module fake_jpeg_18044_n_301 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_301);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_27),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_30),
.Y(n_38)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_0),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_6),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_27),
.Y(n_35)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_17),
.Y(n_45)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_28),
.A2(n_20),
.B1(n_22),
.B2(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_43),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_47),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_48),
.B(n_49),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_27),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_34),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_28),
.A2(n_16),
.B1(n_22),
.B2(n_20),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx24_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_54),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_55),
.A2(n_33),
.B1(n_51),
.B2(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_22),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_61),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_49),
.B(n_22),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_46),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_20),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_41),
.B(n_19),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_47),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_69),
.B(n_46),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_73),
.B(n_75),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_59),
.A2(n_47),
.B1(n_46),
.B2(n_50),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_80),
.A2(n_81),
.B1(n_95),
.B2(n_51),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_59),
.A2(n_43),
.B1(n_52),
.B2(n_40),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_62),
.A2(n_16),
.B1(n_25),
.B2(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_82),
.A2(n_85),
.B1(n_89),
.B2(n_91),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_84),
.B(n_90),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_25),
.B1(n_33),
.B2(n_24),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_31),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_87),
.B(n_74),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_60),
.A2(n_25),
.B1(n_33),
.B2(n_24),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_72),
.B(n_45),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_69),
.A2(n_31),
.B(n_38),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_60),
.A2(n_33),
.B1(n_24),
.B2(n_13),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_51),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_105),
.B1(n_117),
.B2(n_79),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_91),
.B(n_87),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_118),
.Y(n_130)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_111),
.Y(n_138)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_93),
.B(n_19),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_109),
.B(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_19),
.Y(n_110)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_31),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_66),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_112),
.B(n_113),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_73),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_71),
.Y(n_115)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_115),
.Y(n_131)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_19),
.Y(n_119)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_86),
.B(n_21),
.Y(n_121)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_81),
.B1(n_97),
.B2(n_66),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_123),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_100),
.A2(n_94),
.B1(n_29),
.B2(n_30),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_112),
.A2(n_78),
.B1(n_35),
.B2(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_78),
.B1(n_35),
.B2(n_13),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_101),
.C(n_113),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_111),
.C(n_54),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_115),
.B(n_71),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_86),
.B(n_103),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_106),
.A2(n_78),
.B1(n_13),
.B2(n_14),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_137),
.A2(n_140),
.B1(n_117),
.B2(n_23),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_111),
.A2(n_57),
.B1(n_75),
.B2(n_63),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_145),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_116),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_150),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_148),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_132),
.Y(n_150)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_130),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_153),
.B(n_154),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_136),
.Y(n_154)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_159),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_139),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_15),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_133),
.B(n_103),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_173),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_124),
.A2(n_79),
.B1(n_118),
.B2(n_120),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_165),
.B1(n_168),
.B2(n_170),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_53),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_131),
.B(n_54),
.Y(n_164)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_122),
.B1(n_138),
.B2(n_136),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_124),
.B(n_58),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_166),
.B(n_167),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_146),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_142),
.A2(n_125),
.B1(n_129),
.B2(n_135),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_77),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_135),
.A2(n_15),
.B1(n_23),
.B2(n_14),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_129),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_140),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_138),
.B(n_122),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_15),
.B1(n_23),
.B2(n_14),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g173 ( 
.A1(n_126),
.A2(n_1),
.B(n_2),
.Y(n_173)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_176),
.B(n_191),
.C(n_65),
.Y(n_211)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_187),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_58),
.Y(n_187)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_53),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_68),
.Y(n_193)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_193),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_68),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_155),
.A2(n_154),
.B1(n_163),
.B2(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_195),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_120),
.B1(n_118),
.B2(n_1),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_197),
.A2(n_26),
.B1(n_18),
.B2(n_27),
.Y(n_212)
);

INVxp33_ASAP7_75t_L g199 ( 
.A(n_186),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

OAI21xp33_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_153),
.B(n_147),
.Y(n_200)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_188),
.A2(n_156),
.B1(n_173),
.B2(n_151),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_201),
.A2(n_205),
.B1(n_194),
.B2(n_197),
.Y(n_219)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_181),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_185),
.A2(n_182),
.B1(n_179),
.B2(n_183),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_174),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_185),
.A2(n_161),
.B1(n_77),
.B2(n_21),
.Y(n_210)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_217),
.Y(n_236)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_L g215 ( 
.A1(n_196),
.A2(n_77),
.B1(n_65),
.B2(n_1),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_215),
.A2(n_189),
.B1(n_198),
.B2(n_1),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_190),
.Y(n_216)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_216),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_191),
.B(n_9),
.Y(n_217)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_219),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_223),
.B1(n_230),
.B2(n_234),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_208),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_218),
.A2(n_198),
.B1(n_195),
.B2(n_180),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_207),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_180),
.B1(n_176),
.B2(n_2),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_209),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_231),
.A2(n_217),
.B(n_204),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_203),
.B(n_3),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_235),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_214),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_206),
.B(n_4),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g238 ( 
.A(n_223),
.B(n_211),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_238),
.B(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_240),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_236),
.B(n_200),
.C(n_202),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_243),
.C(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_215),
.B1(n_212),
.B2(n_6),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_225),
.B(n_26),
.Y(n_244)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_244),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_21),
.C(n_32),
.Y(n_245)
);

NOR3xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_232),
.C(n_229),
.Y(n_248)
);

BUFx12f_ASAP7_75t_SL g257 ( 
.A(n_248),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_21),
.C(n_32),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_245),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_252),
.B(n_4),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_241),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_254),
.A2(n_259),
.B1(n_249),
.B2(n_5),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_221),
.B1(n_233),
.B2(n_234),
.Y(n_261)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_226),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_251),
.B(n_248),
.Y(n_265)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_264),
.Y(n_271)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_274),
.Y(n_279)
);

FAx1_ASAP7_75t_SL g269 ( 
.A(n_257),
.B(n_5),
.CI(n_7),
.CON(n_269),
.SN(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_269),
.B(n_270),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_32),
.C(n_26),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_255),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_273),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_260),
.B(n_10),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_259),
.A2(n_11),
.B1(n_12),
.B2(n_18),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_275),
.B(n_258),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g276 ( 
.A(n_265),
.B(n_262),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_276),
.A2(n_274),
.B1(n_270),
.B2(n_26),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_266),
.A2(n_256),
.B(n_254),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_283),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_271),
.B(n_267),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_286),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_276),
.A2(n_18),
.B1(n_26),
.B2(n_32),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_290),
.B(n_278),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_18),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_289),
.B(n_280),
.C(n_279),
.Y(n_291)
);

OR2x2_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_282),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_293),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_294),
.A2(n_288),
.B(n_292),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_295),
.Y(n_296)
);

AO21x1_ASAP7_75t_L g297 ( 
.A1(n_296),
.A2(n_32),
.B(n_18),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_298),
.A2(n_18),
.B(n_26),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_32),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_26),
.Y(n_301)
);


endmodule