module fake_ariane_2087_n_800 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_800);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_800;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_584;
wire n_528;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_216;
wire n_540;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_61),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g160 ( 
.A(n_45),
.Y(n_160)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_143),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_51),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_102),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_103),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_154),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_120),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_73),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_4),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_8),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_114),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_13),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_53),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_71),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_7),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_122),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_72),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_6),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_79),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_96),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_60),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_30),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_18),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_129),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_83),
.Y(n_187)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_12),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_113),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_5),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_59),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_148),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_126),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_1),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_115),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_84),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_11),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_107),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_66),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_75),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_141),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_105),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_47),
.Y(n_204)
);

BUFx2_ASAP7_75t_L g205 ( 
.A(n_98),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_16),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_49),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_6),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_23),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_64),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_5),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_112),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_26),
.Y(n_214)
);

OAI21x1_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_77),
.B(n_157),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_163),
.Y(n_216)
);

AND2x4_ASAP7_75t_L g217 ( 
.A(n_163),
.B(n_0),
.Y(n_217)
);

XOR2x2_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_0),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_161),
.B(n_1),
.Y(n_221)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_168),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_178),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_198),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_212),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_172),
.B(n_2),
.Y(n_229)
);

AND2x6_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_200),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_204),
.B(n_2),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

BUFx12f_ASAP7_75t_L g233 ( 
.A(n_162),
.Y(n_233)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_192),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_164),
.B(n_212),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_3),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_185),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_180),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

OAI22x1_ASAP7_75t_R g242 ( 
.A1(n_184),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_9),
.Y(n_243)
);

OAI22x1_ASAP7_75t_R g244 ( 
.A1(n_184),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_244)
);

INVx5_ASAP7_75t_L g245 ( 
.A(n_159),
.Y(n_245)
);

OAI22x1_ASAP7_75t_R g246 ( 
.A1(n_171),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_187),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_193),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_202),
.B(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_180),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_213),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_160),
.Y(n_254)
);

AND2x4_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_15),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_208),
.B(n_16),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_162),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_217),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_251),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_223),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_233),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_233),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_240),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_227),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_227),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_216),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_257),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_235),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_257),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_224),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_216),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_245),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_245),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_245),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_254),
.Y(n_280)
);

BUFx10_ASAP7_75t_L g281 ( 
.A(n_217),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_226),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_254),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_216),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_254),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_254),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_258),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_258),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_216),
.Y(n_289)
);

CKINVDCx6p67_ASAP7_75t_R g290 ( 
.A(n_222),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_220),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_235),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g293 ( 
.A(n_220),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_242),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_225),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_R g297 ( 
.A(n_232),
.B(n_174),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_220),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_222),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_222),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_222),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_225),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_225),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_244),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_237),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_219),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_219),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_268),
.Y(n_308)
);

INVxp67_ASAP7_75t_SL g309 ( 
.A(n_293),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_261),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_221),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_268),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_287),
.B(n_255),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_274),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_293),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_296),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_288),
.B(n_255),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_269),
.B(n_255),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_271),
.B(n_234),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_259),
.Y(n_320)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_298),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_272),
.B(n_234),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_297),
.B(n_221),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_273),
.B(n_229),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_275),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_282),
.Y(n_328)
);

NAND3xp33_ASAP7_75t_L g329 ( 
.A(n_284),
.B(n_249),
.C(n_243),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_259),
.B(n_234),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_266),
.B(n_231),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_239),
.C(n_256),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_296),
.Y(n_333)
);

BUFx6f_ASAP7_75t_SL g334 ( 
.A(n_266),
.Y(n_334)
);

OAI22x1_ASAP7_75t_SL g335 ( 
.A1(n_265),
.A2(n_218),
.B1(n_246),
.B2(n_190),
.Y(n_335)
);

NAND2xp33_ASAP7_75t_L g336 ( 
.A(n_276),
.B(n_256),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_281),
.B(n_248),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_281),
.B(n_165),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_296),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_306),
.B(n_250),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_307),
.B(n_234),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_289),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_260),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_277),
.B(n_166),
.Y(n_344)
);

INVx3_ASAP7_75t_R g345 ( 
.A(n_264),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_305),
.B(n_228),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g347 ( 
.A(n_262),
.B(n_263),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_300),
.Y(n_348)
);

NOR2x1p5_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_175),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_230),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_294),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_301),
.Y(n_354)
);

NAND3xp33_ASAP7_75t_L g355 ( 
.A(n_278),
.B(n_253),
.C(n_252),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_270),
.A2(n_194),
.B1(n_218),
.B2(n_206),
.Y(n_356)
);

BUFx5_ASAP7_75t_L g357 ( 
.A(n_279),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_280),
.Y(n_359)
);

OR2x6_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_228),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_283),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_285),
.B(n_166),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_286),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_267),
.B(n_236),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_304),
.B(n_236),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_297),
.B(n_167),
.Y(n_366)
);

BUFx6f_ASAP7_75t_SL g367 ( 
.A(n_259),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_269),
.B(n_167),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_297),
.B(n_211),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_268),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_261),
.Y(n_371)
);

NAND3xp33_ASAP7_75t_L g372 ( 
.A(n_287),
.B(n_253),
.C(n_252),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_311),
.B(n_211),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_350),
.Y(n_374)
);

BUFx4f_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_325),
.B(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_238),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_313),
.B(n_194),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_360),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_310),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_R g381 ( 
.A(n_334),
.B(n_177),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_337),
.B(n_238),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_313),
.B(n_317),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_318),
.B(n_247),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_357),
.B(n_252),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_308),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_331),
.B(n_247),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_357),
.B(n_252),
.Y(n_389)
);

BUFx2_ASAP7_75t_L g390 ( 
.A(n_360),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_312),
.Y(n_391)
);

NOR3xp33_ASAP7_75t_SL g392 ( 
.A(n_338),
.B(n_199),
.C(n_183),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_253),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_354),
.B(n_253),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_328),
.B(n_371),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_364),
.B(n_241),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_342),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_370),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_357),
.B(n_181),
.Y(n_399)
);

O2A1O1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_336),
.A2(n_197),
.B(n_18),
.C(n_17),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_348),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_357),
.B(n_320),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_352),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_315),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_357),
.B(n_230),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_230),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g410 ( 
.A(n_343),
.B(n_225),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g414 ( 
.A(n_316),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_365),
.B(n_241),
.Y(n_415)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_367),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_L g417 ( 
.A1(n_332),
.A2(n_230),
.B1(n_241),
.B2(n_215),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_L g418 ( 
.A1(n_356),
.A2(n_230),
.B1(n_241),
.B2(n_215),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_309),
.Y(n_419)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_347),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_368),
.A2(n_209),
.B1(n_203),
.B2(n_201),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_367),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_372),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_356),
.A2(n_196),
.B1(n_191),
.B2(n_189),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_316),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_363),
.B(n_17),
.Y(n_426)
);

INVx3_ASAP7_75t_L g427 ( 
.A(n_316),
.Y(n_427)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_372),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_428)
);

BUFx3_ASAP7_75t_L g429 ( 
.A(n_322),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_329),
.A2(n_24),
.B1(n_25),
.B2(n_27),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_329),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_359),
.B(n_158),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_361),
.B(n_28),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_330),
.B(n_29),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_319),
.A2(n_31),
.B(n_32),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_355),
.B(n_358),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_323),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_349),
.Y(n_439)
);

BUFx8_ASAP7_75t_L g440 ( 
.A(n_345),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_SL g441 ( 
.A(n_366),
.B(n_33),
.C(n_34),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_323),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_376),
.A2(n_362),
.B1(n_344),
.B2(n_369),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_384),
.B(n_324),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_377),
.B(n_333),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_420),
.B(n_355),
.Y(n_446)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_414),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_333),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g449 ( 
.A1(n_399),
.A2(n_339),
.B(n_333),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_431),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_399),
.A2(n_339),
.B(n_36),
.Y(n_451)
);

OAI22xp33_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_335),
.B1(n_339),
.B2(n_38),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_378),
.B(n_35),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_378),
.B(n_156),
.Y(n_454)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_429),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_376),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_429),
.B(n_41),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_402),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_436),
.B(n_410),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

OAI21x1_ASAP7_75t_L g461 ( 
.A1(n_408),
.A2(n_42),
.B(n_43),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_386),
.A2(n_44),
.B(n_46),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_383),
.Y(n_463)
);

O2A1O1Ixp5_ASAP7_75t_SL g464 ( 
.A1(n_434),
.A2(n_48),
.B(n_50),
.C(n_52),
.Y(n_464)
);

OAI21x1_ASAP7_75t_L g465 ( 
.A1(n_409),
.A2(n_54),
.B(n_55),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_395),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_386),
.A2(n_62),
.B(n_63),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_389),
.A2(n_65),
.B(n_67),
.Y(n_468)
);

A2O1A1Ixp33_ASAP7_75t_L g469 ( 
.A1(n_400),
.A2(n_68),
.B(n_69),
.C(n_70),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_389),
.A2(n_403),
.B(n_412),
.Y(n_470)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_375),
.B(n_74),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_416),
.Y(n_472)
);

OAI21x1_ASAP7_75t_SL g473 ( 
.A1(n_432),
.A2(n_76),
.B(n_78),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_396),
.B(n_80),
.Y(n_474)
);

O2A1O1Ixp33_ASAP7_75t_L g475 ( 
.A1(n_373),
.A2(n_81),
.B(n_82),
.C(n_85),
.Y(n_475)
);

O2A1O1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_373),
.A2(n_86),
.B(n_87),
.C(n_88),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_403),
.A2(n_89),
.B(n_90),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_414),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_385),
.B(n_91),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_404),
.B(n_92),
.Y(n_480)
);

NOR2x1_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_93),
.Y(n_481)
);

OAI21xp33_ASAP7_75t_SL g482 ( 
.A1(n_397),
.A2(n_94),
.B(n_95),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_413),
.A2(n_433),
.B(n_438),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_442),
.A2(n_97),
.B(n_99),
.Y(n_484)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_393),
.A2(n_100),
.B(n_101),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_375),
.B(n_104),
.Y(n_486)
);

BUFx3_ASAP7_75t_L g487 ( 
.A(n_440),
.Y(n_487)
);

A2O1A1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_388),
.A2(n_106),
.B(n_108),
.C(n_109),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_374),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_424),
.A2(n_111),
.B1(n_116),
.B2(n_117),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_424),
.A2(n_118),
.B1(n_119),
.B2(n_121),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_418),
.A2(n_123),
.B1(n_125),
.B2(n_127),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_388),
.B(n_128),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_405),
.Y(n_494)
);

AO22x1_ASAP7_75t_L g495 ( 
.A1(n_440),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_495)
);

NOR3xp33_ASAP7_75t_L g496 ( 
.A(n_426),
.B(n_439),
.C(n_404),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_418),
.A2(n_401),
.B1(n_423),
.B2(n_430),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g498 ( 
.A(n_419),
.B(n_133),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_390),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_425),
.A2(n_137),
.B(n_138),
.Y(n_500)
);

OAI21x1_ASAP7_75t_L g501 ( 
.A1(n_470),
.A2(n_434),
.B(n_417),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_478),
.Y(n_502)
);

AO21x2_ASAP7_75t_L g503 ( 
.A1(n_497),
.A2(n_394),
.B(n_435),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_460),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_458),
.Y(n_505)
);

AOI22xp33_ASAP7_75t_SL g506 ( 
.A1(n_453),
.A2(n_379),
.B1(n_381),
.B2(n_415),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_489),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_446),
.B(n_422),
.Y(n_508)
);

OAI21x1_ASAP7_75t_L g509 ( 
.A1(n_461),
.A2(n_417),
.B(n_430),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_444),
.A2(n_391),
.B(n_398),
.Y(n_510)
);

AO21x2_ASAP7_75t_L g511 ( 
.A1(n_483),
.A2(n_493),
.B(n_449),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_463),
.Y(n_513)
);

OAI21x1_ASAP7_75t_L g514 ( 
.A1(n_464),
.A2(n_428),
.B(n_427),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_450),
.B(n_387),
.Y(n_515)
);

AO21x2_ASAP7_75t_L g516 ( 
.A1(n_451),
.A2(n_394),
.B(n_407),
.Y(n_516)
);

OAI21x1_ASAP7_75t_L g517 ( 
.A1(n_465),
.A2(n_428),
.B(n_427),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_473),
.A2(n_406),
.B(n_422),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_477),
.A2(n_406),
.B(n_421),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_494),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_479),
.A2(n_414),
.B(n_437),
.Y(n_521)
);

INVx6_ASAP7_75t_SL g522 ( 
.A(n_457),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_447),
.Y(n_524)
);

NOR2x1_ASAP7_75t_L g525 ( 
.A(n_487),
.B(n_414),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_474),
.A2(n_437),
.B(n_441),
.Y(n_526)
);

NAND2x1p5_ASAP7_75t_L g527 ( 
.A(n_455),
.B(n_437),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_447),
.Y(n_528)
);

OAI21x1_ASAP7_75t_L g529 ( 
.A1(n_492),
.A2(n_437),
.B(n_392),
.Y(n_529)
);

OR2x6_ASAP7_75t_L g530 ( 
.A(n_471),
.B(n_381),
.Y(n_530)
);

OAI21x1_ASAP7_75t_L g531 ( 
.A1(n_485),
.A2(n_498),
.B(n_468),
.Y(n_531)
);

BUFx2_ASAP7_75t_L g532 ( 
.A(n_455),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_478),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

BUFx2_ASAP7_75t_L g535 ( 
.A(n_472),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_454),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_478),
.Y(n_537)
);

BUFx12f_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

CKINVDCx14_ASAP7_75t_R g539 ( 
.A(n_480),
.Y(n_539)
);

OAI21x1_ASAP7_75t_L g540 ( 
.A1(n_462),
.A2(n_467),
.B(n_484),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_486),
.B(n_139),
.Y(n_541)
);

CKINVDCx16_ASAP7_75t_R g542 ( 
.A(n_490),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_499),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_445),
.Y(n_544)
);

INVx2_ASAP7_75t_SL g545 ( 
.A(n_481),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_443),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_459),
.Y(n_547)
);

AND2x4_ASAP7_75t_L g548 ( 
.A(n_496),
.B(n_140),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g549 ( 
.A(n_495),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_456),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_518),
.A2(n_476),
.B(n_475),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_491),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_469),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_512),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_518),
.A2(n_500),
.B(n_466),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_546),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_507),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_546),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g559 ( 
.A(n_505),
.B(n_452),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_502),
.Y(n_560)
);

AO21x1_ASAP7_75t_SL g561 ( 
.A1(n_523),
.A2(n_482),
.B(n_488),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_504),
.Y(n_562)
);

INVx3_ASAP7_75t_L g563 ( 
.A(n_533),
.Y(n_563)
);

BUFx4f_ASAP7_75t_L g564 ( 
.A(n_512),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_533),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_513),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_520),
.Y(n_567)
);

OAI21x1_ASAP7_75t_SL g568 ( 
.A1(n_550),
.A2(n_142),
.B(n_144),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_515),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_515),
.Y(n_570)
);

CKINVDCx11_ASAP7_75t_R g571 ( 
.A(n_538),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_543),
.B(n_155),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_538),
.Y(n_573)
);

BUFx2_ASAP7_75t_L g574 ( 
.A(n_522),
.Y(n_574)
);

INVx3_ASAP7_75t_L g575 ( 
.A(n_502),
.Y(n_575)
);

BUFx10_ASAP7_75t_L g576 ( 
.A(n_548),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_542),
.A2(n_146),
.B1(n_147),
.B2(n_149),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_522),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_510),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_508),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_534),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_536),
.A2(n_548),
.B1(n_549),
.B2(n_541),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_547),
.Y(n_583)
);

AOI22xp33_ASAP7_75t_L g584 ( 
.A1(n_536),
.A2(n_548),
.B1(n_541),
.B2(n_506),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_541),
.A2(n_530),
.B1(n_522),
.B2(n_550),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_539),
.A2(n_530),
.B1(n_547),
.B2(n_545),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_530),
.A2(n_532),
.B1(n_544),
.B2(n_527),
.Y(n_588)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_502),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_535),
.B(n_544),
.Y(n_591)
);

BUFx2_ASAP7_75t_L g592 ( 
.A(n_533),
.Y(n_592)
);

INVx6_ASAP7_75t_L g593 ( 
.A(n_533),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_501),
.A2(n_526),
.B(n_519),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_537),
.Y(n_595)
);

AND2x2_ASAP7_75t_SL g596 ( 
.A(n_584),
.B(n_537),
.Y(n_596)
);

BUFx3_ASAP7_75t_L g597 ( 
.A(n_573),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_567),
.Y(n_598)
);

OAI222xp33_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_539),
.B1(n_545),
.B2(n_544),
.C1(n_528),
.C2(n_525),
.Y(n_599)
);

CKINVDCx8_ASAP7_75t_R g600 ( 
.A(n_554),
.Y(n_600)
);

AOI22xp33_ASAP7_75t_SL g601 ( 
.A1(n_552),
.A2(n_509),
.B1(n_503),
.B2(n_501),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_556),
.B(n_528),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_556),
.B(n_537),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_557),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_558),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_571),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_571),
.Y(n_607)
);

AO32x2_ASAP7_75t_L g608 ( 
.A1(n_588),
.A2(n_503),
.A3(n_516),
.B1(n_509),
.B2(n_511),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_558),
.B(n_537),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_562),
.Y(n_610)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_554),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_573),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_R g613 ( 
.A(n_564),
.B(n_527),
.Y(n_613)
);

AND2x2_ASAP7_75t_L g614 ( 
.A(n_572),
.B(n_529),
.Y(n_614)
);

O2A1O1Ixp33_ASAP7_75t_SL g615 ( 
.A1(n_577),
.A2(n_521),
.B(n_526),
.C(n_529),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_564),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_566),
.Y(n_617)
);

CKINVDCx11_ASAP7_75t_R g618 ( 
.A(n_576),
.Y(n_618)
);

OR2x6_ASAP7_75t_L g619 ( 
.A(n_553),
.B(n_519),
.Y(n_619)
);

OAI22xp5_ASAP7_75t_L g620 ( 
.A1(n_584),
.A2(n_559),
.B1(n_585),
.B2(n_553),
.Y(n_620)
);

NOR3xp33_ASAP7_75t_SL g621 ( 
.A(n_591),
.B(n_531),
.C(n_540),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_581),
.Y(n_622)
);

NOR2x1p5_ASAP7_75t_L g623 ( 
.A(n_560),
.B(n_575),
.Y(n_623)
);

INVx3_ASAP7_75t_SL g624 ( 
.A(n_593),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_R g625 ( 
.A(n_576),
.B(n_503),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_555),
.A2(n_517),
.B(n_540),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_569),
.B(n_514),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_570),
.B(n_516),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_574),
.Y(n_629)
);

AOI22xp33_ASAP7_75t_L g630 ( 
.A1(n_576),
.A2(n_516),
.B1(n_514),
.B2(n_511),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_583),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_578),
.B(n_517),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_587),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_586),
.B(n_511),
.Y(n_634)
);

OAI21x1_ASAP7_75t_L g635 ( 
.A1(n_555),
.A2(n_531),
.B(n_551),
.Y(n_635)
);

AOI22xp33_ASAP7_75t_SL g636 ( 
.A1(n_553),
.A2(n_568),
.B1(n_579),
.B2(n_585),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_592),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_560),
.B(n_575),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_589),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_590),
.B(n_595),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_593),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_593),
.Y(n_642)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_580),
.A2(n_589),
.B1(n_563),
.B2(n_565),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_618),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_604),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_639),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_619),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_SL g648 ( 
.A(n_613),
.B(n_563),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_605),
.B(n_594),
.Y(n_649)
);

OR2x2_ASAP7_75t_L g650 ( 
.A(n_605),
.B(n_563),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_602),
.B(n_565),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_622),
.B(n_565),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_631),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_628),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_601),
.B(n_627),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_634),
.B(n_551),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_601),
.B(n_561),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_610),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_633),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_617),
.B(n_619),
.Y(n_660)
);

INVxp67_ASAP7_75t_L g661 ( 
.A(n_609),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_606),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_619),
.Y(n_663)
);

AO21x2_ASAP7_75t_L g664 ( 
.A1(n_625),
.A2(n_589),
.B(n_621),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_598),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_632),
.B(n_614),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_603),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_608),
.B(n_625),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_608),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_608),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_640),
.B(n_638),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_620),
.B(n_630),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_621),
.B(n_596),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_635),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_596),
.B(n_630),
.Y(n_676)
);

CKINVDCx11_ASAP7_75t_R g677 ( 
.A(n_600),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_638),
.B(n_642),
.Y(n_678)
);

INVx4_ASAP7_75t_L g679 ( 
.A(n_639),
.Y(n_679)
);

AND2x4_ASAP7_75t_L g680 ( 
.A(n_623),
.B(n_639),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_626),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_636),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_658),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_658),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_653),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_659),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_666),
.B(n_636),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_667),
.B(n_597),
.Y(n_688)
);

HB1xp67_ASAP7_75t_L g689 ( 
.A(n_650),
.Y(n_689)
);

AND2x2_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_655),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_663),
.B(n_597),
.Y(n_691)
);

INVxp67_ASAP7_75t_SL g692 ( 
.A(n_656),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_659),
.Y(n_693)
);

OR2x2_ASAP7_75t_L g694 ( 
.A(n_661),
.B(n_641),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_655),
.B(n_624),
.Y(n_695)
);

OR2x2_ASAP7_75t_L g696 ( 
.A(n_650),
.B(n_624),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_653),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_665),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_672),
.B(n_639),
.Y(n_699)
);

AND2x4_ASAP7_75t_L g700 ( 
.A(n_663),
.B(n_637),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_651),
.B(n_643),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_673),
.B(n_607),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_665),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_649),
.B(n_611),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_649),
.B(n_611),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_652),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_678),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_647),
.B(n_612),
.Y(n_708)
);

AND2x2_ASAP7_75t_L g709 ( 
.A(n_660),
.B(n_629),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_654),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_660),
.B(n_616),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_646),
.Y(n_712)
);

OAI22xp5_ASAP7_75t_L g713 ( 
.A1(n_682),
.A2(n_657),
.B1(n_673),
.B2(n_674),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_654),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_645),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_682),
.B(n_615),
.C(n_599),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_710),
.Y(n_717)
);

OR2x2_ASAP7_75t_L g718 ( 
.A(n_690),
.B(n_656),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_706),
.B(n_692),
.Y(n_719)
);

BUFx2_ASAP7_75t_L g720 ( 
.A(n_708),
.Y(n_720)
);

OAI33xp33_ASAP7_75t_L g721 ( 
.A1(n_713),
.A2(n_671),
.A3(n_670),
.B1(n_669),
.B2(n_675),
.B3(n_681),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_689),
.B(n_670),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_686),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_714),
.Y(n_724)
);

OR2x2_ASAP7_75t_L g725 ( 
.A(n_690),
.B(n_647),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_689),
.B(n_647),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_683),
.Y(n_727)
);

NAND4xp25_ASAP7_75t_L g728 ( 
.A(n_702),
.B(n_644),
.C(n_657),
.D(n_675),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_684),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_685),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_686),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_693),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_704),
.B(n_644),
.Y(n_733)
);

OR2x2_ASAP7_75t_L g734 ( 
.A(n_695),
.B(n_671),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_669),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_719),
.B(n_687),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_720),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_727),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_718),
.B(n_696),
.Y(n_739)
);

OAI211xp5_ASAP7_75t_L g740 ( 
.A1(n_728),
.A2(n_716),
.B(n_704),
.C(n_705),
.Y(n_740)
);

OAI32xp33_ASAP7_75t_L g741 ( 
.A1(n_728),
.A2(n_674),
.A3(n_701),
.B1(n_695),
.B2(n_688),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_719),
.Y(n_742)
);

OAI22xp33_ASAP7_75t_L g743 ( 
.A1(n_735),
.A2(n_668),
.B1(n_676),
.B2(n_699),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_735),
.B(n_694),
.Y(n_744)
);

OR2x2_ASAP7_75t_L g745 ( 
.A(n_734),
.B(n_705),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_723),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_733),
.B(n_700),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_731),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_742),
.B(n_717),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_747),
.B(n_709),
.Y(n_750)
);

INVx3_ASAP7_75t_L g751 ( 
.A(n_739),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_745),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_740),
.A2(n_707),
.B1(n_700),
.B2(n_725),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_736),
.B(n_722),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_738),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_755),
.Y(n_756)
);

INVxp67_ASAP7_75t_SL g757 ( 
.A(n_753),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_751),
.B(n_737),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_751),
.B(n_736),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_752),
.B(n_753),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_756),
.Y(n_761)
);

AOI221xp5_ASAP7_75t_L g762 ( 
.A1(n_757),
.A2(n_741),
.B1(n_743),
.B2(n_721),
.C(n_740),
.Y(n_762)
);

AOI211xp5_ASAP7_75t_L g763 ( 
.A1(n_760),
.A2(n_754),
.B(n_700),
.C(n_708),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_759),
.B(n_749),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_761),
.Y(n_765)
);

NOR3xp33_ASAP7_75t_L g766 ( 
.A(n_762),
.B(n_760),
.C(n_644),
.Y(n_766)
);

OAI22xp5_ASAP7_75t_L g767 ( 
.A1(n_763),
.A2(n_758),
.B1(n_750),
.B2(n_644),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_765),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_767),
.Y(n_769)
);

XOR2x2_ASAP7_75t_L g770 ( 
.A(n_766),
.B(n_764),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_768),
.B(n_662),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_770),
.A2(n_758),
.B1(n_664),
.B2(n_668),
.Y(n_772)
);

AO22x2_ASAP7_75t_L g773 ( 
.A1(n_769),
.A2(n_709),
.B1(n_711),
.B2(n_708),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_768),
.B(n_677),
.Y(n_774)
);

NAND4xp25_ASAP7_75t_SL g775 ( 
.A(n_769),
.B(n_711),
.C(n_722),
.D(n_726),
.Y(n_775)
);

NOR2x1_ASAP7_75t_L g776 ( 
.A(n_774),
.B(n_724),
.Y(n_776)
);

NAND4xp75_ASAP7_75t_L g777 ( 
.A(n_772),
.B(n_613),
.C(n_730),
.D(n_729),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_771),
.B(n_599),
.C(n_648),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_773),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_775),
.A2(n_712),
.B(n_680),
.Y(n_780)
);

OAI211xp5_ASAP7_75t_SL g781 ( 
.A1(n_774),
.A2(n_712),
.B(n_615),
.C(n_744),
.Y(n_781)
);

CKINVDCx6p67_ASAP7_75t_R g782 ( 
.A(n_779),
.Y(n_782)
);

OAI322xp33_ASAP7_75t_L g783 ( 
.A1(n_776),
.A2(n_679),
.A3(n_748),
.B1(n_746),
.B2(n_697),
.C1(n_681),
.C2(n_646),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_777),
.Y(n_784)
);

OAI211xp5_ASAP7_75t_SL g785 ( 
.A1(n_780),
.A2(n_703),
.B(n_698),
.C(n_732),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_778),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_782),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_786),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_784),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_785),
.A2(n_781),
.B1(n_680),
.B2(n_664),
.Y(n_790)
);

OAI31xp33_ASAP7_75t_L g791 ( 
.A1(n_788),
.A2(n_783),
.A3(n_691),
.B(n_676),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_787),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_789),
.B(n_691),
.Y(n_793)
);

HB1xp67_ASAP7_75t_L g794 ( 
.A(n_792),
.Y(n_794)
);

INVx3_ASAP7_75t_L g795 ( 
.A(n_793),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_794),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_796),
.B(n_795),
.Y(n_797)
);

AOI222xp33_ASAP7_75t_L g798 ( 
.A1(n_797),
.A2(n_791),
.B1(n_790),
.B2(n_691),
.C1(n_680),
.C2(n_715),
.Y(n_798)
);

AOI221xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_646),
.B1(n_680),
.B2(n_679),
.C(n_664),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_799),
.A2(n_679),
.B1(n_646),
.B2(n_693),
.Y(n_800)
);


endmodule