module fake_jpeg_30589_n_434 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_434);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_434;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx11_ASAP7_75t_SL g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_8),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_6),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_6),
.B(n_11),
.Y(n_43)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_8),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_11),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_15),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_48),
.B(n_59),
.Y(n_112)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_49),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_50),
.Y(n_117)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_15),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_53),
.B(n_57),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_54),
.Y(n_124)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx5_ASAP7_75t_SL g143 ( 
.A(n_55),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_56),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_16),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_15),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_63),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_16),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_64),
.B(n_66),
.Y(n_125)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_24),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_67),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g108 ( 
.A(n_70),
.Y(n_108)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

BUFx10_ASAP7_75t_L g113 ( 
.A(n_71),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_72),
.B(n_74),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_14),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_73),
.B(n_44),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_18),
.Y(n_74)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_24),
.Y(n_78)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_81),
.Y(n_153)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_86),
.Y(n_138)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_87),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_33),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_88),
.B(n_94),
.Y(n_141)
);

BUFx5_ASAP7_75t_L g89 ( 
.A(n_17),
.Y(n_89)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_89),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_22),
.Y(n_90)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_29),
.Y(n_91)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_93),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_31),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_96),
.B(n_97),
.Y(n_105)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_84),
.A2(n_19),
.B1(n_37),
.B2(n_35),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_98),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_19),
.B1(n_37),
.B2(n_35),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_90),
.A2(n_45),
.B1(n_26),
.B2(n_21),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_45),
.B1(n_26),
.B2(n_21),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_44),
.B1(n_17),
.B2(n_39),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_115),
.A2(n_78),
.B1(n_65),
.B2(n_80),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_71),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_126),
.B(n_142),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_39),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_130),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_40),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_60),
.B(n_40),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_33),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_82),
.B(n_36),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_62),
.B(n_34),
.C(n_30),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_144),
.A2(n_87),
.B(n_69),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_33),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_67),
.A2(n_30),
.B1(n_34),
.B2(n_44),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_146),
.A2(n_68),
.B1(n_49),
.B2(n_77),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_52),
.A2(n_17),
.B1(n_33),
.B2(n_41),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_150),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_141),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_154),
.B(n_159),
.Y(n_206)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_155),
.Y(n_208)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

INVx6_ASAP7_75t_L g205 ( 
.A(n_157),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_113),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_160),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_133),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_161),
.B(n_167),
.Y(n_210)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_162),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_163),
.A2(n_197),
.B1(n_70),
.B2(n_107),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_125),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_164),
.B(n_179),
.Y(n_225)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_168),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_183),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_143),
.A2(n_55),
.B1(n_95),
.B2(n_58),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_171),
.Y(n_229)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_129),
.Y(n_172)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_172),
.Y(n_236)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_99),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_173),
.Y(n_219)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_136),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_175),
.B(n_181),
.Y(n_227)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_99),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_176),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_182),
.B1(n_132),
.B2(n_124),
.Y(n_224)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

OR2x2_ASAP7_75t_SL g180 ( 
.A(n_112),
.B(n_145),
.Y(n_180)
);

NOR3xp33_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_184),
.C(n_189),
.Y(n_234)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_101),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g182 ( 
.A1(n_100),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_101),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_116),
.B(n_82),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_186),
.B(n_187),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_50),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_144),
.A2(n_83),
.B(n_71),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_188),
.A2(n_149),
.B(n_120),
.Y(n_221)
);

INVx3_ASAP7_75t_SL g189 ( 
.A(n_114),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_112),
.B(n_102),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_190),
.B(n_191),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_127),
.B(n_75),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_151),
.B(n_41),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_192),
.B(n_193),
.Y(n_215)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_134),
.B(n_83),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_195),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_150),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_108),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_196),
.A2(n_198),
.B1(n_107),
.B2(n_152),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_143),
.A2(n_76),
.B1(n_81),
.B2(n_92),
.Y(n_197)
);

BUFx24_ASAP7_75t_L g198 ( 
.A(n_108),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_103),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_199),
.B(n_200),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_151),
.B(n_41),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_103),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_135),
.Y(n_237)
);

OAI22x1_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_115),
.B1(n_153),
.B2(n_120),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_SL g245 ( 
.A1(n_204),
.A2(n_182),
.B(n_187),
.C(n_177),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_209),
.Y(n_270)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_174),
.A2(n_147),
.B(n_138),
.C(n_71),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_214),
.A2(n_221),
.B(n_217),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_216),
.A2(n_111),
.B1(n_135),
.B2(n_113),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_168),
.A2(n_117),
.B1(n_119),
.B2(n_118),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_222),
.B1(n_239),
.B2(n_161),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_118),
.B1(n_114),
.B2(n_119),
.Y(n_222)
);

MAJx2_ASAP7_75t_L g223 ( 
.A(n_169),
.B(n_188),
.C(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_235),
.C(n_172),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_231),
.B1(n_202),
.B2(n_209),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_178),
.A2(n_132),
.B1(n_124),
.B2(n_91),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_180),
.B(n_194),
.C(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_237),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_156),
.A2(n_149),
.B(n_83),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_189),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_195),
.A2(n_93),
.B1(n_96),
.B2(n_153),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_230),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_241),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_206),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_225),
.B(n_154),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_242),
.B(n_249),
.Y(n_285)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_208),
.Y(n_244)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_245),
.A2(n_263),
.B1(n_224),
.B2(n_217),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_232),
.A2(n_179),
.B1(n_162),
.B2(n_171),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_248),
.A2(n_264),
.B1(n_229),
.B2(n_212),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_207),
.B(n_166),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_250),
.B(n_253),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_207),
.B(n_159),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_254),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_252),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_193),
.C(n_181),
.Y(n_253)
);

AOI32xp33_ASAP7_75t_L g254 ( 
.A1(n_204),
.A2(n_189),
.A3(n_165),
.B1(n_175),
.B2(n_198),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_198),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_256),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_185),
.C(n_176),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_213),
.B(n_173),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_257),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_218),
.B(n_201),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_260),
.Y(n_283)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_237),
.Y(n_259)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_199),
.C(n_158),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_227),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_233),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_218),
.A2(n_157),
.B1(n_153),
.B2(n_198),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_262),
.A2(n_266),
.B1(n_267),
.B2(n_239),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_202),
.A2(n_111),
.B1(n_79),
.B2(n_2),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_228),
.Y(n_265)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_265),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_231),
.A2(n_33),
.B1(n_135),
.B2(n_113),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_210),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_268),
.A2(n_271),
.B(n_210),
.Y(n_288)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_228),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_211),
.B1(n_203),
.B2(n_229),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_272),
.A2(n_276),
.B1(n_279),
.B2(n_284),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_274),
.A2(n_278),
.B1(n_281),
.B2(n_289),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_243),
.A2(n_214),
.B1(n_215),
.B2(n_234),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_245),
.A2(n_210),
.B1(n_238),
.B2(n_203),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_243),
.A2(n_215),
.B1(n_233),
.B2(n_213),
.Y(n_284)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_287),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_292),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_245),
.A2(n_219),
.B1(n_212),
.B2(n_226),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_236),
.B1(n_226),
.B2(n_211),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_290),
.A2(n_299),
.B1(n_247),
.B2(n_244),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_260),
.A2(n_236),
.B(n_160),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g293 ( 
.A1(n_270),
.A2(n_160),
.B(n_205),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_297),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_270),
.A2(n_271),
.B(n_268),
.Y(n_297)
);

OAI32xp33_ASAP7_75t_L g298 ( 
.A1(n_245),
.A2(n_160),
.A3(n_205),
.B1(n_2),
.B2(n_3),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_245),
.A2(n_41),
.B1(n_1),
.B2(n_3),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_285),
.B(n_250),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_302),
.B(n_310),
.Y(n_339)
);

AOI22x1_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_263),
.B1(n_252),
.B2(n_240),
.Y(n_303)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_303),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_253),
.C(n_255),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_305),
.B(n_312),
.C(n_282),
.Y(n_338)
);

MAJx2_ASAP7_75t_L g306 ( 
.A(n_288),
.B(n_256),
.C(n_258),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_305),
.Y(n_332)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_309),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_277),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_248),
.C(n_265),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_277),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_321),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_272),
.A2(n_246),
.B1(n_264),
.B2(n_269),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_314),
.A2(n_327),
.B(n_292),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_0),
.Y(n_315)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_315),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_1),
.Y(n_316)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

OA22x2_ASAP7_75t_SL g317 ( 
.A1(n_289),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_273),
.Y(n_318)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_318),
.Y(n_342)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_273),
.Y(n_319)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_319),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_274),
.A2(n_275),
.B1(n_294),
.B2(n_281),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_299),
.A2(n_294),
.B1(n_276),
.B2(n_279),
.Y(n_321)
);

OA21x2_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_4),
.B(n_5),
.Y(n_322)
);

OA21x2_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_301),
.B(n_317),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_287),
.B(n_41),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_324),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_290),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_280),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_326),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_284),
.A2(n_283),
.B1(n_296),
.B2(n_291),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_322),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g370 ( 
.A(n_331),
.B(n_334),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_332),
.B(n_308),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_322),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_337),
.B(n_340),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_346),
.C(n_347),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_327),
.B(n_282),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_L g341 ( 
.A1(n_307),
.A2(n_293),
.B(n_283),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_341),
.A2(n_350),
.B(n_325),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_303),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_312),
.B(n_280),
.C(n_300),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_306),
.B(n_300),
.C(n_285),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_311),
.B(n_278),
.C(n_5),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_349),
.B(n_321),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_325),
.A2(n_4),
.B(n_7),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_339),
.Y(n_352)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_352),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_354),
.B(n_360),
.Y(n_372)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_342),
.Y(n_355)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_355),
.Y(n_375)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_342),
.Y(n_356)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

BUFx24_ASAP7_75t_SL g357 ( 
.A(n_330),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_357),
.B(n_363),
.Y(n_381)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_358),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_332),
.B(n_311),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_364),
.Y(n_373)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_335),
.Y(n_361)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_361),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g386 ( 
.A(n_362),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_308),
.Y(n_364)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_340),
.B(n_304),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_367),
.A2(n_341),
.B(n_333),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_348),
.A2(n_307),
.B1(n_314),
.B2(n_303),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_368),
.A2(n_369),
.B1(n_371),
.B2(n_309),
.Y(n_379)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_343),
.Y(n_369)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_376),
.B(n_364),
.Y(n_399)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_379),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_368),
.A2(n_329),
.B1(n_328),
.B2(n_351),
.Y(n_382)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_362),
.A2(n_370),
.B(n_328),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_383),
.A2(n_344),
.B(n_349),
.Y(n_392)
);

NOR3xp33_ASAP7_75t_SL g384 ( 
.A(n_360),
.B(n_336),
.C(n_350),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_384),
.B(n_334),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_367),
.A2(n_329),
.B1(n_351),
.B2(n_331),
.Y(n_387)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_345),
.Y(n_388)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_388),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_389),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_337),
.B(n_353),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g410 ( 
.A1(n_390),
.A2(n_392),
.B(n_376),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_374),
.B(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_391),
.B(n_395),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_386),
.B(n_354),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_387),
.A2(n_347),
.B1(n_353),
.B2(n_365),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_396),
.B(n_399),
.Y(n_402)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_377),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_380),
.Y(n_404)
);

A2O1A1Ixp33_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_317),
.B(n_315),
.C(n_316),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_400),
.B(n_379),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_401),
.B(n_403),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_365),
.C(n_373),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_404),
.B(n_406),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_393),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_396),
.B(n_381),
.Y(n_408)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_408),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_SL g413 ( 
.A1(n_410),
.A2(n_390),
.B(n_400),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_402),
.B(n_373),
.C(n_395),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_411),
.B(n_416),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_405),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_412),
.B(n_378),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_413),
.A2(n_414),
.B(n_392),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_409),
.A2(n_394),
.B(n_385),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_401),
.Y(n_416)
);

OAI21x1_ASAP7_75t_L g427 ( 
.A1(n_420),
.A2(n_422),
.B(n_319),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_415),
.B(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g428 ( 
.A(n_421),
.B(n_423),
.C(n_372),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_412),
.A2(n_410),
.B1(n_402),
.B2(n_382),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g424 ( 
.A1(n_417),
.A2(n_418),
.B(n_346),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_424),
.A2(n_372),
.B(n_359),
.Y(n_426)
);

NOR2xp67_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_384),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g430 ( 
.A(n_425),
.B(n_427),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_426),
.B(n_428),
.C(n_7),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_429),
.B(n_13),
.C(n_9),
.Y(n_431)
);

O2A1O1Ixp33_ASAP7_75t_SL g432 ( 
.A1(n_431),
.A2(n_430),
.B(n_9),
.C(n_11),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_8),
.B(n_9),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_12),
.B1(n_13),
.B2(n_432),
.Y(n_434)
);


endmodule