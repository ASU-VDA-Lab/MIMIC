module real_jpeg_27902_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_0),
.A2(n_25),
.B1(n_29),
.B2(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_0),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_62),
.B1(n_63),
.B2(n_71),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_1),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_71),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_1),
.A2(n_25),
.B1(n_29),
.B2(n_71),
.Y(n_167)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_2),
.A2(n_103),
.B(n_116),
.Y(n_115)
);

INVx5_ASAP7_75t_L g183 ( 
.A(n_2),
.Y(n_183)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_4),
.A2(n_74),
.B1(n_75),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_4),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_4),
.A2(n_62),
.B1(n_63),
.B2(n_83),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_83),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_83),
.Y(n_182)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_6),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_6),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_55),
.Y(n_126)
);

INVx13_ASAP7_75t_L g75 ( 
.A(n_7),
.Y(n_75)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_8),
.A2(n_11),
.B(n_25),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_9),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_103)
);

OAI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_10),
.A2(n_32),
.B1(n_33),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_10),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_41),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_11),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_11),
.B(n_62),
.Y(n_130)
);

AOI21xp33_ASAP7_75t_L g134 ( 
.A1(n_11),
.A2(n_62),
.B(n_130),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_76),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_11),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_182),
.Y(n_185)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_12),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_13),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_61)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_13),
.Y(n_67)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_15),
.A2(n_69),
.B1(n_74),
.B2(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_69),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_15),
.A2(n_25),
.B1(n_29),
.B2(n_69),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_117),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_19),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_104),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_104),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_84),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_50),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_42),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_31),
.B(n_36),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_39),
.Y(n_38)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_24),
.A2(n_38),
.B1(n_137),
.B2(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_24),
.A2(n_38),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_24),
.A2(n_38),
.B1(n_137),
.B2(n_156),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_24),
.B(n_76),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_24)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_25),
.B(n_44),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp33_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_39)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_28),
.A2(n_33),
.B(n_76),
.C(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_29),
.B(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_32),
.A2(n_33),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_32),
.A2(n_63),
.A3(n_129),
.B1(n_130),
.B2(n_131),
.Y(n_128)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g131 ( 
.A(n_33),
.B(n_66),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_38),
.A2(n_53),
.B(n_56),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_38),
.A2(n_138),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_57),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B(n_47),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_43),
.A2(n_44),
.B1(n_45),
.B2(n_102),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_43),
.B(n_49),
.Y(n_116)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_43),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_43),
.A2(n_167),
.B(n_168),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_43),
.A2(n_174),
.B1(n_182),
.B2(n_183),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_49),
.Y(n_48)
);

INVx11_ASAP7_75t_L g169 ( 
.A(n_44),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_44),
.B(n_76),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_48),
.A2(n_126),
.B(n_127),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_58),
.C(n_72),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_52),
.B1(n_58),
.B2(n_59),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_54),
.B(n_57),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_65),
.B1(n_68),
.B2(n_70),
.Y(n_59)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_60),
.A2(n_65),
.B1(n_68),
.B2(n_112),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_60),
.A2(n_65),
.B1(n_112),
.B2(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_62),
.A2(n_63),
.B1(n_78),
.B2(n_79),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_78),
.Y(n_100)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_63),
.A2(n_73),
.B1(n_80),
.B2(n_100),
.Y(n_99)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_65),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_65),
.Y(n_163)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_72),
.B(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_77),
.B1(n_81),
.B2(n_82),
.Y(n_72)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_76),
.CON(n_73),
.SN(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_74),
.A2(n_78),
.B(n_80),
.C(n_81),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_78),
.Y(n_80)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_76),
.B(n_91),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_82),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_98),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_95),
.B(n_96),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_101),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_99),
.B(n_101),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_108),
.C(n_110),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_105),
.A2(n_106),
.B1(n_201),
.B2(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_113),
.C(n_114),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_111),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_114),
.B1(n_115),
.B2(n_143),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_113),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_198),
.B(n_204),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_149),
.B(n_197),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_139),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_122),
.B(n_139),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_132),
.C(n_135),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_123),
.A2(n_124),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_125),
.B(n_128),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_169),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_127),
.A2(n_169),
.B1(n_173),
.B2(n_175),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_140),
.B(n_146),
.C(n_147),
.Y(n_199)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_191),
.B(n_196),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_170),
.B(n_190),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_159),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_152),
.B(n_159),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_157),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_177),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_166),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_165),
.C(n_166),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_167),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_178),
.B(n_189),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_172),
.B(n_176),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_188),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_181),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_193),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_192),
.B(n_193),
.Y(n_196)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_199),
.B(n_200),
.Y(n_204)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_201),
.Y(n_203)
);


endmodule