module real_aes_11045_n_361 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_350, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_361);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_361;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1744;
wire n_1730;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1940;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_1951;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_1614;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1985;
wire n_1769;
wire n_1812;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_1971;
wire n_731;
wire n_964;
wire n_600;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_365;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_1172;
wire n_459;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_374;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1411;
wire n_1263;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_367;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1986;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1056;
wire n_1592;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1931;
wire n_1721;
wire n_1176;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_362;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_1049;
wire n_1277;
wire n_559;
wire n_1950;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1925;
wire n_1801;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g818 ( .A(n_0), .B(n_819), .Y(n_818) );
CKINVDCx5p33_ASAP7_75t_R g950 ( .A(n_1), .Y(n_950) );
CKINVDCx5p33_ASAP7_75t_R g1473 ( .A(n_2), .Y(n_1473) );
CKINVDCx5p33_ASAP7_75t_R g1516 ( .A(n_3), .Y(n_1516) );
AOI221xp5_ASAP7_75t_L g1334 ( .A1(n_4), .A2(n_248), .B1(n_1088), .B2(n_1126), .C(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1353 ( .A(n_4), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_5), .A2(n_97), .B1(n_452), .B2(n_460), .Y(n_451) );
INVx1_ASAP7_75t_L g553 ( .A(n_5), .Y(n_553) );
INVx1_ASAP7_75t_L g1738 ( .A(n_6), .Y(n_1738) );
OAI22xp5_ASAP7_75t_L g1293 ( .A1(n_7), .A2(n_313), .B1(n_679), .B2(n_682), .Y(n_1293) );
INVx1_ASAP7_75t_L g1313 ( .A(n_7), .Y(n_1313) );
INVx1_ASAP7_75t_L g1943 ( .A(n_8), .Y(n_1943) );
AOI22xp33_ASAP7_75t_L g1967 ( .A1(n_8), .A2(n_143), .B1(n_1374), .B2(n_1968), .Y(n_1967) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_9), .A2(n_209), .B1(n_1125), .B2(n_1126), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_9), .A2(n_209), .B1(n_1139), .B2(n_1141), .Y(n_1138) );
AOI221xp5_ASAP7_75t_L g1269 ( .A1(n_10), .A2(n_201), .B1(n_714), .B2(n_715), .C(n_1088), .Y(n_1269) );
OAI22xp33_ASAP7_75t_L g1274 ( .A1(n_10), .A2(n_316), .B1(n_682), .B2(n_885), .Y(n_1274) );
INVx1_ASAP7_75t_L g1578 ( .A(n_11), .Y(n_1578) );
INVx1_ASAP7_75t_L g701 ( .A(n_12), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_12), .A2(n_107), .B1(n_734), .B2(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g843 ( .A(n_13), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g856 ( .A1(n_13), .A2(n_194), .B1(n_609), .B2(n_615), .Y(n_856) );
OAI22xp33_ASAP7_75t_L g619 ( .A1(n_14), .A2(n_95), .B1(n_620), .B2(n_622), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_14), .A2(n_95), .B1(n_629), .B2(n_641), .C(n_643), .Y(n_640) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_15), .A2(n_114), .B1(n_717), .B2(n_719), .Y(n_716) );
AOI22xp33_ASAP7_75t_SL g727 ( .A1(n_15), .A2(n_114), .B1(n_728), .B2(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g1394 ( .A(n_16), .Y(n_1394) );
OAI211xp5_ASAP7_75t_SL g1412 ( .A1(n_16), .A2(n_622), .B(n_1413), .C(n_1419), .Y(n_1412) );
INVx1_ASAP7_75t_L g1195 ( .A(n_17), .Y(n_1195) );
AOI22xp33_ASAP7_75t_SL g1210 ( .A1(n_17), .A2(n_282), .B1(n_731), .B2(n_1211), .Y(n_1210) );
INVx1_ASAP7_75t_L g1288 ( .A(n_18), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g1389 ( .A(n_19), .Y(n_1389) );
AO221x2_ASAP7_75t_L g1736 ( .A1(n_20), .A2(n_274), .B1(n_1702), .B2(n_1721), .C(n_1737), .Y(n_1736) );
AO22x2_ASAP7_75t_L g1103 ( .A1(n_21), .A2(n_1104), .B1(n_1161), .B2(n_1162), .Y(n_1103) );
INVxp67_ASAP7_75t_SL g1161 ( .A(n_21), .Y(n_1161) );
CKINVDCx16_ASAP7_75t_R g1327 ( .A(n_22), .Y(n_1327) );
AOI21xp5_ASAP7_75t_L g1952 ( .A1(n_23), .A2(n_593), .B(n_594), .Y(n_1952) );
INVx1_ASAP7_75t_L g1955 ( .A(n_23), .Y(n_1955) );
INVx1_ASAP7_75t_L g1643 ( .A(n_24), .Y(n_1643) );
AOI22xp33_ASAP7_75t_L g1673 ( .A1(n_24), .A2(n_120), .B1(n_803), .B2(n_1146), .Y(n_1673) );
AOI22xp33_ASAP7_75t_SL g720 ( .A1(n_25), .A2(n_90), .B1(n_717), .B2(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_SL g755 ( .A(n_25), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_26), .A2(n_358), .B1(n_1148), .B2(n_1238), .Y(n_1237) );
INVxp67_ASAP7_75t_SL g1259 ( .A(n_26), .Y(n_1259) );
OAI222xp33_ASAP7_75t_L g944 ( .A1(n_27), .A2(n_66), .B1(n_145), .B2(n_744), .C1(n_747), .C2(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g960 ( .A(n_27), .Y(n_960) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_28), .Y(n_1027) );
INVx1_ASAP7_75t_L g1344 ( .A(n_29), .Y(n_1344) );
AOI22xp33_ASAP7_75t_SL g1375 ( .A1(n_29), .A2(n_302), .B1(n_1144), .B2(n_1376), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1331 ( .A1(n_30), .A2(n_69), .B1(n_974), .B2(n_1332), .Y(n_1331) );
INVx1_ASAP7_75t_L g1356 ( .A(n_30), .Y(n_1356) );
INVx1_ASAP7_75t_L g1338 ( .A(n_31), .Y(n_1338) );
AOI22xp33_ASAP7_75t_L g1373 ( .A1(n_31), .A2(n_164), .B1(n_1369), .B2(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1441 ( .A(n_32), .Y(n_1441) );
AOI221xp5_ASAP7_75t_L g1484 ( .A1(n_32), .A2(n_155), .B1(n_1485), .B2(n_1486), .C(n_1487), .Y(n_1484) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_33), .B(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g551 ( .A(n_33), .Y(n_551) );
CKINVDCx5p33_ASAP7_75t_R g1391 ( .A(n_34), .Y(n_1391) );
CKINVDCx5p33_ASAP7_75t_R g1174 ( .A(n_35), .Y(n_1174) );
AOI22xp33_ASAP7_75t_L g997 ( .A1(n_36), .A2(n_153), .B1(n_984), .B2(n_998), .Y(n_997) );
AOI22xp33_ASAP7_75t_SL g1017 ( .A1(n_36), .A2(n_153), .B1(n_860), .B2(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1127 ( .A1(n_37), .A2(n_258), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_37), .A2(n_258), .B1(n_803), .B2(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g368 ( .A(n_38), .Y(n_368) );
CKINVDCx5p33_ASAP7_75t_R g1947 ( .A(n_39), .Y(n_1947) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_40), .A2(n_113), .B1(n_880), .B2(n_1340), .Y(n_1339) );
INVx1_ASAP7_75t_L g1364 ( .A(n_40), .Y(n_1364) );
AOI21xp33_ASAP7_75t_L g1941 ( .A1(n_41), .A2(n_531), .B(n_597), .Y(n_1941) );
INVx1_ASAP7_75t_L g1965 ( .A(n_41), .Y(n_1965) );
XOR2xp5_ASAP7_75t_L g1284 ( .A(n_42), .B(n_1285), .Y(n_1284) );
INVxp67_ASAP7_75t_SL g705 ( .A(n_43), .Y(n_705) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_43), .A2(n_176), .B1(n_744), .B2(n_747), .Y(n_743) );
INVx1_ASAP7_75t_L g763 ( .A(n_44), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g799 ( .A1(n_44), .A2(n_221), .B1(n_714), .B2(n_794), .Y(n_799) );
INVx1_ASAP7_75t_L g1591 ( .A(n_45), .Y(n_1591) );
AOI22xp33_ASAP7_75t_L g1612 ( .A1(n_45), .A2(n_285), .B1(n_1131), .B2(n_1134), .Y(n_1612) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_46), .A2(n_148), .B1(n_793), .B2(n_794), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_46), .A2(n_148), .B1(n_629), .B2(n_731), .Y(n_805) );
CKINVDCx5p33_ASAP7_75t_R g1946 ( .A(n_47), .Y(n_1946) );
INVx1_ASAP7_75t_L g1460 ( .A(n_48), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_48), .A2(n_129), .B1(n_738), .B2(n_1146), .Y(n_1505) );
CKINVDCx5p33_ASAP7_75t_R g1652 ( .A(n_49), .Y(n_1652) );
INVx1_ASAP7_75t_L g1552 ( .A(n_50), .Y(n_1552) );
XNOR2xp5_ASAP7_75t_L g1380 ( .A(n_51), .B(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1061 ( .A(n_52), .Y(n_1061) );
OAI221xp5_ASAP7_75t_L g1083 ( .A1(n_52), .A2(n_622), .B1(n_1084), .B2(n_1090), .C(n_1094), .Y(n_1083) );
AOI22xp5_ASAP7_75t_L g1720 ( .A1(n_53), .A2(n_335), .B1(n_1702), .B2(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g1304 ( .A(n_54), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1317 ( .A1(n_54), .A2(n_237), .B1(n_1000), .B2(n_1139), .Y(n_1317) );
INVx1_ASAP7_75t_L g1235 ( .A(n_55), .Y(n_1235) );
INVx1_ASAP7_75t_L g914 ( .A(n_56), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_57), .A2(n_242), .B1(n_1128), .B2(n_1129), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_57), .A2(n_242), .B1(n_803), .B2(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1605 ( .A(n_58), .Y(n_1605) );
AOI22xp33_ASAP7_75t_L g1621 ( .A1(n_58), .A2(n_273), .B1(n_1148), .B2(n_1238), .Y(n_1621) );
INVx1_ASAP7_75t_L g1607 ( .A(n_59), .Y(n_1607) );
AOI22xp33_ASAP7_75t_L g1620 ( .A1(n_59), .A2(n_311), .B1(n_1146), .B2(n_1372), .Y(n_1620) );
INVx1_ASAP7_75t_L g963 ( .A(n_60), .Y(n_963) );
AOI22xp33_ASAP7_75t_SL g986 ( .A1(n_60), .A2(n_112), .B1(n_629), .B2(n_811), .Y(n_986) );
INVx1_ASAP7_75t_L g1299 ( .A(n_61), .Y(n_1299) );
AOI22xp33_ASAP7_75t_L g1318 ( .A1(n_61), .A2(n_197), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
INVx1_ASAP7_75t_L g580 ( .A(n_62), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_62), .A2(n_254), .B1(n_629), .B2(n_631), .C(n_634), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1387 ( .A(n_63), .Y(n_1387) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_64), .A2(n_319), .B1(n_1169), .B2(n_1170), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g1214 ( .A1(n_64), .A2(n_319), .B1(n_502), .B2(n_729), .Y(n_1214) );
INVx1_ASAP7_75t_L g1597 ( .A(n_65), .Y(n_1597) );
OAI22xp5_ASAP7_75t_L g1601 ( .A1(n_65), .A2(n_336), .B1(n_1154), .B2(n_1602), .Y(n_1601) );
AOI22xp33_ASAP7_75t_SL g967 ( .A1(n_66), .A2(n_305), .B1(n_793), .B2(n_968), .Y(n_967) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_67), .A2(n_196), .B1(n_717), .B2(n_791), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_67), .A2(n_196), .B1(n_728), .B2(n_803), .Y(n_802) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_68), .Y(n_1054) );
INVx1_ASAP7_75t_L g1354 ( .A(n_69), .Y(n_1354) );
INVxp33_ASAP7_75t_SL g1531 ( .A(n_70), .Y(n_1531) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_70), .A2(n_350), .B1(n_1566), .B2(n_1568), .Y(n_1565) );
INVx1_ASAP7_75t_L g1295 ( .A(n_71), .Y(n_1295) );
OAI22xp33_ASAP7_75t_L g1401 ( .A1(n_72), .A2(n_351), .B1(n_1066), .B2(n_1067), .Y(n_1401) );
INVx1_ASAP7_75t_L g1421 ( .A(n_72), .Y(n_1421) );
CKINVDCx5p33_ASAP7_75t_R g902 ( .A(n_73), .Y(n_902) );
INVx1_ASAP7_75t_L g1085 ( .A(n_74), .Y(n_1085) );
OAI22xp33_ASAP7_75t_L g1101 ( .A1(n_74), .A2(n_169), .B1(n_679), .B2(n_682), .Y(n_1101) );
CKINVDCx5p33_ASAP7_75t_R g1658 ( .A(n_75), .Y(n_1658) );
INVx1_ASAP7_75t_L g764 ( .A(n_76), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_76), .A2(n_166), .B1(n_717), .B2(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g1437 ( .A(n_77), .Y(n_1437) );
AOI22xp33_ASAP7_75t_L g1489 ( .A1(n_77), .A2(n_229), .B1(n_1144), .B2(n_1490), .Y(n_1489) );
XNOR2xp5_ASAP7_75t_L g1984 ( .A(n_78), .B(n_1985), .Y(n_1984) );
CKINVDCx5p33_ASAP7_75t_R g835 ( .A(n_79), .Y(n_835) );
AOI22xp33_ASAP7_75t_L g1147 ( .A1(n_80), .A2(n_255), .B1(n_803), .B2(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1157 ( .A(n_80), .Y(n_1157) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_81), .Y(n_1541) );
AOI221xp5_ASAP7_75t_L g1572 ( .A1(n_81), .A2(n_353), .B1(n_1319), .B2(n_1573), .C(n_1574), .Y(n_1572) );
INVx1_ASAP7_75t_L g905 ( .A(n_82), .Y(n_905) );
OAI221xp5_ASAP7_75t_L g917 ( .A1(n_82), .A2(n_620), .B1(n_865), .B2(n_918), .C(n_921), .Y(n_917) );
INVx1_ASAP7_75t_L g1113 ( .A(n_83), .Y(n_1113) );
OAI22xp5_ASAP7_75t_L g1153 ( .A1(n_83), .A2(n_195), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
INVx1_ASAP7_75t_L g1400 ( .A(n_84), .Y(n_1400) );
OAI22xp5_ASAP7_75t_L g1405 ( .A1(n_84), .A2(n_296), .B1(n_609), .B2(n_615), .Y(n_1405) );
CKINVDCx20_ASAP7_75t_R g1226 ( .A(n_85), .Y(n_1226) );
XNOR2x2_ASAP7_75t_L g568 ( .A(n_86), .B(n_569), .Y(n_568) );
INVxp67_ASAP7_75t_SL g693 ( .A(n_87), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_87), .A2(n_259), .B1(n_728), .B2(n_738), .Y(n_737) );
OAI221xp5_ASAP7_75t_L g1448 ( .A1(n_88), .A2(n_119), .B1(n_1449), .B2(n_1454), .C(n_1456), .Y(n_1448) );
OAI22xp5_ASAP7_75t_L g1492 ( .A1(n_88), .A2(n_119), .B1(n_1493), .B2(n_1496), .Y(n_1492) );
CKINVDCx5p33_ASAP7_75t_R g596 ( .A(n_89), .Y(n_596) );
INVxp33_ASAP7_75t_L g754 ( .A(n_90), .Y(n_754) );
BUFx2_ASAP7_75t_L g394 ( .A(n_91), .Y(n_394) );
BUFx2_ASAP7_75t_L g492 ( .A(n_91), .Y(n_492) );
INVx1_ASAP7_75t_L g563 ( .A(n_91), .Y(n_563) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_91), .B(n_607), .Y(n_1453) );
INVx1_ASAP7_75t_L g1935 ( .A(n_92), .Y(n_1935) );
AOI22xp33_ASAP7_75t_L g1970 ( .A1(n_92), .A2(n_133), .B1(n_891), .B2(n_1376), .Y(n_1970) );
OAI22xp33_ASAP7_75t_L g912 ( .A1(n_93), .A2(n_102), .B1(n_649), .B2(n_658), .Y(n_912) );
INVx1_ASAP7_75t_L g933 ( .A(n_93), .Y(n_933) );
CKINVDCx5p33_ASAP7_75t_R g1656 ( .A(n_94), .Y(n_1656) );
CKINVDCx5p33_ASAP7_75t_R g1630 ( .A(n_96), .Y(n_1630) );
INVx1_ASAP7_75t_L g431 ( .A(n_97), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g1611 ( .A1(n_98), .A2(n_357), .B1(n_1128), .B2(n_1129), .Y(n_1611) );
AOI22xp33_ASAP7_75t_SL g1617 ( .A1(n_98), .A2(n_357), .B1(n_1500), .B2(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1091 ( .A(n_99), .Y(n_1091) );
OAI22xp33_ASAP7_75t_L g1102 ( .A1(n_99), .A2(n_198), .B1(n_887), .B2(n_889), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g578 ( .A(n_100), .Y(n_578) );
INVx1_ASAP7_75t_L g1064 ( .A(n_101), .Y(n_1064) );
OAI22xp5_ASAP7_75t_L g1071 ( .A1(n_101), .A2(n_108), .B1(n_609), .B2(n_615), .Y(n_1071) );
INVx1_ASAP7_75t_L g932 ( .A(n_102), .Y(n_932) );
OAI221xp5_ASAP7_75t_L g1532 ( .A1(n_103), .A2(n_184), .B1(n_1449), .B2(n_1456), .C(n_1533), .Y(n_1532) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_103), .A2(n_184), .B1(n_1493), .B2(n_1570), .Y(n_1569) );
AOI221xp5_ASAP7_75t_L g1346 ( .A1(n_104), .A2(n_185), .B1(n_531), .B2(n_702), .C(n_1347), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g1368 ( .A1(n_104), .A2(n_185), .B1(n_1369), .B2(n_1372), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_105), .A2(n_205), .B1(n_714), .B2(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_SL g742 ( .A(n_105), .Y(n_742) );
INVx1_ASAP7_75t_L g1593 ( .A(n_106), .Y(n_1593) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_106), .A2(n_125), .B1(n_702), .B2(n_1614), .Y(n_1613) );
INVxp33_ASAP7_75t_L g696 ( .A(n_107), .Y(n_696) );
INVx1_ASAP7_75t_L g1063 ( .A(n_108), .Y(n_1063) );
AO221x1_ASAP7_75t_L g1022 ( .A1(n_109), .A2(n_203), .B1(n_593), .B2(n_594), .C(n_724), .Y(n_1022) );
INVx1_ASAP7_75t_L g1033 ( .A(n_109), .Y(n_1033) );
OAI221xp5_ASAP7_75t_L g1297 ( .A1(n_110), .A2(n_620), .B1(n_865), .B2(n_1298), .C(n_1302), .Y(n_1297) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_110), .A2(n_262), .B1(n_1146), .B2(n_1322), .Y(n_1321) );
INVx1_ASAP7_75t_L g957 ( .A(n_111), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g987 ( .A1(n_111), .A2(n_226), .B1(n_728), .B2(n_984), .Y(n_987) );
INVx1_ASAP7_75t_L g959 ( .A(n_112), .Y(n_959) );
INVx1_ASAP7_75t_L g1363 ( .A(n_113), .Y(n_1363) );
XNOR2x2_ASAP7_75t_L g1583 ( .A(n_115), .B(n_1584), .Y(n_1583) );
INVx1_ASAP7_75t_L g911 ( .A(n_116), .Y(n_911) );
OAI22xp5_ASAP7_75t_L g916 ( .A1(n_116), .A2(n_233), .B1(n_609), .B2(n_615), .Y(n_916) );
CKINVDCx16_ASAP7_75t_R g1716 ( .A(n_117), .Y(n_1716) );
AO22x2_ASAP7_75t_L g939 ( .A1(n_118), .A2(n_940), .B1(n_941), .B2(n_990), .Y(n_939) );
INVxp67_ASAP7_75t_SL g940 ( .A(n_118), .Y(n_940) );
INVx1_ASAP7_75t_L g1648 ( .A(n_120), .Y(n_1648) );
XNOR2xp5_ASAP7_75t_L g892 ( .A(n_121), .B(n_893), .Y(n_892) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_122), .A2(n_278), .B1(n_731), .B2(n_1000), .Y(n_999) );
AOI221xp5_ASAP7_75t_L g1019 ( .A1(n_122), .A2(n_278), .B1(n_531), .B2(n_597), .C(n_873), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_123), .A2(n_204), .B1(n_793), .B2(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_123), .A2(n_204), .B1(n_629), .B2(n_731), .Y(n_981) );
INVx1_ASAP7_75t_L g1058 ( .A(n_124), .Y(n_1058) );
INVx1_ASAP7_75t_L g1587 ( .A(n_125), .Y(n_1587) );
OA22x2_ASAP7_75t_L g391 ( .A1(n_126), .A2(n_392), .B1(n_566), .B2(n_567), .Y(n_391) );
INVxp67_ASAP7_75t_SL g567 ( .A(n_126), .Y(n_567) );
INVx1_ASAP7_75t_L g1265 ( .A(n_127), .Y(n_1265) );
OAI22xp33_ASAP7_75t_L g1275 ( .A1(n_127), .A2(n_201), .B1(n_887), .B2(n_889), .Y(n_1275) );
AOI22xp5_ASAP7_75t_L g1735 ( .A1(n_128), .A2(n_327), .B1(n_1702), .B2(n_1721), .Y(n_1735) );
INVx1_ASAP7_75t_L g1470 ( .A(n_129), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g1145 ( .A1(n_130), .A2(n_161), .B1(n_1141), .B2(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1160 ( .A(n_130), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g1181 ( .A(n_131), .Y(n_1181) );
INVx1_ASAP7_75t_L g1242 ( .A(n_132), .Y(n_1242) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_132), .A2(n_620), .B1(n_1255), .B2(n_1257), .C(n_1260), .Y(n_1254) );
INVx1_ASAP7_75t_L g1936 ( .A(n_133), .Y(n_1936) );
INVx1_ASAP7_75t_L g1292 ( .A(n_134), .Y(n_1292) );
INVx1_ASAP7_75t_L g782 ( .A(n_135), .Y(n_782) );
AOI22xp33_ASAP7_75t_SL g810 ( .A1(n_135), .A2(n_315), .B1(n_629), .B2(n_811), .Y(n_810) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_136), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g1683 ( .A1(n_137), .A2(n_140), .B1(n_1684), .B2(n_1692), .Y(n_1683) );
OAI22xp5_ASAP7_75t_L g1315 ( .A1(n_138), .A2(n_287), .B1(n_1169), .B2(n_1170), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1323 ( .A1(n_138), .A2(n_287), .B1(n_1247), .B2(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1193 ( .A(n_139), .Y(n_1193) );
AOI22xp33_ASAP7_75t_L g1207 ( .A1(n_139), .A2(n_286), .B1(n_1208), .B2(n_1209), .Y(n_1207) );
AOI22xp5_ASAP7_75t_L g1695 ( .A1(n_141), .A2(n_341), .B1(n_1696), .B2(n_1700), .Y(n_1695) );
CKINVDCx5p33_ASAP7_75t_R g432 ( .A(n_142), .Y(n_432) );
INVx1_ASAP7_75t_L g1940 ( .A(n_143), .Y(n_1940) );
CKINVDCx5p33_ASAP7_75t_R g1951 ( .A(n_144), .Y(n_1951) );
INVx1_ASAP7_75t_L g961 ( .A(n_145), .Y(n_961) );
XOR2xp5_ASAP7_75t_L g1521 ( .A(n_146), .B(n_1522), .Y(n_1521) );
AO221x2_ASAP7_75t_L g1755 ( .A1(n_147), .A2(n_215), .B1(n_1696), .B2(n_1702), .C(n_1756), .Y(n_1755) );
INVx1_ASAP7_75t_L g1688 ( .A(n_149), .Y(n_1688) );
INVx1_ASAP7_75t_L g1811 ( .A(n_150), .Y(n_1811) );
AOI22xp5_ASAP7_75t_L g1719 ( .A1(n_151), .A2(n_349), .B1(n_1684), .B2(n_1692), .Y(n_1719) );
INVx1_ASAP7_75t_L g777 ( .A(n_152), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_152), .A2(n_193), .B1(n_674), .B2(n_803), .Y(n_812) );
INVx1_ASAP7_75t_L g1200 ( .A(n_154), .Y(n_1200) );
INVx1_ASAP7_75t_L g1444 ( .A(n_155), .Y(n_1444) );
INVx1_ASAP7_75t_L g697 ( .A(n_156), .Y(n_697) );
INVx1_ASAP7_75t_L g1644 ( .A(n_157), .Y(n_1644) );
AOI221xp5_ASAP7_75t_L g1670 ( .A1(n_157), .A2(n_211), .B1(n_636), .B2(n_1560), .C(n_1671), .Y(n_1670) );
INVx1_ASAP7_75t_L g1689 ( .A(n_158), .Y(n_1689) );
NAND2xp5_ASAP7_75t_L g1694 ( .A(n_158), .B(n_1687), .Y(n_1694) );
AOI221xp5_ASAP7_75t_L g1948 ( .A1(n_159), .A2(n_304), .B1(n_974), .B2(n_1949), .C(n_1950), .Y(n_1948) );
INVx1_ASAP7_75t_L g1958 ( .A(n_159), .Y(n_1958) );
INVx1_ASAP7_75t_L g1109 ( .A(n_160), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_160), .A2(n_189), .B1(n_1131), .B2(n_1134), .Y(n_1130) );
INVx1_ASAP7_75t_L g1151 ( .A(n_161), .Y(n_1151) );
INVx1_ASAP7_75t_L g1632 ( .A(n_162), .Y(n_1632) );
AOI21xp33_ASAP7_75t_L g1667 ( .A1(n_162), .A2(n_1004), .B(n_1668), .Y(n_1667) );
INVx2_ASAP7_75t_L g380 ( .A(n_163), .Y(n_380) );
INVx1_ASAP7_75t_L g1349 ( .A(n_164), .Y(n_1349) );
INVx1_ASAP7_75t_L g1633 ( .A(n_165), .Y(n_1633) );
AOI22xp33_ASAP7_75t_L g1666 ( .A1(n_165), .A2(n_234), .B1(n_804), .B2(n_1051), .Y(n_1666) );
INVx1_ASAP7_75t_L g767 ( .A(n_166), .Y(n_767) );
OAI22xp5_ASAP7_75t_L g1249 ( .A1(n_167), .A2(n_207), .B1(n_1067), .B2(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1271 ( .A(n_167), .Y(n_1271) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_168), .A2(n_266), .B1(n_974), .B2(n_975), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_168), .A2(n_266), .B1(n_983), .B2(n_984), .Y(n_982) );
INVx1_ASAP7_75t_L g1092 ( .A(n_169), .Y(n_1092) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_170), .Y(n_504) );
INVx1_ASAP7_75t_L g450 ( .A(n_171), .Y(n_450) );
BUFx3_ASAP7_75t_L g466 ( .A(n_171), .Y(n_466) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_172), .Y(n_478) );
INVx1_ASAP7_75t_L g1757 ( .A(n_173), .Y(n_1757) );
CKINVDCx5p33_ASAP7_75t_R g1025 ( .A(n_174), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g848 ( .A1(n_175), .A2(n_334), .B1(n_649), .B2(n_658), .Y(n_848) );
INVx1_ASAP7_75t_L g875 ( .A(n_175), .Y(n_875) );
INVx1_ASAP7_75t_L g708 ( .A(n_176), .Y(n_708) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_177), .Y(n_439) );
INVxp33_ASAP7_75t_SL g1528 ( .A(n_178), .Y(n_1528) );
AOI221xp5_ASAP7_75t_L g1559 ( .A1(n_178), .A2(n_297), .B1(n_1146), .B2(n_1560), .C(n_1562), .Y(n_1559) );
AOI221xp5_ASAP7_75t_L g872 ( .A1(n_179), .A2(n_344), .B1(n_593), .B2(n_594), .C(n_873), .Y(n_872) );
OAI22xp33_ASAP7_75t_L g886 ( .A1(n_179), .A2(n_202), .B1(n_887), .B2(n_889), .Y(n_886) );
INVx1_ASAP7_75t_L g927 ( .A(n_180), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g936 ( .A1(n_180), .A2(n_182), .B1(n_887), .B2(n_889), .Y(n_936) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_181), .A2(n_323), .B1(n_609), .B2(n_615), .Y(n_608) );
INVx1_ASAP7_75t_L g647 ( .A(n_181), .Y(n_647) );
AOI221xp5_ASAP7_75t_L g930 ( .A1(n_182), .A2(n_223), .B1(n_593), .B2(n_594), .C(n_704), .Y(n_930) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_183), .A2(n_253), .B1(n_747), .B2(n_769), .C(n_770), .Y(n_768) );
INVx1_ASAP7_75t_L g780 ( .A(n_183), .Y(n_780) );
INVx1_ASAP7_75t_L g1244 ( .A(n_186), .Y(n_1244) );
OAI211xp5_ASAP7_75t_SL g1261 ( .A1(n_186), .A2(n_622), .B(n_1262), .C(n_1270), .Y(n_1261) );
CKINVDCx5p33_ASAP7_75t_R g1010 ( .A(n_187), .Y(n_1010) );
INVx1_ASAP7_75t_L g1809 ( .A(n_188), .Y(n_1809) );
INVx1_ASAP7_75t_L g1119 ( .A(n_189), .Y(n_1119) );
AOI22xp33_ASAP7_75t_SL g1005 ( .A1(n_190), .A2(n_359), .B1(n_674), .B2(n_729), .Y(n_1005) );
INVx1_ASAP7_75t_L g1014 ( .A(n_190), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1475 ( .A(n_191), .Y(n_1475) );
AOI221xp5_ASAP7_75t_L g1418 ( .A1(n_192), .A2(n_360), .B1(n_597), .B2(n_704), .C(n_1088), .Y(n_1418) );
OAI22xp33_ASAP7_75t_L g1424 ( .A1(n_192), .A2(n_291), .B1(n_887), .B2(n_889), .Y(n_1424) );
INVx1_ASAP7_75t_L g778 ( .A(n_193), .Y(n_778) );
INVx1_ASAP7_75t_L g846 ( .A(n_194), .Y(n_846) );
INVx1_ASAP7_75t_L g1116 ( .A(n_195), .Y(n_1116) );
INVx1_ASAP7_75t_L g1301 ( .A(n_197), .Y(n_1301) );
INVx1_ASAP7_75t_L g1086 ( .A(n_198), .Y(n_1086) );
INVx1_ASAP7_75t_L g1758 ( .A(n_199), .Y(n_1758) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_200), .Y(n_1177) );
INVx1_ASAP7_75t_L g869 ( .A(n_202), .Y(n_869) );
INVx1_ASAP7_75t_L g1035 ( .A(n_203), .Y(n_1035) );
INVxp33_ASAP7_75t_L g749 ( .A(n_205), .Y(n_749) );
INVx1_ASAP7_75t_L g490 ( .A(n_206), .Y(n_490) );
INVx1_ASAP7_75t_L g656 ( .A(n_206), .Y(n_656) );
INVx1_ASAP7_75t_L g1272 ( .A(n_207), .Y(n_1272) );
CKINVDCx5p33_ASAP7_75t_R g509 ( .A(n_208), .Y(n_509) );
INVx1_ASAP7_75t_L g1730 ( .A(n_210), .Y(n_1730) );
INVx1_ASAP7_75t_L g1646 ( .A(n_211), .Y(n_1646) );
CKINVDCx5p33_ASAP7_75t_R g1472 ( .A(n_212), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g1183 ( .A(n_213), .Y(n_1183) );
INVx1_ASAP7_75t_L g1554 ( .A(n_214), .Y(n_1554) );
XOR2x2_ASAP7_75t_L g1165 ( .A(n_215), .B(n_1166), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1001 ( .A1(n_216), .A2(n_333), .B1(n_629), .B2(n_1002), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1021 ( .A1(n_216), .A2(n_622), .B1(n_1022), .B2(n_1023), .C(n_1026), .Y(n_1021) );
INVx1_ASAP7_75t_L g1393 ( .A(n_217), .Y(n_1393) );
OAI221xp5_ASAP7_75t_L g1406 ( .A1(n_217), .A2(n_620), .B1(n_865), .B2(n_1407), .C(n_1411), .Y(n_1406) );
CKINVDCx5p33_ASAP7_75t_R g1476 ( .A(n_218), .Y(n_1476) );
CKINVDCx5p33_ASAP7_75t_R g1108 ( .A(n_219), .Y(n_1108) );
XOR2xp5_ASAP7_75t_L g1432 ( .A(n_220), .B(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g771 ( .A(n_221), .Y(n_771) );
INVxp67_ASAP7_75t_SL g1543 ( .A(n_222), .Y(n_1543) );
AOI22xp33_ASAP7_75t_L g1575 ( .A1(n_222), .A2(n_299), .B1(n_1238), .B2(n_1576), .Y(n_1575) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_223), .A2(n_321), .B1(n_682), .B2(n_885), .Y(n_935) );
INVx1_ASAP7_75t_L g1462 ( .A(n_224), .Y(n_1462) );
AOI221xp5_ASAP7_75t_L g1499 ( .A1(n_224), .A2(n_239), .B1(n_1500), .B2(n_1501), .C(n_1502), .Y(n_1499) );
CKINVDCx5p33_ASAP7_75t_R g1932 ( .A(n_225), .Y(n_1932) );
INVx1_ASAP7_75t_L g956 ( .A(n_226), .Y(n_956) );
CKINVDCx5p33_ASAP7_75t_R g601 ( .A(n_227), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g648 ( .A1(n_227), .A2(n_649), .B1(n_657), .B2(n_658), .C(n_661), .Y(n_648) );
CKINVDCx5p33_ASAP7_75t_R g1650 ( .A(n_228), .Y(n_1650) );
INVx1_ASAP7_75t_L g1446 ( .A(n_229), .Y(n_1446) );
CKINVDCx5p33_ASAP7_75t_R g1930 ( .A(n_230), .Y(n_1930) );
INVx1_ASAP7_75t_L g1069 ( .A(n_231), .Y(n_1069) );
AOI22xp5_ASAP7_75t_L g1734 ( .A1(n_232), .A2(n_300), .B1(n_1684), .B2(n_1692), .Y(n_1734) );
INVx1_ASAP7_75t_L g910 ( .A(n_233), .Y(n_910) );
INVx1_ASAP7_75t_L g1628 ( .A(n_234), .Y(n_1628) );
INVx1_ASAP7_75t_L g1291 ( .A(n_235), .Y(n_1291) );
CKINVDCx5p33_ASAP7_75t_R g1180 ( .A(n_236), .Y(n_1180) );
INVx1_ASAP7_75t_L g1303 ( .A(n_237), .Y(n_1303) );
CKINVDCx5p33_ASAP7_75t_R g828 ( .A(n_238), .Y(n_828) );
INVx1_ASAP7_75t_L g1466 ( .A(n_239), .Y(n_1466) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_240), .Y(n_766) );
OAI22xp33_ASAP7_75t_L g1065 ( .A1(n_241), .A2(n_329), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
INVx1_ASAP7_75t_L g1096 ( .A(n_241), .Y(n_1096) );
CKINVDCx5p33_ASAP7_75t_R g1944 ( .A(n_243), .Y(n_1944) );
AOI22xp33_ASAP7_75t_L g1610 ( .A1(n_244), .A2(n_320), .B1(n_1125), .B2(n_1126), .Y(n_1610) );
AOI22xp33_ASAP7_75t_SL g1619 ( .A1(n_244), .A2(n_320), .B1(n_1139), .B2(n_1372), .Y(n_1619) );
CKINVDCx16_ASAP7_75t_R g685 ( .A(n_245), .Y(n_685) );
INVx1_ASAP7_75t_L g837 ( .A(n_246), .Y(n_837) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_246), .A2(n_620), .B1(n_858), .B2(n_861), .C(n_865), .Y(n_857) );
INVx1_ASAP7_75t_L g1060 ( .A(n_247), .Y(n_1060) );
OAI221xp5_ASAP7_75t_L g1072 ( .A1(n_247), .A2(n_620), .B1(n_865), .B2(n_1073), .C(n_1078), .Y(n_1072) );
INVx1_ASAP7_75t_L g1357 ( .A(n_248), .Y(n_1357) );
CKINVDCx5p33_ASAP7_75t_R g832 ( .A(n_249), .Y(n_832) );
INVx1_ASAP7_75t_L g1118 ( .A(n_250), .Y(n_1118) );
AOI22xp33_ASAP7_75t_L g1135 ( .A1(n_250), .A2(n_345), .B1(n_1125), .B2(n_1126), .Y(n_1135) );
CKINVDCx5p33_ASAP7_75t_R g590 ( .A(n_251), .Y(n_590) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_252), .A2(n_268), .B1(n_399), .B2(n_407), .Y(n_398) );
INVx1_ASAP7_75t_L g523 ( .A(n_252), .Y(n_523) );
INVx1_ASAP7_75t_L g781 ( .A(n_253), .Y(n_781) );
AOI21xp33_ASAP7_75t_L g582 ( .A1(n_254), .A2(n_531), .B(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g1158 ( .A(n_255), .Y(n_1158) );
OAI221xp5_ASAP7_75t_L g1171 ( .A1(n_256), .A2(n_622), .B1(n_1172), .B2(n_1178), .C(n_1182), .Y(n_1171) );
AOI22xp33_ASAP7_75t_SL g1213 ( .A1(n_256), .A2(n_332), .B1(n_641), .B2(n_1211), .Y(n_1213) );
OAI211xp5_ASAP7_75t_L g413 ( .A1(n_257), .A2(n_414), .B(n_419), .C(n_426), .Y(n_413) );
INVx1_ASAP7_75t_L g519 ( .A(n_257), .Y(n_519) );
INVx1_ASAP7_75t_L g691 ( .A(n_259), .Y(n_691) );
INVx1_ASAP7_75t_L g1052 ( .A(n_260), .Y(n_1052) );
BUFx3_ASAP7_75t_L g449 ( .A(n_261), .Y(n_449) );
INVx1_ASAP7_75t_L g459 ( .A(n_261), .Y(n_459) );
OAI221xp5_ASAP7_75t_L g1305 ( .A1(n_262), .A2(n_622), .B1(n_1306), .B2(n_1308), .C(n_1314), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g1933 ( .A(n_263), .Y(n_1933) );
INVx1_ASAP7_75t_L g840 ( .A(n_264), .Y(n_840) );
OAI211xp5_ASAP7_75t_L g866 ( .A1(n_264), .A2(n_622), .B(n_867), .C(n_874), .Y(n_866) );
CKINVDCx5p33_ASAP7_75t_R g1008 ( .A(n_265), .Y(n_1008) );
AO22x2_ASAP7_75t_L g758 ( .A1(n_267), .A2(n_759), .B1(n_813), .B2(n_814), .Y(n_758) );
INVxp67_ASAP7_75t_L g813 ( .A(n_267), .Y(n_813) );
INVx1_ASAP7_75t_L g521 ( .A(n_268), .Y(n_521) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_269), .Y(n_376) );
INVx1_ASAP7_75t_L g565 ( .A(n_269), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_269), .B(n_338), .Y(n_607) );
AND2x2_ASAP7_75t_L g611 ( .A(n_269), .B(n_403), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_270), .Y(n_1024) );
INVx1_ASAP7_75t_L g1815 ( .A(n_271), .Y(n_1815) );
AOI21xp33_ASAP7_75t_L g592 ( .A1(n_272), .A2(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g672 ( .A(n_272), .Y(n_672) );
INVx1_ASAP7_75t_L g1604 ( .A(n_273), .Y(n_1604) );
INVx1_ASAP7_75t_L g1731 ( .A(n_275), .Y(n_1731) );
INVx2_ASAP7_75t_L g446 ( .A(n_276), .Y(n_446) );
OR2x2_ASAP7_75t_L g671 ( .A(n_276), .B(n_656), .Y(n_671) );
INVx1_ASAP7_75t_L g1813 ( .A(n_277), .Y(n_1813) );
CKINVDCx16_ASAP7_75t_R g1728 ( .A(n_279), .Y(n_1728) );
INVx1_ASAP7_75t_L g871 ( .A(n_280), .Y(n_871) );
OAI22xp33_ASAP7_75t_L g884 ( .A1(n_280), .A2(n_344), .B1(n_682), .B2(n_885), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g1385 ( .A(n_281), .Y(n_1385) );
INVx1_ASAP7_75t_L g1198 ( .A(n_282), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g575 ( .A(n_283), .Y(n_575) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_284), .Y(n_500) );
INVx1_ASAP7_75t_L g1588 ( .A(n_285), .Y(n_1588) );
INVx1_ASAP7_75t_L g1190 ( .A(n_286), .Y(n_1190) );
INVx1_ASAP7_75t_L g850 ( .A(n_288), .Y(n_850) );
INVx1_ASAP7_75t_L g908 ( .A(n_289), .Y(n_908) );
OAI211xp5_ASAP7_75t_L g925 ( .A1(n_289), .A2(n_622), .B(n_926), .C(n_931), .Y(n_925) );
INVx1_ASAP7_75t_L g1549 ( .A(n_290), .Y(n_1549) );
INVx1_ASAP7_75t_L g1414 ( .A(n_291), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g586 ( .A(n_292), .Y(n_586) );
INVx1_ASAP7_75t_L g1417 ( .A(n_293), .Y(n_1417) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_293), .A2(n_360), .B1(n_679), .B2(n_682), .Y(n_1423) );
INVx1_ASAP7_75t_L g1707 ( .A(n_294), .Y(n_1707) );
INVx1_ASAP7_75t_L g1623 ( .A(n_295), .Y(n_1623) );
INVx1_ASAP7_75t_L g1397 ( .A(n_296), .Y(n_1397) );
INVxp33_ASAP7_75t_L g1530 ( .A(n_297), .Y(n_1530) );
INVx1_ASAP7_75t_L g953 ( .A(n_298), .Y(n_953) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_298), .A2(n_309), .B1(n_717), .B2(n_970), .Y(n_969) );
INVxp33_ASAP7_75t_L g1536 ( .A(n_299), .Y(n_1536) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_301), .Y(n_512) );
INVx1_ASAP7_75t_L g1343 ( .A(n_302), .Y(n_1343) );
AOI22x1_ASAP7_75t_L g992 ( .A1(n_303), .A2(n_993), .B1(n_994), .B2(n_1036), .Y(n_992) );
INVxp67_ASAP7_75t_SL g1036 ( .A(n_303), .Y(n_1036) );
INVx1_ASAP7_75t_L g1956 ( .A(n_304), .Y(n_1956) );
INVx1_ASAP7_75t_L g949 ( .A(n_305), .Y(n_949) );
AOI22xp5_ASAP7_75t_L g1245 ( .A1(n_306), .A2(n_339), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
OAI22xp5_ASAP7_75t_L g1253 ( .A1(n_306), .A2(n_339), .B1(n_609), .B2(n_615), .Y(n_1253) );
INVx1_ASAP7_75t_L g1223 ( .A(n_307), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g713 ( .A1(n_308), .A2(n_354), .B1(n_714), .B2(n_715), .Y(n_713) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_308), .A2(n_354), .B1(n_471), .B2(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g952 ( .A(n_309), .Y(n_952) );
CKINVDCx5p33_ASAP7_75t_R g1655 ( .A(n_310), .Y(n_1655) );
INVx1_ASAP7_75t_L g1600 ( .A(n_311), .Y(n_1600) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_312), .Y(n_898) );
INVx1_ASAP7_75t_L g1307 ( .A(n_313), .Y(n_1307) );
INVx1_ASAP7_75t_L g1739 ( .A(n_314), .Y(n_1739) );
INVx1_ASAP7_75t_L g787 ( .A(n_315), .Y(n_787) );
INVx1_ASAP7_75t_L g1268 ( .A(n_316), .Y(n_1268) );
INVx1_ASAP7_75t_L g1289 ( .A(n_317), .Y(n_1289) );
CKINVDCx5p33_ASAP7_75t_R g1590 ( .A(n_318), .Y(n_1590) );
INVx1_ASAP7_75t_L g929 ( .A(n_321), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_322), .Y(n_899) );
INVx1_ASAP7_75t_L g644 ( .A(n_323), .Y(n_644) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_324), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g1691 ( .A(n_324), .B(n_368), .Y(n_1691) );
AND3x2_ASAP7_75t_L g1699 ( .A(n_324), .B(n_368), .C(n_1688), .Y(n_1699) );
CKINVDCx5p33_ASAP7_75t_R g1403 ( .A(n_325), .Y(n_1403) );
INVx2_ASAP7_75t_L g381 ( .A(n_326), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g1057 ( .A(n_328), .Y(n_1057) );
INVx1_ASAP7_75t_L g1095 ( .A(n_329), .Y(n_1095) );
CKINVDCx5p33_ASAP7_75t_R g830 ( .A(n_330), .Y(n_830) );
INVx1_ASAP7_75t_L g901 ( .A(n_331), .Y(n_901) );
AOI21xp33_ASAP7_75t_L g923 ( .A1(n_331), .A2(n_531), .B(n_924), .Y(n_923) );
OAI221xp5_ASAP7_75t_L g1186 ( .A1(n_332), .A2(n_620), .B1(n_865), .B2(n_1187), .C(n_1194), .Y(n_1186) );
INVx1_ASAP7_75t_L g1020 ( .A(n_333), .Y(n_1020) );
INVx1_ASAP7_75t_L g878 ( .A(n_334), .Y(n_878) );
XNOR2xp5_ASAP7_75t_L g1044 ( .A(n_335), .B(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g1594 ( .A(n_336), .Y(n_1594) );
OAI221xp5_ASAP7_75t_L g1635 ( .A1(n_337), .A2(n_340), .B1(n_1449), .B2(n_1454), .C(n_1636), .Y(n_1635) );
OAI221xp5_ASAP7_75t_L g1661 ( .A1(n_337), .A2(n_340), .B1(n_1496), .B2(n_1662), .C(n_1664), .Y(n_1661) );
INVx1_ASAP7_75t_L g383 ( .A(n_338), .Y(n_383) );
INVx2_ASAP7_75t_L g403 ( .A(n_338), .Y(n_403) );
AO22x2_ASAP7_75t_L g1926 ( .A1(n_341), .A2(n_1927), .B1(n_1971), .B2(n_1972), .Y(n_1926) );
INVxp67_ASAP7_75t_SL g1971 ( .A(n_341), .Y(n_1971) );
AOI22xp33_ASAP7_75t_L g1978 ( .A1(n_341), .A2(n_1979), .B1(n_1983), .B2(n_1986), .Y(n_1978) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_342), .Y(n_397) );
INVx1_ASAP7_75t_L g1555 ( .A(n_343), .Y(n_1555) );
INVx1_ASAP7_75t_L g1111 ( .A(n_345), .Y(n_1111) );
INVx1_ASAP7_75t_L g600 ( .A(n_346), .Y(n_600) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_346), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g468 ( .A1(n_347), .A2(n_469), .B(n_474), .C(n_485), .Y(n_468) );
INVx1_ASAP7_75t_L g558 ( .A(n_347), .Y(n_558) );
INVx1_ASAP7_75t_L g1710 ( .A(n_348), .Y(n_1710) );
INVxp33_ASAP7_75t_SL g1526 ( .A(n_350), .Y(n_1526) );
INVx1_ASAP7_75t_L g1420 ( .A(n_351), .Y(n_1420) );
NOR2xp33_ASAP7_75t_L g1358 ( .A(n_352), .B(n_1359), .Y(n_1358) );
INVxp33_ASAP7_75t_SL g1538 ( .A(n_353), .Y(n_1538) );
CKINVDCx5p33_ASAP7_75t_R g1185 ( .A(n_355), .Y(n_1185) );
INVx1_ASAP7_75t_L g1234 ( .A(n_356), .Y(n_1234) );
INVxp33_ASAP7_75t_SL g1258 ( .A(n_358), .Y(n_1258) );
INVx1_ASAP7_75t_L g1015 ( .A(n_359), .Y(n_1015) );
AOI21xp5_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_384), .B(n_1675), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx3_ASAP7_75t_SL g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_SL g364 ( .A(n_365), .Y(n_364) );
AND2x4_ASAP7_75t_L g365 ( .A(n_366), .B(n_371), .Y(n_365) );
AND2x4_ASAP7_75t_L g1977 ( .A(n_366), .B(n_372), .Y(n_1977) );
NOR2xp33_ASAP7_75t_SL g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVx1_ASAP7_75t_SL g1982 ( .A(n_367), .Y(n_1982) );
NAND2xp5_ASAP7_75t_L g1991 ( .A(n_367), .B(n_369), .Y(n_1991) );
HB1xp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g1981 ( .A(n_369), .B(n_1982), .Y(n_1981) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_377), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g393 ( .A(n_374), .B(n_394), .Y(n_393) );
OR2x6_ASAP7_75t_L g688 ( .A(n_374), .B(n_394), .Y(n_688) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AND2x2_ASAP7_75t_L g712 ( .A(n_375), .B(n_383), .Y(n_712) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
OR2x2_ASAP7_75t_L g531 ( .A(n_376), .B(n_402), .Y(n_531) );
INVx8_ASAP7_75t_L g396 ( .A(n_377), .Y(n_396) );
OR2x6_ASAP7_75t_L g377 ( .A(n_378), .B(n_382), .Y(n_377) );
BUFx6f_ASAP7_75t_L g533 ( .A(n_378), .Y(n_533) );
OR2x6_ASAP7_75t_L g699 ( .A(n_378), .B(n_401), .Y(n_699) );
INVx1_ASAP7_75t_L g863 ( .A(n_378), .Y(n_863) );
INVx2_ASAP7_75t_SL g1080 ( .A(n_378), .Y(n_1080) );
OR2x2_ASAP7_75t_L g1519 ( .A(n_378), .B(n_1453), .Y(n_1519) );
INVx2_ASAP7_75t_SL g1642 ( .A(n_378), .Y(n_1642) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
INVx2_ASAP7_75t_L g406 ( .A(n_380), .Y(n_406) );
AND2x4_ASAP7_75t_L g411 ( .A(n_380), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g418 ( .A(n_380), .Y(n_418) );
INVx1_ASAP7_75t_L g425 ( .A(n_380), .Y(n_425) );
AND2x2_ASAP7_75t_L g430 ( .A(n_380), .B(n_381), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_381), .B(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g412 ( .A(n_381), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_381), .Y(n_417) );
INVx1_ASAP7_75t_L g434 ( .A(n_381), .Y(n_434) );
INVx1_ASAP7_75t_L g614 ( .A(n_381), .Y(n_614) );
AND2x4_ASAP7_75t_L g433 ( .A(n_382), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
OR2x2_ASAP7_75t_L g1155 ( .A(n_383), .B(n_437), .Y(n_1155) );
OR2x2_ASAP7_75t_L g1602 ( .A(n_383), .B(n_437), .Y(n_1602) );
OAI22xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B1(n_1278), .B2(n_1279), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_1037), .B1(n_1038), .B2(n_1277), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
HB1xp67_ASAP7_75t_L g1277 ( .A(n_388), .Y(n_1277) );
XNOR2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_816), .Y(n_388) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_683), .Y(n_389) );
XNOR2x1_ASAP7_75t_L g390 ( .A(n_391), .B(n_568), .Y(n_390) );
INVx1_ASAP7_75t_L g566 ( .A(n_392), .Y(n_566) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B(n_440), .C(n_493), .Y(n_392) );
AOI31xp33_ASAP7_75t_L g1149 ( .A1(n_393), .A2(n_1150), .A3(n_1156), .B(n_1159), .Y(n_1149) );
AND2x4_ASAP7_75t_L g526 ( .A(n_394), .B(n_527), .Y(n_526) );
AND2x4_ASAP7_75t_L g675 ( .A(n_394), .B(n_676), .Y(n_675) );
AND2x4_ASAP7_75t_L g739 ( .A(n_394), .B(n_527), .Y(n_739) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_397), .B(n_398), .C(n_413), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_396), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_396), .A2(n_698), .B1(n_766), .B2(n_787), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g962 ( .A1(n_396), .A2(n_950), .B1(n_963), .B2(n_964), .Y(n_962) );
AOI22xp33_ASAP7_75t_L g1159 ( .A1(n_396), .A2(n_964), .B1(n_1108), .B2(n_1160), .Y(n_1159) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_396), .A2(n_698), .B1(n_1590), .B2(n_1607), .Y(n_1606) );
OAI22xp33_ASAP7_75t_L g516 ( .A1(n_397), .A2(n_510), .B1(n_517), .B2(n_519), .Y(n_516) );
OR2x2_ASAP7_75t_L g399 ( .A(n_400), .B(n_404), .Y(n_399) );
AOI322xp5_ASAP7_75t_L g426 ( .A1(n_400), .A2(n_427), .A3(n_431), .B1(n_432), .B2(n_433), .C1(n_435), .C2(n_439), .Y(n_426) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
AND2x4_ASAP7_75t_L g408 ( .A(n_401), .B(n_409), .Y(n_408) );
AND2x4_ASAP7_75t_L g692 ( .A(n_401), .B(n_612), .Y(n_692) );
AND2x4_ASAP7_75t_L g694 ( .A(n_401), .B(n_409), .Y(n_694) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g423 ( .A(n_403), .Y(n_423) );
INVx2_ASAP7_75t_L g539 ( .A(n_404), .Y(n_539) );
BUFx2_ASAP7_75t_L g1548 ( .A(n_404), .Y(n_1548) );
BUFx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g546 ( .A(n_405), .Y(n_546) );
INVx1_ASAP7_75t_L g574 ( .A(n_405), .Y(n_574) );
INVx1_ASAP7_75t_L g603 ( .A(n_406), .Y(n_603) );
AND2x4_ASAP7_75t_L g612 ( .A(n_406), .B(n_613), .Y(n_612) );
INVx5_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g1156 ( .A1(n_408), .A2(n_692), .B1(n_1157), .B2(n_1158), .Y(n_1156) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
HB1xp67_ASAP7_75t_L g1077 ( .A(n_410), .Y(n_1077) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g542 ( .A(n_411), .Y(n_542) );
INVx3_ASAP7_75t_L g550 ( .A(n_411), .Y(n_550) );
BUFx6f_ASAP7_75t_L g860 ( .A(n_411), .Y(n_860) );
AND2x4_ASAP7_75t_L g424 ( .A(n_412), .B(n_425), .Y(n_424) );
OAI22xp33_ASAP7_75t_L g1640 ( .A1(n_414), .A2(n_1641), .B1(n_1643), .B2(n_1644), .Y(n_1640) );
OAI22xp33_ASAP7_75t_L g1653 ( .A1(n_414), .A2(n_1654), .B1(n_1655), .B2(n_1656), .Y(n_1653) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g1256 ( .A(n_415), .Y(n_1256) );
BUFx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx2_ASAP7_75t_L g536 ( .A(n_416), .Y(n_536) );
INVx3_ASAP7_75t_L g581 ( .A(n_416), .Y(n_581) );
INVx2_ASAP7_75t_L g591 ( .A(n_416), .Y(n_591) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_417), .B(n_418), .Y(n_557) );
INVx1_ASAP7_75t_L g437 ( .A(n_418), .Y(n_437) );
NAND4xp25_ASAP7_75t_SL g689 ( .A(n_419), .B(n_690), .C(n_695), .D(n_700), .Y(n_689) );
NAND4xp25_ASAP7_75t_SL g775 ( .A(n_419), .B(n_776), .C(n_779), .D(n_786), .Y(n_775) );
NAND4xp25_ASAP7_75t_SL g954 ( .A(n_419), .B(n_955), .C(n_958), .D(n_962), .Y(n_954) );
CKINVDCx11_ASAP7_75t_R g419 ( .A(n_420), .Y(n_419) );
AOI211xp5_ASAP7_75t_L g1150 ( .A1(n_420), .A2(n_1151), .B(n_1152), .C(n_1153), .Y(n_1150) );
AOI211xp5_ASAP7_75t_L g1599 ( .A1(n_420), .A2(n_794), .B(n_1600), .C(n_1601), .Y(n_1599) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVxp67_ASAP7_75t_L g438 ( .A(n_422), .Y(n_438) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g564 ( .A(n_423), .B(n_565), .Y(n_564) );
BUFx3_ASAP7_75t_L g624 ( .A(n_424), .Y(n_624) );
BUFx6f_ASAP7_75t_L g704 ( .A(n_424), .Y(n_704) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_424), .Y(n_724) );
BUFx2_ASAP7_75t_L g785 ( .A(n_424), .Y(n_785) );
BUFx3_ASAP7_75t_L g873 ( .A(n_424), .Y(n_873) );
INVx2_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx2_ASAP7_75t_L g793 ( .A(n_428), .Y(n_793) );
INVx2_ASAP7_75t_SL g924 ( .A(n_428), .Y(n_924) );
INVx3_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_429), .Y(n_597) );
AND2x4_ASAP7_75t_L g621 ( .A(n_429), .B(n_611), .Y(n_621) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g584 ( .A(n_430), .Y(n_584) );
AOI322xp5_ASAP7_75t_L g474 ( .A1(n_432), .A2(n_439), .A3(n_475), .B1(n_477), .B2(n_478), .C1(n_479), .C2(n_483), .Y(n_474) );
INVx2_ASAP7_75t_L g707 ( .A(n_433), .Y(n_707) );
AOI222xp33_ASAP7_75t_L g779 ( .A1(n_433), .A2(n_435), .B1(n_780), .B2(n_781), .C1(n_782), .C2(n_783), .Y(n_779) );
INVx2_ASAP7_75t_L g1154 ( .A(n_433), .Y(n_1154) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_434), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_599) );
HB1xp67_ASAP7_75t_L g877 ( .A(n_434), .Y(n_877) );
INVx1_ASAP7_75t_L g1031 ( .A(n_434), .Y(n_1031) );
AOI222xp33_ASAP7_75t_L g700 ( .A1(n_435), .A2(n_701), .B1(n_702), .B2(n_705), .C1(n_706), .C2(n_708), .Y(n_700) );
AOI222xp33_ASAP7_75t_L g958 ( .A1(n_435), .A2(n_702), .B1(n_706), .B2(n_959), .C1(n_960), .C2(n_961), .Y(n_958) );
AND2x4_ASAP7_75t_L g435 ( .A(n_436), .B(n_438), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_436), .A2(n_1008), .B1(n_1010), .B2(n_1030), .Y(n_1029) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI31xp33_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_451), .A3(n_468), .B(n_488), .Y(n_440) );
INVx4_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g752 ( .A1(n_443), .A2(n_753), .B1(n_754), .B2(n_755), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_443), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g951 ( .A1(n_443), .A2(n_753), .B1(n_952), .B2(n_953), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g1107 ( .A1(n_443), .A2(n_461), .B1(n_1108), .B2(n_1109), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g1589 ( .A1(n_443), .A2(n_461), .B1(n_1590), .B2(n_1591), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1957 ( .A1(n_443), .A2(n_461), .B1(n_1930), .B2(n_1958), .Y(n_1957) );
AND2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
AND2x4_ASAP7_75t_L g750 ( .A(n_444), .B(n_751), .Y(n_750) );
AND2x4_ASAP7_75t_L g762 ( .A(n_444), .B(n_751), .Y(n_762) );
INVx1_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
AND2x2_ASAP7_75t_L g745 ( .A(n_445), .B(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g455 ( .A(n_446), .Y(n_455) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_446), .Y(n_463) );
AND2x2_ASAP7_75t_L g497 ( .A(n_446), .B(n_490), .Y(n_497) );
INVx2_ASAP7_75t_L g528 ( .A(n_446), .Y(n_528) );
INVx1_ASAP7_75t_L g524 ( .A(n_447), .Y(n_524) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_447), .Y(n_729) );
BUFx6f_ASAP7_75t_L g738 ( .A(n_447), .Y(n_738) );
BUFx6f_ASAP7_75t_L g845 ( .A(n_447), .Y(n_845) );
INVx2_ASAP7_75t_L g1248 ( .A(n_447), .Y(n_1248) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g507 ( .A(n_448), .Y(n_507) );
INVx1_ASAP7_75t_L g637 ( .A(n_448), .Y(n_637) );
INVx1_ASAP7_75t_L g680 ( .A(n_448), .Y(n_680) );
BUFx6f_ASAP7_75t_L g804 ( .A(n_448), .Y(n_804) );
AND2x4_ASAP7_75t_L g448 ( .A(n_449), .B(n_450), .Y(n_448) );
INVx2_ASAP7_75t_L g467 ( .A(n_449), .Y(n_467) );
AND2x2_ASAP7_75t_L g473 ( .A(n_449), .B(n_466), .Y(n_473) );
INVx1_ASAP7_75t_L g457 ( .A(n_450), .Y(n_457) );
OR2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g477 ( .A(n_453), .Y(n_477) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g470 ( .A(n_454), .B(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g487 ( .A(n_454), .Y(n_487) );
AND2x6_ASAP7_75t_L g753 ( .A(n_454), .B(n_476), .Y(n_753) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AND2x6_ASAP7_75t_L g483 ( .A(n_455), .B(n_484), .Y(n_483) );
INVx2_ASAP7_75t_L g511 ( .A(n_456), .Y(n_511) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_456), .Y(n_1056) );
INVx1_ASAP7_75t_L g1233 ( .A(n_456), .Y(n_1233) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_456), .B(n_671), .Y(n_1513) );
OR2x2_ASAP7_75t_L g456 ( .A(n_457), .B(n_458), .Y(n_456) );
AND2x2_ASAP7_75t_L g515 ( .A(n_457), .B(n_458), .Y(n_515) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x4_ASAP7_75t_L g476 ( .A(n_459), .B(n_466), .Y(n_476) );
INVx4_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_461), .A2(n_697), .B1(n_749), .B2(n_750), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g765 ( .A1(n_461), .A2(n_753), .B1(n_766), .B2(n_767), .C(n_768), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_461), .A2(n_762), .B1(n_949), .B2(n_950), .Y(n_948) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_462), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_462), .B(n_480), .Y(n_1115) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx6_ASAP7_75t_L g633 ( .A(n_464), .Y(n_633) );
INVx2_ASAP7_75t_L g668 ( .A(n_464), .Y(n_668) );
AND2x2_ASAP7_75t_L g676 ( .A(n_464), .B(n_654), .Y(n_676) );
BUFx2_ASAP7_75t_L g734 ( .A(n_464), .Y(n_734) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
INVx1_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g482 ( .A(n_467), .Y(n_482) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AOI211xp5_ASAP7_75t_L g741 ( .A1(n_470), .A2(n_486), .B(n_742), .C(n_743), .Y(n_741) );
HB1xp67_ASAP7_75t_L g1112 ( .A(n_471), .Y(n_1112) );
HB1xp67_ASAP7_75t_L g1486 ( .A(n_471), .Y(n_1486) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x4_ASAP7_75t_L g486 ( .A(n_472), .B(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g630 ( .A(n_472), .Y(n_630) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_472), .Y(n_772) );
INVx1_ASAP7_75t_L g823 ( .A(n_472), .Y(n_823) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g663 ( .A(n_473), .Y(n_663) );
INVx2_ASAP7_75t_L g503 ( .A(n_475), .Y(n_503) );
INVx1_ASAP7_75t_L g842 ( .A(n_475), .Y(n_842) );
INVx2_ASAP7_75t_SL g897 ( .A(n_475), .Y(n_897) );
BUFx6f_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_SL g522 ( .A(n_476), .Y(n_522) );
BUFx6f_ASAP7_75t_L g636 ( .A(n_476), .Y(n_636) );
BUFx2_ASAP7_75t_L g728 ( .A(n_476), .Y(n_728) );
BUFx3_ASAP7_75t_L g827 ( .A(n_476), .Y(n_827) );
BUFx6f_ASAP7_75t_L g891 ( .A(n_476), .Y(n_891) );
BUFx2_ASAP7_75t_L g983 ( .A(n_476), .Y(n_983) );
BUFx6f_ASAP7_75t_L g1051 ( .A(n_476), .Y(n_1051) );
OAI22xp5_ASAP7_75t_L g543 ( .A1(n_478), .A2(n_544), .B1(n_547), .B2(n_551), .Y(n_543) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g746 ( .A(n_481), .Y(n_746) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g651 ( .A(n_482), .Y(n_651) );
INVx3_ASAP7_75t_L g747 ( .A(n_483), .Y(n_747) );
AOI222xp33_ASAP7_75t_L g1110 ( .A1(n_483), .A2(n_1111), .B1(n_1112), .B2(n_1113), .C1(n_1114), .C2(n_1116), .Y(n_1110) );
AOI222xp33_ASAP7_75t_L g1592 ( .A1(n_483), .A2(n_1000), .B1(n_1593), .B2(n_1594), .C1(n_1595), .C2(n_1597), .Y(n_1592) );
AOI222xp33_ASAP7_75t_L g1959 ( .A1(n_483), .A2(n_1114), .B1(n_1946), .B2(n_1947), .C1(n_1951), .C2(n_1960), .Y(n_1959) );
BUFx3_ASAP7_75t_L g660 ( .A(n_484), .Y(n_660) );
CKINVDCx8_ASAP7_75t_R g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g943 ( .A(n_486), .B(n_944), .Y(n_943) );
INVx5_ASAP7_75t_L g1106 ( .A(n_486), .Y(n_1106) );
OAI21xp33_ASAP7_75t_L g770 ( .A1(n_487), .A2(n_771), .B(n_772), .Y(n_770) );
INVx1_ASAP7_75t_SL g756 ( .A(n_488), .Y(n_756) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_491), .Y(n_488) );
AND2x4_ASAP7_75t_L g774 ( .A(n_489), .B(n_491), .Y(n_774) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
AND2x4_ASAP7_75t_L g527 ( .A(n_490), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g882 ( .A(n_491), .Y(n_882) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g498 ( .A(n_492), .Y(n_498) );
OR2x6_ASAP7_75t_L g530 ( .A(n_492), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_494), .B(n_529), .Y(n_493) );
OAI33xp33_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_499), .A3(n_508), .B1(n_516), .B2(n_520), .B3(n_525), .Y(n_494) );
INVx1_ASAP7_75t_SL g726 ( .A(n_495), .Y(n_726) );
OAI33xp33_ASAP7_75t_L g824 ( .A1(n_495), .A2(n_825), .A3(n_831), .B1(n_836), .B2(n_841), .B3(n_847), .Y(n_824) );
OAI33xp33_ASAP7_75t_L g895 ( .A1(n_495), .A2(n_847), .A3(n_896), .B1(n_900), .B2(n_903), .B3(n_909), .Y(n_895) );
OAI33xp33_ASAP7_75t_L g1048 ( .A1(n_495), .A2(n_525), .A3(n_1049), .B1(n_1055), .B2(n_1059), .B3(n_1062), .Y(n_1048) );
OAI33xp33_ASAP7_75t_L g1383 ( .A1(n_495), .A2(n_525), .A3(n_1384), .B1(n_1388), .B2(n_1392), .B3(n_1395), .Y(n_1383) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_498), .Y(n_495) );
OR2x6_ASAP7_75t_L g639 ( .A(n_496), .B(n_498), .Y(n_639) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx1_ASAP7_75t_L g808 ( .A(n_497), .Y(n_808) );
INVx2_ASAP7_75t_SL g1504 ( .A(n_497), .Y(n_1504) );
INVx1_ASAP7_75t_L g1574 ( .A(n_497), .Y(n_1574) );
BUFx3_ASAP7_75t_L g1672 ( .A(n_497), .Y(n_1672) );
INVx2_ASAP7_75t_L g626 ( .A(n_498), .Y(n_626) );
AND2x4_ASAP7_75t_L g711 ( .A(n_498), .B(n_712), .Y(n_711) );
OR2x2_ASAP7_75t_L g807 ( .A(n_498), .B(n_808), .Y(n_807) );
BUFx2_ASAP7_75t_L g1099 ( .A(n_498), .Y(n_1099) );
AND2x4_ASAP7_75t_L g1123 ( .A(n_498), .B(n_712), .Y(n_1123) );
OAI31xp33_ASAP7_75t_L g1167 ( .A1(n_498), .A2(n_1168), .A3(n_1171), .B(n_1186), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_501), .B1(n_504), .B2(n_505), .Y(n_499) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_500), .A2(n_504), .B1(n_538), .B2(n_540), .Y(n_537) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
OAI22xp5_ASAP7_75t_L g643 ( .A1(n_503), .A2(n_644), .B1(n_645), .B2(n_647), .Y(n_643) );
INVx2_ASAP7_75t_SL g1324 ( .A(n_503), .Y(n_1324) );
INVx1_ASAP7_75t_L g1968 ( .A(n_503), .Y(n_1968) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g646 ( .A(n_507), .Y(n_646) );
OR2x2_ASAP7_75t_L g1515 ( .A(n_507), .B(n_671), .Y(n_1515) );
OAI22xp33_ASAP7_75t_SL g508 ( .A1(n_509), .A2(n_510), .B1(n_512), .B2(n_513), .Y(n_508) );
OAI22xp33_ASAP7_75t_L g532 ( .A1(n_509), .A2(n_512), .B1(n_533), .B2(n_534), .Y(n_532) );
OAI22xp33_ASAP7_75t_L g831 ( .A1(n_510), .A2(n_832), .B1(n_833), .B2(n_835), .Y(n_831) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_510), .A2(n_837), .B1(n_838), .B2(n_840), .Y(n_836) );
OAI22xp33_ASAP7_75t_L g900 ( .A1(n_510), .A2(n_833), .B1(n_901), .B2(n_902), .Y(n_900) );
OAI22xp33_ASAP7_75t_L g1059 ( .A1(n_510), .A2(n_517), .B1(n_1060), .B2(n_1061), .Y(n_1059) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g888 ( .A(n_511), .Y(n_888) );
INVx2_ASAP7_75t_L g904 ( .A(n_511), .Y(n_904) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g907 ( .A(n_514), .Y(n_907) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx2_ASAP7_75t_L g518 ( .A(n_515), .Y(n_518) );
BUFx2_ASAP7_75t_L g834 ( .A(n_515), .Y(n_834) );
BUFx4f_ASAP7_75t_L g839 ( .A(n_515), .Y(n_839) );
INVx1_ASAP7_75t_L g947 ( .A(n_515), .Y(n_947) );
OAI22xp33_ASAP7_75t_L g1055 ( .A1(n_517), .A2(n_1056), .B1(n_1057), .B2(n_1058), .Y(n_1055) );
BUFx3_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
OR2x6_ASAP7_75t_L g682 ( .A(n_518), .B(n_670), .Y(n_682) );
OAI22xp33_ASAP7_75t_L g1392 ( .A1(n_518), .A2(n_1232), .B1(n_1393), .B2(n_1394), .Y(n_1392) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_521), .A2(n_522), .B1(n_523), .B2(n_524), .Y(n_520) );
INVx2_ASAP7_75t_L g674 ( .A(n_522), .Y(n_674) );
INVx1_ASAP7_75t_L g998 ( .A(n_522), .Y(n_998) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_526), .A2(n_628), .B1(n_638), .B2(n_640), .C(n_648), .Y(n_627) );
AOI33xp33_ASAP7_75t_L g1136 ( .A1(n_526), .A2(n_1137), .A3(n_1138), .B1(n_1143), .B2(n_1145), .B3(n_1147), .Y(n_1136) );
BUFx4f_ASAP7_75t_L g1240 ( .A(n_526), .Y(n_1240) );
BUFx4f_ASAP7_75t_L g1377 ( .A(n_526), .Y(n_1377) );
INVx2_ASAP7_75t_L g1488 ( .A(n_527), .Y(n_1488) );
INVx2_ASAP7_75t_SL g1564 ( .A(n_527), .Y(n_1564) );
CKINVDCx5p33_ASAP7_75t_R g1668 ( .A(n_527), .Y(n_1668) );
AND2x4_ASAP7_75t_L g654 ( .A(n_528), .B(n_655), .Y(n_654) );
OAI33xp33_ASAP7_75t_L g529 ( .A1(n_530), .A2(n_532), .A3(n_537), .B1(n_543), .B2(n_552), .B3(n_559), .Y(n_529) );
OAI33xp33_ASAP7_75t_L g1458 ( .A1(n_530), .A2(n_1459), .A3(n_1465), .B1(n_1471), .B2(n_1474), .B3(n_1477), .Y(n_1458) );
OAI33xp33_ASAP7_75t_L g1534 ( .A1(n_530), .A2(n_1477), .A3(n_1535), .B1(n_1540), .B2(n_1547), .B3(n_1553), .Y(n_1534) );
INVx1_ASAP7_75t_L g1639 ( .A(n_530), .Y(n_1639) );
OAI22xp33_ASAP7_75t_L g552 ( .A1(n_533), .A2(n_553), .B1(n_554), .B2(n_558), .Y(n_552) );
INVx1_ASAP7_75t_L g1176 ( .A(n_533), .Y(n_1176) );
INVx1_ASAP7_75t_L g1197 ( .A(n_533), .Y(n_1197) );
OAI221xp5_ASAP7_75t_L g1302 ( .A1(n_533), .A2(n_556), .B1(n_864), .B2(n_1303), .C(n_1304), .Y(n_1302) );
OAI221xp5_ASAP7_75t_L g1306 ( .A1(n_533), .A2(n_581), .B1(n_1087), .B2(n_1292), .C(n_1307), .Y(n_1306) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_533), .A2(n_556), .B1(n_1081), .B2(n_1389), .C(n_1391), .Y(n_1411) );
BUFx2_ASAP7_75t_L g1654 ( .A(n_533), .Y(n_1654) );
OAI221xp5_ASAP7_75t_L g1194 ( .A1(n_534), .A2(n_1081), .B1(n_1195), .B2(n_1196), .C(n_1198), .Y(n_1194) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_536), .B(n_599), .Y(n_598) );
OR2x6_ASAP7_75t_L g865 ( .A(n_536), .B(n_605), .Y(n_865) );
OR2x2_ASAP7_75t_L g1260 ( .A(n_536), .B(n_605), .Y(n_1260) );
HB1xp67_ASAP7_75t_L g1539 ( .A(n_536), .Y(n_1539) );
OAI22xp5_ASAP7_75t_L g918 ( .A1(n_538), .A2(n_898), .B1(n_899), .B2(n_919), .Y(n_918) );
OAI221xp5_ASAP7_75t_L g1413 ( .A1(n_538), .A2(n_1414), .B1(n_1415), .B2(n_1417), .C(n_1418), .Y(n_1413) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g1267 ( .A(n_540), .Y(n_1267) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x4_ASAP7_75t_L g616 ( .A(n_541), .B(n_617), .Y(n_616) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
OAI22xp5_ASAP7_75t_L g858 ( .A1(n_544), .A2(n_828), .B1(n_830), .B2(n_859), .Y(n_858) );
OAI22xp5_ASAP7_75t_L g1298 ( .A1(n_544), .A2(n_1299), .B1(n_1300), .B2(n_1301), .Y(n_1298) );
INVx2_ASAP7_75t_SL g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g1074 ( .A(n_545), .Y(n_1074) );
INVx2_ASAP7_75t_L g1469 ( .A(n_545), .Y(n_1469) );
INVx2_ASAP7_75t_L g1542 ( .A(n_545), .Y(n_1542) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g1189 ( .A(n_546), .Y(n_1189) );
OAI22xp5_ASAP7_75t_L g1645 ( .A1(n_547), .A2(n_1646), .B1(n_1647), .B2(n_1648), .Y(n_1645) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g798 ( .A(n_549), .Y(n_798) );
INVx2_ASAP7_75t_L g1192 ( .A(n_549), .Y(n_1192) );
INVx3_ASAP7_75t_L g1312 ( .A(n_549), .Y(n_1312) );
INVx2_ASAP7_75t_L g1416 ( .A(n_549), .Y(n_1416) );
INVx2_ASAP7_75t_L g1551 ( .A(n_549), .Y(n_1551) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
INVx3_ASAP7_75t_L g577 ( .A(n_550), .Y(n_577) );
INVx3_ASAP7_75t_L g920 ( .A(n_550), .Y(n_920) );
OAI221xp5_ASAP7_75t_L g1084 ( .A1(n_554), .A2(n_862), .B1(n_1085), .B2(n_1086), .C(n_1087), .Y(n_1084) );
OAI22xp33_ASAP7_75t_L g1553 ( .A1(n_554), .A2(n_1537), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx2_ASAP7_75t_L g1173 ( .A(n_555), .Y(n_1173) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_556), .A2(n_832), .B1(n_835), .B2(n_862), .C(n_864), .Y(n_861) );
BUFx3_ASAP7_75t_L g922 ( .A(n_556), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_556), .B(n_1029), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1464 ( .A(n_556), .Y(n_1464) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AOI33xp33_ASAP7_75t_L g710 ( .A1(n_560), .A2(n_711), .A3(n_713), .B1(n_716), .B2(n_720), .B3(n_722), .Y(n_710) );
AOI33xp33_ASAP7_75t_L g1121 ( .A1(n_560), .A2(n_1122), .A3(n_1124), .B1(n_1127), .B2(n_1130), .B3(n_1135), .Y(n_1121) );
AOI33xp33_ASAP7_75t_L g1609 ( .A1(n_560), .A2(n_1122), .A3(n_1610), .B1(n_1611), .B2(n_1612), .B3(n_1613), .Y(n_1609) );
INVx6_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx5_ASAP7_75t_L g800 ( .A(n_561), .Y(n_800) );
OR2x6_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NAND2x1p5_ASAP7_75t_L g653 ( .A(n_562), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
OR2x2_ASAP7_75t_L g670 ( .A(n_563), .B(n_671), .Y(n_670) );
AND2x4_ASAP7_75t_L g1440 ( .A(n_563), .B(n_611), .Y(n_1440) );
BUFx2_ASAP7_75t_L g594 ( .A(n_564), .Y(n_594) );
INVx2_ASAP7_75t_L g1089 ( .A(n_564), .Y(n_1089) );
NAND4xp25_ASAP7_75t_L g569 ( .A(n_570), .B(n_627), .C(n_665), .D(n_677), .Y(n_569) );
OAI31xp33_ASAP7_75t_L g570 ( .A1(n_571), .A2(n_608), .A3(n_619), .B(n_625), .Y(n_570) );
OAI221xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_579), .B1(n_585), .B2(n_589), .C(n_595), .Y(n_571) );
OAI22xp5_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B1(n_576), .B2(n_578), .Y(n_572) );
OAI22xp5_ASAP7_75t_L g585 ( .A1(n_573), .A2(n_586), .B1(n_587), .B2(n_588), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_573), .A2(n_587), .B1(n_1024), .B2(n_1025), .Y(n_1023) );
BUFx2_ASAP7_75t_L g1179 ( .A(n_573), .Y(n_1179) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_573), .A2(n_859), .B1(n_1258), .B2(n_1259), .Y(n_1257) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g868 ( .A(n_574), .Y(n_868) );
INVx1_ASAP7_75t_L g1310 ( .A(n_574), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1409 ( .A(n_574), .Y(n_1409) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_575), .A2(n_578), .B1(n_635), .B2(n_637), .Y(n_634) );
INVx2_ASAP7_75t_L g721 ( .A(n_576), .Y(n_721) );
INVx2_ASAP7_75t_SL g791 ( .A(n_576), .Y(n_791) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx2_ASAP7_75t_L g587 ( .A(n_577), .Y(n_587) );
INVx2_ASAP7_75t_L g971 ( .A(n_577), .Y(n_971) );
INVx1_ASAP7_75t_L g1546 ( .A(n_577), .Y(n_1546) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B(n_582), .Y(n_579) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_581), .A2(n_1057), .B1(n_1058), .B2(n_1079), .C(n_1081), .Y(n_1078) );
BUFx2_ASAP7_75t_L g714 ( .A(n_583), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_583), .B(n_854), .Y(n_853) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx2_ASAP7_75t_L g593 ( .A(n_584), .Y(n_593) );
INVx2_ASAP7_75t_SL g1337 ( .A(n_584), .Y(n_1337) );
AOI222xp33_ASAP7_75t_L g665 ( .A1(n_586), .A2(n_596), .B1(n_666), .B2(n_672), .C1(n_673), .C2(n_675), .Y(n_665) );
INVx1_ASAP7_75t_L g719 ( .A(n_587), .Y(n_719) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_588), .A2(n_590), .B1(n_678), .B2(n_681), .Y(n_677) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B(n_592), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g1474 ( .A1(n_591), .A2(n_862), .B1(n_1475), .B2(n_1476), .Y(n_1474) );
OAI21xp5_ASAP7_75t_SL g1950 ( .A1(n_591), .A2(n_1951), .B(n_1952), .Y(n_1950) );
BUFx3_ASAP7_75t_L g1125 ( .A(n_593), .Y(n_1125) );
A2O1A1Ixp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_597), .B(n_598), .C(n_604), .Y(n_595) );
INVx1_ASAP7_75t_L g1615 ( .A(n_597), .Y(n_1615) );
NAND2x1p5_ASAP7_75t_L g1455 ( .A(n_602), .B(n_1452), .Y(n_1455) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x6_ASAP7_75t_L g880 ( .A(n_603), .B(n_605), .Y(n_880) );
A2O1A1Ixp33_ASAP7_75t_L g1026 ( .A1(n_604), .A2(n_793), .B(n_1027), .C(n_1028), .Y(n_1026) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g854 ( .A(n_605), .Y(n_854) );
INVx1_ASAP7_75t_L g1341 ( .A(n_605), .Y(n_1341) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx3_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_610), .A2(n_616), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
INVx3_ASAP7_75t_L g1169 ( .A(n_610), .Y(n_1169) );
AOI22xp33_ASAP7_75t_L g1342 ( .A1(n_610), .A2(n_616), .B1(n_1343), .B2(n_1344), .Y(n_1342) );
AOI22xp33_ASAP7_75t_L g1934 ( .A1(n_610), .A2(n_616), .B1(n_1935), .B2(n_1936), .Y(n_1934) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g618 ( .A(n_611), .Y(n_618) );
INVx1_ASAP7_75t_L g718 ( .A(n_612), .Y(n_718) );
BUFx2_ASAP7_75t_L g974 ( .A(n_612), .Y(n_974) );
BUFx6f_ASAP7_75t_L g1018 ( .A(n_612), .Y(n_1018) );
BUFx2_ASAP7_75t_L g1128 ( .A(n_612), .Y(n_1128) );
BUFx6f_ASAP7_75t_L g1133 ( .A(n_612), .Y(n_1133) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx3_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx3_ASAP7_75t_L g1170 ( .A(n_616), .Y(n_1170) );
AND2x4_ASAP7_75t_L g623 ( .A(n_617), .B(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
CKINVDCx6p67_ASAP7_75t_R g620 ( .A(n_621), .Y(n_620) );
AOI22xp5_ASAP7_75t_L g1016 ( .A1(n_621), .A2(n_1017), .B1(n_1019), .B2(n_1020), .Y(n_1016) );
AOI221xp5_ASAP7_75t_L g1345 ( .A1(n_621), .A2(n_1346), .B1(n_1348), .B2(n_1349), .C(n_1350), .Y(n_1345) );
AOI222xp33_ASAP7_75t_L g1929 ( .A1(n_621), .A2(n_623), .B1(n_1930), .B2(n_1931), .C1(n_1932), .C2(n_1933), .Y(n_1929) );
INVx8_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI221xp5_ASAP7_75t_L g1330 ( .A1(n_623), .A2(n_1331), .B1(n_1334), .B2(n_1338), .C(n_1339), .Y(n_1330) );
INVx1_ASAP7_75t_L g979 ( .A(n_624), .Y(n_979) );
OAI31xp33_ASAP7_75t_L g1252 ( .A1(n_625), .A2(n_1253), .A3(n_1254), .B(n_1261), .Y(n_1252) );
OAI31xp33_ASAP7_75t_L g1404 ( .A1(n_625), .A2(n_1405), .A3(n_1406), .B(n_1412), .Y(n_1404) );
INVx1_ASAP7_75t_L g1479 ( .A(n_625), .Y(n_1479) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
NOR2xp67_ASAP7_75t_L g852 ( .A(n_626), .B(n_853), .Y(n_852) );
INVx3_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx6f_ASAP7_75t_L g642 ( .A(n_633), .Y(n_642) );
INVx2_ASAP7_75t_L g732 ( .A(n_633), .Y(n_732) );
INVx2_ASAP7_75t_L g751 ( .A(n_633), .Y(n_751) );
INVx1_ASAP7_75t_L g811 ( .A(n_633), .Y(n_811) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_633), .Y(n_1004) );
INVx2_ASAP7_75t_L g1140 ( .A(n_633), .Y(n_1140) );
INVx1_ASAP7_75t_L g1371 ( .A(n_633), .Y(n_1371) );
INVx1_ASAP7_75t_L g1319 ( .A(n_635), .Y(n_1319) );
INVx2_ASAP7_75t_SL g635 ( .A(n_636), .Y(n_635) );
BUFx3_ASAP7_75t_L g1144 ( .A(n_636), .Y(n_1144) );
AND2x4_ASAP7_75t_L g1482 ( .A(n_636), .B(n_1483), .Y(n_1482) );
INVx1_ASAP7_75t_L g1567 ( .A(n_636), .Y(n_1567) );
OAI22xp33_ASAP7_75t_L g896 ( .A1(n_637), .A2(n_897), .B1(n_898), .B2(n_899), .Y(n_896) );
INVx1_ASAP7_75t_L g1238 ( .A(n_637), .Y(n_1238) );
INVx1_ASAP7_75t_L g1376 ( .A(n_637), .Y(n_1376) );
INVx1_ASAP7_75t_L g1399 ( .A(n_637), .Y(n_1399) );
INVx2_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g1137 ( .A(n_639), .Y(n_1137) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_639), .Y(n_1206) );
OAI22xp5_ASAP7_75t_SL g1229 ( .A1(n_639), .A2(n_1230), .B1(n_1239), .B2(n_1241), .Y(n_1229) );
OAI22xp5_ASAP7_75t_L g1963 ( .A1(n_639), .A2(n_1239), .B1(n_1964), .B2(n_1969), .Y(n_1963) );
INVx4_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g1485 ( .A(n_642), .Y(n_1485) );
INVx1_ASAP7_75t_L g984 ( .A(n_645), .Y(n_984) );
INVx2_ASAP7_75t_SL g1209 ( .A(n_645), .Y(n_1209) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
BUFx2_ASAP7_75t_L g1568 ( .A(n_646), .Y(n_1568) );
INVx2_ASAP7_75t_L g1007 ( .A(n_649), .Y(n_1007) );
INVx1_ASAP7_75t_L g1204 ( .A(n_649), .Y(n_1204) );
INVx1_ASAP7_75t_L g1251 ( .A(n_649), .Y(n_1251) );
INVx2_ASAP7_75t_L g1362 ( .A(n_649), .Y(n_1362) );
NAND2x1p5_ASAP7_75t_L g649 ( .A(n_650), .B(n_652), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g1495 ( .A(n_651), .Y(n_1495) );
INVx2_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
OR2x6_ASAP7_75t_L g658 ( .A(n_653), .B(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g664 ( .A(n_653), .Y(n_664) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_653), .B(n_659), .Y(n_1067) );
AND2x4_ASAP7_75t_L g1494 ( .A(n_654), .B(n_1495), .Y(n_1494) );
AND2x2_ASAP7_75t_L g1497 ( .A(n_654), .B(n_660), .Y(n_1497) );
INVx1_ASAP7_75t_L g1510 ( .A(n_654), .Y(n_1510) );
AND2x4_ASAP7_75t_L g1663 ( .A(n_654), .B(n_1495), .Y(n_1663) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g1009 ( .A(n_658), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1570 ( .A(n_659), .B(n_1510), .Y(n_1570) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
INVx1_ASAP7_75t_L g1216 ( .A(n_661), .Y(n_1216) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_662), .B(n_664), .Y(n_661) );
HB1xp67_ASAP7_75t_L g1374 ( .A(n_662), .Y(n_1374) );
BUFx2_ASAP7_75t_SL g1573 ( .A(n_662), .Y(n_1573) );
BUFx6f_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g736 ( .A(n_663), .Y(n_736) );
BUFx4f_ASAP7_75t_L g1000 ( .A(n_663), .Y(n_1000) );
INVx2_ASAP7_75t_SL g1212 ( .A(n_663), .Y(n_1212) );
BUFx3_ASAP7_75t_L g1322 ( .A(n_663), .Y(n_1322) );
AND2x4_ASAP7_75t_L g1507 ( .A(n_663), .B(n_1483), .Y(n_1507) );
INVx1_ASAP7_75t_L g1961 ( .A(n_663), .Y(n_1961) );
AND2x2_ASAP7_75t_L g821 ( .A(n_664), .B(n_822), .Y(n_821) );
AOI222xp33_ASAP7_75t_L g1032 ( .A1(n_666), .A2(n_675), .B1(n_678), .B2(n_1024), .C1(n_1027), .C2(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1219 ( .A1(n_666), .A2(n_673), .B1(n_1177), .B2(n_1180), .Y(n_1219) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_666), .A2(n_673), .B1(n_1291), .B2(n_1292), .C(n_1293), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_666), .A2(n_673), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_669), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g1146 ( .A(n_668), .Y(n_1146) );
AND2x2_ASAP7_75t_L g673 ( .A(n_669), .B(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OR2x6_ASAP7_75t_L g679 ( .A(n_670), .B(n_680), .Y(n_679) );
OR2x2_ASAP7_75t_L g885 ( .A(n_670), .B(n_680), .Y(n_885) );
OR2x2_ASAP7_75t_L g887 ( .A(n_670), .B(n_888), .Y(n_887) );
OR2x2_ASAP7_75t_L g889 ( .A(n_670), .B(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g1483 ( .A(n_671), .Y(n_1483) );
AOI22xp5_ASAP7_75t_L g1034 ( .A1(n_673), .A2(n_681), .B1(n_1025), .B2(n_1035), .Y(n_1034) );
OR2x6_ASAP7_75t_L g851 ( .A(n_675), .B(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g1520 ( .A(n_675), .Y(n_1520) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_678), .A2(n_681), .B1(n_1174), .B2(n_1181), .Y(n_1218) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_678), .A2(n_681), .B1(n_1356), .B2(n_1357), .Y(n_1355) );
CKINVDCx6p67_ASAP7_75t_R g678 ( .A(n_679), .Y(n_678) );
OAI22xp5_ASAP7_75t_L g1062 ( .A1(n_680), .A2(n_826), .B1(n_1063), .B2(n_1064), .Y(n_1062) );
INVx2_ASAP7_75t_L g1491 ( .A(n_680), .Y(n_1491) );
CKINVDCx6p67_ASAP7_75t_R g681 ( .A(n_682), .Y(n_681) );
OA22x2_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_757), .B1(n_758), .B2(n_815), .Y(n_683) );
INVx1_ASAP7_75t_L g815 ( .A(n_684), .Y(n_815) );
XNOR2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g1726 ( .A1(n_685), .A2(n_1717), .B1(n_1727), .B2(n_1728), .Y(n_1726) );
AOI211xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_709), .C(n_740), .Y(n_686) );
AOI221x1_ASAP7_75t_L g759 ( .A1(n_687), .A2(n_760), .B1(n_773), .B2(n_775), .C(n_788), .Y(n_759) );
AOI221x1_ASAP7_75t_L g941 ( .A1(n_687), .A2(n_773), .B1(n_942), .B2(n_954), .C(n_965), .Y(n_941) );
CKINVDCx16_ASAP7_75t_R g687 ( .A(n_688), .Y(n_687) );
AOI31xp33_ASAP7_75t_L g1598 ( .A1(n_688), .A2(n_1599), .A3(n_1603), .B(n_1606), .Y(n_1598) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_692), .B1(n_693), .B2(n_694), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g776 ( .A1(n_692), .A2(n_694), .B1(n_777), .B2(n_778), .Y(n_776) );
AOI22xp33_ASAP7_75t_L g955 ( .A1(n_692), .A2(n_694), .B1(n_956), .B2(n_957), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1603 ( .A1(n_692), .A2(n_694), .B1(n_1604), .B2(n_1605), .Y(n_1603) );
INVx4_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx5_ASAP7_75t_L g964 ( .A(n_699), .Y(n_964) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_SL g1126 ( .A(n_703), .Y(n_1126) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
BUFx6f_ASAP7_75t_L g715 ( .A(n_704), .Y(n_715) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g709 ( .A(n_710), .B(n_725), .Y(n_709) );
NAND3xp33_ASAP7_75t_L g789 ( .A(n_711), .B(n_790), .C(n_792), .Y(n_789) );
NAND3xp33_ASAP7_75t_L g972 ( .A(n_711), .B(n_973), .C(n_977), .Y(n_972) );
BUFx2_ASAP7_75t_SL g864 ( .A(n_712), .Y(n_864) );
INVx1_ASAP7_75t_L g1082 ( .A(n_712), .Y(n_1082) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g795 ( .A(n_724), .Y(n_795) );
HB1xp67_ASAP7_75t_L g968 ( .A(n_724), .Y(n_968) );
AOI33xp33_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_727), .A3(n_730), .B1(n_733), .B2(n_737), .B3(n_739), .Y(n_725) );
AOI33xp33_ASAP7_75t_L g996 ( .A1(n_726), .A2(n_739), .A3(n_997), .B1(n_999), .B2(n_1001), .B3(n_1005), .Y(n_996) );
BUFx6f_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
NAND3xp33_ASAP7_75t_L g809 ( .A(n_739), .B(n_810), .C(n_812), .Y(n_809) );
INVx1_ASAP7_75t_L g847 ( .A(n_739), .Y(n_847) );
INVx1_ASAP7_75t_L g989 ( .A(n_739), .Y(n_989) );
AOI31xp33_ASAP7_75t_SL g740 ( .A1(n_741), .A2(n_748), .A3(n_752), .B(n_756), .Y(n_740) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g769 ( .A(n_745), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1117 ( .A1(n_753), .A2(n_762), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_753), .A2(n_762), .B1(n_1587), .B2(n_1588), .Y(n_1586) );
AOI22xp33_ASAP7_75t_L g1954 ( .A1(n_753), .A2(n_762), .B1(n_1955), .B2(n_1956), .Y(n_1954) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g814 ( .A(n_759), .Y(n_814) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_765), .Y(n_760) );
INVx1_ASAP7_75t_L g1142 ( .A(n_772), .Y(n_1142) );
AND2x4_ASAP7_75t_L g1508 ( .A(n_772), .B(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1561 ( .A(n_772), .Y(n_1561) );
AOI211x1_ASAP7_75t_L g1584 ( .A1(n_773), .A2(n_1585), .B(n_1598), .C(n_1608), .Y(n_1584) );
AOI221x1_ASAP7_75t_SL g1927 ( .A1(n_773), .A2(n_1099), .B1(n_1928), .B2(n_1953), .C(n_1963), .Y(n_1927) );
BUFx6f_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AOI211x1_ASAP7_75t_SL g1104 ( .A1(n_774), .A2(n_1105), .B(n_1120), .C(n_1149), .Y(n_1104) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NAND4xp25_ASAP7_75t_L g788 ( .A(n_789), .B(n_796), .C(n_801), .D(n_809), .Y(n_788) );
INVx1_ASAP7_75t_L g1093 ( .A(n_791), .Y(n_1093) );
INVx2_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
NAND3xp33_ASAP7_75t_L g796 ( .A(n_797), .B(n_799), .C(n_800), .Y(n_796) );
NAND3xp33_ASAP7_75t_L g966 ( .A(n_800), .B(n_967), .C(n_969), .Y(n_966) );
CKINVDCx8_ASAP7_75t_R g1477 ( .A(n_800), .Y(n_1477) );
NAND3xp33_ASAP7_75t_L g801 ( .A(n_802), .B(n_805), .C(n_806), .Y(n_801) );
BUFx6f_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g829 ( .A(n_804), .Y(n_829) );
INVx1_ASAP7_75t_L g1053 ( .A(n_804), .Y(n_1053) );
NAND3xp33_ASAP7_75t_L g980 ( .A(n_806), .B(n_981), .C(n_982), .Y(n_980) );
INVx3_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_937), .Y(n_816) );
XOR2xp5_ASAP7_75t_L g817 ( .A(n_818), .B(n_892), .Y(n_817) );
AND4x1_ASAP7_75t_L g819 ( .A(n_820), .B(n_849), .C(n_855), .D(n_883), .Y(n_819) );
NOR3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_824), .C(n_848), .Y(n_820) );
NOR3xp33_ASAP7_75t_L g894 ( .A(n_821), .B(n_895), .C(n_912), .Y(n_894) );
AOI221xp5_ASAP7_75t_L g1006 ( .A1(n_821), .A2(n_1007), .B1(n_1008), .B2(n_1009), .C(n_1010), .Y(n_1006) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_821), .Y(n_1047) );
BUFx2_ASAP7_75t_L g1228 ( .A(n_821), .Y(n_1228) );
AOI221xp5_ASAP7_75t_L g1287 ( .A1(n_821), .A2(n_1009), .B1(n_1251), .B2(n_1288), .C(n_1289), .Y(n_1287) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1501 ( .A(n_823), .Y(n_1501) );
OAI22xp33_ASAP7_75t_L g825 ( .A1(n_826), .A2(n_828), .B1(n_829), .B2(n_830), .Y(n_825) );
OAI22xp33_ASAP7_75t_L g1384 ( .A1(n_826), .A2(n_1385), .B1(n_1386), .B2(n_1387), .Y(n_1384) );
INVx2_ASAP7_75t_SL g826 ( .A(n_827), .Y(n_826) );
BUFx3_ASAP7_75t_L g1246 ( .A(n_827), .Y(n_1246) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_829), .A2(n_842), .B1(n_910), .B2(n_911), .Y(n_909) );
INVx2_ASAP7_75t_SL g833 ( .A(n_834), .Y(n_833) );
BUFx2_ASAP7_75t_L g1236 ( .A(n_838), .Y(n_1236) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g1243 ( .A(n_839), .Y(n_1243) );
INVx2_ASAP7_75t_SL g1665 ( .A(n_839), .Y(n_1665) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B1(n_844), .B2(n_846), .Y(n_841) );
INVx2_ASAP7_75t_SL g844 ( .A(n_845), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g849 ( .A(n_850), .B(n_851), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_851), .B(n_914), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_851), .B(n_1069), .Y(n_1068) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_851), .B(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1225 ( .A(n_851), .B(n_1226), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1294 ( .A(n_851), .B(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1359 ( .A(n_851), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_851), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1931 ( .A(n_853), .Y(n_1931) );
AND2x2_ASAP7_75t_L g876 ( .A(n_854), .B(n_877), .Y(n_876) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_854), .B(n_877), .Y(n_1184) );
OAI31xp33_ASAP7_75t_L g855 ( .A1(n_856), .A2(n_857), .A3(n_866), .B(n_881), .Y(n_855) );
INVx2_ASAP7_75t_SL g1129 ( .A(n_859), .Y(n_1129) );
INVx2_ASAP7_75t_L g1949 ( .A(n_859), .Y(n_1949) );
INVx4_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_SL g870 ( .A(n_860), .Y(n_870) );
INVx2_ASAP7_75t_SL g928 ( .A(n_860), .Y(n_928) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_860), .Y(n_1134) );
INVx2_ASAP7_75t_SL g1300 ( .A(n_860), .Y(n_1300) );
INVx2_ASAP7_75t_SL g1333 ( .A(n_860), .Y(n_1333) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g1461 ( .A(n_863), .Y(n_1461) );
INVx2_ASAP7_75t_L g1350 ( .A(n_865), .Y(n_1350) );
OAI221xp5_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_870), .B2(n_871), .C(n_872), .Y(n_867) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_868), .A2(n_927), .B1(n_928), .B2(n_929), .C(n_930), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1178 ( .A1(n_870), .A2(n_1179), .B1(n_1180), .B2(n_1181), .Y(n_1178) );
OAI22xp5_ASAP7_75t_L g1471 ( .A1(n_870), .A2(n_1467), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
AND2x6_ASAP7_75t_L g1442 ( .A(n_873), .B(n_1440), .Y(n_1442) );
NAND2x1p5_ASAP7_75t_L g1457 ( .A(n_873), .B(n_1452), .Y(n_1457) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_875), .A2(n_876), .B1(n_878), .B2(n_879), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g931 ( .A1(n_876), .A2(n_879), .B1(n_932), .B2(n_933), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_876), .A2(n_879), .B1(n_1095), .B2(n_1096), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_879), .A2(n_1183), .B1(n_1184), .B2(n_1185), .Y(n_1182) );
AOI22xp33_ASAP7_75t_L g1270 ( .A1(n_879), .A2(n_1184), .B1(n_1271), .B2(n_1272), .Y(n_1270) );
AOI22xp5_ASAP7_75t_L g1314 ( .A1(n_879), .A2(n_1184), .B1(n_1288), .B2(n_1289), .Y(n_1314) );
AOI22xp33_ASAP7_75t_L g1419 ( .A1(n_879), .A2(n_1184), .B1(n_1420), .B2(n_1421), .Y(n_1419) );
AOI22xp5_ASAP7_75t_L g1945 ( .A1(n_879), .A2(n_1184), .B1(n_1946), .B2(n_1947), .Y(n_1945) );
CKINVDCx11_ASAP7_75t_R g879 ( .A(n_880), .Y(n_879) );
OAI31xp33_ASAP7_75t_L g915 ( .A1(n_881), .A2(n_916), .A3(n_917), .B(n_925), .Y(n_915) );
OAI21xp5_ASAP7_75t_L g1011 ( .A1(n_881), .A2(n_1012), .B(n_1021), .Y(n_1011) );
OAI31xp33_ASAP7_75t_L g1296 ( .A1(n_881), .A2(n_1297), .A3(n_1305), .B(n_1315), .Y(n_1296) );
BUFx8_ASAP7_75t_SL g881 ( .A(n_882), .Y(n_881) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .Y(n_883) );
INVx1_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
BUFx2_ASAP7_75t_L g1148 ( .A(n_891), .Y(n_1148) );
BUFx4f_ASAP7_75t_L g1208 ( .A(n_891), .Y(n_1208) );
AND4x1_ASAP7_75t_L g893 ( .A(n_894), .B(n_913), .C(n_915), .D(n_934), .Y(n_893) );
OAI21xp33_ASAP7_75t_SL g921 ( .A1(n_902), .A2(n_922), .B(n_923), .Y(n_921) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_905), .B1(n_906), .B2(n_908), .Y(n_903) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_904), .A2(n_1242), .B1(n_1243), .B2(n_1244), .C(n_1245), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1969 ( .A1(n_906), .A2(n_1232), .B1(n_1932), .B2(n_1933), .C(n_1970), .Y(n_1969) );
INVx2_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g1942 ( .A1(n_919), .A2(n_1548), .B1(n_1943), .B2(n_1944), .Y(n_1942) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_L g976 ( .A(n_920), .Y(n_976) );
AND2x4_ASAP7_75t_L g1439 ( .A(n_920), .B(n_1440), .Y(n_1439) );
NOR2xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_936), .Y(n_934) );
OAI22x1_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_939), .B1(n_991), .B2(n_992), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_939), .Y(n_938) );
INVx1_ASAP7_75t_L g990 ( .A(n_941), .Y(n_990) );
NAND3xp33_ASAP7_75t_L g942 ( .A(n_943), .B(n_948), .C(n_951), .Y(n_942) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
HB1xp67_ASAP7_75t_L g1390 ( .A(n_947), .Y(n_1390) );
NAND4xp25_ASAP7_75t_L g965 ( .A(n_966), .B(n_972), .C(n_980), .D(n_985), .Y(n_965) );
INVx1_ASAP7_75t_L g1410 ( .A(n_970), .Y(n_1410) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
INVx1_ASAP7_75t_L g975 ( .A(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx1_ASAP7_75t_L g1152 ( .A(n_979), .Y(n_1152) );
NAND3xp33_ASAP7_75t_L g985 ( .A(n_986), .B(n_987), .C(n_988), .Y(n_985) );
AOI33xp33_ASAP7_75t_L g1205 ( .A1(n_988), .A2(n_1206), .A3(n_1207), .B1(n_1210), .B2(n_1213), .B3(n_1214), .Y(n_1205) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx2_ASAP7_75t_SL g991 ( .A(n_992), .Y(n_991) );
INVx2_ASAP7_75t_L g993 ( .A(n_994), .Y(n_993) );
NAND4xp75_ASAP7_75t_L g994 ( .A(n_995), .B(n_1011), .C(n_1032), .D(n_1034), .Y(n_994) );
AND2x2_ASAP7_75t_L g995 ( .A(n_996), .B(n_1006), .Y(n_995) );
INVx2_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1007), .Y(n_1066) );
AOI22xp5_ASAP7_75t_L g1203 ( .A1(n_1009), .A2(n_1183), .B1(n_1185), .B2(n_1204), .Y(n_1203) );
AOI22xp5_ASAP7_75t_L g1361 ( .A1(n_1009), .A2(n_1362), .B1(n_1363), .B2(n_1364), .Y(n_1361) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1016), .Y(n_1012) );
NAND2x1p5_ASAP7_75t_L g1340 ( .A(n_1030), .B(n_1341), .Y(n_1340) );
NAND2x1_ASAP7_75t_SL g1451 ( .A(n_1030), .B(n_1452), .Y(n_1451) );
INVx2_ASAP7_75t_L g1030 ( .A(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1038), .Y(n_1037) );
XNOR2xp5_ASAP7_75t_L g1038 ( .A(n_1039), .B(n_1164), .Y(n_1038) );
AOI22xp5_ASAP7_75t_L g1039 ( .A1(n_1040), .A2(n_1041), .B1(n_1103), .B2(n_1163), .Y(n_1039) );
INVx1_ASAP7_75t_L g1040 ( .A(n_1041), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_1044), .Y(n_1043) );
AND4x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1068), .C(n_1070), .D(n_1100), .Y(n_1045) );
NOR3xp33_ASAP7_75t_SL g1046 ( .A(n_1047), .B(n_1048), .C(n_1065), .Y(n_1046) );
NOR3xp33_ASAP7_75t_L g1382 ( .A(n_1047), .B(n_1383), .C(n_1401), .Y(n_1382) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_1050), .A2(n_1052), .B1(n_1053), .B2(n_1054), .Y(n_1049) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
BUFx2_ASAP7_75t_L g1367 ( .A(n_1051), .Y(n_1367) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1051), .Y(n_1396) );
BUFx3_ASAP7_75t_L g1500 ( .A(n_1051), .Y(n_1500) );
OAI22xp5_ASAP7_75t_L g1073 ( .A1(n_1052), .A2(n_1054), .B1(n_1074), .B2(n_1075), .Y(n_1073) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1053), .Y(n_1320) );
OAI22xp33_ASAP7_75t_L g1388 ( .A1(n_1056), .A2(n_1389), .B1(n_1390), .B2(n_1391), .Y(n_1388) );
OAI31xp33_ASAP7_75t_L g1070 ( .A1(n_1071), .A2(n_1072), .A3(n_1083), .B(n_1097), .Y(n_1070) );
OAI22xp5_ASAP7_75t_SL g1090 ( .A1(n_1074), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
OAI22xp5_ASAP7_75t_L g1465 ( .A1(n_1075), .A2(n_1466), .B1(n_1467), .B2(n_1470), .Y(n_1465) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx1_ASAP7_75t_L g1076 ( .A(n_1077), .Y(n_1076) );
BUFx2_ASAP7_75t_L g1537 ( .A(n_1079), .Y(n_1537) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1255 ( .A1(n_1081), .A2(n_1175), .B1(n_1234), .B2(n_1235), .C(n_1256), .Y(n_1255) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_1087), .A2(n_1173), .B1(n_1174), .B2(n_1175), .C(n_1177), .Y(n_1172) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
INVx2_ASAP7_75t_SL g1088 ( .A(n_1089), .Y(n_1088) );
AOI31xp33_ASAP7_75t_L g1659 ( .A1(n_1097), .A2(n_1660), .A3(n_1669), .B(n_1674), .Y(n_1659) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
AOI31xp33_ASAP7_75t_SL g1329 ( .A1(n_1098), .A2(n_1330), .A3(n_1342), .B(n_1345), .Y(n_1329) );
CKINVDCx8_ASAP7_75t_R g1098 ( .A(n_1099), .Y(n_1098) );
NOR2xp33_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1102), .Y(n_1100) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1103), .Y(n_1163) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1104), .Y(n_1162) );
NAND4xp25_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .C(n_1110), .D(n_1117), .Y(n_1105) );
NAND4xp25_ASAP7_75t_SL g1585 ( .A(n_1106), .B(n_1586), .C(n_1589), .D(n_1592), .Y(n_1585) );
BUFx2_ASAP7_75t_L g1962 ( .A(n_1106), .Y(n_1962) );
BUFx4f_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1115), .Y(n_1596) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1121), .B(n_1136), .Y(n_1120) );
BUFx3_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx3_ASAP7_75t_L g1131 ( .A(n_1132), .Y(n_1131) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_1133), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1133), .B(n_1440), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1634 ( .A(n_1133), .B(n_1440), .Y(n_1634) );
INVx1_ASAP7_75t_L g1651 ( .A(n_1134), .Y(n_1651) );
AOI33xp33_ASAP7_75t_L g1365 ( .A1(n_1137), .A2(n_1366), .A3(n_1368), .B1(n_1373), .B2(n_1375), .B3(n_1377), .Y(n_1365) );
AOI33xp33_ASAP7_75t_L g1616 ( .A1(n_1137), .A2(n_1377), .A3(n_1617), .B1(n_1619), .B2(n_1620), .B3(n_1621), .Y(n_1616) );
BUFx3_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1576 ( .A(n_1140), .Y(n_1576) );
INVx1_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
AOI22xp5_ASAP7_75t_L g1164 ( .A1(n_1165), .A2(n_1220), .B1(n_1221), .B2(n_1276), .Y(n_1164) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1165), .Y(n_1276) );
NAND3xp33_ASAP7_75t_L g1166 ( .A(n_1167), .B(n_1199), .C(n_1201), .Y(n_1166) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_1188), .A2(n_1190), .B1(n_1191), .B2(n_1193), .Y(n_1187) );
BUFx2_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
INVx2_ASAP7_75t_L g1264 ( .A(n_1189), .Y(n_1264) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
NOR2xp33_ASAP7_75t_SL g1201 ( .A(n_1202), .B(n_1217), .Y(n_1201) );
NAND3xp33_ASAP7_75t_SL g1202 ( .A(n_1203), .B(n_1205), .C(n_1215), .Y(n_1202) );
AOI33xp33_ASAP7_75t_L g1316 ( .A1(n_1206), .A2(n_1240), .A3(n_1317), .B1(n_1318), .B2(n_1321), .B3(n_1323), .Y(n_1316) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1209), .Y(n_1386) );
INVx1_ASAP7_75t_L g1211 ( .A(n_1212), .Y(n_1211) );
INVx2_ASAP7_75t_L g1372 ( .A(n_1212), .Y(n_1372) );
NAND3xp33_ASAP7_75t_SL g1360 ( .A(n_1215), .B(n_1361), .C(n_1365), .Y(n_1360) );
INVx1_ASAP7_75t_L g1215 ( .A(n_1216), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1217 ( .A(n_1218), .B(n_1219), .Y(n_1217) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
XNOR2xp5_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1224), .Y(n_1222) );
AND4x1_ASAP7_75t_L g1224 ( .A(n_1225), .B(n_1227), .C(n_1252), .D(n_1273), .Y(n_1224) );
NOR3xp33_ASAP7_75t_SL g1227 ( .A(n_1228), .B(n_1229), .C(n_1249), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1230 ( .A1(n_1231), .A2(n_1234), .B1(n_1235), .B2(n_1236), .C(n_1237), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1964 ( .A1(n_1231), .A2(n_1944), .B1(n_1965), .B2(n_1966), .C(n_1967), .Y(n_1964) );
BUFx2_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1966 ( .A(n_1238), .Y(n_1966) );
CKINVDCx5p33_ASAP7_75t_R g1239 ( .A(n_1240), .Y(n_1239) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
INVx1_ASAP7_75t_L g1618 ( .A(n_1248), .Y(n_1618) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
OAI221xp5_ASAP7_75t_L g1262 ( .A1(n_1263), .A2(n_1265), .B1(n_1266), .B2(n_1268), .C(n_1269), .Y(n_1262) );
INVx2_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
INVx2_ASAP7_75t_L g1647 ( .A(n_1264), .Y(n_1647) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
NOR2xp33_ASAP7_75t_L g1273 ( .A(n_1274), .B(n_1275), .Y(n_1273) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
XNOR2xp5_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1428), .Y(n_1279) );
AOI22xp5_ASAP7_75t_L g1280 ( .A1(n_1281), .A2(n_1378), .B1(n_1425), .B2(n_1426), .Y(n_1280) );
HB1xp67_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1282), .Y(n_1427) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_1283), .A2(n_1284), .B1(n_1325), .B2(n_1326), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
NAND4xp75_ASAP7_75t_SL g1285 ( .A(n_1286), .B(n_1294), .C(n_1296), .D(n_1316), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1287), .B(n_1290), .Y(n_1286) );
OAI22xp5_ASAP7_75t_L g1308 ( .A1(n_1291), .A2(n_1309), .B1(n_1311), .B2(n_1313), .Y(n_1308) );
BUFx2_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
XNOR2xp5_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
OAI22xp5_ASAP7_75t_L g1714 ( .A1(n_1327), .A2(n_1715), .B1(n_1716), .B2(n_1717), .Y(n_1714) );
NOR4xp75_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1351), .C(n_1358), .D(n_1360), .Y(n_1328) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1333), .Y(n_1332) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
BUFx2_ASAP7_75t_L g1347 ( .A(n_1337), .Y(n_1347) );
AND2x4_ASAP7_75t_L g1445 ( .A(n_1337), .B(n_1440), .Y(n_1445) );
NOR3xp33_ASAP7_75t_L g1937 ( .A(n_1350), .B(n_1938), .C(n_1948), .Y(n_1937) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1352), .B(n_1355), .Y(n_1351) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
INVx1_ASAP7_75t_L g1425 ( .A(n_1378), .Y(n_1425) );
HB1xp67_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx1_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
AND4x1_ASAP7_75t_L g1381 ( .A(n_1382), .B(n_1402), .C(n_1404), .D(n_1422), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g1407 ( .A1(n_1385), .A2(n_1387), .B1(n_1408), .B2(n_1410), .Y(n_1407) );
OAI22xp5_ASAP7_75t_L g1395 ( .A1(n_1396), .A2(n_1397), .B1(n_1398), .B2(n_1400), .Y(n_1395) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1424), .Y(n_1422) );
HB1xp67_ASAP7_75t_L g1426 ( .A(n_1427), .Y(n_1426) );
XNOR2xp5_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1580), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1430), .Y(n_1429) );
AO22x2_ASAP7_75t_L g1430 ( .A1(n_1431), .A2(n_1432), .B1(n_1521), .B2(n_1579), .Y(n_1430) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1478), .Y(n_1433) );
NOR3xp33_ASAP7_75t_L g1434 ( .A(n_1435), .B(n_1448), .C(n_1458), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1435 ( .A(n_1436), .B(n_1443), .Y(n_1435) );
AOI22xp33_ASAP7_75t_L g1436 ( .A1(n_1437), .A2(n_1438), .B1(n_1441), .B2(n_1442), .Y(n_1436) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
BUFx2_ASAP7_75t_L g1527 ( .A(n_1439), .Y(n_1527) );
BUFx2_ASAP7_75t_L g1629 ( .A(n_1439), .Y(n_1629) );
AOI22xp33_ASAP7_75t_L g1525 ( .A1(n_1442), .A2(n_1526), .B1(n_1527), .B2(n_1528), .Y(n_1525) );
AOI22xp33_ASAP7_75t_L g1627 ( .A1(n_1442), .A2(n_1628), .B1(n_1629), .B2(n_1630), .Y(n_1627) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_1444), .A2(n_1445), .B1(n_1446), .B2(n_1447), .Y(n_1443) );
AOI22xp33_ASAP7_75t_L g1529 ( .A1(n_1445), .A2(n_1447), .B1(n_1530), .B2(n_1531), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1631 ( .A1(n_1445), .A2(n_1632), .B1(n_1633), .B2(n_1634), .Y(n_1631) );
INVx2_ASAP7_75t_SL g1449 ( .A(n_1450), .Y(n_1449) );
INVx2_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx3_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
BUFx4f_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
BUFx4f_ASAP7_75t_L g1533 ( .A(n_1455), .Y(n_1533) );
BUFx2_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
BUFx2_ASAP7_75t_L g1636 ( .A(n_1457), .Y(n_1636) );
OAI22xp33_ASAP7_75t_L g1459 ( .A1(n_1460), .A2(n_1461), .B1(n_1462), .B2(n_1463), .Y(n_1459) );
BUFx3_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
OAI21xp5_ASAP7_75t_L g1939 ( .A1(n_1464), .A2(n_1940), .B(n_1941), .Y(n_1939) );
INVx2_ASAP7_75t_L g1467 ( .A(n_1468), .Y(n_1467) );
INVx2_ASAP7_75t_L g1468 ( .A(n_1469), .Y(n_1468) );
AOI221xp5_ASAP7_75t_L g1481 ( .A1(n_1472), .A2(n_1482), .B1(n_1484), .B2(n_1489), .C(n_1492), .Y(n_1481) );
AOI22xp33_ASAP7_75t_L g1511 ( .A1(n_1473), .A2(n_1475), .B1(n_1512), .B2(n_1514), .Y(n_1511) );
AOI221xp5_ASAP7_75t_L g1498 ( .A1(n_1476), .A2(n_1499), .B1(n_1505), .B2(n_1506), .C(n_1508), .Y(n_1498) );
OAI33xp33_ASAP7_75t_L g1637 ( .A1(n_1477), .A2(n_1638), .A3(n_1640), .B1(n_1645), .B2(n_1649), .B3(n_1653), .Y(n_1637) );
AOI22xp33_ASAP7_75t_L g1478 ( .A1(n_1479), .A2(n_1480), .B1(n_1516), .B2(n_1517), .Y(n_1478) );
AOI22xp33_ASAP7_75t_L g1556 ( .A1(n_1479), .A2(n_1517), .B1(n_1557), .B2(n_1578), .Y(n_1556) );
NAND3xp33_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1498), .C(n_1511), .Y(n_1480) );
AOI221xp5_ASAP7_75t_L g1558 ( .A1(n_1482), .A2(n_1549), .B1(n_1559), .B2(n_1565), .C(n_1569), .Y(n_1558) );
AOI21xp5_ASAP7_75t_L g1660 ( .A1(n_1482), .A2(n_1650), .B(n_1661), .Y(n_1660) );
BUFx2_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
BUFx2_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
INVx2_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
INVx2_ASAP7_75t_SL g1496 ( .A(n_1497), .Y(n_1496) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1504), .Y(n_1503) );
AOI221xp5_ASAP7_75t_L g1571 ( .A1(n_1506), .A2(n_1508), .B1(n_1555), .B2(n_1572), .C(n_1575), .Y(n_1571) );
AOI221xp5_ASAP7_75t_L g1669 ( .A1(n_1506), .A2(n_1508), .B1(n_1656), .B2(n_1670), .C(n_1673), .Y(n_1669) );
BUFx6f_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx1_ASAP7_75t_SL g1509 ( .A(n_1510), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_1512), .A2(n_1514), .B1(n_1552), .B2(n_1554), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1674 ( .A1(n_1512), .A2(n_1514), .B1(n_1652), .B2(n_1655), .Y(n_1674) );
INVx6_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
INVx4_ASAP7_75t_L g1514 ( .A(n_1515), .Y(n_1514) );
AOI21xp33_ASAP7_75t_L g1657 ( .A1(n_1517), .A2(n_1658), .B(n_1659), .Y(n_1657) );
INVx5_ASAP7_75t_L g1517 ( .A(n_1518), .Y(n_1517) );
AND2x4_ASAP7_75t_L g1518 ( .A(n_1519), .B(n_1520), .Y(n_1518) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1521), .Y(n_1579) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1556), .Y(n_1522) );
NOR3xp33_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1532), .C(n_1534), .Y(n_1523) );
NAND2xp5_ASAP7_75t_L g1524 ( .A(n_1525), .B(n_1529), .Y(n_1524) );
OAI22xp33_ASAP7_75t_L g1535 ( .A1(n_1536), .A2(n_1537), .B1(n_1538), .B2(n_1539), .Y(n_1535) );
OAI22xp5_ASAP7_75t_L g1540 ( .A1(n_1541), .A2(n_1542), .B1(n_1543), .B2(n_1544), .Y(n_1540) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
INVx1_ASAP7_75t_L g1545 ( .A(n_1546), .Y(n_1545) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_1548), .A2(n_1549), .B1(n_1550), .B2(n_1552), .Y(n_1547) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1551), .Y(n_1550) );
NAND3xp33_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1571), .C(n_1577), .Y(n_1557) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx1_ASAP7_75t_L g1562 ( .A(n_1563), .Y(n_1562) );
INVx1_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1567), .Y(n_1566) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
XNOR2xp5_ASAP7_75t_L g1582 ( .A(n_1583), .B(n_1622), .Y(n_1582) );
INVx1_ASAP7_75t_L g1595 ( .A(n_1596), .Y(n_1595) );
NAND2xp5_ASAP7_75t_L g1608 ( .A(n_1609), .B(n_1616), .Y(n_1608) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1615), .Y(n_1614) );
XNOR2x1_ASAP7_75t_L g1622 ( .A(n_1623), .B(n_1624), .Y(n_1622) );
AND2x2_ASAP7_75t_L g1624 ( .A(n_1625), .B(n_1657), .Y(n_1624) );
NOR3xp33_ASAP7_75t_SL g1625 ( .A(n_1626), .B(n_1635), .C(n_1637), .Y(n_1625) );
NAND2xp5_ASAP7_75t_L g1626 ( .A(n_1627), .B(n_1631), .Y(n_1626) );
OAI211xp5_ASAP7_75t_L g1664 ( .A1(n_1630), .A2(n_1665), .B(n_1666), .C(n_1667), .Y(n_1664) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx3_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
OAI22xp5_ASAP7_75t_L g1649 ( .A1(n_1647), .A2(n_1650), .B1(n_1651), .B2(n_1652), .Y(n_1649) );
INVx1_ASAP7_75t_SL g1662 ( .A(n_1663), .Y(n_1662) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1672), .Y(n_1671) );
OAI221xp5_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1922), .B1(n_1925), .B2(n_1973), .C(n_1978), .Y(n_1675) );
NOR3xp33_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1892), .C(n_1919), .Y(n_1676) );
AOI33xp33_ASAP7_75t_L g1677 ( .A1(n_1678), .A2(n_1772), .A3(n_1817), .B1(n_1844), .B2(n_1863), .B3(n_1879), .Y(n_1677) );
AOI211xp5_ASAP7_75t_L g1678 ( .A1(n_1679), .A2(n_1722), .B(n_1744), .C(n_1761), .Y(n_1678) );
NOR2xp33_ASAP7_75t_L g1679 ( .A(n_1680), .B(n_1703), .Y(n_1679) );
OR2x2_ASAP7_75t_L g1770 ( .A(n_1680), .B(n_1771), .Y(n_1770) );
NOR2x1_ASAP7_75t_R g1803 ( .A(n_1680), .B(n_1804), .Y(n_1803) );
AND2x2_ASAP7_75t_L g1819 ( .A(n_1680), .B(n_1759), .Y(n_1819) );
NAND2xp5_ASAP7_75t_L g1884 ( .A(n_1680), .B(n_1866), .Y(n_1884) );
AOI211xp5_ASAP7_75t_SL g1895 ( .A1(n_1680), .A2(n_1743), .B(n_1896), .C(n_1897), .Y(n_1895) );
INVx2_ASAP7_75t_L g1680 ( .A(n_1681), .Y(n_1680) );
NAND2xp5_ASAP7_75t_L g1751 ( .A(n_1681), .B(n_1752), .Y(n_1751) );
INVx2_ASAP7_75t_L g1681 ( .A(n_1682), .Y(n_1681) );
INVx4_ASAP7_75t_L g1768 ( .A(n_1682), .Y(n_1768) );
NAND2xp5_ASAP7_75t_L g1774 ( .A(n_1682), .B(n_1775), .Y(n_1774) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1682), .B(n_1743), .Y(n_1798) );
NAND2xp5_ASAP7_75t_L g1824 ( .A(n_1682), .B(n_1732), .Y(n_1824) );
OR2x2_ASAP7_75t_L g1835 ( .A(n_1682), .B(n_1769), .Y(n_1835) );
NOR2xp33_ASAP7_75t_L g1849 ( .A(n_1682), .B(n_1743), .Y(n_1849) );
NAND2xp5_ASAP7_75t_L g1858 ( .A(n_1682), .B(n_1753), .Y(n_1858) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1682), .B(n_1705), .Y(n_1886) );
AND2x2_ASAP7_75t_L g1891 ( .A(n_1682), .B(n_1787), .Y(n_1891) );
AND2x2_ASAP7_75t_L g1894 ( .A(n_1682), .B(n_1741), .Y(n_1894) );
AOI21xp5_ASAP7_75t_L g1906 ( .A1(n_1682), .A2(n_1794), .B(n_1803), .Y(n_1906) );
NAND2xp5_ASAP7_75t_L g1910 ( .A(n_1682), .B(n_1754), .Y(n_1910) );
AND2x6_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1695), .Y(n_1682) );
AND2x4_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1690), .Y(n_1684) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
OR2x2_ASAP7_75t_L g1709 ( .A(n_1686), .B(n_1691), .Y(n_1709) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1689), .Y(n_1686) );
HB1xp67_ASAP7_75t_L g1989 ( .A(n_1687), .Y(n_1989) );
INVx1_ASAP7_75t_L g1687 ( .A(n_1688), .Y(n_1687) );
INVx1_ASAP7_75t_L g1698 ( .A(n_1689), .Y(n_1698) );
AND2x4_ASAP7_75t_L g1692 ( .A(n_1690), .B(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1690 ( .A(n_1691), .Y(n_1690) );
OR2x2_ASAP7_75t_L g1713 ( .A(n_1691), .B(n_1694), .Y(n_1713) );
INVx1_ASAP7_75t_L g1693 ( .A(n_1694), .Y(n_1693) );
INVx1_ASAP7_75t_L g1715 ( .A(n_1696), .Y(n_1715) );
INVx1_ASAP7_75t_L g1810 ( .A(n_1696), .Y(n_1810) );
BUFx3_ASAP7_75t_L g1924 ( .A(n_1696), .Y(n_1924) );
AND2x4_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1699), .Y(n_1696) );
AND2x2_ASAP7_75t_L g1721 ( .A(n_1697), .B(n_1699), .Y(n_1721) );
HB1xp67_ASAP7_75t_L g1990 ( .A(n_1697), .Y(n_1990) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
AND2x4_ASAP7_75t_L g1702 ( .A(n_1698), .B(n_1699), .Y(n_1702) );
INVx2_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
OAI22xp5_ASAP7_75t_L g1808 ( .A1(n_1701), .A2(n_1809), .B1(n_1810), .B2(n_1811), .Y(n_1808) );
INVx2_ASAP7_75t_L g1701 ( .A(n_1702), .Y(n_1701) );
INVx1_ASAP7_75t_SL g1717 ( .A(n_1702), .Y(n_1717) );
OAI222xp33_ASAP7_75t_L g1773 ( .A1(n_1703), .A2(n_1774), .B1(n_1778), .B2(n_1781), .C1(n_1784), .C2(n_1786), .Y(n_1773) );
OAI321xp33_ASAP7_75t_L g1909 ( .A1(n_1703), .A2(n_1837), .A3(n_1865), .B1(n_1910), .B2(n_1911), .C(n_1913), .Y(n_1909) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_1704), .B(n_1753), .Y(n_1826) );
AOI221xp5_ASAP7_75t_L g1844 ( .A1(n_1704), .A2(n_1749), .B1(n_1845), .B2(n_1854), .C(n_1855), .Y(n_1844) );
AND2x2_ASAP7_75t_L g1704 ( .A(n_1705), .B(n_1718), .Y(n_1704) );
INVx3_ASAP7_75t_L g1748 ( .A(n_1705), .Y(n_1748) );
OR2x2_ASAP7_75t_L g1762 ( .A(n_1705), .B(n_1763), .Y(n_1762) );
OR2x2_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1714), .Y(n_1705) );
OAI22xp33_ASAP7_75t_L g1706 ( .A1(n_1707), .A2(n_1708), .B1(n_1710), .B2(n_1711), .Y(n_1706) );
OAI22xp5_ASAP7_75t_L g1729 ( .A1(n_1708), .A2(n_1713), .B1(n_1730), .B2(n_1731), .Y(n_1729) );
OAI22xp33_ASAP7_75t_L g1756 ( .A1(n_1708), .A2(n_1713), .B1(n_1757), .B2(n_1758), .Y(n_1756) );
BUFx3_ASAP7_75t_L g1814 ( .A(n_1708), .Y(n_1814) );
BUFx6f_ASAP7_75t_L g1708 ( .A(n_1709), .Y(n_1708) );
OAI22xp5_ASAP7_75t_L g1737 ( .A1(n_1709), .A2(n_1713), .B1(n_1738), .B2(n_1739), .Y(n_1737) );
HB1xp67_ASAP7_75t_L g1816 ( .A(n_1711), .Y(n_1816) );
INVx1_ASAP7_75t_L g1711 ( .A(n_1712), .Y(n_1711) );
INVx1_ASAP7_75t_L g1712 ( .A(n_1713), .Y(n_1712) );
OR2x2_ASAP7_75t_L g1763 ( .A(n_1718), .B(n_1755), .Y(n_1763) );
OR2x2_ASAP7_75t_L g1771 ( .A(n_1718), .B(n_1754), .Y(n_1771) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1718), .B(n_1754), .Y(n_1787) );
AND2x2_ASAP7_75t_L g1796 ( .A(n_1718), .B(n_1748), .Y(n_1796) );
INVx2_ASAP7_75t_L g1802 ( .A(n_1718), .Y(n_1802) );
OAI22xp5_ASAP7_75t_L g1869 ( .A1(n_1718), .A2(n_1842), .B1(n_1870), .B2(n_1872), .Y(n_1869) );
AND2x2_ASAP7_75t_L g1877 ( .A(n_1718), .B(n_1755), .Y(n_1877) );
AOI221xp5_ASAP7_75t_L g1893 ( .A1(n_1718), .A2(n_1877), .B1(n_1894), .B2(n_1895), .C(n_1899), .Y(n_1893) );
AND2x4_ASAP7_75t_L g1718 ( .A(n_1719), .B(n_1720), .Y(n_1718) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1721), .Y(n_1727) );
NAND2xp5_ASAP7_75t_L g1722 ( .A(n_1723), .B(n_1740), .Y(n_1722) );
OAI22xp33_ASAP7_75t_L g1875 ( .A1(n_1723), .A2(n_1846), .B1(n_1876), .B2(n_1878), .Y(n_1875) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
AND2x2_ASAP7_75t_L g1724 ( .A(n_1725), .B(n_1732), .Y(n_1724) );
CKINVDCx6p67_ASAP7_75t_R g1743 ( .A(n_1725), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1759 ( .A(n_1725), .B(n_1760), .Y(n_1759) );
NAND2xp5_ASAP7_75t_L g1766 ( .A(n_1725), .B(n_1767), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1775 ( .A(n_1725), .B(n_1776), .Y(n_1775) );
OR2x2_ASAP7_75t_L g1780 ( .A(n_1725), .B(n_1742), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1725), .B(n_1785), .Y(n_1784) );
OR2x2_ASAP7_75t_L g1829 ( .A(n_1725), .B(n_1769), .Y(n_1829) );
AND2x2_ASAP7_75t_L g1868 ( .A(n_1725), .B(n_1742), .Y(n_1868) );
AND2x2_ASAP7_75t_L g1912 ( .A(n_1725), .B(n_1790), .Y(n_1912) );
OR2x6_ASAP7_75t_SL g1725 ( .A(n_1726), .B(n_1729), .Y(n_1725) );
AND2x2_ASAP7_75t_L g1785 ( .A(n_1732), .B(n_1768), .Y(n_1785) );
NAND2xp5_ASAP7_75t_L g1797 ( .A(n_1732), .B(n_1798), .Y(n_1797) );
AND2x2_ASAP7_75t_L g1841 ( .A(n_1732), .B(n_1743), .Y(n_1841) );
INVx1_ASAP7_75t_L g1896 ( .A(n_1732), .Y(n_1896) );
AND2x2_ASAP7_75t_L g1732 ( .A(n_1733), .B(n_1736), .Y(n_1732) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1733), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1769 ( .A(n_1733), .B(n_1736), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1776 ( .A(n_1733), .B(n_1777), .Y(n_1776) );
AND2x2_ASAP7_75t_L g1733 ( .A(n_1734), .B(n_1735), .Y(n_1733) );
AND2x2_ASAP7_75t_L g1760 ( .A(n_1736), .B(n_1742), .Y(n_1760) );
INVx1_ASAP7_75t_L g1777 ( .A(n_1736), .Y(n_1777) );
NOR2xp33_ASAP7_75t_L g1838 ( .A(n_1736), .B(n_1743), .Y(n_1838) );
OAI22xp5_ASAP7_75t_L g1761 ( .A1(n_1740), .A2(n_1762), .B1(n_1764), .B2(n_1770), .Y(n_1761) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
AND2x2_ASAP7_75t_L g1741 ( .A(n_1742), .B(n_1743), .Y(n_1741) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1743), .B(n_1776), .Y(n_1794) );
AND2x2_ASAP7_75t_L g1853 ( .A(n_1743), .B(n_1760), .Y(n_1853) );
AND2x2_ASAP7_75t_L g1871 ( .A(n_1743), .B(n_1785), .Y(n_1871) );
AND2x2_ASAP7_75t_L g1880 ( .A(n_1743), .B(n_1777), .Y(n_1880) );
OAI322xp33_ASAP7_75t_L g1883 ( .A1(n_1743), .A2(n_1829), .A3(n_1833), .B1(n_1884), .B2(n_1885), .C1(n_1887), .C2(n_1888), .Y(n_1883) );
NAND2xp5_ASAP7_75t_L g1885 ( .A(n_1743), .B(n_1886), .Y(n_1885) );
OR2x2_ASAP7_75t_L g1898 ( .A(n_1743), .B(n_1777), .Y(n_1898) );
NOR2xp33_ASAP7_75t_L g1908 ( .A(n_1743), .B(n_1824), .Y(n_1908) );
INVxp67_ASAP7_75t_L g1744 ( .A(n_1745), .Y(n_1744) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1746), .B(n_1749), .Y(n_1745) );
O2A1O1Ixp33_ASAP7_75t_L g1836 ( .A1(n_1746), .A2(n_1770), .B(n_1837), .C(n_1839), .Y(n_1836) );
INVx1_ASAP7_75t_SL g1746 ( .A(n_1747), .Y(n_1746) );
AND2x2_ASAP7_75t_L g1818 ( .A(n_1747), .B(n_1819), .Y(n_1818) );
INVx3_ASAP7_75t_L g1747 ( .A(n_1748), .Y(n_1747) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1748), .B(n_1802), .Y(n_1801) );
INVx1_ASAP7_75t_L g1833 ( .A(n_1748), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1854 ( .A(n_1748), .B(n_1754), .Y(n_1854) );
AND2x2_ASAP7_75t_L g1862 ( .A(n_1748), .B(n_1753), .Y(n_1862) );
O2A1O1Ixp33_ASAP7_75t_SL g1919 ( .A1(n_1748), .A2(n_1763), .B(n_1920), .C(n_1921), .Y(n_1919) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1759), .Y(n_1749) );
NOR2xp33_ASAP7_75t_L g1795 ( .A(n_1750), .B(n_1796), .Y(n_1795) );
INVx1_ASAP7_75t_L g1750 ( .A(n_1751), .Y(n_1750) );
INVx1_ASAP7_75t_L g1752 ( .A(n_1753), .Y(n_1752) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1753), .Y(n_1799) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1753), .Y(n_1832) );
INVx2_ASAP7_75t_SL g1753 ( .A(n_1754), .Y(n_1753) );
INVx2_ASAP7_75t_SL g1754 ( .A(n_1755), .Y(n_1754) );
HB1xp67_ASAP7_75t_L g1823 ( .A(n_1755), .Y(n_1823) );
NOR2xp33_ASAP7_75t_L g1778 ( .A(n_1759), .B(n_1779), .Y(n_1778) );
INVx1_ASAP7_75t_L g1804 ( .A(n_1760), .Y(n_1804) );
OAI22xp5_ASAP7_75t_L g1905 ( .A1(n_1762), .A2(n_1882), .B1(n_1906), .B2(n_1907), .Y(n_1905) );
INVx1_ASAP7_75t_L g1783 ( .A(n_1763), .Y(n_1783) );
INVxp67_ASAP7_75t_SL g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1766), .Y(n_1765) );
AOI22xp33_ASAP7_75t_L g1859 ( .A1(n_1767), .A2(n_1831), .B1(n_1860), .B2(n_1862), .Y(n_1859) );
NOR2xp33_ASAP7_75t_L g1767 ( .A(n_1768), .B(n_1769), .Y(n_1767) );
AND2x2_ASAP7_75t_L g1782 ( .A(n_1768), .B(n_1783), .Y(n_1782) );
NAND2xp5_ASAP7_75t_L g1852 ( .A(n_1768), .B(n_1853), .Y(n_1852) );
INVx1_ASAP7_75t_L g1861 ( .A(n_1768), .Y(n_1861) );
AND2x2_ASAP7_75t_L g1867 ( .A(n_1768), .B(n_1868), .Y(n_1867) );
O2A1O1Ixp33_ASAP7_75t_L g1917 ( .A1(n_1768), .A2(n_1804), .B(n_1825), .C(n_1918), .Y(n_1917) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1769), .Y(n_1790) );
INVx1_ASAP7_75t_L g1791 ( .A(n_1770), .Y(n_1791) );
AOI221xp5_ASAP7_75t_L g1863 ( .A1(n_1771), .A2(n_1864), .B1(n_1867), .B2(n_1869), .C(n_1875), .Y(n_1863) );
INVx2_ASAP7_75t_L g1866 ( .A(n_1771), .Y(n_1866) );
NOR3xp33_ASAP7_75t_L g1772 ( .A(n_1773), .B(n_1788), .C(n_1792), .Y(n_1772) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1774), .Y(n_1904) );
AND2x2_ASAP7_75t_L g1860 ( .A(n_1776), .B(n_1861), .Y(n_1860) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1776), .Y(n_1873) );
NAND3xp33_ASAP7_75t_L g1913 ( .A(n_1779), .B(n_1866), .C(n_1886), .Y(n_1913) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1780), .Y(n_1779) );
INVx1_ASAP7_75t_L g1781 ( .A(n_1782), .Y(n_1781) );
INVx1_ASAP7_75t_L g1786 ( .A(n_1787), .Y(n_1786) );
AOI211xp5_ASAP7_75t_SL g1903 ( .A1(n_1787), .A2(n_1904), .B(n_1905), .C(n_1909), .Y(n_1903) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
NAND2xp5_ASAP7_75t_L g1789 ( .A(n_1790), .B(n_1791), .Y(n_1789) );
NAND2xp5_ASAP7_75t_L g1848 ( .A(n_1790), .B(n_1849), .Y(n_1848) );
NAND3xp33_ASAP7_75t_L g1856 ( .A(n_1790), .B(n_1802), .C(n_1857), .Y(n_1856) );
NAND2xp5_ASAP7_75t_L g1902 ( .A(n_1790), .B(n_1798), .Y(n_1902) );
OAI221xp5_ASAP7_75t_L g1792 ( .A1(n_1793), .A2(n_1795), .B1(n_1797), .B2(n_1799), .C(n_1800), .Y(n_1792) );
INVx1_ASAP7_75t_L g1793 ( .A(n_1794), .Y(n_1793) );
AOI221xp5_ASAP7_75t_L g1914 ( .A1(n_1796), .A2(n_1840), .B1(n_1847), .B2(n_1915), .C(n_1917), .Y(n_1914) );
NAND2xp5_ASAP7_75t_L g1916 ( .A(n_1796), .B(n_1799), .Y(n_1916) );
AND2x2_ASAP7_75t_L g1821 ( .A(n_1797), .B(n_1822), .Y(n_1821) );
A2O1A1Ixp33_ASAP7_75t_SL g1839 ( .A1(n_1799), .A2(n_1840), .B(n_1841), .C(n_1842), .Y(n_1839) );
AOI21xp5_ASAP7_75t_L g1800 ( .A1(n_1801), .A2(n_1803), .B(n_1805), .Y(n_1800) );
NOR2xp33_ASAP7_75t_L g1830 ( .A(n_1801), .B(n_1823), .Y(n_1830) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1801), .Y(n_1878) );
NAND2xp5_ASAP7_75t_L g1882 ( .A(n_1801), .B(n_1823), .Y(n_1882) );
OAI321xp33_ASAP7_75t_L g1820 ( .A1(n_1802), .A2(n_1804), .A3(n_1821), .B1(n_1824), .B2(n_1825), .C(n_1827), .Y(n_1820) );
INVx1_ASAP7_75t_L g1843 ( .A(n_1802), .Y(n_1843) );
AND2x2_ASAP7_75t_L g1887 ( .A(n_1804), .B(n_1873), .Y(n_1887) );
CKINVDCx14_ASAP7_75t_R g1805 ( .A(n_1806), .Y(n_1805) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
NAND3xp33_ASAP7_75t_SL g1855 ( .A(n_1807), .B(n_1856), .C(n_1859), .Y(n_1855) );
OR2x6_ASAP7_75t_SL g1807 ( .A(n_1808), .B(n_1812), .Y(n_1807) );
OAI22xp5_ASAP7_75t_L g1812 ( .A1(n_1813), .A2(n_1814), .B1(n_1815), .B2(n_1816), .Y(n_1812) );
NOR3xp33_ASAP7_75t_SL g1817 ( .A(n_1818), .B(n_1820), .C(n_1836), .Y(n_1817) );
INVxp67_ASAP7_75t_L g1921 ( .A(n_1818), .Y(n_1921) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
INVx1_ASAP7_75t_L g1901 ( .A(n_1823), .Y(n_1901) );
INVx1_ASAP7_75t_L g1840 ( .A(n_1824), .Y(n_1840) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1826), .Y(n_1825) );
AOI22xp33_ASAP7_75t_L g1827 ( .A1(n_1828), .A2(n_1830), .B1(n_1831), .B2(n_1834), .Y(n_1827) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_1832), .B(n_1833), .Y(n_1831) );
NAND2xp5_ASAP7_75t_L g1865 ( .A(n_1833), .B(n_1866), .Y(n_1865) );
OAI211xp5_ASAP7_75t_L g1892 ( .A1(n_1833), .A2(n_1893), .B(n_1903), .C(n_1914), .Y(n_1892) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1835), .Y(n_1834) );
NOR2xp33_ASAP7_75t_L g1889 ( .A(n_1837), .B(n_1890), .Y(n_1889) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
INVx1_ASAP7_75t_L g1920 ( .A(n_1841), .Y(n_1920) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
NAND2xp5_ASAP7_75t_L g1845 ( .A(n_1846), .B(n_1850), .Y(n_1845) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1847 ( .A(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g1874 ( .A(n_1849), .Y(n_1874) );
INVx1_ASAP7_75t_L g1850 ( .A(n_1851), .Y(n_1850) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1852), .Y(n_1851) );
INVx1_ASAP7_75t_L g1918 ( .A(n_1853), .Y(n_1918) );
INVx1_ASAP7_75t_L g1857 ( .A(n_1858), .Y(n_1857) );
INVx1_ASAP7_75t_L g1888 ( .A(n_1862), .Y(n_1888) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1865), .Y(n_1864) );
INVx1_ASAP7_75t_L g1870 ( .A(n_1871), .Y(n_1870) );
OR2x2_ASAP7_75t_L g1872 ( .A(n_1873), .B(n_1874), .Y(n_1872) );
INVx1_ASAP7_75t_L g1876 ( .A(n_1877), .Y(n_1876) );
AOI211xp5_ASAP7_75t_L g1879 ( .A1(n_1880), .A2(n_1881), .B(n_1883), .C(n_1889), .Y(n_1879) );
INVx1_ASAP7_75t_L g1881 ( .A(n_1882), .Y(n_1881) );
INVx1_ASAP7_75t_L g1890 ( .A(n_1891), .Y(n_1890) );
INVx1_ASAP7_75t_L g1897 ( .A(n_1898), .Y(n_1897) );
INVx1_ASAP7_75t_L g1899 ( .A(n_1900), .Y(n_1899) );
OR2x2_ASAP7_75t_L g1900 ( .A(n_1901), .B(n_1902), .Y(n_1900) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
INVx1_ASAP7_75t_L g1911 ( .A(n_1912), .Y(n_1911) );
INVx1_ASAP7_75t_L g1915 ( .A(n_1916), .Y(n_1915) );
HB1xp67_ASAP7_75t_L g1922 ( .A(n_1923), .Y(n_1922) );
INVx1_ASAP7_75t_L g1923 ( .A(n_1924), .Y(n_1923) );
INVx2_ASAP7_75t_SL g1925 ( .A(n_1926), .Y(n_1925) );
INVx1_ASAP7_75t_L g1972 ( .A(n_1927), .Y(n_1972) );
HB1xp67_ASAP7_75t_L g1985 ( .A(n_1927), .Y(n_1985) );
NAND3xp33_ASAP7_75t_L g1928 ( .A(n_1929), .B(n_1934), .C(n_1937), .Y(n_1928) );
OAI21xp5_ASAP7_75t_SL g1938 ( .A1(n_1939), .A2(n_1942), .B(n_1945), .Y(n_1938) );
NAND4xp25_ASAP7_75t_SL g1953 ( .A(n_1954), .B(n_1957), .C(n_1959), .D(n_1962), .Y(n_1953) );
INVx1_ASAP7_75t_L g1960 ( .A(n_1961), .Y(n_1960) );
CKINVDCx14_ASAP7_75t_R g1973 ( .A(n_1974), .Y(n_1973) );
BUFx2_ASAP7_75t_L g1974 ( .A(n_1975), .Y(n_1974) );
INVx1_ASAP7_75t_L g1975 ( .A(n_1976), .Y(n_1975) );
INVx1_ASAP7_75t_L g1976 ( .A(n_1977), .Y(n_1976) );
INVx1_ASAP7_75t_L g1979 ( .A(n_1980), .Y(n_1979) );
CKINVDCx5p33_ASAP7_75t_R g1980 ( .A(n_1981), .Y(n_1980) );
A2O1A1Ixp33_ASAP7_75t_L g1987 ( .A1(n_1982), .A2(n_1988), .B(n_1990), .C(n_1991), .Y(n_1987) );
INVxp33_ASAP7_75t_SL g1983 ( .A(n_1984), .Y(n_1983) );
HB1xp67_ASAP7_75t_L g1986 ( .A(n_1987), .Y(n_1986) );
INVx1_ASAP7_75t_L g1988 ( .A(n_1989), .Y(n_1988) );
endmodule