module fake_ariane_2266_n_1706 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_1706);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1706;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_137;
wire n_1298;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_136;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_149;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_209;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_159;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_144;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_155;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_145;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_451;
wire n_745;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_157;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1524;
wire n_1476;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_140;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_152;
wire n_169;
wire n_1288;
wire n_1201;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_161;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_139;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_153;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1670;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_52),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_30),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_4),
.Y(n_140)
);

BUFx10_ASAP7_75t_L g141 ( 
.A(n_6),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_81),
.Y(n_142)
);

CKINVDCx5p33_ASAP7_75t_R g143 ( 
.A(n_29),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_105),
.Y(n_144)
);

CKINVDCx5p33_ASAP7_75t_R g145 ( 
.A(n_57),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_38),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_42),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_50),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_44),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_55),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_63),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_96),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_104),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_36),
.Y(n_154)
);

CKINVDCx5p33_ASAP7_75t_R g155 ( 
.A(n_25),
.Y(n_155)
);

BUFx10_ASAP7_75t_L g156 ( 
.A(n_129),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_52),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_117),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_27),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_76),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_10),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_58),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_83),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_75),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_43),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_90),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_1),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g170 ( 
.A(n_30),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_116),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_119),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_29),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_22),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_120),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_89),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_13),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_13),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_60),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_103),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_42),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_134),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_80),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_91),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_17),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_84),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_132),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_94),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_6),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_109),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_28),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_125),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_47),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_12),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_20),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_2),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_22),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_88),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_32),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_48),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_71),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_12),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_59),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_61),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_47),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_78),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_5),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_25),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_56),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_102),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_43),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_54),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_17),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_107),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_123),
.Y(n_221)
);

BUFx2_ASAP7_75t_SL g222 ( 
.A(n_72),
.Y(n_222)
);

BUFx8_ASAP7_75t_SL g223 ( 
.A(n_69),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_5),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_24),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g226 ( 
.A(n_40),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_1),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_130),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_4),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_113),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_23),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_49),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_35),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_55),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_34),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_100),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_131),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_62),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_26),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_122),
.Y(n_243)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_82),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_135),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_11),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_20),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_0),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_32),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_18),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_35),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_41),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_44),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_7),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_73),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_24),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_23),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_87),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_97),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_37),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_124),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_68),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_54),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_112),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

BUFx3_ASAP7_75t_L g269 ( 
.A(n_15),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_67),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_151),
.Y(n_271)
);

INVxp67_ASAP7_75t_SL g272 ( 
.A(n_137),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_223),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_149),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_210),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_175),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_185),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_226),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_0),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_136),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_158),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_199),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_139),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_139),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_163),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_138),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_140),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_163),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_165),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_165),
.Y(n_292)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_137),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_143),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_150),
.B(n_157),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_167),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_201),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_167),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_205),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_225),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

INVxp67_ASAP7_75t_SL g302 ( 
.A(n_154),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_232),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_145),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_154),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_146),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_147),
.Y(n_308)
);

INVxp33_ASAP7_75t_SL g309 ( 
.A(n_148),
.Y(n_309)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_185),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_155),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_188),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_252),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_210),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_159),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_261),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_188),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_210),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_152),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_220),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_190),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_156),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_156),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_L g325 ( 
.A(n_234),
.B(n_3),
.Y(n_325)
);

INVxp67_ASAP7_75t_SL g326 ( 
.A(n_160),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_190),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_195),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_156),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_195),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_160),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_156),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_206),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_206),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_166),
.Y(n_335)
);

INVxp33_ASAP7_75t_L g336 ( 
.A(n_173),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_169),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_210),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_208),
.B(n_3),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_208),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_211),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_246),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_173),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_210),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_174),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_211),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_275),
.B(n_218),
.Y(n_347)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_275),
.B(n_218),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_277),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_323),
.B(n_141),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_277),
.Y(n_352)
);

AND2x4_ASAP7_75t_L g353 ( 
.A(n_279),
.B(n_228),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_279),
.B(n_310),
.Y(n_354)
);

AND2x6_ASAP7_75t_L g355 ( 
.A(n_282),
.B(n_161),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_277),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_314),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_279),
.B(n_231),
.Y(n_358)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_310),
.B(n_228),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g360 ( 
.A(n_310),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_282),
.B(n_269),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g362 ( 
.A(n_274),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_314),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_314),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_318),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_318),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_338),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_338),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_338),
.Y(n_370)
);

AND2x4_ASAP7_75t_L g371 ( 
.A(n_285),
.B(n_286),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_344),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_344),
.Y(n_373)
);

INVx4_ASAP7_75t_L g374 ( 
.A(n_344),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_285),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_286),
.B(n_231),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_323),
.B(n_230),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_324),
.B(n_141),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_287),
.B(n_238),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_287),
.B(n_238),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_290),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_290),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_291),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_291),
.B(n_245),
.Y(n_384)
);

CKINVDCx14_ASAP7_75t_R g385 ( 
.A(n_319),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_292),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_292),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_296),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_296),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_298),
.Y(n_390)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_298),
.B(n_269),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_312),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_312),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_317),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_317),
.Y(n_395)
);

INVx4_ASAP7_75t_L g396 ( 
.A(n_322),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_309),
.B(n_288),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_322),
.B(n_247),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_327),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_327),
.B(n_247),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_328),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_328),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_330),
.Y(n_403)
);

BUFx2_ASAP7_75t_L g404 ( 
.A(n_276),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_330),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_333),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_333),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_334),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_334),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_230),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_340),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_346),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_397),
.B(n_278),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_387),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_377),
.B(n_324),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_387),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_387),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_387),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_387),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_354),
.B(n_278),
.Y(n_424)
);

NAND2x1p5_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_245),
.Y(n_425)
);

NAND3xp33_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_281),
.C(n_289),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_387),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_354),
.B(n_294),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_387),
.Y(n_430)
);

OA22x2_ASAP7_75t_L g431 ( 
.A1(n_362),
.A2(n_297),
.B1(n_274),
.B2(n_272),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_348),
.Y(n_432)
);

NAND3xp33_ASAP7_75t_L g433 ( 
.A(n_396),
.B(n_307),
.C(n_304),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_348),
.Y(n_435)
);

BUFx4f_ASAP7_75t_L g436 ( 
.A(n_388),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_351),
.B(n_308),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_388),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_388),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_377),
.B(n_311),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_388),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_388),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_388),
.Y(n_443)
);

INVx4_ASAP7_75t_L g444 ( 
.A(n_371),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_388),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_351),
.B(n_315),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_360),
.B(n_320),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_385),
.Y(n_449)
);

INVxp33_ASAP7_75t_L g450 ( 
.A(n_362),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_399),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_378),
.B(n_335),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_381),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_354),
.B(n_337),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_399),
.Y(n_457)
);

NOR3xp33_ASAP7_75t_L g458 ( 
.A(n_404),
.B(n_339),
.C(n_345),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_414),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_378),
.A2(n_316),
.B1(n_325),
.B2(n_280),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_399),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_354),
.B(n_272),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_414),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_360),
.B(n_321),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_354),
.B(n_293),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_399),
.Y(n_468)
);

INVx5_ASAP7_75t_L g469 ( 
.A(n_355),
.Y(n_469)
);

OR2x6_ASAP7_75t_L g470 ( 
.A(n_404),
.B(n_325),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_361),
.Y(n_471)
);

OR2x6_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_400),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g473 ( 
.A(n_361),
.Y(n_473)
);

OAI22xp33_ASAP7_75t_L g474 ( 
.A1(n_347),
.A2(n_336),
.B1(n_297),
.B2(n_178),
.Y(n_474)
);

INVxp33_ASAP7_75t_L g475 ( 
.A(n_398),
.Y(n_475)
);

NAND3xp33_ASAP7_75t_L g476 ( 
.A(n_396),
.B(n_331),
.C(n_306),
.Y(n_476)
);

INVx4_ASAP7_75t_SL g477 ( 
.A(n_355),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_360),
.B(n_329),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_371),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_371),
.B(n_293),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_399),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_402),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

BUFx4f_ASAP7_75t_L g484 ( 
.A(n_402),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_R g485 ( 
.A(n_353),
.B(n_273),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_402),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_385),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g488 ( 
.A1(n_396),
.A2(n_250),
.B1(n_182),
.B2(n_183),
.Y(n_488)
);

NAND3xp33_ASAP7_75t_L g489 ( 
.A(n_396),
.B(n_358),
.C(n_414),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g490 ( 
.A(n_361),
.B(n_306),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_353),
.A2(n_302),
.B1(n_326),
.B2(n_332),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_391),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_389),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_390),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_407),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_391),
.B(n_331),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_396),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_392),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_392),
.B(n_394),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_402),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_407),
.B(n_326),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_402),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_402),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_411),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_407),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_395),
.B(n_343),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_355),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g512 ( 
.A(n_395),
.B(n_343),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_407),
.B(n_301),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_411),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_411),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_411),
.Y(n_516)
);

AND2x2_ASAP7_75t_SL g517 ( 
.A(n_410),
.B(n_264),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_411),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_411),
.Y(n_520)
);

INVx2_ASAP7_75t_SL g521 ( 
.A(n_353),
.Y(n_521)
);

INVx1_ASAP7_75t_SL g522 ( 
.A(n_391),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_353),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_401),
.B(n_301),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_411),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_353),
.B(n_141),
.Y(n_526)
);

BUFx10_ASAP7_75t_L g527 ( 
.A(n_359),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_413),
.Y(n_528)
);

AOI22xp33_ASAP7_75t_L g529 ( 
.A1(n_359),
.A2(n_196),
.B1(n_268),
.B2(n_187),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_413),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_413),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g533 ( 
.A(n_398),
.B(n_342),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_359),
.B(n_141),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_359),
.B(n_407),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_413),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_413),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_413),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_413),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_347),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_356),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_359),
.B(n_295),
.Y(n_542)
);

BUFx8_ASAP7_75t_SL g543 ( 
.A(n_400),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_375),
.Y(n_544)
);

BUFx6f_ASAP7_75t_SL g545 ( 
.A(n_410),
.Y(n_545)
);

BUFx4f_ASAP7_75t_L g546 ( 
.A(n_355),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_401),
.B(n_342),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_374),
.Y(n_548)
);

INVx4_ASAP7_75t_L g549 ( 
.A(n_410),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_403),
.B(n_266),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_403),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_356),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_405),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_374),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_400),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_358),
.B(n_187),
.Y(n_556)
);

OAI22xp33_ASAP7_75t_L g557 ( 
.A1(n_349),
.A2(n_236),
.B1(n_177),
.B2(n_198),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_356),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_410),
.A2(n_196),
.B1(n_217),
.B2(n_202),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_405),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_409),
.B(n_271),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_356),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g563 ( 
.A(n_409),
.B(n_283),
.Y(n_563)
);

BUFx8_ASAP7_75t_SL g564 ( 
.A(n_410),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_540),
.B(n_412),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_448),
.B(n_415),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_517),
.B(n_415),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_517),
.B(n_375),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_444),
.B(n_375),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_467),
.B(n_440),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_449),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_541),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_479),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_467),
.B(n_375),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_444),
.B(n_382),
.Y(n_576)
);

OAI22xp33_ASAP7_75t_L g577 ( 
.A1(n_472),
.A2(n_349),
.B1(n_376),
.B2(n_379),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_467),
.B(n_382),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_425),
.B(n_382),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_429),
.Y(n_580)
);

AOI22xp33_ASAP7_75t_L g581 ( 
.A1(n_431),
.A2(n_408),
.B1(n_406),
.B2(n_393),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_432),
.B(n_284),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_418),
.B(n_382),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_504),
.B(n_383),
.Y(n_584)
);

AOI22xp33_ASAP7_75t_L g585 ( 
.A1(n_431),
.A2(n_408),
.B1(n_406),
.B2(n_393),
.Y(n_585)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_480),
.A2(n_379),
.B1(n_376),
.B2(n_380),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_425),
.B(n_383),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_459),
.Y(n_589)
);

NOR2xp67_ASAP7_75t_L g590 ( 
.A(n_478),
.B(n_380),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_425),
.B(n_383),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_424),
.B(n_384),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_475),
.B(n_384),
.Y(n_593)
);

NOR2xp67_ASAP7_75t_L g594 ( 
.A(n_426),
.B(n_386),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_428),
.B(n_386),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_541),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_456),
.B(n_386),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_552),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_513),
.B(n_393),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_454),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_465),
.B(n_393),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_454),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_460),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_492),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g606 ( 
.A(n_555),
.B(n_406),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_545),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_510),
.B(n_406),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_464),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_512),
.B(n_408),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_471),
.B(n_374),
.Y(n_611)
);

BUFx6f_ASAP7_75t_SL g612 ( 
.A(n_470),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_473),
.B(n_374),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_435),
.B(n_295),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_522),
.B(n_374),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_558),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_524),
.B(n_189),
.Y(n_618)
);

OR2x2_ASAP7_75t_SL g619 ( 
.A(n_542),
.B(n_299),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_493),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_494),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_556),
.B(n_364),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_495),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_527),
.B(n_465),
.Y(n_624)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_466),
.B(n_364),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_L g626 ( 
.A1(n_463),
.A2(n_248),
.B(n_192),
.C(n_194),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_465),
.B(n_257),
.Y(n_627)
);

AO221x1_ASAP7_75t_L g628 ( 
.A1(n_474),
.A2(n_230),
.B1(n_192),
.B2(n_194),
.C(n_197),
.Y(n_628)
);

BUFx8_ASAP7_75t_L g629 ( 
.A(n_542),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_556),
.B(n_364),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_558),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_562),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_562),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_496),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_465),
.B(n_257),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_500),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_556),
.B(n_364),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_544),
.Y(n_638)
);

AND2x4_ASAP7_75t_L g639 ( 
.A(n_472),
.B(n_197),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_514),
.B(n_497),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_514),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_544),
.Y(n_643)
);

NAND2x1p5_ASAP7_75t_L g644 ( 
.A(n_549),
.B(n_364),
.Y(n_644)
);

NOR3xp33_ASAP7_75t_L g645 ( 
.A(n_416),
.B(n_202),
.C(n_200),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_501),
.B(n_551),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_553),
.B(n_366),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_549),
.B(n_204),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_422),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_560),
.B(n_366),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_497),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_533),
.B(n_366),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_533),
.B(n_366),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_514),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_509),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_509),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_490),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_437),
.B(n_446),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_450),
.B(n_300),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_422),
.Y(n_660)
);

NAND2xp33_ASAP7_75t_L g661 ( 
.A(n_514),
.B(n_355),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_431),
.A2(n_253),
.B1(n_200),
.B2(n_268),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_521),
.B(n_350),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_514),
.B(n_144),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_521),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_453),
.B(n_207),
.Y(n_666)
);

BUFx6f_ASAP7_75t_SL g667 ( 
.A(n_470),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_523),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_545),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_SL g670 ( 
.A(n_490),
.B(n_212),
.Y(n_670)
);

AOI22xp5_ASAP7_75t_L g671 ( 
.A1(n_523),
.A2(n_144),
.B1(n_244),
.B2(n_176),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_472),
.A2(n_244),
.B1(n_222),
.B2(n_270),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_423),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_548),
.B(n_350),
.Y(n_674)
);

INVx2_ASAP7_75t_SL g675 ( 
.A(n_498),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_535),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_472),
.Y(n_677)
);

BUFx5_ASAP7_75t_L g678 ( 
.A(n_417),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_561),
.B(n_303),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_548),
.B(n_264),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_548),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_554),
.B(n_161),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_554),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_554),
.B(n_352),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_436),
.B(n_161),
.Y(n_685)
);

AOI22xp5_ASAP7_75t_L g686 ( 
.A1(n_458),
.A2(n_222),
.B1(n_209),
.B2(n_267),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_476),
.B(n_213),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_547),
.Y(n_688)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_545),
.A2(n_563),
.B1(n_492),
.B2(n_470),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_499),
.B(n_489),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_436),
.A2(n_373),
.B(n_372),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_499),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_499),
.B(n_529),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_557),
.B(n_352),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_559),
.B(n_357),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_433),
.B(n_357),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_423),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_526),
.B(n_363),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_534),
.B(n_363),
.Y(n_699)
);

NOR3xp33_ASAP7_75t_L g700 ( 
.A(n_488),
.B(n_550),
.C(n_487),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_470),
.B(n_214),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_491),
.B(n_216),
.Y(n_702)
);

BUFx6f_ASAP7_75t_SL g703 ( 
.A(n_449),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_419),
.B(n_370),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_417),
.Y(n_705)
);

AOI22xp5_ASAP7_75t_L g706 ( 
.A1(n_485),
.A2(n_180),
.B1(n_186),
.B2(n_184),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_546),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_419),
.B(n_372),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_421),
.B(n_372),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_564),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_427),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_421),
.B(n_373),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_421),
.B(n_373),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_441),
.B(n_217),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_461),
.B(n_219),
.Y(n_715)
);

BUFx3_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_436),
.B(n_161),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_546),
.Y(n_718)
);

INVx8_ASAP7_75t_L g719 ( 
.A(n_543),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_441),
.B(n_219),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_484),
.B(n_161),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_420),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_441),
.B(n_227),
.Y(n_723)
);

INVx3_ASAP7_75t_L g724 ( 
.A(n_442),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_442),
.B(n_227),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_420),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_442),
.B(n_233),
.Y(n_727)
);

NOR3xp33_ASAP7_75t_L g728 ( 
.A(n_487),
.B(n_253),
.C(n_248),
.Y(n_728)
);

OAI221xp5_ASAP7_75t_L g729 ( 
.A1(n_438),
.A2(n_233),
.B1(n_237),
.B2(n_239),
.C(n_242),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_462),
.B(n_237),
.Y(n_730)
);

INVx6_ASAP7_75t_L g731 ( 
.A(n_607),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_620),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_577),
.B(n_484),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_571),
.B(n_543),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_582),
.B(n_313),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_621),
.Y(n_736)
);

AOI21xp5_ASAP7_75t_L g737 ( 
.A1(n_567),
.A2(n_484),
.B(n_439),
.Y(n_737)
);

BUFx6f_ASAP7_75t_L g738 ( 
.A(n_707),
.Y(n_738)
);

AND2x6_ASAP7_75t_L g739 ( 
.A(n_677),
.B(n_438),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_690),
.A2(n_447),
.B(n_439),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_577),
.B(n_590),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_596),
.Y(n_742)
);

AOI21xp5_ASAP7_75t_L g743 ( 
.A1(n_646),
.A2(n_451),
.B(n_447),
.Y(n_743)
);

AND2x2_ASAP7_75t_SL g744 ( 
.A(n_607),
.B(n_546),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_593),
.B(n_592),
.Y(n_745)
);

AOI21xp5_ASAP7_75t_L g746 ( 
.A1(n_584),
.A2(n_452),
.B(n_451),
.Y(n_746)
);

NOR2xp67_ASAP7_75t_L g747 ( 
.A(n_572),
.B(n_600),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_677),
.B(n_477),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_593),
.B(n_462),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_598),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_707),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_623),
.Y(n_752)
);

OAI21xp5_ASAP7_75t_L g753 ( 
.A1(n_592),
.A2(n_483),
.B(n_452),
.Y(n_753)
);

NOR2xp33_ASAP7_75t_L g754 ( 
.A(n_688),
.B(n_462),
.Y(n_754)
);

AOI22xp33_ASAP7_75t_L g755 ( 
.A1(n_702),
.A2(n_662),
.B1(n_628),
.B2(n_715),
.Y(n_755)
);

AO21x1_ASAP7_75t_L g756 ( 
.A1(n_583),
.A2(n_597),
.B(n_595),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_606),
.B(n_468),
.Y(n_757)
);

INVx3_ASAP7_75t_L g758 ( 
.A(n_707),
.Y(n_758)
);

NOR2xp67_ASAP7_75t_L g759 ( 
.A(n_602),
.B(n_468),
.Y(n_759)
);

O2A1O1Ixp33_ASAP7_75t_SL g760 ( 
.A1(n_579),
.A2(n_505),
.B(n_538),
.C(n_483),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_566),
.A2(n_468),
.B1(n_518),
.B2(n_486),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_598),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_606),
.B(n_486),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_657),
.B(n_266),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_659),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_675),
.B(n_266),
.Y(n_766)
);

INVx3_ASAP7_75t_L g767 ( 
.A(n_707),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_674),
.A2(n_505),
.B(n_503),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_618),
.B(n_518),
.Y(n_769)
);

BUFx12f_ASAP7_75t_L g770 ( 
.A(n_629),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_702),
.A2(n_648),
.B1(n_568),
.B2(n_666),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_638),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_684),
.A2(n_507),
.B(n_503),
.Y(n_773)
);

O2A1O1Ixp33_ASAP7_75t_L g774 ( 
.A1(n_652),
.A2(n_239),
.B(n_242),
.C(n_538),
.Y(n_774)
);

OAI22xp5_ASAP7_75t_L g775 ( 
.A1(n_586),
.A2(n_519),
.B1(n_508),
.B2(n_515),
.Y(n_775)
);

AOI21xp5_ASAP7_75t_L g776 ( 
.A1(n_599),
.A2(n_508),
.B(n_507),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_608),
.B(n_610),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_575),
.B(n_519),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_578),
.B(n_427),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_708),
.A2(n_516),
.B(n_515),
.Y(n_780)
);

INVx3_ASAP7_75t_L g781 ( 
.A(n_718),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_648),
.B(n_634),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_638),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_636),
.B(n_430),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_669),
.B(n_477),
.Y(n_785)
);

NOR2x1p5_ASAP7_75t_L g786 ( 
.A(n_710),
.B(n_224),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_641),
.B(n_430),
.Y(n_787)
);

AOI21xp33_ASAP7_75t_L g788 ( 
.A1(n_687),
.A2(n_516),
.B(n_525),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_710),
.Y(n_789)
);

OAI21xp33_ASAP7_75t_L g790 ( 
.A1(n_687),
.A2(n_254),
.B(n_235),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_665),
.A2(n_525),
.B1(n_530),
.B2(n_531),
.Y(n_791)
);

AOI22xp5_ASAP7_75t_L g792 ( 
.A1(n_666),
.A2(n_530),
.B1(n_531),
.B2(n_532),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_580),
.Y(n_793)
);

AND2x4_ASAP7_75t_L g794 ( 
.A(n_669),
.B(n_477),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_709),
.A2(n_532),
.B(n_537),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_629),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_595),
.B(n_434),
.Y(n_797)
);

HB1xp67_ASAP7_75t_L g798 ( 
.A(n_605),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_565),
.B(n_434),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_643),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_597),
.B(n_443),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_716),
.Y(n_802)
);

AOI21x1_ASAP7_75t_L g803 ( 
.A1(n_685),
.A2(n_539),
.B(n_537),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_676),
.B(n_443),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_653),
.B(n_445),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_643),
.Y(n_806)
);

AND2x4_ASAP7_75t_L g807 ( 
.A(n_639),
.B(n_477),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_712),
.A2(n_539),
.B(n_536),
.Y(n_808)
);

AOI21xp5_ASAP7_75t_L g809 ( 
.A1(n_713),
.A2(n_536),
.B(n_528),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_574),
.B(n_445),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_SL g811 ( 
.A(n_679),
.B(n_266),
.Y(n_811)
);

OAI21xp5_ASAP7_75t_L g812 ( 
.A1(n_570),
.A2(n_528),
.B(n_520),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_704),
.A2(n_520),
.B(n_506),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_588),
.B(n_457),
.Y(n_814)
);

OR2x6_ASAP7_75t_L g815 ( 
.A(n_719),
.B(n_457),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_589),
.B(n_481),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_604),
.B(n_481),
.Y(n_817)
);

HB1xp67_ASAP7_75t_L g818 ( 
.A(n_639),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_609),
.B(n_482),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_611),
.B(n_482),
.Y(n_820)
);

AOI21x1_ASAP7_75t_L g821 ( 
.A1(n_685),
.A2(n_369),
.B(n_367),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_678),
.B(n_469),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_615),
.B(n_249),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_R g824 ( 
.A(n_719),
.B(n_469),
.Y(n_824)
);

AO21x1_ASAP7_75t_L g825 ( 
.A1(n_658),
.A2(n_367),
.B(n_369),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_613),
.B(n_251),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_718),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_718),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_640),
.A2(n_153),
.B(n_265),
.Y(n_829)
);

INVx4_ASAP7_75t_L g830 ( 
.A(n_719),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_640),
.A2(n_142),
.B(n_262),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_579),
.A2(n_591),
.B(n_587),
.Y(n_832)
);

INVxp67_ASAP7_75t_L g833 ( 
.A(n_569),
.Y(n_833)
);

AO21x2_ASAP7_75t_L g834 ( 
.A1(n_664),
.A2(n_367),
.B(n_369),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_573),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_616),
.B(n_658),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_647),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_718),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_603),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_644),
.Y(n_840)
);

INVx1_ASAP7_75t_SL g841 ( 
.A(n_619),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_587),
.A2(n_229),
.B(n_168),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_581),
.B(n_255),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_689),
.B(n_256),
.Y(n_844)
);

O2A1O1Ixp33_ASAP7_75t_SL g845 ( 
.A1(n_591),
.A2(n_367),
.B(n_369),
.C(n_11),
.Y(n_845)
);

OAI22xp5_ASAP7_75t_L g846 ( 
.A1(n_668),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_846)
);

OAI21xp5_ASAP7_75t_L g847 ( 
.A1(n_570),
.A2(n_355),
.B(n_469),
.Y(n_847)
);

BUFx4f_ASAP7_75t_L g848 ( 
.A(n_715),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_585),
.B(n_263),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_614),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_576),
.A2(n_355),
.B(n_511),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_585),
.B(n_230),
.Y(n_852)
);

AOI21xp33_ASAP7_75t_L g853 ( 
.A1(n_701),
.A2(n_215),
.B(n_171),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_693),
.B(n_625),
.Y(n_854)
);

O2A1O1Ixp33_ASAP7_75t_L g855 ( 
.A1(n_576),
.A2(n_8),
.B(n_9),
.C(n_14),
.Y(n_855)
);

OAI21xp5_ASAP7_75t_L g856 ( 
.A1(n_681),
.A2(n_355),
.B(n_511),
.Y(n_856)
);

NAND3xp33_ASAP7_75t_L g857 ( 
.A(n_728),
.B(n_230),
.C(n_164),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_622),
.B(n_172),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_L g859 ( 
.A1(n_630),
.A2(n_9),
.B(n_14),
.C(n_15),
.Y(n_859)
);

NOR2x2_ASAP7_75t_L g860 ( 
.A(n_703),
.B(n_16),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_637),
.B(n_179),
.Y(n_861)
);

AOI22x1_ASAP7_75t_L g862 ( 
.A1(n_683),
.A2(n_365),
.B1(n_368),
.B2(n_181),
.Y(n_862)
);

NOR2xp33_ASAP7_75t_L g863 ( 
.A(n_651),
.B(n_655),
.Y(n_863)
);

OAI22xp5_ASAP7_75t_L g864 ( 
.A1(n_594),
.A2(n_241),
.B1(n_193),
.B2(n_203),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_603),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_617),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_662),
.B(n_365),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_670),
.B(n_16),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_612),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_650),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_645),
.B(n_191),
.Y(n_871)
);

INVx3_ASAP7_75t_L g872 ( 
.A(n_644),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_656),
.B(n_221),
.Y(n_873)
);

A2O1A1Ixp33_ASAP7_75t_L g874 ( 
.A1(n_729),
.A2(n_368),
.B(n_365),
.C(n_243),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_678),
.B(n_511),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_706),
.B(n_240),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_672),
.B(n_18),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_680),
.A2(n_726),
.B(n_722),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_686),
.B(n_671),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_680),
.A2(n_511),
.B(n_469),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_631),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_705),
.A2(n_511),
.B(n_469),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_724),
.B(n_19),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_632),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_633),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_714),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_724),
.B(n_19),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_692),
.A2(n_365),
.B(n_368),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_720),
.Y(n_889)
);

INVx3_ASAP7_75t_L g890 ( 
.A(n_603),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_700),
.B(n_368),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_SL g892 ( 
.A(n_678),
.B(n_368),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_612),
.A2(n_667),
.B1(n_624),
.B2(n_694),
.Y(n_893)
);

AND2x2_ASAP7_75t_SL g894 ( 
.A(n_661),
.B(n_368),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_667),
.B(n_21),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_649),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_603),
.Y(n_897)
);

INVx4_ASAP7_75t_L g898 ( 
.A(n_703),
.Y(n_898)
);

BUFx3_ASAP7_75t_L g899 ( 
.A(n_642),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_601),
.A2(n_624),
.B(n_711),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_723),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_725),
.B(n_21),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_642),
.A2(n_654),
.B1(n_663),
.B2(n_730),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_727),
.B(n_26),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_626),
.B(n_27),
.Y(n_905)
);

O2A1O1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_696),
.A2(n_28),
.B(n_31),
.C(n_33),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_698),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_745),
.B(n_673),
.Y(n_908)
);

BUFx12f_ASAP7_75t_L g909 ( 
.A(n_770),
.Y(n_909)
);

OAI22xp5_ASAP7_75t_L g910 ( 
.A1(n_782),
.A2(n_654),
.B1(n_642),
.B2(n_699),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_732),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_734),
.A2(n_627),
.B1(n_635),
.B2(n_721),
.Y(n_912)
);

BUFx8_ASAP7_75t_SL g913 ( 
.A(n_789),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_783),
.Y(n_914)
);

BUFx4f_ASAP7_75t_L g915 ( 
.A(n_796),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_798),
.Y(n_916)
);

NOR2xp67_ASAP7_75t_L g917 ( 
.A(n_898),
.B(n_627),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_833),
.B(n_660),
.Y(n_918)
);

OAI22xp5_ASAP7_75t_L g919 ( 
.A1(n_777),
.A2(n_654),
.B1(n_682),
.B2(n_695),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_789),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_833),
.B(n_836),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_734),
.B(n_654),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_783),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_797),
.A2(n_682),
.B(n_717),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_907),
.B(n_697),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_L g926 ( 
.A(n_811),
.B(n_721),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_844),
.B(n_678),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_741),
.A2(n_691),
.B(n_368),
.C(n_365),
.Y(n_928)
);

AO32x2_ASAP7_75t_L g929 ( 
.A1(n_903),
.A2(n_678),
.A3(n_368),
.B1(n_365),
.B2(n_39),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_879),
.A2(n_33),
.B(n_36),
.C(n_37),
.Y(n_930)
);

INVx3_ASAP7_75t_L g931 ( 
.A(n_785),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_736),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_877),
.A2(n_40),
.B(n_41),
.C(n_45),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_800),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_844),
.A2(n_678),
.B1(n_355),
.B2(n_365),
.Y(n_935)
);

AOI22xp5_ASAP7_75t_L g936 ( 
.A1(n_747),
.A2(n_355),
.B1(n_365),
.B2(n_48),
.Y(n_936)
);

AND2x2_ASAP7_75t_SL g937 ( 
.A(n_755),
.B(n_45),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_848),
.B(n_46),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_752),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_765),
.B(n_50),
.Y(n_940)
);

OAI22xp5_ASAP7_75t_L g941 ( 
.A1(n_755),
.A2(n_733),
.B1(n_793),
.B2(n_749),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_SL g942 ( 
.A(n_848),
.B(n_51),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_823),
.A2(n_51),
.B1(n_53),
.B2(n_56),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_772),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_SL g945 ( 
.A1(n_895),
.A2(n_53),
.B1(n_64),
.B2(n_65),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_748),
.B(n_70),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_735),
.B(n_74),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_798),
.B(n_818),
.Y(n_948)
);

OR2x2_ASAP7_75t_L g949 ( 
.A(n_818),
.B(n_841),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_754),
.A2(n_77),
.B(n_79),
.C(n_85),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_764),
.B(n_86),
.Y(n_951)
);

INVx1_ASAP7_75t_SL g952 ( 
.A(n_824),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_739),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_806),
.Y(n_954)
);

OR2x6_ASAP7_75t_L g955 ( 
.A(n_807),
.B(n_133),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_866),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_750),
.Y(n_957)
);

OAI22xp5_ASAP7_75t_L g958 ( 
.A1(n_733),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_837),
.B(n_99),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_790),
.B(n_101),
.Y(n_960)
);

OR2x6_ASAP7_75t_SL g961 ( 
.A(n_868),
.B(n_106),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_748),
.B(n_110),
.Y(n_962)
);

AOI22x1_ASAP7_75t_L g963 ( 
.A1(n_737),
.A2(n_115),
.B1(n_118),
.B2(n_121),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_766),
.B(n_126),
.Y(n_964)
);

OAI22xp5_ASAP7_75t_L g965 ( 
.A1(n_757),
.A2(n_763),
.B1(n_754),
.B2(n_870),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_895),
.B(n_802),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_886),
.B(n_889),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_802),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_824),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_881),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_785),
.Y(n_971)
);

A2O1A1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_832),
.A2(n_788),
.B(n_901),
.C(n_855),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_801),
.A2(n_753),
.B(n_892),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_807),
.B(n_840),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_756),
.B(n_750),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_884),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_830),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_762),
.B(n_739),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_840),
.B(n_738),
.Y(n_979)
);

OAI21xp33_ASAP7_75t_SL g980 ( 
.A1(n_894),
.A2(n_792),
.B(n_887),
.Y(n_980)
);

BUFx3_ASAP7_75t_L g981 ( 
.A(n_830),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_762),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_898),
.Y(n_983)
);

BUFx3_ASAP7_75t_L g984 ( 
.A(n_815),
.Y(n_984)
);

BUFx4f_ASAP7_75t_L g985 ( 
.A(n_731),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_905),
.A2(n_904),
.B1(n_902),
.B2(n_819),
.Y(n_986)
);

OAI22x1_ASAP7_75t_L g987 ( 
.A1(n_893),
.A2(n_786),
.B1(n_869),
.B2(n_857),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_835),
.Y(n_988)
);

OAI21xp33_ASAP7_75t_L g989 ( 
.A1(n_826),
.A2(n_853),
.B(n_846),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_803),
.A2(n_825),
.B(n_821),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_835),
.Y(n_991)
);

NOR2xp67_ASAP7_75t_L g992 ( 
.A(n_869),
.B(n_876),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_739),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_815),
.B(n_867),
.Y(n_994)
);

INVx6_ASAP7_75t_L g995 ( 
.A(n_815),
.Y(n_995)
);

A2O1A1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_874),
.A2(n_906),
.B(n_863),
.C(n_774),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_738),
.B(n_751),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_892),
.A2(n_769),
.B(n_805),
.Y(n_998)
);

A2O1A1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_874),
.A2(n_863),
.B(n_878),
.C(n_799),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_871),
.B(n_843),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_814),
.A2(n_817),
.B1(n_816),
.B2(n_787),
.Y(n_1001)
);

O2A1O1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_859),
.A2(n_861),
.B(n_858),
.C(n_883),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_740),
.A2(n_776),
.B(n_813),
.Y(n_1003)
);

BUFx12f_ASAP7_75t_L g1004 ( 
.A(n_731),
.Y(n_1004)
);

OR2x2_ASAP7_75t_L g1005 ( 
.A(n_849),
.B(n_873),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_746),
.A2(n_808),
.B(n_809),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_743),
.A2(n_820),
.B(n_795),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_759),
.B(n_731),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_742),
.Y(n_1009)
);

OAI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_768),
.A2(n_773),
.B(n_780),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_779),
.B(n_850),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_896),
.Y(n_1012)
);

O2A1O1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_845),
.A2(n_760),
.B(n_791),
.C(n_775),
.Y(n_1013)
);

AO32x2_ASAP7_75t_L g1014 ( 
.A1(n_761),
.A2(n_838),
.A3(n_864),
.B1(n_845),
.B2(n_760),
.Y(n_1014)
);

AOI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_900),
.A2(n_778),
.B(n_784),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_812),
.A2(n_875),
.B(n_822),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_896),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_885),
.B(n_854),
.Y(n_1018)
);

AND2x4_ASAP7_75t_L g1019 ( 
.A(n_794),
.B(n_872),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_804),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_899),
.Y(n_1021)
);

AO32x2_ASAP7_75t_L g1022 ( 
.A1(n_838),
.A2(n_834),
.A3(n_852),
.B1(n_891),
.B2(n_862),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_799),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_899),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_834),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_822),
.A2(n_875),
.B(n_894),
.Y(n_1026)
);

OAI22xp5_ASAP7_75t_L g1027 ( 
.A1(n_810),
.A2(n_839),
.B1(n_865),
.B2(n_890),
.Y(n_1027)
);

A2O1A1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_810),
.A2(n_781),
.B(n_828),
.C(n_767),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_738),
.B(n_751),
.Y(n_1029)
);

INVx2_ASAP7_75t_SL g1030 ( 
.A(n_744),
.Y(n_1030)
);

NAND2x1_ASAP7_75t_L g1031 ( 
.A(n_758),
.B(n_767),
.Y(n_1031)
);

A2O1A1Ixp33_ASAP7_75t_L g1032 ( 
.A1(n_758),
.A2(n_828),
.B(n_781),
.C(n_842),
.Y(n_1032)
);

OAI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_839),
.A2(n_865),
.B1(n_890),
.B2(n_897),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_839),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_865),
.Y(n_1035)
);

OAI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_865),
.A2(n_897),
.B1(n_744),
.B2(n_751),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_R g1037 ( 
.A(n_738),
.B(n_751),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_827),
.B(n_847),
.Y(n_1038)
);

AO31x2_ASAP7_75t_L g1039 ( 
.A1(n_888),
.A2(n_882),
.A3(n_880),
.B(n_831),
.Y(n_1039)
);

INVxp67_ASAP7_75t_L g1040 ( 
.A(n_829),
.Y(n_1040)
);

NOR2xp33_ASAP7_75t_L g1041 ( 
.A(n_827),
.B(n_851),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_827),
.B(n_856),
.Y(n_1042)
);

INVxp67_ASAP7_75t_L g1043 ( 
.A(n_860),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_860),
.A2(n_702),
.B1(n_755),
.B2(n_615),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_R g1045 ( 
.A(n_830),
.B(n_449),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_783),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_783),
.Y(n_1047)
);

OA21x2_ASAP7_75t_L g1048 ( 
.A1(n_1006),
.A2(n_1003),
.B(n_1010),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_989),
.A2(n_996),
.B(n_986),
.C(n_938),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_965),
.A2(n_927),
.B(n_1007),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_965),
.A2(n_973),
.B(n_986),
.Y(n_1051)
);

AOI221xp5_ASAP7_75t_L g1052 ( 
.A1(n_1044),
.A2(n_941),
.B1(n_940),
.B2(n_943),
.C(n_933),
.Y(n_1052)
);

OAI21x1_ASAP7_75t_L g1053 ( 
.A1(n_990),
.A2(n_1015),
.B(n_1010),
.Y(n_1053)
);

BUFx6f_ASAP7_75t_L g1054 ( 
.A(n_985),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_999),
.A2(n_941),
.B(n_972),
.Y(n_1055)
);

INVx5_ASAP7_75t_L g1056 ( 
.A(n_913),
.Y(n_1056)
);

AO31x2_ASAP7_75t_L g1057 ( 
.A1(n_1025),
.A2(n_975),
.A3(n_1001),
.B(n_928),
.Y(n_1057)
);

AOI221xp5_ASAP7_75t_SL g1058 ( 
.A1(n_930),
.A2(n_1013),
.B1(n_916),
.B2(n_1002),
.C(n_980),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_1001),
.A2(n_998),
.B(n_908),
.Y(n_1059)
);

AO31x2_ASAP7_75t_L g1060 ( 
.A1(n_975),
.A2(n_919),
.A3(n_910),
.B(n_1016),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_1019),
.B(n_931),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_968),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_SL g1063 ( 
.A1(n_908),
.A2(n_1026),
.B(n_921),
.Y(n_1063)
);

BUFx12f_ASAP7_75t_L g1064 ( 
.A(n_909),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_920),
.Y(n_1065)
);

AO31x2_ASAP7_75t_L g1066 ( 
.A1(n_919),
.A2(n_910),
.A3(n_1027),
.B(n_1018),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_921),
.B(n_967),
.Y(n_1067)
);

AOI22xp5_ASAP7_75t_L g1068 ( 
.A1(n_937),
.A2(n_945),
.B1(n_948),
.B2(n_926),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1000),
.A2(n_942),
.B1(n_1023),
.B2(n_966),
.Y(n_1069)
);

AO31x2_ASAP7_75t_L g1070 ( 
.A1(n_1027),
.A2(n_1018),
.A3(n_924),
.B(n_1011),
.Y(n_1070)
);

INVx3_ASAP7_75t_L g1071 ( 
.A(n_953),
.Y(n_1071)
);

AO31x2_ASAP7_75t_L g1072 ( 
.A1(n_1011),
.A2(n_978),
.A3(n_959),
.B(n_1028),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_967),
.A2(n_1040),
.B(n_1036),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_1020),
.B(n_918),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_SL g1075 ( 
.A1(n_922),
.A2(n_1032),
.B(n_950),
.C(n_1031),
.Y(n_1075)
);

OAI21x1_ASAP7_75t_L g1076 ( 
.A1(n_963),
.A2(n_1042),
.B(n_1033),
.Y(n_1076)
);

OAI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_935),
.A2(n_1005),
.B(n_912),
.Y(n_1077)
);

AO21x1_ASAP7_75t_L g1078 ( 
.A1(n_960),
.A2(n_958),
.B(n_1041),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_1043),
.B(n_947),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_983),
.Y(n_1080)
);

BUFx3_ASAP7_75t_L g1081 ( 
.A(n_915),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_911),
.B(n_932),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_953),
.A2(n_993),
.B(n_1033),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_918),
.B(n_925),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_964),
.A2(n_951),
.B(n_992),
.C(n_917),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_925),
.B(n_1030),
.Y(n_1086)
);

INVx3_ASAP7_75t_SL g1087 ( 
.A(n_977),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_997),
.A2(n_1029),
.B(n_979),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_952),
.B(n_969),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_939),
.A2(n_961),
.B1(n_955),
.B2(n_962),
.Y(n_1090)
);

BUFx4f_ASAP7_75t_SL g1091 ( 
.A(n_1004),
.Y(n_1091)
);

BUFx2_ASAP7_75t_L g1092 ( 
.A(n_1024),
.Y(n_1092)
);

OAI22xp5_ASAP7_75t_L g1093 ( 
.A1(n_955),
.A2(n_946),
.B1(n_962),
.B2(n_952),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1038),
.A2(n_955),
.B(n_985),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_L g1095 ( 
.A(n_936),
.B(n_1034),
.C(n_1035),
.Y(n_1095)
);

OAI21x1_ASAP7_75t_L g1096 ( 
.A1(n_1047),
.A2(n_914),
.B(n_1046),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1034),
.A2(n_946),
.B(n_1035),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_915),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1037),
.Y(n_1099)
);

BUFx3_ASAP7_75t_L g1100 ( 
.A(n_981),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_1019),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_987),
.A2(n_991),
.B1(n_988),
.B2(n_944),
.C(n_994),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_949),
.B(n_970),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_956),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_976),
.Y(n_1105)
);

AOI221x1_ASAP7_75t_L g1106 ( 
.A1(n_923),
.A2(n_934),
.B1(n_954),
.B2(n_1021),
.C(n_957),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1009),
.B(n_982),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_931),
.B(n_971),
.Y(n_1108)
);

BUFx2_ASAP7_75t_L g1109 ( 
.A(n_1045),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1034),
.A2(n_974),
.B(n_971),
.Y(n_1110)
);

AOI21x1_ASAP7_75t_L g1111 ( 
.A1(n_1008),
.A2(n_1017),
.B(n_1012),
.Y(n_1111)
);

AO31x2_ASAP7_75t_L g1112 ( 
.A1(n_1022),
.A2(n_929),
.A3(n_1014),
.B(n_1039),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_995),
.B(n_984),
.Y(n_1113)
);

AOI22xp33_ASAP7_75t_L g1114 ( 
.A1(n_995),
.A2(n_929),
.B1(n_1014),
.B2(n_1022),
.Y(n_1114)
);

AO21x2_ASAP7_75t_L g1115 ( 
.A1(n_1022),
.A2(n_1014),
.B(n_1039),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1039),
.A2(n_990),
.B(n_1006),
.Y(n_1116)
);

OAI22x1_ASAP7_75t_L g1117 ( 
.A1(n_961),
.A2(n_689),
.B1(n_844),
.B2(n_771),
.Y(n_1117)
);

OAI21x1_ASAP7_75t_L g1118 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1003),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_921),
.B(n_745),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_921),
.B(n_745),
.Y(n_1120)
);

AND2x2_ASAP7_75t_L g1121 ( 
.A(n_948),
.B(n_615),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_948),
.B(n_615),
.Y(n_1123)
);

AOI221x1_ASAP7_75t_L g1124 ( 
.A1(n_958),
.A2(n_986),
.B1(n_941),
.B2(n_989),
.C(n_910),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_911),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_915),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_999),
.A2(n_741),
.B(n_771),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_937),
.A2(n_745),
.B1(n_771),
.B2(n_927),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_989),
.A2(n_745),
.B(n_741),
.C(n_416),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1003),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_913),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_948),
.B(n_615),
.Y(n_1134)
);

OA21x2_ASAP7_75t_L g1135 ( 
.A1(n_1006),
.A2(n_1003),
.B(n_1010),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1136)
);

O2A1O1Ixp33_ASAP7_75t_SL g1137 ( 
.A1(n_927),
.A2(n_745),
.B(n_741),
.C(n_782),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1138)
);

AO22x2_ASAP7_75t_L g1139 ( 
.A1(n_941),
.A2(n_986),
.B1(n_679),
.B2(n_741),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_913),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_989),
.A2(n_745),
.B(n_741),
.C(n_416),
.Y(n_1141)
);

O2A1O1Ixp33_ASAP7_75t_SL g1142 ( 
.A1(n_927),
.A2(n_745),
.B(n_741),
.C(n_782),
.Y(n_1142)
);

BUFx6f_ASAP7_75t_L g1143 ( 
.A(n_985),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_985),
.Y(n_1144)
);

OAI22xp33_ASAP7_75t_L g1145 ( 
.A1(n_961),
.A2(n_771),
.B1(n_811),
.B2(n_351),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1146)
);

OR2x2_ASAP7_75t_L g1147 ( 
.A(n_949),
.B(n_600),
.Y(n_1147)
);

HB1xp67_ASAP7_75t_L g1148 ( 
.A(n_948),
.Y(n_1148)
);

AOI221x1_ASAP7_75t_L g1149 ( 
.A1(n_958),
.A2(n_986),
.B1(n_941),
.B2(n_989),
.C(n_910),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_921),
.B(n_745),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_911),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_911),
.Y(n_1153)
);

AOI22xp33_ASAP7_75t_SL g1154 ( 
.A1(n_937),
.A2(n_378),
.B1(n_351),
.B2(n_811),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_920),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_911),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1003),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_948),
.B(n_615),
.Y(n_1158)
);

AOI21x1_ASAP7_75t_L g1159 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1003),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_989),
.A2(n_771),
.B(n_927),
.C(n_745),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1162)
);

INVxp67_ASAP7_75t_L g1163 ( 
.A(n_948),
.Y(n_1163)
);

NAND2x1p5_ASAP7_75t_L g1164 ( 
.A(n_952),
.B(n_969),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_999),
.A2(n_741),
.B(n_771),
.Y(n_1165)
);

AND2x2_ASAP7_75t_L g1166 ( 
.A(n_948),
.B(n_615),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1012),
.Y(n_1167)
);

AOI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_937),
.A2(n_771),
.B1(n_745),
.B2(n_1044),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_SL g1169 ( 
.A(n_920),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_911),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_921),
.B(n_745),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_915),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_L g1173 ( 
.A1(n_999),
.A2(n_741),
.B(n_771),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_990),
.A2(n_1006),
.B(n_1003),
.Y(n_1174)
);

OAI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_999),
.A2(n_741),
.B(n_771),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1176)
);

AO22x2_ASAP7_75t_L g1177 ( 
.A1(n_941),
.A2(n_986),
.B1(n_679),
.B2(n_741),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1019),
.B(n_677),
.Y(n_1178)
);

NOR2x1_ASAP7_75t_L g1179 ( 
.A(n_920),
.B(n_898),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_965),
.A2(n_777),
.B(n_927),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_921),
.B(n_745),
.Y(n_1181)
);

AND2x2_ASAP7_75t_SL g1182 ( 
.A(n_937),
.B(n_1044),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_1019),
.B(n_677),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_909),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_913),
.Y(n_1185)
);

NAND2xp5_ASAP7_75t_SL g1186 ( 
.A(n_927),
.B(n_771),
.Y(n_1186)
);

INVx5_ASAP7_75t_L g1187 ( 
.A(n_913),
.Y(n_1187)
);

HB1xp67_ASAP7_75t_L g1188 ( 
.A(n_1148),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1182),
.A2(n_1154),
.B1(n_1145),
.B2(n_1168),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1082),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1119),
.B(n_1151),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_1126),
.Y(n_1192)
);

INVx6_ASAP7_75t_L g1193 ( 
.A(n_1054),
.Y(n_1193)
);

AOI21xp33_ASAP7_75t_L g1194 ( 
.A1(n_1049),
.A2(n_1177),
.B(n_1139),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1168),
.A2(n_1052),
.B1(n_1129),
.B2(n_1117),
.Y(n_1195)
);

BUFx3_ASAP7_75t_L g1196 ( 
.A(n_1099),
.Y(n_1196)
);

CKINVDCx11_ASAP7_75t_R g1197 ( 
.A(n_1184),
.Y(n_1197)
);

OAI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1068),
.A2(n_1129),
.B1(n_1124),
.B2(n_1149),
.Y(n_1198)
);

INVx5_ASAP7_75t_L g1199 ( 
.A(n_1071),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1054),
.Y(n_1200)
);

CKINVDCx11_ASAP7_75t_R g1201 ( 
.A(n_1080),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1171),
.B(n_1181),
.Y(n_1202)
);

INVx6_ASAP7_75t_L g1203 ( 
.A(n_1054),
.Y(n_1203)
);

INVx4_ASAP7_75t_L g1204 ( 
.A(n_1091),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1139),
.A2(n_1177),
.B1(n_1090),
.B2(n_1186),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1090),
.A2(n_1093),
.B1(n_1077),
.B2(n_1165),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1068),
.A2(n_1128),
.B1(n_1175),
.B2(n_1165),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1120),
.B(n_1067),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_1160),
.A2(n_1120),
.B1(n_1133),
.B2(n_1136),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1092),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_1147),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1093),
.A2(n_1158),
.B1(n_1166),
.B2(n_1121),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1067),
.B(n_1163),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_SL g1214 ( 
.A1(n_1077),
.A2(n_1175),
.B1(n_1128),
.B2(n_1173),
.Y(n_1214)
);

CKINVDCx20_ASAP7_75t_R g1215 ( 
.A(n_1062),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1143),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1123),
.A2(n_1134),
.B1(n_1173),
.B2(n_1078),
.Y(n_1217)
);

INVx1_ASAP7_75t_SL g1218 ( 
.A(n_1155),
.Y(n_1218)
);

AOI22x1_ASAP7_75t_SL g1219 ( 
.A1(n_1140),
.A2(n_1185),
.B1(n_1098),
.B2(n_1056),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1079),
.B(n_1061),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_1056),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1152),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1153),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1132),
.Y(n_1224)
);

AOI22xp33_ASAP7_75t_L g1225 ( 
.A1(n_1055),
.A2(n_1162),
.B1(n_1125),
.B2(n_1122),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1055),
.A2(n_1161),
.B1(n_1176),
.B2(n_1146),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1156),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1138),
.A2(n_1150),
.B(n_1180),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1170),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1061),
.B(n_1178),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1056),
.Y(n_1231)
);

CKINVDCx6p67_ASAP7_75t_R g1232 ( 
.A(n_1187),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1143),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1104),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1105),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1107),
.Y(n_1236)
);

NAND2x1p5_ASAP7_75t_L g1237 ( 
.A(n_1071),
.B(n_1143),
.Y(n_1237)
);

AOI22xp33_ASAP7_75t_L g1238 ( 
.A1(n_1084),
.A2(n_1074),
.B1(n_1069),
.B2(n_1086),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1130),
.A2(n_1141),
.B(n_1051),
.Y(n_1239)
);

BUFx2_ASAP7_75t_L g1240 ( 
.A(n_1065),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1107),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1084),
.B(n_1069),
.Y(n_1242)
);

BUFx10_ASAP7_75t_L g1243 ( 
.A(n_1144),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1086),
.A2(n_1103),
.B1(n_1114),
.B2(n_1063),
.Y(n_1244)
);

CKINVDCx11_ASAP7_75t_R g1245 ( 
.A(n_1109),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1096),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1089),
.Y(n_1247)
);

BUFx4f_ASAP7_75t_SL g1248 ( 
.A(n_1081),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1073),
.A2(n_1094),
.B1(n_1167),
.B2(n_1183),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_1144),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1089),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1164),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1101),
.B(n_1164),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1169),
.A2(n_1050),
.B1(n_1101),
.B2(n_1095),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1100),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1187),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1101),
.A2(n_1059),
.B1(n_1115),
.B2(n_1113),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1106),
.Y(n_1258)
);

BUFx2_ASAP7_75t_L g1259 ( 
.A(n_1179),
.Y(n_1259)
);

INVx3_ASAP7_75t_L g1260 ( 
.A(n_1088),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1115),
.A2(n_1108),
.B1(n_1083),
.B2(n_1127),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1070),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1070),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1070),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_1172),
.Y(n_1265)
);

INVx6_ASAP7_75t_L g1266 ( 
.A(n_1097),
.Y(n_1266)
);

INVx6_ASAP7_75t_L g1267 ( 
.A(n_1110),
.Y(n_1267)
);

AOI211xp5_ASAP7_75t_L g1268 ( 
.A1(n_1085),
.A2(n_1058),
.B(n_1142),
.C(n_1137),
.Y(n_1268)
);

BUFx12f_ASAP7_75t_L g1269 ( 
.A(n_1102),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1111),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1058),
.A2(n_1048),
.B1(n_1135),
.B2(n_1159),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1066),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1066),
.B(n_1112),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1048),
.Y(n_1274)
);

BUFx6f_ASAP7_75t_L g1275 ( 
.A(n_1076),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1135),
.A2(n_1053),
.B1(n_1116),
.B2(n_1066),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1072),
.B(n_1060),
.Y(n_1277)
);

CKINVDCx14_ASAP7_75t_R g1278 ( 
.A(n_1075),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1057),
.Y(n_1279)
);

AOI22x1_ASAP7_75t_L g1280 ( 
.A1(n_1118),
.A2(n_1131),
.B1(n_1157),
.B2(n_1174),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1057),
.Y(n_1281)
);

BUFx2_ASAP7_75t_L g1282 ( 
.A(n_1060),
.Y(n_1282)
);

INVx6_ASAP7_75t_L g1283 ( 
.A(n_1060),
.Y(n_1283)
);

INVx4_ASAP7_75t_L g1284 ( 
.A(n_1057),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1112),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1112),
.A2(n_1168),
.B1(n_1068),
.B2(n_1129),
.Y(n_1286)
);

NAND2x1p5_ASAP7_75t_L g1287 ( 
.A(n_1099),
.B(n_952),
.Y(n_1287)
);

INVx3_ASAP7_75t_L g1288 ( 
.A(n_1061),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1091),
.Y(n_1289)
);

OAI22xp33_ASAP7_75t_L g1290 ( 
.A1(n_1168),
.A2(n_1068),
.B1(n_1129),
.B2(n_771),
.Y(n_1290)
);

INVx8_ASAP7_75t_L g1291 ( 
.A(n_1064),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1168),
.A2(n_1068),
.B1(n_1129),
.B2(n_771),
.Y(n_1292)
);

CKINVDCx11_ASAP7_75t_R g1293 ( 
.A(n_1064),
.Y(n_1293)
);

INVx8_ASAP7_75t_L g1294 ( 
.A(n_1064),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1064),
.Y(n_1295)
);

BUFx3_ASAP7_75t_L g1296 ( 
.A(n_1099),
.Y(n_1296)
);

AOI22xp33_ASAP7_75t_SL g1297 ( 
.A1(n_1182),
.A2(n_937),
.B1(n_811),
.B2(n_1090),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1082),
.Y(n_1298)
);

INVx2_ASAP7_75t_SL g1299 ( 
.A(n_1091),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1082),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1082),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1082),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1082),
.Y(n_1303)
);

INVx1_ASAP7_75t_SL g1304 ( 
.A(n_1087),
.Y(n_1304)
);

CKINVDCx6p67_ASAP7_75t_R g1305 ( 
.A(n_1056),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1082),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1182),
.A2(n_937),
.B1(n_1154),
.B2(n_1145),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1082),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1263),
.Y(n_1309)
);

AOI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1290),
.A2(n_1292),
.B1(n_1297),
.B2(n_1307),
.Y(n_1310)
);

OAI21x1_ASAP7_75t_L g1311 ( 
.A1(n_1280),
.A2(n_1228),
.B(n_1239),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1264),
.Y(n_1312)
);

BUFx5_ASAP7_75t_L g1313 ( 
.A(n_1272),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1307),
.A2(n_1189),
.B1(n_1290),
.B2(n_1292),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1188),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1273),
.B(n_1192),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1189),
.A2(n_1206),
.B1(n_1195),
.B2(n_1207),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1260),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1213),
.B(n_1208),
.Y(n_1319)
);

BUFx2_ASAP7_75t_L g1320 ( 
.A(n_1260),
.Y(n_1320)
);

AND2x4_ASAP7_75t_SL g1321 ( 
.A(n_1254),
.B(n_1249),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1285),
.Y(n_1322)
);

HB1xp67_ASAP7_75t_L g1323 ( 
.A(n_1210),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1247),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1277),
.A2(n_1276),
.B(n_1226),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1191),
.B(n_1202),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1274),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1285),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1272),
.B(n_1251),
.Y(n_1329)
);

BUFx2_ASAP7_75t_L g1330 ( 
.A(n_1274),
.Y(n_1330)
);

AOI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1209),
.A2(n_1225),
.B(n_1226),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1285),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1252),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1271),
.A2(n_1276),
.B(n_1225),
.Y(n_1334)
);

BUFx4f_ASAP7_75t_SL g1335 ( 
.A(n_1215),
.Y(n_1335)
);

BUFx6f_ASAP7_75t_L g1336 ( 
.A(n_1283),
.Y(n_1336)
);

AO21x2_ASAP7_75t_L g1337 ( 
.A1(n_1198),
.A2(n_1258),
.B(n_1194),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1248),
.B(n_1240),
.Y(n_1338)
);

HB1xp67_ASAP7_75t_L g1339 ( 
.A(n_1222),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1223),
.B(n_1227),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1229),
.B(n_1214),
.Y(n_1341)
);

AOI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1282),
.A2(n_1262),
.B(n_1281),
.Y(n_1342)
);

INVxp67_ASAP7_75t_L g1343 ( 
.A(n_1265),
.Y(n_1343)
);

AOI222xp33_ASAP7_75t_L g1344 ( 
.A1(n_1195),
.A2(n_1207),
.B1(n_1198),
.B2(n_1286),
.C1(n_1217),
.C2(n_1205),
.Y(n_1344)
);

AO21x1_ASAP7_75t_L g1345 ( 
.A1(n_1286),
.A2(n_1268),
.B(n_1242),
.Y(n_1345)
);

INVx5_ASAP7_75t_L g1346 ( 
.A(n_1283),
.Y(n_1346)
);

INVx2_ASAP7_75t_SL g1347 ( 
.A(n_1266),
.Y(n_1347)
);

OA21x2_ASAP7_75t_L g1348 ( 
.A1(n_1262),
.A2(n_1279),
.B(n_1257),
.Y(n_1348)
);

AO211x2_ASAP7_75t_L g1349 ( 
.A1(n_1217),
.A2(n_1269),
.B(n_1205),
.C(n_1278),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1234),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1257),
.A2(n_1261),
.B(n_1254),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1248),
.B(n_1304),
.Y(n_1352)
);

BUFx2_ASAP7_75t_L g1353 ( 
.A(n_1283),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1235),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1246),
.A2(n_1270),
.B(n_1241),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_1218),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1236),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1212),
.B(n_1261),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1284),
.B(n_1256),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1190),
.B(n_1308),
.Y(n_1360)
);

NOR2xp33_ASAP7_75t_L g1361 ( 
.A(n_1196),
.B(n_1296),
.Y(n_1361)
);

OA21x2_ASAP7_75t_L g1362 ( 
.A1(n_1244),
.A2(n_1238),
.B(n_1303),
.Y(n_1362)
);

INVx2_ASAP7_75t_L g1363 ( 
.A(n_1275),
.Y(n_1363)
);

AND2x2_ASAP7_75t_L g1364 ( 
.A(n_1298),
.B(n_1300),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1301),
.B(n_1302),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1275),
.Y(n_1366)
);

HB1xp67_ASAP7_75t_L g1367 ( 
.A(n_1306),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1211),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1253),
.A2(n_1269),
.B(n_1259),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1287),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1266),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1220),
.B(n_1288),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1266),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1237),
.A2(n_1288),
.B(n_1230),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1199),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1199),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1199),
.A2(n_1237),
.B(n_1299),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1199),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1200),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1200),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_1255),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1200),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1200),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1233),
.A2(n_1256),
.B(n_1216),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1233),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1255),
.B(n_1233),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1233),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1216),
.A2(n_1289),
.B(n_1204),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1221),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1232),
.B(n_1305),
.Y(n_1391)
);

NOR2xp33_ASAP7_75t_L g1392 ( 
.A(n_1335),
.B(n_1201),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1315),
.B(n_1291),
.Y(n_1393)
);

OAI21xp33_ASAP7_75t_SL g1394 ( 
.A1(n_1310),
.A2(n_1289),
.B(n_1204),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1319),
.B(n_1367),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1352),
.B(n_1219),
.Y(n_1396)
);

AND2x4_ASAP7_75t_L g1397 ( 
.A(n_1329),
.B(n_1231),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1341),
.B(n_1193),
.Y(n_1398)
);

OAI211xp5_ASAP7_75t_L g1399 ( 
.A1(n_1314),
.A2(n_1197),
.B(n_1245),
.C(n_1224),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1341),
.B(n_1203),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1373),
.B(n_1224),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1387),
.Y(n_1402)
);

NAND2xp5_ASAP7_75t_L g1403 ( 
.A(n_1368),
.B(n_1291),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1345),
.A2(n_1243),
.B(n_1250),
.C(n_1294),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1329),
.B(n_1295),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_SL g1406 ( 
.A(n_1331),
.B(n_1295),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1326),
.B(n_1293),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1339),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1345),
.B(n_1351),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_SL g1410 ( 
.A1(n_1389),
.A2(n_1343),
.B(n_1382),
.C(n_1323),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1317),
.A2(n_1344),
.B(n_1356),
.C(n_1337),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1350),
.Y(n_1412)
);

AOI211xp5_ASAP7_75t_L g1413 ( 
.A1(n_1358),
.A2(n_1334),
.B(n_1351),
.C(n_1349),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1358),
.A2(n_1349),
.B1(n_1321),
.B2(n_1362),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1338),
.B(n_1361),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1378),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1350),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1364),
.B(n_1365),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1378),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_SL g1420 ( 
.A1(n_1378),
.A2(n_1385),
.B(n_1379),
.Y(n_1420)
);

AO32x2_ASAP7_75t_L g1421 ( 
.A1(n_1333),
.A2(n_1347),
.A3(n_1362),
.B1(n_1316),
.B2(n_1337),
.Y(n_1421)
);

INVx4_ASAP7_75t_L g1422 ( 
.A(n_1378),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1340),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1316),
.B(n_1324),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1329),
.B(n_1359),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1359),
.B(n_1324),
.Y(n_1426)
);

NAND2xp33_ASAP7_75t_R g1427 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1354),
.Y(n_1428)
);

A2O1A1Ixp33_ASAP7_75t_L g1429 ( 
.A1(n_1321),
.A2(n_1371),
.B(n_1311),
.C(n_1375),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1347),
.A2(n_1362),
.B(n_1374),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1391),
.Y(n_1431)
);

O2A1O1Ixp33_ASAP7_75t_SL g1432 ( 
.A1(n_1390),
.A2(n_1376),
.B(n_1377),
.C(n_1379),
.Y(n_1432)
);

AOI221xp5_ASAP7_75t_L g1433 ( 
.A1(n_1337),
.A2(n_1360),
.B1(n_1357),
.B2(n_1354),
.C(n_1312),
.Y(n_1433)
);

OAI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1390),
.A2(n_1376),
.B1(n_1377),
.B2(n_1380),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1369),
.B(n_1383),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1309),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1369),
.B(n_1383),
.Y(n_1438)
);

AO21x1_ASAP7_75t_L g1439 ( 
.A1(n_1381),
.A2(n_1384),
.B(n_1386),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1369),
.B(n_1388),
.Y(n_1440)
);

AO32x2_ASAP7_75t_L g1441 ( 
.A1(n_1325),
.A2(n_1355),
.A3(n_1342),
.B1(n_1348),
.B2(n_1330),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1384),
.A2(n_1386),
.B1(n_1325),
.B2(n_1372),
.Y(n_1442)
);

OA21x2_ASAP7_75t_L g1443 ( 
.A1(n_1330),
.A2(n_1363),
.B(n_1366),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1437),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1412),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1417),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1422),
.B(n_1359),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1428),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1414),
.A2(n_1322),
.B1(n_1332),
.B2(n_1328),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1443),
.Y(n_1450)
);

OR2x2_ASAP7_75t_L g1451 ( 
.A(n_1423),
.B(n_1309),
.Y(n_1451)
);

NAND2xp5_ASAP7_75t_L g1452 ( 
.A(n_1395),
.B(n_1370),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1418),
.B(n_1312),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1408),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1439),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1426),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1424),
.B(n_1320),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1436),
.Y(n_1458)
);

NOR2x1_ASAP7_75t_L g1459 ( 
.A(n_1434),
.B(n_1318),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1435),
.Y(n_1460)
);

OR2x2_ASAP7_75t_L g1461 ( 
.A(n_1402),
.B(n_1320),
.Y(n_1461)
);

AND2x4_ASAP7_75t_L g1462 ( 
.A(n_1425),
.B(n_1346),
.Y(n_1462)
);

OAI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1406),
.A2(n_1375),
.B(n_1366),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1438),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1442),
.B(n_1327),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_R g1467 ( 
.A(n_1431),
.B(n_1353),
.Y(n_1467)
);

AND2x2_ASAP7_75t_SL g1468 ( 
.A(n_1419),
.B(n_1353),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1420),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1398),
.B(n_1355),
.Y(n_1470)
);

AND2x6_ASAP7_75t_L g1471 ( 
.A(n_1397),
.B(n_1336),
.Y(n_1471)
);

INVxp67_ASAP7_75t_L g1472 ( 
.A(n_1455),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1455),
.Y(n_1473)
);

NOR3xp33_ASAP7_75t_L g1474 ( 
.A(n_1459),
.B(n_1411),
.C(n_1399),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1450),
.Y(n_1475)
);

AND2x4_ASAP7_75t_L g1476 ( 
.A(n_1447),
.B(n_1416),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_1459),
.Y(n_1477)
);

BUFx3_ASAP7_75t_L g1478 ( 
.A(n_1471),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1444),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1460),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1444),
.Y(n_1481)
);

NAND4xp25_ASAP7_75t_L g1482 ( 
.A(n_1454),
.B(n_1413),
.C(n_1393),
.D(n_1403),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1449),
.A2(n_1409),
.B1(n_1414),
.B2(n_1433),
.Y(n_1483)
);

AOI211x1_ASAP7_75t_L g1484 ( 
.A1(n_1452),
.A2(n_1407),
.B(n_1401),
.C(n_1400),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1461),
.Y(n_1485)
);

AO21x2_ASAP7_75t_L g1486 ( 
.A1(n_1470),
.A2(n_1430),
.B(n_1429),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1464),
.B(n_1421),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1458),
.B(n_1413),
.Y(n_1488)
);

AND2x2_ASAP7_75t_SL g1489 ( 
.A(n_1468),
.B(n_1416),
.Y(n_1489)
);

NOR3xp33_ASAP7_75t_L g1490 ( 
.A(n_1469),
.B(n_1404),
.C(n_1394),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1445),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1458),
.B(n_1410),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1454),
.B(n_1432),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1466),
.B(n_1421),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1468),
.B(n_1441),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1463),
.A2(n_1394),
.B1(n_1313),
.B2(n_1405),
.Y(n_1496)
);

INVx4_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1468),
.B(n_1441),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1456),
.B(n_1441),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1477),
.B(n_1456),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1477),
.B(n_1469),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1475),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1479),
.Y(n_1503)
);

INVx4_ASAP7_75t_L g1504 ( 
.A(n_1489),
.Y(n_1504)
);

INVxp67_ASAP7_75t_SL g1505 ( 
.A(n_1472),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1478),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1479),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1479),
.Y(n_1508)
);

AND2x2_ASAP7_75t_SL g1509 ( 
.A(n_1489),
.B(n_1462),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1495),
.B(n_1457),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1497),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1481),
.Y(n_1512)
);

INVx1_ASAP7_75t_SL g1513 ( 
.A(n_1492),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1497),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1480),
.B(n_1451),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1480),
.B(n_1453),
.Y(n_1516)
);

AND2x4_ASAP7_75t_SL g1517 ( 
.A(n_1497),
.B(n_1462),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1472),
.B(n_1446),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1495),
.B(n_1447),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1481),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1498),
.B(n_1447),
.Y(n_1522)
);

INVx2_ASAP7_75t_SL g1523 ( 
.A(n_1478),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1475),
.Y(n_1524)
);

AND3x2_ASAP7_75t_L g1525 ( 
.A(n_1474),
.B(n_1396),
.C(n_1405),
.Y(n_1525)
);

NAND2x1p5_ASAP7_75t_L g1526 ( 
.A(n_1489),
.B(n_1497),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1498),
.B(n_1465),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1473),
.B(n_1448),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1475),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1498),
.B(n_1465),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1507),
.Y(n_1531)
);

AO22x1_ASAP7_75t_L g1532 ( 
.A1(n_1505),
.A2(n_1474),
.B1(n_1490),
.B2(n_1488),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1507),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1509),
.B(n_1489),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1502),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1502),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1503),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1503),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1509),
.B(n_1485),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1508),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1502),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1484),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1516),
.B(n_1492),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1509),
.B(n_1485),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1508),
.Y(n_1546)
);

INVxp67_ASAP7_75t_L g1547 ( 
.A(n_1513),
.Y(n_1547)
);

NOR2x1_ASAP7_75t_L g1548 ( 
.A(n_1504),
.B(n_1497),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1505),
.B(n_1484),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1508),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1512),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1509),
.B(n_1478),
.Y(n_1552)
);

HB1xp67_ASAP7_75t_L g1553 ( 
.A(n_1518),
.Y(n_1553)
);

BUFx2_ASAP7_75t_L g1554 ( 
.A(n_1504),
.Y(n_1554)
);

NAND2xp33_ASAP7_75t_L g1555 ( 
.A(n_1526),
.B(n_1490),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1512),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1527),
.B(n_1530),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1516),
.B(n_1491),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1517),
.B(n_1478),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1504),
.B(n_1496),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1512),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1527),
.B(n_1493),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1502),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1524),
.Y(n_1565)
);

OR2x2_ASAP7_75t_L g1566 ( 
.A(n_1516),
.B(n_1491),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1517),
.B(n_1476),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1521),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1515),
.B(n_1491),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1530),
.B(n_1488),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1521),
.Y(n_1571)
);

INVx2_ASAP7_75t_SL g1572 ( 
.A(n_1517),
.Y(n_1572)
);

NAND2x1p5_ASAP7_75t_L g1573 ( 
.A(n_1548),
.B(n_1504),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1534),
.B(n_1517),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1531),
.Y(n_1575)
);

INVx3_ASAP7_75t_L g1576 ( 
.A(n_1534),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1552),
.B(n_1530),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1531),
.Y(n_1578)
);

OAI22xp33_ASAP7_75t_L g1579 ( 
.A1(n_1549),
.A2(n_1482),
.B1(n_1504),
.B2(n_1427),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1532),
.Y(n_1580)
);

INVx1_ASAP7_75t_SL g1581 ( 
.A(n_1532),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1552),
.B(n_1506),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1558),
.B(n_1518),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1553),
.B(n_1520),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1547),
.B(n_1520),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1533),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1548),
.B(n_1506),
.Y(n_1587)
);

INVx6_ASAP7_75t_L g1588 ( 
.A(n_1560),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1533),
.Y(n_1589)
);

HB1xp67_ASAP7_75t_L g1590 ( 
.A(n_1537),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1540),
.B(n_1526),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1535),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1535),
.Y(n_1593)
);

NAND3xp33_ASAP7_75t_L g1594 ( 
.A(n_1543),
.B(n_1525),
.C(n_1482),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1537),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1572),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1570),
.B(n_1544),
.Y(n_1597)
);

NOR3xp33_ASAP7_75t_L g1598 ( 
.A(n_1555),
.B(n_1528),
.C(n_1501),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1538),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1544),
.B(n_1556),
.Y(n_1600)
);

INVx2_ASAP7_75t_SL g1601 ( 
.A(n_1572),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1563),
.B(n_1528),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1538),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1560),
.B(n_1506),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1567),
.B(n_1523),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1567),
.B(n_1523),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1540),
.B(n_1523),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1580),
.A2(n_1561),
.B1(n_1483),
.B2(n_1486),
.Y(n_1608)
);

OAI21xp5_ASAP7_75t_SL g1609 ( 
.A1(n_1580),
.A2(n_1525),
.B(n_1554),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1590),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1590),
.Y(n_1611)
);

AOI32xp33_ASAP7_75t_L g1612 ( 
.A1(n_1581),
.A2(n_1545),
.A3(n_1554),
.B1(n_1499),
.B2(n_1500),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1599),
.Y(n_1613)
);

INVxp67_ASAP7_75t_L g1614 ( 
.A(n_1581),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1597),
.B(n_1510),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1604),
.B(n_1545),
.Y(n_1616)
);

INVx1_ASAP7_75t_SL g1617 ( 
.A(n_1588),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1604),
.B(n_1519),
.Y(n_1618)
);

INVxp67_ASAP7_75t_L g1619 ( 
.A(n_1596),
.Y(n_1619)
);

NAND2x1_ASAP7_75t_L g1620 ( 
.A(n_1588),
.B(n_1500),
.Y(n_1620)
);

AOI31xp33_ASAP7_75t_L g1621 ( 
.A1(n_1573),
.A2(n_1526),
.A3(n_1392),
.B(n_1500),
.Y(n_1621)
);

OAI22xp5_ASAP7_75t_L g1622 ( 
.A1(n_1594),
.A2(n_1579),
.B1(n_1588),
.B2(n_1598),
.Y(n_1622)
);

OAI21xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1587),
.A2(n_1522),
.B(n_1519),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1594),
.A2(n_1526),
.B1(n_1483),
.B2(n_1514),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1597),
.B(n_1510),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1599),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1595),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1579),
.A2(n_1486),
.B1(n_1494),
.B2(n_1487),
.Y(n_1628)
);

AOI21xp33_ASAP7_75t_L g1629 ( 
.A1(n_1576),
.A2(n_1535),
.B(n_1536),
.Y(n_1629)
);

AOI22xp33_ASAP7_75t_SL g1630 ( 
.A1(n_1576),
.A2(n_1499),
.B1(n_1486),
.B2(n_1526),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1595),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1603),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1608),
.A2(n_1598),
.B1(n_1576),
.B2(n_1577),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1630),
.A2(n_1588),
.B1(n_1576),
.B2(n_1573),
.Y(n_1634)
);

INVxp67_ASAP7_75t_SL g1635 ( 
.A(n_1614),
.Y(n_1635)
);

CKINVDCx14_ASAP7_75t_R g1636 ( 
.A(n_1622),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1627),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1631),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1614),
.B(n_1600),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1630),
.A2(n_1585),
.B1(n_1573),
.B2(n_1600),
.C(n_1584),
.Y(n_1640)
);

OAI21xp5_ASAP7_75t_L g1641 ( 
.A1(n_1609),
.A2(n_1573),
.B(n_1587),
.Y(n_1641)
);

OAI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1612),
.A2(n_1582),
.B(n_1607),
.Y(n_1642)
);

AOI221xp5_ASAP7_75t_L g1643 ( 
.A1(n_1628),
.A2(n_1585),
.B1(n_1584),
.B2(n_1586),
.C(n_1589),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1632),
.Y(n_1644)
);

INVx1_ASAP7_75t_SL g1645 ( 
.A(n_1617),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1610),
.Y(n_1646)
);

AOI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1624),
.A2(n_1577),
.B1(n_1588),
.B2(n_1607),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1611),
.Y(n_1648)
);

OAI32xp33_ASAP7_75t_L g1649 ( 
.A1(n_1623),
.A2(n_1591),
.A3(n_1602),
.B1(n_1587),
.B2(n_1583),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1619),
.B(n_1616),
.Y(n_1650)
);

OAI22xp5_ASAP7_75t_L g1651 ( 
.A1(n_1621),
.A2(n_1574),
.B1(n_1596),
.B2(n_1601),
.Y(n_1651)
);

INVx1_ASAP7_75t_SL g1652 ( 
.A(n_1645),
.Y(n_1652)
);

XOR2x2_ASAP7_75t_L g1653 ( 
.A(n_1640),
.B(n_1620),
.Y(n_1653)
);

OAI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1640),
.A2(n_1619),
.B(n_1629),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1635),
.B(n_1613),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1650),
.B(n_1626),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1636),
.B(n_1596),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1637),
.Y(n_1658)
);

AOI21xp5_ASAP7_75t_L g1659 ( 
.A1(n_1649),
.A2(n_1601),
.B(n_1615),
.Y(n_1659)
);

XOR2x2_ASAP7_75t_L g1660 ( 
.A(n_1633),
.B(n_1625),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1651),
.B(n_1601),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1638),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1643),
.A2(n_1582),
.B1(n_1592),
.B2(n_1593),
.Y(n_1663)
);

NAND3xp33_ASAP7_75t_L g1664 ( 
.A(n_1654),
.B(n_1634),
.C(n_1639),
.Y(n_1664)
);

NAND4xp75_ASAP7_75t_L g1665 ( 
.A(n_1657),
.B(n_1641),
.C(n_1647),
.D(n_1646),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1652),
.B(n_1642),
.Y(n_1666)
);

INVx2_ASAP7_75t_SL g1667 ( 
.A(n_1652),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1661),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1663),
.A2(n_1644),
.B1(n_1648),
.B2(n_1592),
.C(n_1593),
.Y(n_1669)
);

OAI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1659),
.A2(n_1575),
.B(n_1578),
.C(n_1586),
.Y(n_1670)
);

NOR3xp33_ASAP7_75t_L g1671 ( 
.A(n_1655),
.B(n_1593),
.C(n_1592),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1658),
.B(n_1618),
.Y(n_1672)
);

NAND3xp33_ASAP7_75t_SL g1673 ( 
.A(n_1656),
.B(n_1662),
.C(n_1653),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1660),
.Y(n_1674)
);

AOI222xp33_ASAP7_75t_L g1675 ( 
.A1(n_1674),
.A2(n_1575),
.B1(n_1578),
.B2(n_1589),
.C1(n_1603),
.C2(n_1542),
.Y(n_1675)
);

OAI211xp5_ASAP7_75t_SL g1676 ( 
.A1(n_1664),
.A2(n_1602),
.B(n_1583),
.C(n_1511),
.Y(n_1676)
);

AOI221xp5_ASAP7_75t_L g1677 ( 
.A1(n_1673),
.A2(n_1542),
.B1(n_1565),
.B2(n_1536),
.C(n_1564),
.Y(n_1677)
);

A2O1A1Ixp33_ASAP7_75t_L g1678 ( 
.A1(n_1669),
.A2(n_1574),
.B(n_1536),
.C(n_1542),
.Y(n_1678)
);

OAI211xp5_ASAP7_75t_L g1679 ( 
.A1(n_1668),
.A2(n_1606),
.B(n_1605),
.C(n_1511),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1675),
.Y(n_1680)
);

AO21x1_ASAP7_75t_L g1681 ( 
.A1(n_1676),
.A2(n_1666),
.B(n_1671),
.Y(n_1681)
);

AOI22xp5_ASAP7_75t_L g1682 ( 
.A1(n_1677),
.A2(n_1667),
.B1(n_1665),
.B2(n_1670),
.Y(n_1682)
);

NAND3xp33_ASAP7_75t_L g1683 ( 
.A(n_1679),
.B(n_1672),
.C(n_1606),
.Y(n_1683)
);

AOI221xp5_ASAP7_75t_L g1684 ( 
.A1(n_1678),
.A2(n_1565),
.B1(n_1564),
.B2(n_1539),
.C(n_1568),
.Y(n_1684)
);

OAI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1677),
.A2(n_1565),
.B1(n_1605),
.B2(n_1511),
.C(n_1514),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1681),
.Y(n_1686)
);

XNOR2xp5_ASAP7_75t_L g1687 ( 
.A(n_1682),
.B(n_1501),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1683),
.B(n_1519),
.Y(n_1688)
);

OAI22x1_ASAP7_75t_L g1689 ( 
.A1(n_1680),
.A2(n_1571),
.B1(n_1539),
.B2(n_1568),
.Y(n_1689)
);

NOR2xp67_ASAP7_75t_L g1690 ( 
.A(n_1685),
.B(n_1559),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1689),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1686),
.A2(n_1684),
.B(n_1571),
.Y(n_1692)
);

AOI322xp5_ASAP7_75t_L g1693 ( 
.A1(n_1688),
.A2(n_1689),
.A3(n_1687),
.B1(n_1690),
.B2(n_1499),
.C1(n_1487),
.C2(n_1494),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1693),
.B(n_1501),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1694),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_SL g1696 ( 
.A1(n_1695),
.A2(n_1691),
.B1(n_1692),
.B2(n_1546),
.Y(n_1696)
);

INVx1_ASAP7_75t_SL g1697 ( 
.A(n_1695),
.Y(n_1697)
);

OAI22xp5_ASAP7_75t_SL g1698 ( 
.A1(n_1697),
.A2(n_1550),
.B1(n_1541),
.B2(n_1562),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1696),
.A2(n_1541),
.B1(n_1546),
.B2(n_1562),
.Y(n_1699)
);

OAI22xp5_ASAP7_75t_L g1700 ( 
.A1(n_1699),
.A2(n_1566),
.B1(n_1559),
.B2(n_1569),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1698),
.A2(n_1557),
.B(n_1551),
.Y(n_1701)
);

AOI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1700),
.A2(n_1701),
.B1(n_1550),
.B2(n_1557),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1702),
.A2(n_1551),
.B(n_1566),
.Y(n_1703)
);

OAI21xp5_ASAP7_75t_L g1704 ( 
.A1(n_1703),
.A2(n_1529),
.B(n_1524),
.Y(n_1704)
);

OAI221xp5_ASAP7_75t_R g1705 ( 
.A1(n_1704),
.A2(n_1467),
.B1(n_1569),
.B2(n_1511),
.C(n_1514),
.Y(n_1705)
);

AOI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1705),
.A2(n_1415),
.B(n_1511),
.C(n_1514),
.Y(n_1706)
);


endmodule