module fake_jpeg_24380_n_318 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx8_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_19),
.B(n_0),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_20),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_20),
.Y(n_55)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g42 ( 
.A1(n_35),
.A2(n_14),
.B1(n_25),
.B2(n_26),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_53),
.B1(n_35),
.B2(n_34),
.Y(n_69)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_50),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_29),
.Y(n_49)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_33),
.B(n_22),
.Y(n_52)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_52),
.B(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_35),
.A2(n_23),
.B1(n_22),
.B2(n_26),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_55),
.B(n_31),
.Y(n_66)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_35),
.B(n_14),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_56),
.B(n_36),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_SL g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_59),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_49),
.A2(n_34),
.B1(n_26),
.B2(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_77),
.B1(n_69),
.B2(n_59),
.Y(n_80)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_69),
.B1(n_72),
.B2(n_44),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_32),
.Y(n_62)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_66),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_52),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_35),
.B1(n_34),
.B2(n_17),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_29),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_74),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_45),
.B(n_31),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_75),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_32),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_68),
.Y(n_79)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_62),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_82),
.A2(n_98),
.B1(n_99),
.B2(n_72),
.Y(n_113)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_64),
.A2(n_40),
.B1(n_44),
.B2(n_51),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_91),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_57),
.Y(n_89)
);

INVx13_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_93),
.B(n_95),
.Y(n_118)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_68),
.Y(n_95)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_74),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_47),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_59),
.A2(n_56),
.B1(n_36),
.B2(n_47),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_64),
.A2(n_51),
.B1(n_47),
.B2(n_27),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_94),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_105),
.Y(n_131)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_89),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_104),
.Y(n_146)
);

NAND2x1_ASAP7_75t_SL g103 ( 
.A(n_98),
.B(n_58),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_103),
.A2(n_115),
.B(n_77),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_100),
.B(n_65),
.Y(n_105)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_110),
.Y(n_142)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_112),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_113),
.A2(n_65),
.B1(n_62),
.B2(n_70),
.Y(n_136)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_79),
.Y(n_114)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_114),
.Y(n_139)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_83),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_116),
.Y(n_138)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_84),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_120),
.Y(n_127)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_119),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_87),
.B(n_66),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_93),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_123),
.Y(n_132)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_96),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

INVx13_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_91),
.B1(n_92),
.B2(n_78),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_126),
.B1(n_136),
.B2(n_141),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_78),
.B1(n_92),
.B2(n_94),
.Y(n_126)
);

OAI21xp33_ASAP7_75t_SL g173 ( 
.A1(n_129),
.A2(n_36),
.B(n_30),
.Y(n_173)
);

AO22x1_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_98),
.B1(n_80),
.B2(n_58),
.Y(n_130)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_130),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_73),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_101),
.B(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_135),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_77),
.C(n_70),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_137),
.B(n_36),
.C(n_63),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_115),
.A2(n_58),
.B1(n_39),
.B2(n_54),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_121),
.A2(n_103),
.B1(n_115),
.B2(n_117),
.Y(n_144)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_144),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_118),
.B(n_45),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_58),
.Y(n_147)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_103),
.A2(n_61),
.B1(n_76),
.B2(n_88),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_148),
.A2(n_61),
.B1(n_76),
.B2(n_106),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_110),
.Y(n_151)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_108),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_163),
.C(n_137),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_106),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_158),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_142),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_160),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_114),
.Y(n_157)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_157),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_143),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_31),
.B(n_16),
.C(n_24),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_159),
.B(n_27),
.Y(n_189)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_124),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_162),
.B(n_171),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_146),
.B(n_112),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_128),
.Y(n_181)
);

HAxp5_ASAP7_75t_SL g167 ( 
.A(n_147),
.B(n_48),
.CON(n_167),
.SN(n_167)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_167),
.A2(n_172),
.B(n_145),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_95),
.B1(n_139),
.B2(n_138),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_128),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_170),
.Y(n_185)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_146),
.Y(n_171)
);

OAI21xp33_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_13),
.B(n_12),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_173),
.A2(n_141),
.B1(n_61),
.B2(n_76),
.Y(n_199)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_174),
.B(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_135),
.Y(n_175)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_144),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_196),
.Y(n_204)
);

OAI22x1_ASAP7_75t_L g179 ( 
.A1(n_150),
.A2(n_130),
.B1(n_148),
.B2(n_126),
.Y(n_179)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_195),
.B1(n_174),
.B2(n_159),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_180),
.B(n_189),
.Y(n_219)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_181),
.Y(n_222)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_188),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_190),
.B(n_194),
.C(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_193),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_199),
.B1(n_201),
.B2(n_200),
.Y(n_210)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_149),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_136),
.C(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_165),
.A2(n_127),
.B(n_134),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_116),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_150),
.A2(n_133),
.B1(n_138),
.B2(n_43),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_200),
.A2(n_171),
.B1(n_168),
.B2(n_170),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g201 ( 
.A1(n_165),
.A2(n_133),
.B(n_48),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_218),
.C(n_199),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_168),
.C(n_175),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_214),
.C(n_221),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_156),
.Y(n_208)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_216),
.B(n_220),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_210),
.A2(n_213),
.B1(n_182),
.B2(n_183),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_184),
.B1(n_191),
.B2(n_193),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_153),
.C(n_164),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_215),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_160),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_158),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_153),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_194),
.B(n_164),
.C(n_161),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_149),
.C(n_143),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_223),
.B(n_187),
.C(n_182),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_205),
.B(n_201),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_234),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_226),
.B(n_229),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g230 ( 
.A(n_204),
.B(n_179),
.Y(n_230)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_230),
.A2(n_231),
.B(n_240),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_186),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_242),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_219),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_196),
.C(n_143),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_213),
.A2(n_102),
.B1(n_50),
.B2(n_74),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_236),
.A2(n_209),
.B1(n_211),
.B2(n_206),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_71),
.C(n_17),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_239),
.B(n_241),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_214),
.B(n_21),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_223),
.B(n_71),
.C(n_24),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_71),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_202),
.A2(n_71),
.B(n_109),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_243),
.B(n_244),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_222),
.B(n_71),
.C(n_38),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_236),
.Y(n_247)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_247),
.Y(n_269)
);

A2O1A1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_231),
.A2(n_220),
.B(n_203),
.C(n_202),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_257),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_262),
.B1(n_38),
.B2(n_30),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_225),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_251),
.B(n_259),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_238),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_255),
.Y(n_273)
);

BUFx12_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_235),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_256),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_206),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_18),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_260),
.B(n_18),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_229),
.A2(n_81),
.B1(n_38),
.B2(n_30),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_249),
.B(n_228),
.C(n_234),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_266),
.C(n_271),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_262),
.B(n_228),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_264),
.B(n_265),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_258),
.A2(n_246),
.B(n_251),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_240),
.C(n_230),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_270),
.B1(n_38),
.B2(n_30),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_250),
.A2(n_21),
.B1(n_28),
.B2(n_15),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_81),
.C(n_11),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_255),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_274),
.B(n_13),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_81),
.C(n_38),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_276),
.B(n_257),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_0),
.Y(n_290)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_278),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_266),
.B(n_248),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_281),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_272),
.B(n_254),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_13),
.Y(n_282)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_282),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_276),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_12),
.C(n_11),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_288),
.B(n_289),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_11),
.B1(n_21),
.B2(n_15),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_290),
.C(n_285),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_28),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_274),
.B(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_291),
.B(n_292),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_280),
.B(n_268),
.C(n_28),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_268),
.C(n_15),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_294),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_1),
.B(n_2),
.Y(n_298)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_298),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.C1(n_5),
.C2(n_6),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_295),
.A2(n_284),
.B1(n_2),
.B2(n_3),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_304),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_18),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g305 ( 
.A(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_306),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_297),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_306)
);

AOI31xp33_ASAP7_75t_L g311 ( 
.A1(n_307),
.A2(n_296),
.A3(n_291),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_302),
.B(n_299),
.Y(n_308)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_311),
.A3(n_301),
.B1(n_293),
.B2(n_305),
.C1(n_7),
.C2(n_1),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_309),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_5),
.B(n_6),
.Y(n_313)
);

NAND2xp33_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_9),
.Y(n_315)
);

NAND4xp25_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_5),
.C(n_6),
.D(n_7),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_7),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_8),
.Y(n_318)
);


endmodule