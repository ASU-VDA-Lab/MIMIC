module real_jpeg_12986_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_249;
wire n_286;
wire n_292;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_244;
wire n_128;
wire n_202;
wire n_179;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

BUFx2_ASAP7_75t_L g75 ( 
.A(n_0),
.Y(n_75)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_3),
.A2(n_63),
.B1(n_66),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_3),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_3),
.A2(n_49),
.B1(n_51),
.B2(n_78),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_78),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_78),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_4),
.A2(n_25),
.B1(n_29),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_4),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_4),
.A2(n_40),
.B1(n_49),
.B2(n_51),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_4),
.A2(n_40),
.B1(n_63),
.B2(n_66),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_5),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_5),
.A2(n_29),
.B(n_32),
.C(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_5),
.B(n_38),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_5),
.A2(n_28),
.B1(n_49),
.B2(n_51),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_5),
.A2(n_87),
.B1(n_116),
.B2(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_53),
.Y(n_188)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_35),
.B1(n_36),
.B2(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_25),
.B1(n_29),
.B2(n_44),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_10),
.A2(n_44),
.B1(n_49),
.B2(n_51),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_10),
.A2(n_44),
.B1(n_63),
.B2(n_66),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_11),
.A2(n_63),
.B1(n_66),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_11),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_49),
.B1(n_51),
.B2(n_80),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_80),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_12),
.A2(n_49),
.B1(n_51),
.B2(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_12),
.A2(n_63),
.B1(n_66),
.B2(n_71),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_12),
.A2(n_35),
.B1(n_36),
.B2(n_71),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_12),
.A2(n_25),
.B1(n_29),
.B2(n_71),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_13),
.A2(n_49),
.B1(n_51),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_68),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_13),
.A2(n_63),
.B1(n_66),
.B2(n_68),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_68),
.Y(n_246)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_15),
.A2(n_35),
.B1(n_36),
.B2(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_15),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_49),
.B1(n_51),
.B2(n_55),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_15),
.A2(n_55),
.B1(n_63),
.B2(n_66),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_15),
.A2(n_25),
.B1(n_29),
.B2(n_55),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_273),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_251),
.B(n_272),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_224),
.B(n_250),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_125),
.B(n_203),
.C(n_223),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_98),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_21),
.B(n_98),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_72),
.C(n_85),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_22),
.B(n_200),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_41),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_42),
.C(n_56),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_38),
.B2(n_39),
.Y(n_23)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g82 ( 
.A1(n_28),
.A2(n_33),
.B(n_35),
.Y(n_82)
);

HAxp5_ASAP7_75t_SL g135 ( 
.A(n_28),
.B(n_36),
.CON(n_135),
.SN(n_135)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_28),
.B(n_60),
.C(n_66),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_28),
.B(n_87),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_28),
.B(n_62),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_30),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_30),
.A2(n_38),
.B1(n_107),
.B2(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_30),
.B(n_269),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_34),
.A2(n_104),
.B1(n_105),
.B2(n_106),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g287 ( 
.A1(n_34),
.A2(n_288),
.B(n_289),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_35),
.A2(n_36),
.B1(n_47),
.B2(n_48),
.Y(n_52)
);

NOR3xp33_ASAP7_75t_L g136 ( 
.A(n_35),
.B(n_48),
.C(n_49),
.Y(n_136)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_38),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_38),
.B(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_39),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_56),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_53),
.B2(n_54),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_45),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_45),
.A2(n_53),
.B1(n_95),
.B2(n_135),
.Y(n_150)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_45),
.A2(n_111),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_45),
.B(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_45),
.A2(n_53),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_52),
.Y(n_45)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_94),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_46),
.B(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_46),
.A2(n_240),
.B(n_241),
.Y(n_239)
);

OA22x2_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_46)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_47),
.A2(n_51),
.B(n_134),
.C(n_136),
.Y(n_133)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_49),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_51),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_51),
.B(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_53),
.B(n_111),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g109 ( 
.A(n_54),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_67),
.B(n_69),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_57),
.B(n_123),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_57),
.A2(n_142),
.B1(n_144),
.B2(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_57),
.A2(n_144),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_57),
.A2(n_144),
.B1(n_152),
.B2(n_162),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_57),
.A2(n_144),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_57),
.A2(n_69),
.B(n_212),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_57),
.A2(n_67),
.B(n_144),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_60),
.B1(n_63),
.B2(n_66),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_SL g59 ( 
.A(n_60),
.Y(n_59)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_121),
.B(n_122),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

CKINVDCx6p67_ASAP7_75t_R g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_66),
.B(n_75),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_66),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_67),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_72),
.B(n_85),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_72)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_76),
.B2(n_79),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_74),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_74),
.A2(n_119),
.B(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_75),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_75),
.B(n_138),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_79),
.Y(n_117)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_83),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_91),
.C(n_93),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_86),
.A2(n_91),
.B1(n_92),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_86),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_90),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_87),
.A2(n_116),
.B1(n_167),
.B2(n_175),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_87),
.A2(n_116),
.B(n_231),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_88),
.B(n_185),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_93),
.B(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g282 ( 
.A1(n_96),
.A2(n_283),
.B(n_284),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_113),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_99),
.B(n_114),
.C(n_124),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_102),
.B2(n_112),
.Y(n_99)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_108),
.C(n_112),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_104),
.A2(n_244),
.B(n_245),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_104),
.A2(n_267),
.B(n_268),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_124),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_120),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_115),
.B(n_120),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_116),
.A2(n_169),
.B(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_121),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_122),
.B(n_143),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_198),
.B(n_202),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_153),
.B(n_197),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_148),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_130),
.B(n_148),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_145),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_139),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_132),
.B(n_139),
.C(n_145),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_133),
.B(n_137),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_138),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_141),
.B(n_143),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_150),
.C(n_151),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_149),
.B(n_194),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_151),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_154),
.A2(n_192),
.B(n_196),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_181),
.B(n_191),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_170),
.B(n_180),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_157),
.B(n_165),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_157)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_158),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_163),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_176),
.B(n_179),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_183),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_183),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_184),
.B(n_187),
.C(n_190),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_189),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_195),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_193),
.B(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_199),
.B(n_201),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_204),
.B(n_222),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_207),
.C(n_214),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_210),
.B2(n_213),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_208),
.B(n_213),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_210),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_215),
.B(n_217),
.C(n_220),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_220),
.Y(n_216)
);

INVxp33_ASAP7_75t_L g284 ( 
.A(n_218),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_219),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_225),
.B(n_226),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_249),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_234),
.B1(n_247),
.B2(n_248),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_248),
.C(n_249),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_233),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_229),
.A2(n_230),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_232),
.Y(n_263)
);

AOI21xp33_ASAP7_75t_L g277 ( 
.A1(n_230),
.A2(n_263),
.B(n_265),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_239),
.C(n_243),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_243),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_271),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_271),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_255),
.B2(n_270),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_256),
.C(n_262),
.Y(n_275)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_255),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_262),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_260),
.B(n_261),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_257),
.B(n_260),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_259),
.Y(n_283)
);

FAx1_ASAP7_75t_SL g276 ( 
.A(n_261),
.B(n_277),
.CI(n_278),
.CON(n_276),
.SN(n_276)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_291),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_275),
.B(n_276),
.Y(n_292)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_276),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_287),
.B2(n_290),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_282),
.B1(n_285),
.B2(n_286),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_287),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);


endmodule