module fake_jpeg_11151_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx5_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_8),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_9),
.Y(n_71)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_51),
.B(n_0),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_62),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_87),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_82),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g100 ( 
.A(n_88),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_71),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_91),
.B(n_96),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_SL g93 ( 
.A(n_82),
.Y(n_93)
);

INVx13_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_70),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_6),
.Y(n_117)
);

INVx13_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

INVx13_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_85),
.A2(n_67),
.B(n_69),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_99),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_89),
.A2(n_60),
.B1(n_56),
.B2(n_69),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_104),
.B1(n_105),
.B2(n_110),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_55),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_103),
.B(n_111),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_56),
.B1(n_68),
.B2(n_66),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_83),
.A2(n_61),
.B1(n_53),
.B2(n_58),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_63),
.B1(n_72),
.B2(n_67),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_109),
.B1(n_113),
.B2(n_88),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_72),
.B1(n_65),
.B2(n_50),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_29),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_94),
.A2(n_65),
.B1(n_2),
.B2(n_3),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_1),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_4),
.B(n_5),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_112),
.A2(n_102),
.B(n_109),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_90),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_115),
.Y(n_123)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_118),
.Y(n_139)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_120),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_121),
.A2(n_125),
.B(n_131),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_124),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_110),
.B(n_7),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_99),
.B(n_90),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_10),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_132),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_25),
.B1(n_27),
.B2(n_33),
.Y(n_150)
);

AO22x1_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_98),
.B1(n_30),
.B2(n_32),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_10),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_133),
.B(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_11),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_137),
.B(n_34),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_12),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_15),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_13),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_14),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_147),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_119),
.B(n_48),
.C(n_21),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_38),
.C(n_40),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_128),
.A2(n_119),
.B1(n_130),
.B2(n_131),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_146),
.A2(n_149),
.B1(n_150),
.B2(n_47),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_122),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_130),
.A2(n_17),
.B1(n_22),
.B2(n_23),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_152),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_37),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_154),
.Y(n_164)
);

OAI21xp33_ASAP7_75t_SL g156 ( 
.A1(n_139),
.A2(n_128),
.B(n_129),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_158),
.B1(n_162),
.B2(n_151),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_161),
.C(n_149),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_41),
.C(n_43),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_163),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_160),
.B(n_145),
.C(n_142),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_165),
.A2(n_166),
.B1(n_155),
.B2(n_157),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_160),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_169),
.B(n_167),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_153),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_141),
.C(n_143),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_172),
.A2(n_140),
.B(n_164),
.Y(n_173)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_173),
.Y(n_174)
);


endmodule