module fake_jpeg_20111_n_146 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_3),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_10),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_43),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_1),
.B(n_14),
.Y(n_57)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_32),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_21),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_15),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_5),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_4),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_75),
.B(n_49),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_77),
.B(n_64),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_78),
.Y(n_86)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_79),
.A2(n_56),
.B1(n_51),
.B2(n_47),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g87 ( 
.A(n_80),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_78),
.Y(n_82)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_79),
.A2(n_46),
.B1(n_58),
.B2(n_59),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_83),
.A2(n_91),
.B1(n_66),
.B2(n_64),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_88),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_53),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_47),
.B1(n_71),
.B2(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_81),
.B(n_70),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_95),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_2),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_69),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_99),
.B(n_2),
.Y(n_119)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_101),
.Y(n_106)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_66),
.B1(n_72),
.B2(n_67),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_84),
.A2(n_61),
.B(n_63),
.C(n_65),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_103),
.B(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_104),
.B(n_86),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_116),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_97),
.B(n_65),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_108),
.B(n_6),
.C(n_7),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_102),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_109),
.B(n_114),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_110),
.A2(n_72),
.B1(n_68),
.B2(n_7),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_113),
.B(n_105),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_96),
.B(n_60),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_96),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_117),
.Y(n_129)
);

BUFx8_ASAP7_75t_L g116 ( 
.A(n_103),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_96),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_118),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_119),
.B(n_22),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_120),
.A2(n_123),
.B1(n_109),
.B2(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_44),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_3),
.B(n_6),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_126),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_131),
.B(n_132),
.Y(n_135)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_128),
.A2(n_116),
.A3(n_117),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_16),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_8),
.B1(n_9),
.B2(n_17),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_136),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_123),
.C(n_129),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_134),
.C(n_135),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_139),
.B(n_130),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_24),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_27),
.C(n_29),
.Y(n_144)
);

OAI221xp5_ASAP7_75t_L g145 ( 
.A1(n_144),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.C(n_38),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_42),
.Y(n_146)
);


endmodule