module fake_jpeg_29194_n_547 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_547);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_547;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

CKINVDCx14_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_9),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_4),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

BUFx12_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_14),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_22),
.B(n_54),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_55),
.B(n_101),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_56),
.Y(n_128)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_58),
.Y(n_145)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_60),
.Y(n_143)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_61),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_62),
.Y(n_148)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_35),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_63),
.B(n_65),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_64),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_7),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_35),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_66),
.B(n_72),
.Y(n_154)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_67),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g140 ( 
.A(n_68),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_69),
.Y(n_166)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_71),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_16),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_26),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_77),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_23),
.Y(n_79)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_33),
.A2(n_15),
.B1(n_5),
.B2(n_2),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_80),
.A2(n_53),
.B1(n_50),
.B2(n_28),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx5_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_83),
.Y(n_178)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_86),
.Y(n_160)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_51),
.B(n_8),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_88),
.B(n_48),
.Y(n_174)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_91),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_25),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_92),
.B(n_97),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_93),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_17),
.Y(n_94)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_94),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_96),
.Y(n_127)
);

INVx6_ASAP7_75t_SL g97 ( 
.A(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_49),
.Y(n_99)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_18),
.Y(n_100)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_22),
.B(n_8),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_40),
.Y(n_102)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_102),
.Y(n_150)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_103),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_40),
.Y(n_104)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_104),
.Y(n_155)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_42),
.Y(n_105)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_106),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_107),
.Y(n_113)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_25),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_52),
.Y(n_175)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_16),
.Y(n_109)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_49),
.Y(n_111)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_65),
.B(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_121),
.B(n_130),
.Y(n_208)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_88),
.A2(n_48),
.B(n_39),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_122),
.B(n_129),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_84),
.A2(n_32),
.B1(n_18),
.B2(n_30),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_125),
.A2(n_126),
.B1(n_139),
.B2(n_147),
.Y(n_181)
);

OAI22xp33_ASAP7_75t_L g126 ( 
.A1(n_64),
.A2(n_32),
.B1(n_18),
.B2(n_36),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g129 ( 
.A(n_80),
.B(n_25),
.CON(n_129),
.SN(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_94),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_137),
.A2(n_10),
.B(n_15),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_69),
.A2(n_53),
.B1(n_50),
.B2(n_46),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_92),
.B(n_41),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_142),
.B(n_173),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_71),
.A2(n_28),
.B1(n_46),
.B2(n_43),
.Y(n_147)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_162),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_63),
.B(n_43),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_169),
.B(n_176),
.Y(n_197)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_61),
.Y(n_171)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_92),
.B(n_37),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_39),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_66),
.B(n_37),
.Y(n_176)
);

INVx5_ASAP7_75t_L g179 ( 
.A(n_178),
.Y(n_179)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_124),
.B(n_38),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_180),
.B(n_189),
.Y(n_248)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_165),
.Y(n_182)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_182),
.Y(n_256)
);

INVx8_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_183),
.Y(n_270)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_157),
.Y(n_184)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_184),
.Y(n_258)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_140),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_128),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_186),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_34),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_209),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_188),
.B(n_192),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_117),
.B(n_38),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_119),
.Y(n_190)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_190),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_174),
.A2(n_34),
.B1(n_41),
.B2(n_111),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_193),
.B(n_195),
.Y(n_262)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_161),
.Y(n_194)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_120),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_128),
.Y(n_196)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_131),
.A2(n_27),
.B(n_21),
.Y(n_198)
);

A2O1A1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_198),
.A2(n_126),
.B(n_164),
.C(n_52),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_129),
.A2(n_32),
.B1(n_70),
.B2(n_75),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_199),
.A2(n_216),
.B1(n_225),
.B2(n_116),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_114),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_192),
.Y(n_236)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_202),
.Y(n_265)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_205),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_125),
.A2(n_77),
.B1(n_73),
.B2(n_81),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_206),
.A2(n_223),
.B1(n_159),
.B2(n_143),
.Y(n_254)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_133),
.Y(n_207)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_207),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_163),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_136),
.A2(n_85),
.B1(n_93),
.B2(n_104),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_210),
.A2(n_166),
.B1(n_106),
.B2(n_143),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g211 ( 
.A(n_140),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_115),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_134),
.Y(n_214)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_214),
.Y(n_274)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_113),
.Y(n_215)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_215),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_32),
.B1(n_79),
.B2(n_36),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_154),
.B(n_21),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_217),
.B(n_224),
.Y(n_250)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_218),
.Y(n_269)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_219),
.Y(n_272)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_123),
.Y(n_220)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_220),
.Y(n_273)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_226),
.Y(n_247)
);

BUFx12f_ASAP7_75t_L g222 ( 
.A(n_132),
.Y(n_222)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_222),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_136),
.A2(n_102),
.B1(n_95),
.B2(n_62),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_175),
.B(n_27),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_151),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_83),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_229),
.B1(n_151),
.B2(n_166),
.Y(n_237)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_150),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_228),
.B(n_230),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_L g229 ( 
.A1(n_118),
.A2(n_60),
.B1(n_56),
.B2(n_107),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_146),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_232),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_167),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_146),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_148),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_197),
.B(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_235),
.B(n_183),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_236),
.B(n_191),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_243),
.B1(n_266),
.B2(n_229),
.Y(n_276)
);

NAND2x1_ASAP7_75t_SL g239 ( 
.A(n_181),
.B(n_156),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_239),
.A2(n_184),
.B(n_218),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_153),
.C(n_170),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_241),
.B(n_207),
.C(n_182),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_188),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_254),
.A2(n_225),
.B1(n_141),
.B2(n_233),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

AOI32xp33_ASAP7_75t_L g263 ( 
.A1(n_201),
.A2(n_112),
.A3(n_145),
.B1(n_158),
.B2(n_160),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_263),
.B(n_208),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_204),
.A2(n_198),
.B1(n_227),
.B2(n_224),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_268),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_200),
.B(n_148),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_212),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g275 ( 
.A(n_250),
.B(n_188),
.C(n_200),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_275),
.B(n_278),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_276),
.A2(n_280),
.B1(n_244),
.B2(n_249),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_277),
.A2(n_282),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_287),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_237),
.A2(n_168),
.B1(n_203),
.B2(n_190),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_260),
.Y(n_281)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_281),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_283),
.B(n_288),
.C(n_291),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g284 ( 
.A(n_271),
.B(n_205),
.Y(n_284)
);

OAI21xp33_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_269),
.B(n_267),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_286),
.B(n_296),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_230),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_194),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_289),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_250),
.B(n_202),
.C(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_220),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_293),
.B(n_257),
.Y(n_330)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_247),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_294),
.B(n_299),
.Y(n_313)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_255),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_235),
.B(n_248),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_272),
.Y(n_297)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_297),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_239),
.A2(n_141),
.B1(n_196),
.B2(n_186),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_298),
.A2(n_303),
.B1(n_243),
.B2(n_258),
.Y(n_312)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_272),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_257),
.B(n_219),
.C(n_149),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_263),
.Y(n_315)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_302),
.B(n_304),
.Y(n_333)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_246),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_239),
.A2(n_179),
.B(n_127),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_258),
.B(n_244),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_273),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_311),
.A2(n_329),
.B1(n_336),
.B2(n_303),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_312),
.A2(n_326),
.B1(n_328),
.B2(n_242),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_314),
.A2(n_285),
.B(n_293),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_283),
.C(n_291),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_290),
.B(n_253),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_318),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_325),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_286),
.B(n_245),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_330),
.Y(n_339)
);

OAI21xp33_ASAP7_75t_L g359 ( 
.A1(n_324),
.A2(n_256),
.B(n_265),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_279),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_301),
.A2(n_238),
.B1(n_270),
.B2(n_269),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_302),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_327),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_301),
.A2(n_238),
.B1(n_270),
.B2(n_242),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_281),
.A2(n_270),
.B1(n_274),
.B2(n_264),
.Y(n_329)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_300),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_331),
.B(n_335),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_287),
.B(n_257),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_276),
.A2(n_231),
.B1(n_258),
.B2(n_264),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_288),
.B(n_274),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_337),
.B(n_234),
.Y(n_357)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_334),
.Y(n_340)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_340),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_318),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_341),
.B(n_346),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_342),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_345),
.B(n_322),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_318),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_348),
.A2(n_355),
.B(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_334),
.Y(n_350)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_311),
.A2(n_292),
.B1(n_285),
.B2(n_289),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_356),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_332),
.B(n_278),
.C(n_275),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_354),
.C(n_364),
.Y(n_374)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_338),
.Y(n_353)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_353),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_306),
.C(n_297),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_318),
.A2(n_280),
.B(n_299),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_336),
.A2(n_295),
.B1(n_307),
.B2(n_255),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_357),
.B(n_358),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_315),
.A2(n_240),
.B1(n_256),
.B2(n_234),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g381 ( 
.A1(n_359),
.A2(n_326),
.B(n_328),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g360 ( 
.A1(n_314),
.A2(n_335),
.B(n_308),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_361),
.A2(n_362),
.B1(n_347),
.B2(n_359),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_325),
.A2(n_240),
.B1(n_265),
.B2(n_304),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_362),
.A2(n_329),
.B1(n_323),
.B2(n_327),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_333),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_363),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_322),
.B(n_252),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_313),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_365),
.B(n_368),
.Y(n_382)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_315),
.A2(n_259),
.B1(n_252),
.B2(n_144),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_367),
.B(n_337),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_313),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_340),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_370),
.B(n_379),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_372),
.A2(n_387),
.B1(n_392),
.B2(n_342),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_376),
.B(n_351),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_339),
.B(n_320),
.Y(n_380)
);

CKINVDCx14_ASAP7_75t_R g412 ( 
.A(n_380),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_381),
.A2(n_396),
.B(n_356),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_350),
.B(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_385),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_343),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_386),
.B(n_394),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_361),
.A2(n_317),
.B1(n_310),
.B2(n_321),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_SL g388 ( 
.A(n_339),
.B(n_316),
.Y(n_388)
);

NAND3xp33_ASAP7_75t_L g414 ( 
.A(n_388),
.B(n_357),
.C(n_344),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_389),
.B(n_393),
.C(n_354),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_SL g390 ( 
.A(n_345),
.B(n_309),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_352),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_364),
.B(n_309),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_349),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_363),
.B(n_310),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_395),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_347),
.A2(n_308),
.B(n_330),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_348),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_360),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_349),
.B(n_317),
.Y(n_399)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_399),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_401),
.A2(n_397),
.B1(n_391),
.B2(n_375),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_403),
.B(n_404),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_405),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_406),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_388),
.B(n_395),
.Y(n_407)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_407),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_374),
.B(n_389),
.C(n_364),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_409),
.B(n_419),
.C(n_393),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_385),
.B(n_316),
.Y(n_410)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_399),
.Y(n_413)
);

INVxp67_ASAP7_75t_L g450 ( 
.A(n_413),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_414),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_394),
.Y(n_416)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_417),
.B1(n_426),
.B2(n_427),
.Y(n_440)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_397),
.A2(n_347),
.B1(n_355),
.B2(n_358),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_418),
.A2(n_425),
.B1(n_392),
.B2(n_387),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_374),
.B(n_367),
.C(n_344),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_381),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_379),
.B(n_353),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_422),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_366),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_383),
.B(n_333),
.Y(n_423)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_424),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_380),
.B(n_323),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_397),
.A2(n_312),
.B1(n_152),
.B2(n_91),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_383),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_382),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_371),
.B(n_259),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_428),
.B(n_396),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_370),
.B(n_222),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_429),
.B(n_373),
.Y(n_453)
);

XOR2x1_ASAP7_75t_SL g430 ( 
.A(n_406),
.B(n_391),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_430),
.B(n_441),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_434),
.B(n_447),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_435),
.A2(n_418),
.B1(n_425),
.B2(n_369),
.Y(n_457)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_438),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_401),
.A2(n_412),
.B1(n_408),
.B2(n_375),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_439),
.A2(n_442),
.B1(n_446),
.B2(n_426),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_408),
.A2(n_382),
.B1(n_384),
.B2(n_378),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_409),
.B(n_390),
.Y(n_443)
);

XOR2xp5_ASAP7_75t_L g470 ( 
.A(n_443),
.B(n_444),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_427),
.A2(n_384),
.B1(n_378),
.B2(n_377),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_419),
.B(n_376),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_403),
.B(n_373),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_448),
.B(n_451),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_404),
.B(n_420),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_415),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_434),
.B(n_421),
.C(n_422),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_459),
.C(n_460),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_455),
.B(n_457),
.Y(n_474)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_440),
.Y(n_458)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_458),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_451),
.B(n_411),
.C(n_402),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_411),
.C(n_402),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_436),
.A2(n_413),
.B1(n_369),
.B2(n_423),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_472),
.B1(n_433),
.B2(n_410),
.Y(n_485)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_449),
.Y(n_464)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_465),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_430),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_466),
.B(n_473),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_468),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_445),
.B(n_416),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_447),
.B(n_448),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_469),
.B(n_211),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_432),
.A2(n_407),
.B1(n_372),
.B2(n_417),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_437),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_441),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_475),
.B(n_484),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_459),
.A2(n_450),
.B1(n_415),
.B2(n_400),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_477),
.B(n_485),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_460),
.A2(n_450),
.B(n_400),
.Y(n_481)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_481),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_466),
.A2(n_438),
.B(n_433),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_482),
.B(n_11),
.Y(n_505)
);

MAJx2_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_377),
.C(n_431),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_443),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_486),
.B(n_487),
.C(n_470),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_428),
.C(n_157),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_461),
.B(n_222),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_488),
.B(n_490),
.Y(n_502)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_454),
.B(n_211),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_491),
.B(n_52),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_478),
.A2(n_462),
.B(n_469),
.Y(n_492)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_492),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_507),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_478),
.B(n_470),
.C(n_463),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_494),
.B(n_501),
.C(n_29),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_476),
.B(n_479),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_496),
.B(n_500),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_480),
.A2(n_463),
.B(n_457),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_499),
.B(n_504),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_45),
.Y(n_500)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_474),
.B(n_36),
.C(n_211),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_483),
.B(n_11),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_503),
.B(n_506),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_474),
.B(n_52),
.C(n_31),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_505),
.B(n_10),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_29),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_497),
.A2(n_491),
.B1(n_475),
.B2(n_482),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_509),
.B(n_510),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_500),
.A2(n_486),
.B1(n_484),
.B2(n_31),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_31),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_511),
.B(n_516),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_513),
.B(n_3),
.Y(n_527)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_514),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_498),
.B(n_29),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_493),
.B(n_52),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_517),
.B(n_519),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_505),
.B(n_5),
.Y(n_519)
);

AOI321xp33_ASAP7_75t_L g521 ( 
.A1(n_495),
.A2(n_10),
.A3(n_14),
.B1(n_3),
.B2(n_4),
.C(n_15),
.Y(n_521)
);

NOR2xp67_ASAP7_75t_L g528 ( 
.A(n_521),
.B(n_520),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_518),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_523),
.B(n_527),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g524 ( 
.A1(n_512),
.A2(n_502),
.B1(n_495),
.B2(n_501),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_524),
.B(n_529),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_528),
.B(n_508),
.Y(n_536)
);

CKINVDCx14_ASAP7_75t_R g529 ( 
.A(n_513),
.Y(n_529)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_530),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_531),
.B(n_534),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_SL g533 ( 
.A1(n_529),
.A2(n_511),
.B(n_508),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_SL g537 ( 
.A1(n_533),
.A2(n_535),
.B(n_532),
.Y(n_537)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_522),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_536),
.B(n_526),
.C(n_4),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_537),
.B(n_539),
.Y(n_541)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_535),
.B(n_525),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_540),
.B(n_10),
.C(n_11),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_538),
.B(n_0),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_543),
.B(n_541),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g545 ( 
.A1(n_544),
.A2(n_0),
.B(n_1),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_545),
.B(n_1),
.Y(n_546)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_546),
.A2(n_1),
.B(n_415),
.Y(n_547)
);


endmodule