module real_aes_7202_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_502;
wire n_434;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_756;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g514 ( .A1(n_0), .A2(n_179), .B(n_515), .C(n_518), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_1), .B(n_510), .Y(n_519) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g128 ( .A(n_2), .Y(n_128) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_3), .A2(n_105), .B1(n_117), .B2(n_777), .Y(n_104) );
INVx1_ASAP7_75t_L g177 ( .A(n_4), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g583 ( .A(n_5), .B(n_180), .Y(n_583) );
OAI22xp5_ASAP7_75t_SL g132 ( .A1(n_6), .A2(n_133), .B1(n_136), .B2(n_137), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g137 ( .A(n_6), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g553 ( .A1(n_7), .A2(n_478), .B(n_554), .Y(n_553) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_8), .A2(n_187), .B(n_533), .Y(n_532) );
AOI22xp33_ASAP7_75t_L g233 ( .A1(n_9), .A2(n_39), .B1(n_167), .B2(n_215), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_10), .B(n_187), .Y(n_195) );
AND2x6_ASAP7_75t_L g182 ( .A(n_11), .B(n_183), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_12), .A2(n_182), .B(n_483), .C(n_527), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g133 ( .A1(n_13), .A2(n_43), .B1(n_134), .B2(n_135), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_13), .Y(n_134) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g129 ( .A(n_14), .B(n_40), .Y(n_129) );
INVx1_ASAP7_75t_L g161 ( .A(n_15), .Y(n_161) );
INVx1_ASAP7_75t_L g158 ( .A(n_16), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_17), .B(n_163), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_18), .B(n_180), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_19), .B(n_154), .Y(n_261) );
AO32x2_ASAP7_75t_L g231 ( .A1(n_20), .A2(n_153), .A3(n_187), .B1(n_206), .B2(n_232), .Y(n_231) );
AOI222xp33_ASAP7_75t_SL g131 ( .A1(n_21), .A2(n_132), .B1(n_138), .B2(n_756), .C1(n_757), .C2(n_759), .Y(n_131) );
NAND2xp5_ASAP7_75t_SL g228 ( .A(n_22), .B(n_167), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_23), .B(n_154), .Y(n_184) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_24), .A2(n_58), .B1(n_167), .B2(n_215), .Y(n_234) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_25), .Y(n_130) );
AOI22xp33_ASAP7_75t_SL g217 ( .A1(n_26), .A2(n_84), .B1(n_163), .B2(n_167), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_27), .B(n_167), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_28), .A2(n_206), .B(n_483), .C(n_501), .Y(n_500) );
A2O1A1Ixp33_ASAP7_75t_L g535 ( .A1(n_29), .A2(n_206), .B(n_483), .C(n_536), .Y(n_535) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_30), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_31), .B(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_32), .A2(n_478), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_33), .B(n_208), .Y(n_249) );
INVx2_ASAP7_75t_L g165 ( .A(n_34), .Y(n_165) );
A2O1A1Ixp33_ASAP7_75t_L g480 ( .A1(n_35), .A2(n_481), .B(n_485), .C(n_491), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_36), .B(n_167), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_37), .B(n_208), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_38), .B(n_226), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_40), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_41), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g531 ( .A(n_42), .Y(n_531) );
INVx1_ASAP7_75t_L g135 ( .A(n_43), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_44), .B(n_180), .Y(n_548) );
OAI22xp5_ASAP7_75t_SL g769 ( .A1(n_45), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_769) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_45), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_46), .B(n_478), .Y(n_534) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_47), .A2(n_141), .B1(n_142), .B2(n_463), .Y(n_140) );
INVx1_ASAP7_75t_L g463 ( .A(n_47), .Y(n_463) );
OAI22xp5_ASAP7_75t_SL g770 ( .A1(n_47), .A2(n_49), .B1(n_463), .B2(n_771), .Y(n_770) );
A2O1A1Ixp33_ASAP7_75t_L g545 ( .A1(n_48), .A2(n_481), .B(n_491), .C(n_546), .Y(n_545) );
CKINVDCx20_ASAP7_75t_R g771 ( .A(n_49), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_50), .B(n_167), .Y(n_190) );
INVx1_ASAP7_75t_L g516 ( .A(n_51), .Y(n_516) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_52), .A2(n_93), .B1(n_215), .B2(n_216), .Y(n_214) );
INVx1_ASAP7_75t_L g547 ( .A(n_53), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_54), .B(n_167), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_55), .B(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_56), .B(n_478), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_57), .B(n_175), .Y(n_194) );
AOI22xp33_ASAP7_75t_SL g259 ( .A1(n_59), .A2(n_63), .B1(n_163), .B2(n_167), .Y(n_259) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_60), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_61), .B(n_167), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_62), .B(n_167), .Y(n_223) );
INVx1_ASAP7_75t_L g183 ( .A(n_64), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_65), .B(n_478), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_66), .B(n_510), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g556 ( .A1(n_67), .A2(n_169), .B(n_175), .C(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_68), .B(n_167), .Y(n_178) );
INVx1_ASAP7_75t_L g157 ( .A(n_69), .Y(n_157) );
OAI22xp33_ASAP7_75t_SL g766 ( .A1(n_70), .A2(n_767), .B1(n_774), .B2(n_775), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_70), .Y(n_774) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_71), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_72), .B(n_180), .Y(n_489) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_73), .A2(n_187), .A3(n_206), .B1(n_213), .B2(n_218), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_74), .B(n_181), .Y(n_528) );
INVx1_ASAP7_75t_L g202 ( .A(n_75), .Y(n_202) );
INVx1_ASAP7_75t_L g244 ( .A(n_76), .Y(n_244) );
CKINVDCx16_ASAP7_75t_R g513 ( .A(n_77), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_78), .B(n_488), .Y(n_502) );
A2O1A1Ixp33_ASAP7_75t_L g580 ( .A1(n_79), .A2(n_483), .B(n_491), .C(n_581), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_80), .B(n_163), .Y(n_245) );
CKINVDCx16_ASAP7_75t_R g555 ( .A(n_81), .Y(n_555) );
INVx1_ASAP7_75t_L g116 ( .A(n_82), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_83), .B(n_487), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_85), .B(n_215), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_86), .Y(n_494) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_87), .B(n_163), .Y(n_248) );
INVx2_ASAP7_75t_L g155 ( .A(n_88), .Y(n_155) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_89), .Y(n_587) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_90), .B(n_205), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_91), .B(n_163), .Y(n_191) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
OR2x2_ASAP7_75t_L g125 ( .A(n_92), .B(n_126), .Y(n_125) );
OR2x2_ASAP7_75t_L g466 ( .A(n_92), .B(n_127), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g258 ( .A1(n_94), .A2(n_103), .B1(n_163), .B2(n_164), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_95), .B(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g486 ( .A(n_96), .Y(n_486) );
INVxp67_ASAP7_75t_L g558 ( .A(n_97), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_98), .B(n_163), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g524 ( .A(n_100), .Y(n_524) );
INVx1_ASAP7_75t_L g582 ( .A(n_101), .Y(n_582) );
AND2x2_ASAP7_75t_L g549 ( .A(n_102), .B(n_208), .Y(n_549) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx2_ASAP7_75t_SL g777 ( .A(n_107), .Y(n_777) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g469 ( .A(n_113), .B(n_127), .Y(n_469) );
NOR2x2_ASAP7_75t_L g761 ( .A(n_113), .B(n_126), .Y(n_761) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx3_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
AOI22xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_131), .B1(n_762), .B2(n_765), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g764 ( .A(n_122), .Y(n_764) );
AOI21xp5_ASAP7_75t_L g765 ( .A1(n_123), .A2(n_766), .B(n_776), .Y(n_765) );
NOR2xp33_ASAP7_75t_SL g123 ( .A(n_124), .B(n_130), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
HB1xp67_ASAP7_75t_L g776 ( .A(n_125), .Y(n_776) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
INVx1_ASAP7_75t_L g756 ( .A(n_132), .Y(n_756) );
CKINVDCx14_ASAP7_75t_R g136 ( .A(n_133), .Y(n_136) );
OAI22x1_ASAP7_75t_SL g138 ( .A1(n_139), .A2(n_464), .B1(n_467), .B2(n_470), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g757 ( .A1(n_140), .A2(n_464), .B1(n_469), .B2(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_141), .A2(n_142), .B1(n_768), .B2(n_769), .Y(n_767) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_SL g142 ( .A(n_143), .B(n_429), .Y(n_142) );
NOR3xp33_ASAP7_75t_L g143 ( .A(n_144), .B(n_333), .C(n_417), .Y(n_143) );
NAND4xp25_ASAP7_75t_L g144 ( .A(n_145), .B(n_276), .C(n_298), .D(n_314), .Y(n_144) );
AOI221xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_209), .B1(n_235), .B2(n_254), .C(n_262), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_185), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g288 ( .A(n_148), .B(n_254), .Y(n_288) );
NAND4xp25_ASAP7_75t_L g328 ( .A(n_148), .B(n_316), .C(n_329), .D(n_331), .Y(n_328) );
INVxp67_ASAP7_75t_L g445 ( .A(n_148), .Y(n_445) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OR2x2_ASAP7_75t_L g327 ( .A(n_149), .B(n_265), .Y(n_327) );
AND2x2_ASAP7_75t_L g351 ( .A(n_149), .B(n_185), .Y(n_351) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x2_ASAP7_75t_L g318 ( .A(n_150), .B(n_253), .Y(n_318) );
AND2x2_ASAP7_75t_L g358 ( .A(n_150), .B(n_339), .Y(n_358) );
AND2x2_ASAP7_75t_L g375 ( .A(n_150), .B(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_150), .B(n_186), .Y(n_399) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x2_ASAP7_75t_L g252 ( .A(n_151), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g270 ( .A(n_151), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g282 ( .A(n_151), .B(n_186), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_151), .B(n_196), .Y(n_304) );
OA21x2_ASAP7_75t_L g151 ( .A1(n_152), .A2(n_159), .B(n_184), .Y(n_151) );
OA21x2_ASAP7_75t_L g196 ( .A1(n_152), .A2(n_197), .B(n_207), .Y(n_196) );
INVx2_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_153), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_154), .Y(n_187) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
AND2x2_ASAP7_75t_SL g208 ( .A(n_155), .B(n_156), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
OAI21xp5_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_173), .B(n_182), .Y(n_159) );
O2A1O1Ixp33_ASAP7_75t_L g160 ( .A1(n_161), .A2(n_162), .B(n_166), .C(n_169), .Y(n_160) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_162), .A2(n_528), .B(n_529), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g536 ( .A1(n_162), .A2(n_537), .B(n_538), .Y(n_536) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
INVx2_ASAP7_75t_L g168 ( .A(n_165), .Y(n_168) );
INVx1_ASAP7_75t_L g176 ( .A(n_165), .Y(n_176) );
INVx3_ASAP7_75t_L g243 ( .A(n_167), .Y(n_243) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_167), .Y(n_584) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx1_ASAP7_75t_L g215 ( .A(n_168), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_168), .Y(n_216) );
AND2x6_ASAP7_75t_L g483 ( .A(n_168), .B(n_484), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g581 ( .A1(n_169), .A2(n_582), .B(n_583), .C(n_584), .Y(n_581) );
INVx1_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_170), .A2(n_247), .B(n_248), .Y(n_246) );
INVx4_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g488 ( .A(n_171), .Y(n_488) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx3_ASAP7_75t_L g181 ( .A(n_172), .Y(n_181) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_172), .Y(n_205) );
INVx1_ASAP7_75t_L g226 ( .A(n_172), .Y(n_226) );
AND2x2_ASAP7_75t_L g479 ( .A(n_172), .B(n_176), .Y(n_479) );
INVx1_ASAP7_75t_L g484 ( .A(n_172), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_177), .B(n_178), .C(n_179), .Y(n_173) );
O2A1O1Ixp5_ASAP7_75t_L g201 ( .A1(n_174), .A2(n_202), .B(n_203), .C(n_204), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_174), .A2(n_502), .B(n_503), .Y(n_501) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_179), .A2(n_193), .B(n_194), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g232 ( .A1(n_179), .A2(n_205), .B1(n_233), .B2(n_234), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_179), .A2(n_205), .B1(n_258), .B2(n_259), .Y(n_257) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_180), .A2(n_190), .B(n_191), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_180), .A2(n_199), .B(n_200), .Y(n_198) );
O2A1O1Ixp5_ASAP7_75t_SL g242 ( .A1(n_180), .A2(n_243), .B(n_244), .C(n_245), .Y(n_242) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_180), .B(n_558), .Y(n_557) );
INVx5_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g213 ( .A1(n_181), .A2(n_205), .B1(n_214), .B2(n_217), .Y(n_213) );
OAI21xp5_ASAP7_75t_L g188 ( .A1(n_182), .A2(n_189), .B(n_192), .Y(n_188) );
BUFx3_ASAP7_75t_L g206 ( .A(n_182), .Y(n_206) );
OAI21xp5_ASAP7_75t_L g221 ( .A1(n_182), .A2(n_222), .B(n_227), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g241 ( .A1(n_182), .A2(n_242), .B(n_246), .Y(n_241) );
AND2x4_ASAP7_75t_L g478 ( .A(n_182), .B(n_479), .Y(n_478) );
INVx4_ASAP7_75t_SL g492 ( .A(n_182), .Y(n_492) );
NAND2x1p5_ASAP7_75t_L g525 ( .A(n_182), .B(n_479), .Y(n_525) );
AND2x2_ASAP7_75t_L g285 ( .A(n_185), .B(n_286), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g334 ( .A1(n_185), .A2(n_335), .B1(n_338), .B2(n_340), .C(n_344), .Y(n_334) );
AND2x2_ASAP7_75t_L g393 ( .A(n_185), .B(n_358), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_185), .B(n_375), .Y(n_427) );
AND2x2_ASAP7_75t_L g185 ( .A(n_186), .B(n_196), .Y(n_185) );
INVx3_ASAP7_75t_L g253 ( .A(n_186), .Y(n_253) );
AND2x2_ASAP7_75t_L g302 ( .A(n_186), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g356 ( .A(n_186), .B(n_271), .Y(n_356) );
AND2x2_ASAP7_75t_L g414 ( .A(n_186), .B(n_415), .Y(n_414) );
OA21x2_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_195), .Y(n_186) );
INVx4_ASAP7_75t_L g256 ( .A(n_187), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_187), .A2(n_534), .B(n_535), .Y(n_533) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_187), .Y(n_552) );
AND2x2_ASAP7_75t_L g254 ( .A(n_196), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g271 ( .A(n_196), .Y(n_271) );
INVx1_ASAP7_75t_L g326 ( .A(n_196), .Y(n_326) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_196), .Y(n_332) );
AND2x2_ASAP7_75t_L g377 ( .A(n_196), .B(n_253), .Y(n_377) );
OR2x2_ASAP7_75t_L g416 ( .A(n_196), .B(n_255), .Y(n_416) );
OAI21xp5_ASAP7_75t_L g197 ( .A1(n_198), .A2(n_201), .B(n_206), .Y(n_197) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_204), .A2(n_228), .B(n_229), .Y(n_227) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
INVx4_ASAP7_75t_L g517 ( .A(n_205), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g275 ( .A(n_206), .B(n_256), .C(n_257), .Y(n_275) );
INVx2_ASAP7_75t_L g218 ( .A(n_208), .Y(n_218) );
OA21x2_ASAP7_75t_L g220 ( .A1(n_208), .A2(n_221), .B(n_230), .Y(n_220) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_208), .A2(n_241), .B(n_249), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_208), .A2(n_477), .B(n_480), .Y(n_476) );
INVx1_ASAP7_75t_L g507 ( .A(n_208), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g543 ( .A1(n_208), .A2(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_209), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
AND2x2_ASAP7_75t_L g412 ( .A(n_210), .B(n_409), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_210), .B(n_394), .Y(n_444) );
BUFx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g343 ( .A(n_211), .B(n_267), .Y(n_343) );
AND2x2_ASAP7_75t_L g392 ( .A(n_211), .B(n_238), .Y(n_392) );
INVx1_ASAP7_75t_L g438 ( .A(n_211), .Y(n_438) );
INVx1_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
BUFx6f_ASAP7_75t_L g251 ( .A(n_212), .Y(n_251) );
AND2x2_ASAP7_75t_L g293 ( .A(n_212), .B(n_267), .Y(n_293) );
INVx1_ASAP7_75t_L g310 ( .A(n_212), .Y(n_310) );
AND2x2_ASAP7_75t_L g316 ( .A(n_212), .B(n_231), .Y(n_316) );
HB1xp67_ASAP7_75t_L g490 ( .A(n_216), .Y(n_490) );
INVx2_ASAP7_75t_L g518 ( .A(n_216), .Y(n_518) );
INVx1_ASAP7_75t_L g504 ( .A(n_218), .Y(n_504) );
AND2x2_ASAP7_75t_L g384 ( .A(n_219), .B(n_292), .Y(n_384) );
INVx2_ASAP7_75t_L g449 ( .A(n_219), .Y(n_449) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_231), .Y(n_219) );
AND2x2_ASAP7_75t_L g266 ( .A(n_220), .B(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g279 ( .A(n_220), .B(n_239), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_220), .B(n_238), .Y(n_307) );
INVx1_ASAP7_75t_L g313 ( .A(n_220), .Y(n_313) );
INVx1_ASAP7_75t_L g330 ( .A(n_220), .Y(n_330) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_220), .Y(n_342) );
INVx2_ASAP7_75t_L g410 ( .A(n_220), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_223), .A2(n_224), .B(n_225), .Y(n_222) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
INVx2_ASAP7_75t_L g267 ( .A(n_231), .Y(n_267) );
BUFx2_ASAP7_75t_L g364 ( .A(n_231), .Y(n_364) );
AND2x2_ASAP7_75t_L g409 ( .A(n_231), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_237), .B(n_346), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g432 ( .A1(n_237), .A2(n_408), .B(n_422), .Y(n_432) );
AND2x2_ASAP7_75t_L g457 ( .A(n_237), .B(n_343), .Y(n_457) );
BUFx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g379 ( .A(n_239), .Y(n_379) );
AND2x2_ASAP7_75t_L g408 ( .A(n_239), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_240), .Y(n_292) );
INVx2_ASAP7_75t_L g311 ( .A(n_240), .Y(n_311) );
OR2x2_ASAP7_75t_L g312 ( .A(n_240), .B(n_313), .Y(n_312) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx2_ASAP7_75t_L g265 ( .A(n_251), .Y(n_265) );
OR2x2_ASAP7_75t_L g278 ( .A(n_251), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g346 ( .A(n_251), .B(n_342), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_251), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g447 ( .A(n_251), .B(n_448), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_251), .B(n_384), .Y(n_459) );
AND2x2_ASAP7_75t_L g338 ( .A(n_252), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g361 ( .A(n_252), .B(n_254), .Y(n_361) );
INVx2_ASAP7_75t_L g273 ( .A(n_253), .Y(n_273) );
AND2x2_ASAP7_75t_L g301 ( .A(n_253), .B(n_274), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_253), .B(n_326), .Y(n_382) );
AND2x2_ASAP7_75t_L g296 ( .A(n_254), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g443 ( .A(n_254), .Y(n_443) );
AND2x2_ASAP7_75t_L g455 ( .A(n_254), .B(n_318), .Y(n_455) );
AND2x2_ASAP7_75t_L g281 ( .A(n_255), .B(n_271), .Y(n_281) );
INVx1_ASAP7_75t_L g376 ( .A(n_255), .Y(n_376) );
AO21x1_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_257), .B(n_260), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_256), .B(n_494), .Y(n_493) );
INVx3_ASAP7_75t_L g510 ( .A(n_256), .Y(n_510) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_256), .A2(n_523), .B(n_530), .Y(n_522) );
AO21x2_ASAP7_75t_L g578 ( .A1(n_256), .A2(n_579), .B(n_586), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g586 ( .A(n_256), .B(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x4_ASAP7_75t_L g274 ( .A(n_261), .B(n_275), .Y(n_274) );
INVxp67_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_264), .B(n_268), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_265), .B(n_312), .Y(n_321) );
OR2x2_ASAP7_75t_L g453 ( .A(n_265), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g370 ( .A(n_266), .B(n_311), .Y(n_370) );
AND2x2_ASAP7_75t_L g378 ( .A(n_266), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g437 ( .A(n_266), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g461 ( .A(n_266), .B(n_308), .Y(n_461) );
NOR2xp67_ASAP7_75t_L g419 ( .A(n_267), .B(n_420), .Y(n_419) );
OR2x2_ASAP7_75t_L g448 ( .A(n_267), .B(n_311), .Y(n_448) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g269 ( .A(n_270), .B(n_272), .Y(n_269) );
AND2x2_ASAP7_75t_L g300 ( .A(n_270), .B(n_301), .Y(n_300) );
INVxp67_ASAP7_75t_L g462 ( .A(n_270), .Y(n_462) );
NOR2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g297 ( .A(n_273), .Y(n_297) );
AND2x2_ASAP7_75t_L g348 ( .A(n_273), .B(n_281), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_273), .B(n_416), .Y(n_442) );
INVx2_ASAP7_75t_L g287 ( .A(n_274), .Y(n_287) );
INVx3_ASAP7_75t_L g339 ( .A(n_274), .Y(n_339) );
OR2x2_ASAP7_75t_L g367 ( .A(n_274), .B(n_368), .Y(n_367) );
AOI311xp33_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_280), .A3(n_282), .B(n_283), .C(n_294), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g314 ( .A1(n_277), .A2(n_315), .B(n_317), .C(n_319), .Y(n_314) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_SL g299 ( .A(n_279), .Y(n_299) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g317 ( .A(n_281), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_281), .B(n_297), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_281), .B(n_282), .Y(n_450) );
AND2x2_ASAP7_75t_L g372 ( .A(n_282), .B(n_286), .Y(n_372) );
AOI21xp33_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_288), .B(n_289), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g430 ( .A(n_286), .B(n_318), .Y(n_430) );
INVx2_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g303 ( .A(n_287), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g324 ( .A(n_287), .Y(n_324) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
AND2x2_ASAP7_75t_L g315 ( .A(n_291), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g360 ( .A(n_293), .Y(n_360) );
AND2x4_ASAP7_75t_L g422 ( .A(n_293), .B(n_391), .Y(n_422) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AOI222xp33_ASAP7_75t_L g373 ( .A1(n_296), .A2(n_362), .B1(n_374), .B2(n_378), .C1(n_380), .C2(n_384), .Y(n_373) );
A2O1A1Ixp33_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_302), .C(n_305), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_299), .B(n_343), .Y(n_366) );
INVx1_ASAP7_75t_L g388 ( .A(n_301), .Y(n_388) );
INVx1_ASAP7_75t_L g322 ( .A(n_303), .Y(n_322) );
OR2x2_ASAP7_75t_L g387 ( .A(n_304), .B(n_388), .Y(n_387) );
OAI21xp33_ASAP7_75t_SL g305 ( .A1(n_306), .A2(n_308), .B(n_312), .Y(n_305) );
NAND3xp33_ASAP7_75t_L g323 ( .A(n_306), .B(n_324), .C(n_325), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_306), .A2(n_343), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_310), .Y(n_363) );
AND2x2_ASAP7_75t_SL g329 ( .A(n_311), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g420 ( .A(n_311), .Y(n_420) );
HB1xp67_ASAP7_75t_L g436 ( .A(n_311), .Y(n_436) );
INVx2_ASAP7_75t_L g394 ( .A(n_312), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_316), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g368 ( .A(n_318), .Y(n_368) );
OAI221xp5_ASAP7_75t_L g319 ( .A1(n_320), .A2(n_322), .B1(n_323), .B2(n_327), .C(n_328), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp5_ASAP7_75t_SL g401 ( .A(n_322), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_SL g456 ( .A(n_322), .Y(n_456) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVx2_ASAP7_75t_L g337 ( .A(n_329), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_329), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g395 ( .A(n_329), .B(n_343), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_329), .B(n_405), .Y(n_404) );
AND2x2_ASAP7_75t_L g428 ( .A(n_329), .B(n_363), .Y(n_428) );
BUFx3_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND5xp2_ASAP7_75t_L g333 ( .A(n_334), .B(n_352), .C(n_373), .D(n_385), .E(n_400), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI32xp33_ASAP7_75t_L g425 ( .A1(n_337), .A2(n_364), .A3(n_380), .B1(n_426), .B2(n_428), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_339), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_343), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_SL g349 ( .A(n_343), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_349), .B2(n_350), .Y(n_344) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI221xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_359), .B1(n_361), .B2(n_362), .C(n_365), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_357), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g424 ( .A(n_356), .B(n_375), .Y(n_424) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
AOI221xp5_ASAP7_75t_L g439 ( .A1(n_361), .A2(n_422), .B1(n_440), .B2(n_445), .C(n_446), .Y(n_439) );
AND2x2_ASAP7_75t_L g362 ( .A(n_363), .B(n_364), .Y(n_362) );
INVx2_ASAP7_75t_L g405 ( .A(n_364), .Y(n_405) );
OAI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_367), .B1(n_369), .B2(n_371), .Y(n_365) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g383 ( .A(n_375), .Y(n_383) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AOI222xp33_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_389), .B1(n_393), .B2(n_394), .C1(n_395), .C2(n_396), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g389 ( .A(n_390), .B(n_392), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
OAI22xp33_ASAP7_75t_L g440 ( .A1(n_394), .A2(n_441), .B1(n_443), .B2(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_SL g398 ( .A(n_399), .Y(n_398) );
AOI21xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_406), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g406 ( .A1(n_407), .A2(n_411), .B(n_413), .Y(n_406) );
INVx2_ASAP7_75t_SL g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g454 ( .A(n_409), .Y(n_454) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
A2O1A1Ixp33_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_421), .B(n_423), .C(n_425), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AOI211xp5_ASAP7_75t_L g429 ( .A1(n_430), .A2(n_431), .B(n_433), .C(n_458), .Y(n_429) );
CKINVDCx16_ASAP7_75t_R g434 ( .A(n_430), .Y(n_434) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
OAI211xp5_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_435), .B(n_439), .C(n_451), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_437), .Y(n_435) );
AOI21xp33_ASAP7_75t_L g446 ( .A1(n_447), .A2(n_449), .B(n_450), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_455), .B1(n_456), .B2(n_457), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
AOI21xp33_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_462), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g758 ( .A(n_470), .Y(n_758) );
OR3x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_670), .C(n_713), .Y(n_470) );
NAND5xp2_ASAP7_75t_L g471 ( .A(n_472), .B(n_597), .C(n_627), .D(n_644), .E(n_659), .Y(n_471) );
AOI221xp5_ASAP7_75t_SL g472 ( .A1(n_473), .A2(n_520), .B1(n_560), .B2(n_566), .C(n_570), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_495), .Y(n_473) );
OR2x2_ASAP7_75t_L g575 ( .A(n_474), .B(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g614 ( .A(n_474), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g632 ( .A(n_474), .B(n_633), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_474), .B(n_568), .Y(n_649) );
OR2x2_ASAP7_75t_L g661 ( .A(n_474), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_474), .B(n_620), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_474), .B(n_694), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_474), .B(n_598), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_474), .B(n_606), .Y(n_712) );
AND2x2_ASAP7_75t_L g744 ( .A(n_474), .B(n_508), .Y(n_744) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_474), .Y(n_752) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_475), .B(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g572 ( .A(n_475), .B(n_550), .Y(n_572) );
BUFx2_ASAP7_75t_L g594 ( .A(n_475), .Y(n_594) );
AND2x2_ASAP7_75t_L g623 ( .A(n_475), .B(n_496), .Y(n_623) );
AND2x2_ASAP7_75t_L g678 ( .A(n_475), .B(n_576), .Y(n_678) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_493), .Y(n_475) );
BUFx2_ASAP7_75t_L g499 ( .A(n_478), .Y(n_499) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_SL g512 ( .A1(n_482), .A2(n_492), .B(n_513), .C(n_514), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g554 ( .A1(n_482), .A2(n_492), .B(n_555), .C(n_556), .Y(n_554) );
INVx5_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
O2A1O1Ixp33_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_487), .B(n_489), .C(n_490), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g546 ( .A1(n_487), .A2(n_490), .B(n_547), .C(n_548), .Y(n_546) );
INVx2_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_495), .B(n_632), .Y(n_641) );
OAI32xp33_ASAP7_75t_L g655 ( .A1(n_495), .A2(n_591), .A3(n_656), .B1(n_657), .B2(n_658), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_495), .B(n_657), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_495), .B(n_575), .Y(n_698) );
INVx1_ASAP7_75t_SL g727 ( .A(n_495), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g736 ( .A(n_495), .B(n_522), .C(n_678), .D(n_737), .Y(n_736) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_508), .Y(n_495) );
INVx5_ASAP7_75t_L g569 ( .A(n_496), .Y(n_569) );
AND2x2_ASAP7_75t_L g598 ( .A(n_496), .B(n_509), .Y(n_598) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_496), .Y(n_677) );
AND2x2_ASAP7_75t_L g747 ( .A(n_496), .B(n_694), .Y(n_747) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_505), .Y(n_496) );
AOI21xp5_ASAP7_75t_SL g497 ( .A1(n_498), .A2(n_500), .B(n_504), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
AND2x4_ASAP7_75t_L g620 ( .A(n_508), .B(n_569), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_508), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g654 ( .A(n_508), .B(n_576), .Y(n_654) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AND2x2_ASAP7_75t_L g568 ( .A(n_509), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g606 ( .A(n_509), .B(n_578), .Y(n_606) );
AND2x2_ASAP7_75t_L g615 ( .A(n_509), .B(n_577), .Y(n_615) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_519), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_517), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_520), .A2(n_684), .B1(n_686), .B2(n_688), .C1(n_691), .C2(n_692), .Y(n_683) );
AND2x4_ASAP7_75t_L g520 ( .A(n_521), .B(n_539), .Y(n_520) );
AND2x2_ASAP7_75t_L g616 ( .A(n_521), .B(n_617), .Y(n_616) );
NAND3xp33_ASAP7_75t_L g733 ( .A(n_521), .B(n_594), .C(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g521 ( .A(n_522), .B(n_532), .Y(n_521) );
INVx5_ASAP7_75t_SL g565 ( .A(n_522), .Y(n_565) );
OAI322xp33_ASAP7_75t_L g570 ( .A1(n_522), .A2(n_571), .A3(n_573), .B1(n_574), .B2(n_588), .C1(n_591), .C2(n_593), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_522), .B(n_563), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_522), .B(n_551), .Y(n_742) );
OAI21xp5_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_525), .B(n_526), .Y(n_523) );
INVx2_ASAP7_75t_L g563 ( .A(n_532), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_532), .B(n_541), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_539), .B(n_601), .Y(n_656) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g635 ( .A(n_540), .B(n_636), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_541), .B(n_550), .Y(n_540) );
OR2x2_ASAP7_75t_L g564 ( .A(n_541), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_541), .B(n_572), .Y(n_571) );
OR2x2_ASAP7_75t_L g603 ( .A(n_541), .B(n_551), .Y(n_603) );
AND2x2_ASAP7_75t_L g626 ( .A(n_541), .B(n_563), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_541), .B(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g642 ( .A(n_541), .B(n_601), .Y(n_642) );
AND2x2_ASAP7_75t_L g650 ( .A(n_541), .B(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_541), .B(n_610), .Y(n_700) );
INVx5_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g590 ( .A(n_542), .B(n_565), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_542), .B(n_592), .Y(n_591) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_551), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_542), .B(n_664), .Y(n_705) );
OR2x2_ASAP7_75t_L g721 ( .A(n_542), .B(n_665), .Y(n_721) );
AND2x2_ASAP7_75t_SL g728 ( .A(n_542), .B(n_682), .Y(n_728) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_542), .Y(n_735) );
OR2x6_ASAP7_75t_L g542 ( .A(n_543), .B(n_549), .Y(n_542) );
AND2x2_ASAP7_75t_L g589 ( .A(n_550), .B(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g639 ( .A(n_550), .B(n_563), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_550), .B(n_565), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_550), .B(n_601), .Y(n_723) );
INVx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_551), .B(n_565), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_551), .B(n_563), .Y(n_611) );
OR2x2_ASAP7_75t_L g665 ( .A(n_551), .B(n_563), .Y(n_665) );
AND2x2_ASAP7_75t_L g682 ( .A(n_551), .B(n_562), .Y(n_682) );
INVxp67_ASAP7_75t_L g704 ( .A(n_551), .Y(n_704) );
AND2x2_ASAP7_75t_L g731 ( .A(n_551), .B(n_601), .Y(n_731) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_551), .Y(n_738) );
OA21x2_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_559), .Y(n_551) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_564), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_562), .B(n_612), .Y(n_685) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g601 ( .A(n_563), .B(n_565), .Y(n_601) );
OR2x2_ASAP7_75t_L g668 ( .A(n_563), .B(n_669), .Y(n_668) );
INVx2_ASAP7_75t_L g612 ( .A(n_564), .Y(n_612) );
OR2x2_ASAP7_75t_L g673 ( .A(n_564), .B(n_665), .Y(n_673) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx1_ASAP7_75t_L g573 ( .A(n_568), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_568), .B(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g574 ( .A(n_569), .B(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_569), .B(n_596), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_569), .B(n_576), .Y(n_608) );
INVx2_ASAP7_75t_L g653 ( .A(n_569), .Y(n_653) );
AND2x2_ASAP7_75t_L g666 ( .A(n_569), .B(n_606), .Y(n_666) );
AND2x2_ASAP7_75t_L g691 ( .A(n_569), .B(n_615), .Y(n_691) );
INVx1_ASAP7_75t_L g643 ( .A(n_574), .Y(n_643) );
INVx2_ASAP7_75t_SL g630 ( .A(n_575), .Y(n_630) );
INVx1_ASAP7_75t_L g633 ( .A(n_576), .Y(n_633) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
HB1xp67_ASAP7_75t_L g596 ( .A(n_577), .Y(n_596) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g694 ( .A(n_578), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_585), .Y(n_579) );
INVx1_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
AND2x2_ASAP7_75t_L g663 ( .A(n_590), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g669 ( .A(n_590), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g671 ( .A1(n_590), .A2(n_672), .B1(n_674), .B2(n_679), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_590), .B(n_682), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_591), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_SL g625 ( .A(n_592), .Y(n_625) );
OR2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
OR2x2_ASAP7_75t_L g607 ( .A(n_594), .B(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_594), .B(n_598), .Y(n_658) );
AND2x2_ASAP7_75t_L g681 ( .A(n_594), .B(n_682), .Y(n_681) );
BUFx2_ASAP7_75t_L g657 ( .A(n_596), .Y(n_657) );
AOI211xp5_ASAP7_75t_L g597 ( .A1(n_598), .A2(n_599), .B(n_604), .C(n_618), .Y(n_597) );
INVx1_ASAP7_75t_L g621 ( .A(n_598), .Y(n_621) );
OAI221xp5_ASAP7_75t_SL g729 ( .A1(n_598), .A2(n_730), .B1(n_732), .B2(n_733), .C(n_736), .Y(n_729) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
INVx1_ASAP7_75t_L g748 ( .A(n_601), .Y(n_748) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g697 ( .A(n_603), .B(n_636), .Y(n_697) );
A2O1A1Ixp33_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_607), .B(n_609), .C(n_613), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_612), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
OAI32xp33_ASAP7_75t_L g722 ( .A1(n_611), .A2(n_612), .A3(n_675), .B1(n_712), .B2(n_723), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
AND2x2_ASAP7_75t_L g754 ( .A(n_614), .B(n_653), .Y(n_754) );
AND2x2_ASAP7_75t_L g701 ( .A(n_615), .B(n_653), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_615), .B(n_623), .Y(n_719) );
AOI31xp33_ASAP7_75t_SL g618 ( .A1(n_619), .A2(n_621), .A3(n_622), .B(n_624), .Y(n_618) );
INVxp67_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_620), .B(n_632), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_620), .B(n_630), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_620), .A2(n_650), .B1(n_740), .B2(n_743), .C(n_745), .Y(n_739) );
CKINVDCx16_ASAP7_75t_R g622 ( .A(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
AND2x2_ASAP7_75t_L g645 ( .A(n_625), .B(n_646), .Y(n_645) );
AOI222xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_634), .B1(n_637), .B2(n_640), .C1(n_642), .C2(n_643), .Y(n_627) );
NAND2xp5_ASAP7_75t_SL g628 ( .A(n_629), .B(n_631), .Y(n_628) );
INVx1_ASAP7_75t_L g710 ( .A(n_629), .Y(n_710) );
INVx1_ASAP7_75t_L g732 ( .A(n_632), .Y(n_732) );
INVx2_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_635), .A2(n_746), .B1(n_748), .B2(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g651 ( .A(n_636), .Y(n_651) );
INVx1_ASAP7_75t_SL g638 ( .A(n_639), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_648), .B1(n_650), .B2(n_652), .C(n_655), .Y(n_644) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g689 ( .A(n_647), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g741 ( .A(n_647), .B(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g716 ( .A(n_652), .Y(n_716) );
AND2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g680 ( .A(n_653), .Y(n_680) );
INVx1_ASAP7_75t_L g662 ( .A(n_654), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_657), .B(n_744), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_660), .A2(n_663), .B1(n_666), .B2(n_667), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_SL g753 ( .A(n_666), .Y(n_753) );
INVxp33_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_668), .B(n_712), .Y(n_711) );
OAI32xp33_ASAP7_75t_L g702 ( .A1(n_669), .A2(n_703), .A3(n_704), .B1(n_705), .B2(n_706), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g670 ( .A(n_671), .B(n_683), .C(n_695), .D(n_707), .Y(n_670) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
NAND2xp33_ASAP7_75t_SL g674 ( .A(n_675), .B(n_676), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_678), .B(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
CKINVDCx16_ASAP7_75t_R g688 ( .A(n_689), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_692), .A2(n_708), .B1(n_725), .B2(n_728), .C(n_729), .Y(n_724) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g743 ( .A(n_694), .B(n_744), .Y(n_743) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_698), .B1(n_699), .B2(n_701), .C(n_702), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g734 ( .A(n_704), .B(n_735), .Y(n_734) );
AOI21xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_710), .B(n_711), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NAND4xp25_ASAP7_75t_L g713 ( .A(n_714), .B(n_724), .C(n_739), .D(n_750), .Y(n_713) );
O2A1O1Ixp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_718), .B(n_720), .C(n_722), .Y(n_714) );
NAND2xp5_ASAP7_75t_SL g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
INVxp67_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_L g755 ( .A(n_742), .Y(n_755) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_754), .B(n_755), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g759 ( .A(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
BUFx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g775 ( .A(n_767), .Y(n_775) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g773 ( .A(n_770), .Y(n_773) );
endmodule