module fake_jpeg_21383_n_174 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_174);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_174;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx11_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx16f_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_34),
.Y(n_55)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_32),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_0),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_7),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_31),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_5),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_15),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_43),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_52),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_76),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_81),
.Y(n_90)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_82),
.Y(n_89)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

CKINVDCx6p67_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_97),
.Y(n_100)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_78),
.Y(n_93)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_91),
.A2(n_71),
.B1(n_63),
.B2(n_66),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_98),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_95),
.B(n_64),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_109),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_87),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_102),
.B(n_106),
.Y(n_119)
);

NAND3xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_58),
.C(n_70),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_103),
.B(n_50),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_94),
.A2(n_56),
.B1(n_52),
.B2(n_70),
.Y(n_108)
);

AOI32xp33_ASAP7_75t_L g127 ( 
.A1(n_108),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_64),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_84),
.B1(n_85),
.B2(n_62),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_110),
.A2(n_111),
.B1(n_62),
.B2(n_53),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_48),
.B1(n_53),
.B2(n_75),
.Y(n_111)
);

AO22x1_ASAP7_75t_L g112 ( 
.A1(n_91),
.A2(n_65),
.B1(n_67),
.B2(n_73),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_114),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_75),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_126),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_55),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_118),
.B(n_121),
.Y(n_129)
);

NAND2xp33_ASAP7_75t_SL g140 ( 
.A(n_120),
.B(n_124),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_112),
.B(n_74),
.C(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_113),
.Y(n_123)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_104),
.A2(n_61),
.B1(n_65),
.B2(n_51),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_110),
.A2(n_72),
.B1(n_68),
.B2(n_22),
.Y(n_126)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_100),
.B(n_18),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_128),
.Y(n_136)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_132),
.Y(n_150)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_125),
.B(n_103),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_134),
.B(n_129),
.C(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_135),
.A2(n_117),
.B(n_118),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_141),
.B(n_144),
.C(n_146),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_148),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_111),
.C(n_107),
.Y(n_146)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_105),
.B(n_2),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_147),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_150),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_152),
.B(n_154),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_142),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_145),
.B(n_24),
.C(n_41),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_28),
.B(n_40),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_159),
.C(n_158),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_153),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_160),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g161 ( 
.A(n_158),
.B(n_151),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_162),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_161),
.C(n_153),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_155),
.C(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_149),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_166),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_168),
.B(n_23),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_19),
.B(n_30),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_170),
.A2(n_17),
.B(n_29),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_171),
.A2(n_130),
.B1(n_11),
.B2(n_39),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_8),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_173),
.A2(n_6),
.B1(n_25),
.B2(n_37),
.Y(n_174)
);


endmodule