module fake_netlist_1_3950_n_537 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_537);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_537;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_357;
wire n_90;
wire n_245;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_159;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_99;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_71), .Y(n_76) );
CKINVDCx5p33_ASAP7_75t_R g77 ( .A(n_17), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_34), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_18), .Y(n_79) );
CKINVDCx16_ASAP7_75t_R g80 ( .A(n_44), .Y(n_80) );
INVx2_ASAP7_75t_L g81 ( .A(n_17), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_65), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_64), .Y(n_84) );
INVx3_ASAP7_75t_L g85 ( .A(n_50), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_25), .Y(n_86) );
INVxp33_ASAP7_75t_SL g87 ( .A(n_13), .Y(n_87) );
BUFx3_ASAP7_75t_L g88 ( .A(n_8), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_58), .Y(n_89) );
BUFx2_ASAP7_75t_L g90 ( .A(n_18), .Y(n_90) );
CKINVDCx16_ASAP7_75t_R g91 ( .A(n_30), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_70), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_43), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_37), .Y(n_94) );
INVx2_ASAP7_75t_L g95 ( .A(n_68), .Y(n_95) );
INVx1_ASAP7_75t_SL g96 ( .A(n_15), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_48), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_5), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_10), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_23), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_16), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_5), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_74), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_26), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_63), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_19), .Y(n_106) );
INVxp33_ASAP7_75t_L g107 ( .A(n_57), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_59), .Y(n_109) );
CKINVDCx14_ASAP7_75t_R g110 ( .A(n_60), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_88), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_85), .B(n_0), .Y(n_112) );
NOR2x1_ASAP7_75t_L g113 ( .A(n_88), .B(n_0), .Y(n_113) );
AND2x2_ASAP7_75t_SL g114 ( .A(n_80), .B(n_35), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_80), .Y(n_115) );
AND2x4_ASAP7_75t_L g116 ( .A(n_85), .B(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_88), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_85), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_85), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_84), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_102), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_102), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_91), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g124 ( .A(n_90), .B(n_1), .Y(n_124) );
NAND2xp5_ASAP7_75t_SL g125 ( .A(n_91), .B(n_2), .Y(n_125) );
CKINVDCx16_ASAP7_75t_R g126 ( .A(n_110), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_84), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_90), .B(n_2), .Y(n_128) );
CKINVDCx20_ASAP7_75t_R g129 ( .A(n_109), .Y(n_129) );
NOR2xp67_ASAP7_75t_L g130 ( .A(n_103), .B(n_3), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_84), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_95), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_129), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_118), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g136 ( .A(n_122), .B(n_107), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_122), .B(n_107), .Y(n_137) );
CKINVDCx16_ASAP7_75t_R g138 ( .A(n_126), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_118), .Y(n_139) );
INVx4_ASAP7_75t_L g140 ( .A(n_112), .Y(n_140) );
BUFx8_ASAP7_75t_SL g141 ( .A(n_123), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_119), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_119), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_126), .B(n_103), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_122), .B(n_76), .Y(n_145) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_114), .B(n_94), .Y(n_146) );
NAND2xp33_ASAP7_75t_R g147 ( .A(n_115), .B(n_87), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_119), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_118), .Y(n_149) );
INVx2_ASAP7_75t_SL g150 ( .A(n_112), .Y(n_150) );
BUFx6f_ASAP7_75t_SL g151 ( .A(n_114), .Y(n_151) );
INVxp67_ASAP7_75t_SL g152 ( .A(n_124), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_128), .B(n_110), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_118), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_118), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_122), .B(n_76), .Y(n_156) );
AND2x2_ASAP7_75t_L g157 ( .A(n_128), .B(n_102), .Y(n_157) );
AND2x6_ASAP7_75t_L g158 ( .A(n_112), .B(n_78), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_132), .Y(n_159) );
CKINVDCx5p33_ASAP7_75t_R g160 ( .A(n_141), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g161 ( .A(n_153), .B(n_114), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_142), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g163 ( .A1(n_145), .A2(n_112), .B(n_116), .C(n_117), .Y(n_163) );
NOR2xp67_ASAP7_75t_L g164 ( .A(n_146), .B(n_116), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g165 ( .A(n_138), .Y(n_165) );
NOR2xp33_ASAP7_75t_R g166 ( .A(n_138), .B(n_128), .Y(n_166) );
BUFx8_ASAP7_75t_L g167 ( .A(n_151), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_153), .B(n_116), .Y(n_168) );
AOI22xp33_ASAP7_75t_L g169 ( .A1(n_151), .A2(n_116), .B1(n_125), .B2(n_124), .Y(n_169) );
AOI22xp33_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_113), .B1(n_118), .B2(n_117), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_142), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_158), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
INVx2_ASAP7_75t_SL g174 ( .A(n_153), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_140), .B(n_130), .Y(n_176) );
NAND3xp33_ASAP7_75t_SL g177 ( .A(n_134), .B(n_77), .C(n_108), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_152), .B(n_130), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_144), .B(n_104), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_148), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_157), .B(n_113), .Y(n_182) );
INVx6_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
A2O1A1Ixp33_ASAP7_75t_L g185 ( .A1(n_145), .A2(n_111), .B(n_121), .C(n_131), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_157), .B(n_79), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_136), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_140), .Y(n_189) );
INVx5_ASAP7_75t_L g190 ( .A(n_158), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_157), .B(n_111), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_140), .Y(n_192) );
NOR2xp67_ASAP7_75t_L g193 ( .A(n_156), .B(n_121), .Y(n_193) );
BUFx2_ASAP7_75t_L g194 ( .A(n_184), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_175), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_183), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_188), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_174), .B(n_136), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_181), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_181), .Y(n_200) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
BUFx10_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_191), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_165), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_168), .A2(n_150), .B(n_140), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_172), .Y(n_206) );
NAND2x1_ASAP7_75t_L g207 ( .A(n_183), .B(n_158), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_189), .Y(n_208) );
BUFx8_ASAP7_75t_L g209 ( .A(n_172), .Y(n_209) );
AND2x2_ASAP7_75t_L g210 ( .A(n_174), .B(n_137), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_190), .B(n_150), .Y(n_211) );
AO32x2_ASAP7_75t_L g212 ( .A1(n_185), .A2(n_150), .A3(n_151), .B1(n_158), .B2(n_132), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_165), .Y(n_213) );
AND2x6_ASAP7_75t_L g214 ( .A(n_172), .B(n_158), .Y(n_214) );
NAND2x1p5_ASAP7_75t_L g215 ( .A(n_184), .B(n_137), .Y(n_215) );
BUFx12f_ASAP7_75t_L g216 ( .A(n_160), .Y(n_216) );
AND2x6_ASAP7_75t_L g217 ( .A(n_172), .B(n_158), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_187), .Y(n_218) );
OAI21x1_ASAP7_75t_L g219 ( .A1(n_162), .A2(n_156), .B(n_135), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_189), .Y(n_220) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_161), .A2(n_158), .B1(n_101), .B2(n_79), .Y(n_221) );
INVx1_ASAP7_75t_SL g222 ( .A(n_187), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_182), .B(n_158), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_163), .A2(n_131), .B(n_133), .C(n_127), .Y(n_224) );
INVxp67_ASAP7_75t_L g225 ( .A(n_187), .Y(n_225) );
INVx6_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_224), .A2(n_164), .B(n_178), .C(n_193), .Y(n_227) );
AOI22xp5_ASAP7_75t_L g228 ( .A1(n_197), .A2(n_147), .B1(n_179), .B2(n_169), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_209), .Y(n_229) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_219), .A2(n_176), .B(n_170), .Y(n_230) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_224), .A2(n_182), .B(n_192), .C(n_180), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_199), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g233 ( .A1(n_218), .A2(n_171), .B1(n_162), .B2(n_180), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_203), .B(n_187), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_210), .B(n_190), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_209), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_199), .Y(n_237) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_219), .A2(n_192), .B(n_173), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_213), .Y(n_239) );
INVx2_ASAP7_75t_L g240 ( .A(n_200), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_200), .Y(n_241) );
OAI21x1_ASAP7_75t_SL g242 ( .A1(n_221), .A2(n_171), .B(n_186), .Y(n_242) );
OR2x6_ASAP7_75t_L g243 ( .A(n_207), .B(n_167), .Y(n_243) );
OAI21x1_ASAP7_75t_L g244 ( .A1(n_205), .A2(n_186), .B(n_173), .Y(n_244) );
NAND2x1p5_ASAP7_75t_L g245 ( .A(n_206), .B(n_190), .Y(n_245) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_211), .A2(n_133), .B(n_120), .Y(n_246) );
AOI221xp5_ASAP7_75t_L g247 ( .A1(n_225), .A2(n_177), .B1(n_160), .B2(n_96), .C(n_99), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_210), .B(n_167), .Y(n_248) );
OAI21x1_ASAP7_75t_L g249 ( .A1(n_211), .A2(n_215), .B(n_139), .Y(n_249) );
AND2x4_ASAP7_75t_L g250 ( .A(n_195), .B(n_190), .Y(n_250) );
AND2x4_ASAP7_75t_L g251 ( .A(n_208), .B(n_190), .Y(n_251) );
OAI22xp5_ASAP7_75t_SL g252 ( .A1(n_201), .A2(n_216), .B1(n_204), .B2(n_222), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_234), .A2(n_198), .B1(n_215), .B2(n_223), .Y(n_253) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_232), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_232), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_238), .A2(n_206), .B(n_220), .Y(n_257) );
BUFx8_ASAP7_75t_L g258 ( .A(n_229), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_234), .B(n_228), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_227), .A2(n_206), .B(n_196), .Y(n_260) );
AOI221xp5_ASAP7_75t_L g261 ( .A1(n_247), .A2(n_96), .B1(n_106), .B2(n_99), .C(n_101), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_237), .Y(n_262) );
AOI22xp33_ASAP7_75t_L g263 ( .A1(n_248), .A2(n_167), .B1(n_216), .B2(n_196), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_237), .Y(n_264) );
AOI22xp33_ASAP7_75t_L g265 ( .A1(n_252), .A2(n_167), .B1(n_194), .B2(n_214), .Y(n_265) );
NAND4xp25_ASAP7_75t_L g266 ( .A(n_231), .B(n_147), .C(n_106), .D(n_98), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_240), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_240), .B(n_209), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_242), .A2(n_206), .B(n_154), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g270 ( .A1(n_236), .A2(n_217), .B1(n_214), .B2(n_194), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_241), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g272 ( .A1(n_239), .A2(n_235), .B1(n_236), .B2(n_243), .Y(n_272) );
AND2x4_ASAP7_75t_L g273 ( .A(n_236), .B(n_214), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_254), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_255), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_271), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_255), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_256), .B(n_241), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_256), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_262), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_271), .Y(n_281) );
AND2x2_ASAP7_75t_L g282 ( .A(n_262), .B(n_212), .Y(n_282) );
AO31x2_ASAP7_75t_L g283 ( .A1(n_257), .A2(n_233), .A3(n_133), .B(n_131), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_264), .Y(n_284) );
AND2x2_ASAP7_75t_L g285 ( .A(n_267), .B(n_212), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_259), .B(n_212), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_268), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_269), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_253), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_272), .B(n_212), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_273), .B(n_212), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_273), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_260), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_243), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_273), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_282), .B(n_78), .Y(n_296) );
HB1xp67_ASAP7_75t_L g297 ( .A(n_276), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_276), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_281), .Y(n_299) );
AND2x4_ASAP7_75t_L g300 ( .A(n_292), .B(n_249), .Y(n_300) );
AND2x2_ASAP7_75t_L g301 ( .A(n_282), .B(n_82), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_278), .B(n_82), .Y(n_302) );
OR2x2_ASAP7_75t_L g303 ( .A(n_275), .B(n_265), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_275), .Y(n_304) );
AND2x2_ASAP7_75t_L g305 ( .A(n_278), .B(n_83), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_283), .Y(n_307) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_294), .B(n_270), .Y(n_308) );
AND2x4_ASAP7_75t_SL g309 ( .A(n_292), .B(n_243), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_277), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_277), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_279), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_279), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_285), .B(n_83), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_280), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_285), .B(n_86), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_286), .B(n_86), .Y(n_317) );
AND2x2_ASAP7_75t_L g318 ( .A(n_291), .B(n_89), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_288), .Y(n_319) );
OAI33xp33_ASAP7_75t_L g320 ( .A1(n_287), .A2(n_97), .A3(n_89), .B1(n_92), .B2(n_93), .B3(n_105), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_280), .B(n_263), .Y(n_321) );
INVx2_ASAP7_75t_SL g322 ( .A(n_292), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_284), .Y(n_323) );
NAND3xp33_ASAP7_75t_L g324 ( .A(n_288), .B(n_258), .C(n_261), .Y(n_324) );
AND2x4_ASAP7_75t_L g325 ( .A(n_291), .B(n_249), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_286), .B(n_290), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_323), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_318), .B(n_284), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_304), .Y(n_329) );
NOR4xp25_ASAP7_75t_SL g330 ( .A(n_323), .B(n_287), .C(n_258), .D(n_293), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_326), .B(n_289), .Y(n_331) );
AOI322xp5_ASAP7_75t_L g332 ( .A1(n_318), .A2(n_274), .A3(n_81), .B1(n_98), .B2(n_290), .C1(n_289), .C2(n_93), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_326), .B(n_283), .Y(n_333) );
AND2x2_ASAP7_75t_L g334 ( .A(n_325), .B(n_283), .Y(n_334) );
NOR2x1_ASAP7_75t_L g335 ( .A(n_324), .B(n_294), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_325), .B(n_283), .Y(n_336) );
AND2x2_ASAP7_75t_L g337 ( .A(n_325), .B(n_283), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_283), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_325), .B(n_293), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_297), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_302), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_304), .B(n_295), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_319), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_310), .B(n_295), .Y(n_344) );
AOI211xp5_ASAP7_75t_L g345 ( .A1(n_324), .A2(n_81), .B(n_98), .C(n_105), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_302), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_319), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_310), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_311), .B(n_81), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
OR2x2_ASAP7_75t_L g351 ( .A(n_311), .B(n_120), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_312), .B(n_95), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_321), .B(n_258), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_305), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_317), .B(n_92), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_298), .Y(n_357) );
NOR3xp33_ASAP7_75t_L g358 ( .A(n_320), .B(n_97), .C(n_120), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_312), .B(n_313), .Y(n_359) );
CKINVDCx5p33_ASAP7_75t_R g360 ( .A(n_309), .Y(n_360) );
NAND2xp67_ASAP7_75t_L g361 ( .A(n_309), .B(n_127), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
OAI33xp33_ASAP7_75t_L g363 ( .A1(n_321), .A2(n_127), .A3(n_4), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_317), .B(n_3), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_313), .B(n_132), .Y(n_365) );
AND2x4_ASAP7_75t_SL g366 ( .A(n_298), .B(n_243), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_315), .B(n_132), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_322), .B(n_243), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_315), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_322), .B(n_132), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_322), .B(n_132), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_331), .B(n_308), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_331), .B(n_308), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_346), .B(n_308), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_359), .B(n_296), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_359), .Y(n_376) );
XNOR2x2_ASAP7_75t_L g377 ( .A(n_335), .B(n_303), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_340), .B(n_299), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_329), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_317), .A3(n_296), .B1(n_301), .B2(n_314), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_329), .Y(n_381) );
OR2x2_ASAP7_75t_L g382 ( .A(n_333), .B(n_341), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_327), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_333), .B(n_299), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_354), .B(n_296), .Y(n_385) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_354), .B(n_301), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_350), .B(n_299), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_339), .B(n_307), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
NAND2x1p5_ASAP7_75t_L g390 ( .A(n_368), .B(n_306), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_369), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_342), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_344), .Y(n_395) );
INVxp33_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
NAND2xp33_ASAP7_75t_L g397 ( .A(n_360), .B(n_303), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_344), .B(n_301), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_352), .B(n_314), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_352), .B(n_314), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_360), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_339), .B(n_307), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_334), .B(n_316), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_328), .B(n_306), .Y(n_404) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_330), .A2(n_320), .B(n_306), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_357), .B(n_316), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_356), .B(n_316), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_332), .B(n_300), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_364), .B(n_4), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_349), .B(n_300), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_349), .B(n_300), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_365), .Y(n_412) );
INVx1_ASAP7_75t_SL g413 ( .A(n_366), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_365), .Y(n_414) );
OAI32xp33_ASAP7_75t_L g415 ( .A1(n_338), .A2(n_104), .A3(n_309), .B1(n_9), .B2(n_10), .Y(n_415) );
AOI211xp5_ASAP7_75t_SL g416 ( .A1(n_368), .A2(n_300), .B(n_242), .C(n_235), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_367), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_334), .B(n_6), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_343), .B(n_7), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_343), .B(n_9), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_366), .Y(n_421) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_367), .A2(n_11), .B(n_12), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_338), .B(n_11), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_388), .B(n_336), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_376), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_393), .B(n_336), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_383), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g428 ( .A1(n_380), .A2(n_368), .B(n_337), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g429 ( .A(n_409), .B(n_423), .C(n_386), .D(n_418), .Y(n_429) );
NOR2xp33_ASAP7_75t_L g430 ( .A(n_396), .B(n_363), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g431 ( .A1(n_401), .A2(n_351), .B1(n_337), .B2(n_355), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_389), .Y(n_432) );
AOI322xp5_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_372), .A3(n_373), .B1(n_385), .B2(n_374), .C1(n_407), .C2(n_375), .Y(n_433) );
AOI32xp33_ASAP7_75t_L g434 ( .A1(n_416), .A2(n_358), .A3(n_370), .B1(n_371), .B2(n_361), .Y(n_434) );
NOR2x1_ASAP7_75t_L g435 ( .A(n_405), .B(n_351), .Y(n_435) );
OAI21xp5_ASAP7_75t_L g436 ( .A1(n_422), .A2(n_371), .B(n_370), .Y(n_436) );
OAI322xp33_ASAP7_75t_L g437 ( .A1(n_377), .A2(n_362), .A3(n_347), .B1(n_355), .B2(n_361), .C1(n_16), .C2(n_19), .Y(n_437) );
OAI322xp33_ASAP7_75t_L g438 ( .A1(n_382), .A2(n_362), .A3(n_347), .B1(n_14), .B2(n_15), .C1(n_20), .C2(n_13), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_388), .B(n_402), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_391), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_402), .B(n_12), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_379), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_394), .B(n_20), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_381), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_403), .B(n_244), .Y(n_445) );
AOI32xp33_ASAP7_75t_L g446 ( .A1(n_416), .A2(n_235), .A3(n_250), .B1(n_251), .B2(n_230), .Y(n_446) );
AOI322xp5_ASAP7_75t_L g447 ( .A1(n_375), .A2(n_235), .A3(n_250), .B1(n_251), .B2(n_100), .C1(n_159), .C2(n_149), .Y(n_447) );
OAI22xp33_ASAP7_75t_L g448 ( .A1(n_413), .A2(n_246), .B1(n_245), .B2(n_250), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_415), .A2(n_159), .B1(n_250), .B2(n_149), .C(n_135), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_408), .A2(n_244), .B1(n_230), .B2(n_251), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_395), .B(n_159), .Y(n_452) );
INVxp67_ASAP7_75t_SL g453 ( .A(n_378), .Y(n_453) );
OAI22xp5_ASAP7_75t_L g454 ( .A1(n_413), .A2(n_246), .B1(n_251), .B2(n_245), .Y(n_454) );
XNOR2xp5_ASAP7_75t_L g455 ( .A(n_421), .B(n_245), .Y(n_455) );
INVxp67_ASAP7_75t_L g456 ( .A(n_387), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_406), .Y(n_457) );
OAI21xp33_ASAP7_75t_L g458 ( .A1(n_398), .A2(n_159), .B(n_155), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_384), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_398), .B(n_159), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g461 ( .A1(n_422), .A2(n_217), .B(n_214), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_419), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_419), .Y(n_463) );
AOI22xp5_ASAP7_75t_L g464 ( .A1(n_399), .A2(n_159), .B1(n_217), .B2(n_214), .Y(n_464) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_399), .A2(n_159), .B1(n_217), .B2(n_214), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_390), .B(n_21), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_412), .B(n_155), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_433), .B(n_417), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_462), .B(n_414), .Y(n_469) );
INVxp67_ASAP7_75t_L g470 ( .A(n_430), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_427), .Y(n_471) );
AOI32xp33_ASAP7_75t_L g472 ( .A1(n_441), .A2(n_400), .A3(n_420), .B1(n_410), .B2(n_411), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_428), .A2(n_390), .B1(n_400), .B2(n_420), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_432), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_446), .B(n_392), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_440), .Y(n_476) );
OAI21xp5_ASAP7_75t_L g477 ( .A1(n_428), .A2(n_217), .B(n_155), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_442), .Y(n_478) );
BUFx2_ASAP7_75t_SL g479 ( .A(n_453), .Y(n_479) );
OAI211xp5_ASAP7_75t_L g480 ( .A1(n_429), .A2(n_154), .B(n_139), .C(n_135), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_444), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_439), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_463), .B(n_22), .Y(n_483) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_435), .A2(n_217), .B(n_154), .Y(n_484) );
NOR2xp33_ASAP7_75t_L g485 ( .A(n_429), .B(n_24), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_450), .Y(n_486) );
NOR3xp33_ASAP7_75t_L g487 ( .A(n_437), .B(n_139), .C(n_29), .Y(n_487) );
OAI221xp5_ASAP7_75t_L g488 ( .A1(n_434), .A2(n_226), .B1(n_183), .B2(n_32), .C(n_33), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_425), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_457), .B(n_28), .Y(n_490) );
O2A1O1Ixp5_ASAP7_75t_L g491 ( .A1(n_438), .A2(n_31), .B(n_36), .C(n_38), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_431), .B(n_202), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_426), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_456), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g495 ( .A1(n_443), .A2(n_39), .B1(n_40), .B2(n_41), .C(n_42), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g496 ( .A1(n_424), .A2(n_226), .B1(n_202), .B2(n_183), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_470), .A2(n_459), .B(n_445), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_479), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_473), .A2(n_455), .B1(n_436), .B2(n_451), .Y(n_499) );
AOI21xp33_ASAP7_75t_L g500 ( .A1(n_485), .A2(n_460), .B(n_452), .Y(n_500) );
XNOR2x1_ASAP7_75t_L g501 ( .A(n_468), .B(n_436), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_478), .Y(n_502) );
NAND2xp33_ASAP7_75t_L g503 ( .A(n_477), .B(n_461), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_471), .Y(n_504) );
BUFx2_ASAP7_75t_L g505 ( .A(n_482), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_481), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_485), .A2(n_447), .B(n_461), .C(n_449), .Y(n_507) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_480), .A2(n_458), .B(n_466), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_475), .A2(n_448), .B(n_454), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_474), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_476), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_472), .A2(n_467), .B1(n_465), .B2(n_464), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_494), .B(n_45), .Y(n_513) );
AO22x1_ASAP7_75t_SL g514 ( .A1(n_498), .A2(n_486), .B1(n_493), .B2(n_489), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_505), .A2(n_475), .B(n_491), .Y(n_515) );
OAI211xp5_ASAP7_75t_L g516 ( .A1(n_509), .A2(n_488), .B(n_487), .C(n_490), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g517 ( .A1(n_499), .A2(n_469), .B1(n_492), .B2(n_490), .C(n_483), .Y(n_517) );
OAI21xp5_ASAP7_75t_L g518 ( .A1(n_501), .A2(n_484), .B(n_495), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_503), .A2(n_496), .B(n_47), .Y(n_519) );
OAI22xp33_ASAP7_75t_SL g520 ( .A1(n_504), .A2(n_226), .B1(n_49), .B2(n_51), .Y(n_520) );
OAI22xp33_ASAP7_75t_SL g521 ( .A1(n_504), .A2(n_502), .B1(n_506), .B2(n_511), .Y(n_521) );
OAI211xp5_ASAP7_75t_SL g522 ( .A1(n_507), .A2(n_46), .B(n_52), .C(n_53), .Y(n_522) );
NAND2xp33_ASAP7_75t_L g523 ( .A(n_515), .B(n_497), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g524 ( .A1(n_516), .A2(n_513), .B(n_500), .C(n_508), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_521), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_517), .B(n_510), .Y(n_526) );
NAND4xp75_ASAP7_75t_L g527 ( .A(n_518), .B(n_513), .C(n_512), .D(n_56), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_526), .B(n_519), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_525), .A2(n_514), .B1(n_520), .B2(n_522), .Y(n_529) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_524), .B(n_54), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_528), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_530), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_531), .Y(n_533) );
AOI222xp33_ASAP7_75t_SL g534 ( .A1(n_533), .A2(n_532), .B1(n_529), .B2(n_523), .C1(n_527), .C2(n_67), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_534), .Y(n_535) );
AOI322xp5_ASAP7_75t_L g536 ( .A1(n_535), .A2(n_55), .A3(n_61), .B1(n_62), .B2(n_66), .C1(n_69), .C2(n_72), .Y(n_536) );
AOI221xp5_ASAP7_75t_L g537 ( .A1(n_536), .A2(n_73), .B1(n_75), .B2(n_226), .C(n_202), .Y(n_537) );
endmodule