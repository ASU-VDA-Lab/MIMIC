module fake_jpeg_13759_n_146 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_146);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_146;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_61),
.A2(n_49),
.B1(n_52),
.B2(n_45),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_63),
.A2(n_61),
.B1(n_60),
.B2(n_53),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_65),
.Y(n_74)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_50),
.Y(n_73)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_71),
.Y(n_84)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_72),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_50),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_77),
.A2(n_64),
.B1(n_62),
.B2(n_58),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_83),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_57),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_82),
.B(n_1),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_54),
.Y(n_83)
);

BUFx10_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_73),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_43),
.Y(n_111)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g116 ( 
.A(n_88),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_78),
.B(n_46),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_90),
.C(n_99),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_82),
.B(n_59),
.C(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_56),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_93),
.B(n_97),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_94),
.Y(n_106)
);

AND2x6_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_24),
.Y(n_95)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_18),
.A3(n_21),
.B1(n_25),
.B2(n_26),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_96),
.A2(n_8),
.B(n_10),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_0),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_22),
.C(n_41),
.Y(n_99)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_100),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_75),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_6),
.B(n_7),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_107)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_107),
.B(n_110),
.C(n_114),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_93),
.B(n_7),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_109),
.B(n_115),
.Y(n_124)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_32),
.B(n_34),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_11),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_118),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_97),
.B(n_14),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_16),
.Y(n_115)
);

XOR2x1_ASAP7_75t_L g117 ( 
.A(n_102),
.B(n_17),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_117),
.B(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_92),
.B(n_27),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_29),
.C(n_31),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_129),
.C(n_112),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_104),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_105),
.B(n_36),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_128),
.B(n_130),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_38),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g131 ( 
.A1(n_117),
.A2(n_40),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_128),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_133),
.B(n_134),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_126),
.Y(n_137)
);

MAJx2_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_138),
.C(n_136),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_132),
.A2(n_127),
.B(n_131),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_139),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_124),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_135),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_143),
.A2(n_107),
.B(n_123),
.C(n_122),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_116),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_145),
.B(n_112),
.Y(n_146)
);


endmodule