module fake_jpeg_13755_n_254 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_254);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_254;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_228;
wire n_178;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

BUFx4f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_1),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_46),
.Y(n_47)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_15),
.B(n_9),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_51),
.B(n_56),
.Y(n_95)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_52),
.Y(n_98)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_16),
.Y(n_53)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_53),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_20),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_16),
.B(n_4),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_17),
.B(n_4),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_60),
.B(n_61),
.Y(n_100)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_26),
.B(n_10),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_75),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_64),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_65),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_70),
.Y(n_132)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_71),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_37),
.Y(n_72)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_72),
.Y(n_134)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_37),
.Y(n_74)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_74),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_17),
.B(n_4),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_78),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_27),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_79),
.B(n_81),
.Y(n_120)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

BUFx4f_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_32),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_46),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_85),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_86),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g85 ( 
.A(n_39),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_46),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_87),
.B(n_90),
.Y(n_127)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_89),
.Y(n_123)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_19),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_25),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_32),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_21),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_56),
.A2(n_41),
.B1(n_22),
.B2(n_28),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_97),
.A2(n_95),
.B1(n_117),
.B2(n_106),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_51),
.B(n_36),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_102),
.B(n_111),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_62),
.B(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_28),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_117),
.B(n_124),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_41),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_128),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_21),
.Y(n_125)
);

NOR2x1_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_65),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_77),
.B(n_29),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_78),
.B(n_29),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_131),
.B(n_133),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_38),
.Y(n_133)
);

AOI32xp33_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_47),
.A3(n_81),
.B1(n_69),
.B2(n_48),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_138),
.B(n_144),
.Y(n_188)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_94),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_95),
.B(n_38),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_141),
.B(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_82),
.C(n_25),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_145),
.B(n_150),
.Y(n_181)
);

BUFx16f_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_146),
.B(n_153),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_95),
.B(n_123),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_123),
.C(n_100),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_148),
.B(n_152),
.Y(n_191)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_130),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_133),
.Y(n_150)
);

AO21x1_ASAP7_75t_L g151 ( 
.A1(n_100),
.A2(n_122),
.B(n_124),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_112),
.B(n_119),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_121),
.Y(n_154)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_101),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_155),
.A2(n_165),
.B(n_167),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_106),
.B(n_99),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_156),
.B(n_159),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_92),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_169),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_115),
.B1(n_104),
.B2(n_116),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_158),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_127),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_103),
.A2(n_105),
.B1(n_109),
.B2(n_129),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_94),
.A2(n_126),
.B1(n_136),
.B2(n_107),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_162),
.A2(n_173),
.B1(n_167),
.B2(n_174),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_93),
.B(n_96),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_163),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_98),
.B(n_126),
.C(n_136),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_164),
.A2(n_168),
.B(n_173),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_134),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_135),
.Y(n_166)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_166),
.Y(n_199)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_122),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_123),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_170),
.B(n_171),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_128),
.B(n_131),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_114),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_161),
.B(n_165),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_182),
.A2(n_187),
.B1(n_192),
.B2(n_196),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_147),
.A2(n_151),
.B1(n_169),
.B2(n_148),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_157),
.A2(n_168),
.B1(n_144),
.B2(n_141),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_195),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_142),
.B1(n_164),
.B2(n_137),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_174),
.B1(n_149),
.B2(n_145),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_139),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_193),
.B(n_198),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_200),
.B(n_203),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_177),
.B(n_155),
.Y(n_201)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_201),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_172),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_205),
.Y(n_219)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_199),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_140),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_210),
.Y(n_227)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_207),
.Y(n_220)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_208),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_165),
.B(n_146),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_209),
.B(n_213),
.C(n_195),
.Y(n_226)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_184),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_211),
.A2(n_214),
.B1(n_215),
.B2(n_186),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_197),
.B1(n_185),
.B2(n_189),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_146),
.B(n_181),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_179),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

NOR4xp25_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_198),
.C(n_180),
.D(n_190),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_217),
.B(n_226),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_202),
.A2(n_185),
.B1(n_180),
.B2(n_190),
.Y(n_218)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_218),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_221),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_212),
.Y(n_229)
);

MAJx2_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_192),
.C(n_194),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_231),
.C(n_234),
.Y(n_236)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_229),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_194),
.C(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_183),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_232),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_188),
.C(n_201),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_235),
.A2(n_216),
.B1(n_178),
.B2(n_220),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_237),
.B(n_239),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_231),
.B(n_201),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_238),
.B(n_234),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_233),
.B(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_240),
.B(n_219),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_243),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_245),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_241),
.B(n_227),
.Y(n_245)
);

OAI31xp33_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_230),
.A3(n_228),
.B(n_239),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_246),
.B(n_236),
.C(n_238),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_248),
.B(n_244),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_249),
.B(n_250),
.Y(n_251)
);

AOI21x1_ASAP7_75t_SL g252 ( 
.A1(n_251),
.A2(n_247),
.B(n_209),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_252),
.A2(n_226),
.B(n_216),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_236),
.Y(n_254)
);


endmodule