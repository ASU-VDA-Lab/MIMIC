module fake_aes_3225_n_46 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_46);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_46;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx1_ASAP7_75t_L g16 ( .A(n_3), .Y(n_16) );
CKINVDCx5p33_ASAP7_75t_R g17 ( .A(n_3), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_6), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_5), .Y(n_19) );
INVx2_ASAP7_75t_L g20 ( .A(n_8), .Y(n_20) );
NOR2x1_ASAP7_75t_L g21 ( .A(n_11), .B(n_15), .Y(n_21) );
CKINVDCx20_ASAP7_75t_R g22 ( .A(n_2), .Y(n_22) );
INVx2_ASAP7_75t_L g23 ( .A(n_20), .Y(n_23) );
OR2x2_ASAP7_75t_SL g24 ( .A(n_16), .B(n_0), .Y(n_24) );
INVxp67_ASAP7_75t_L g25 ( .A(n_18), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_17), .Y(n_26) );
OAI21xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_20), .B(n_21), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_25), .B(n_17), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_26), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
NAND4xp25_ASAP7_75t_SL g31 ( .A(n_29), .B(n_22), .C(n_24), .D(n_27), .Y(n_31) );
OAI33xp33_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_23), .A3(n_19), .B1(n_28), .B2(n_4), .B3(n_5), .Y(n_32) );
AOI221xp5_ASAP7_75t_L g33 ( .A1(n_31), .A2(n_29), .B1(n_30), .B2(n_19), .C(n_4), .Y(n_33) );
OAI21xp33_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_29), .B(n_1), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_34), .Y(n_35) );
OAI322xp33_ASAP7_75t_SL g36 ( .A1(n_33), .A2(n_0), .A3(n_1), .B1(n_2), .B2(n_6), .C1(n_7), .C2(n_9), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
NOR2x1_ASAP7_75t_L g38 ( .A(n_35), .B(n_7), .Y(n_38) );
INVx1_ASAP7_75t_SL g39 ( .A(n_35), .Y(n_39) );
OAI221xp5_ASAP7_75t_L g40 ( .A1(n_37), .A2(n_10), .B1(n_12), .B2(n_13), .C(n_14), .Y(n_40) );
INVx1_ASAP7_75t_L g41 ( .A(n_39), .Y(n_41) );
INVx3_ASAP7_75t_L g42 ( .A(n_38), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_40), .Y(n_43) );
OAI22xp5_ASAP7_75t_L g44 ( .A1(n_42), .A2(n_36), .B1(n_43), .B2(n_41), .Y(n_44) );
BUFx2_ASAP7_75t_L g45 ( .A(n_41), .Y(n_45) );
NAND3xp33_ASAP7_75t_L g46 ( .A(n_44), .B(n_42), .C(n_45), .Y(n_46) );
endmodule