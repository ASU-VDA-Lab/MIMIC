module real_jpeg_31215_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_237;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_0),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_0),
.B(n_92),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_1),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_2),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_2),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_2),
.B(n_75),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_2),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_2),
.Y(n_220)
);

NAND2x1_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_3),
.B(n_62),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_3),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_3),
.B(n_24),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_4),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_4),
.B(n_55),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_6),
.Y(n_122)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_7),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g74 ( 
.A(n_8),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_8),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_8),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_8),
.B(n_140),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_8),
.B(n_176),
.Y(n_175)
);

NAND2xp33_ASAP7_75t_R g40 ( 
.A(n_9),
.B(n_41),
.Y(n_40)
);

AO22x1_ASAP7_75t_L g51 ( 
.A1(n_9),
.A2(n_13),
.B1(n_41),
.B2(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_9),
.B(n_99),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_9),
.B(n_117),
.Y(n_116)
);

NAND2x1_ASAP7_75t_L g159 ( 
.A(n_9),
.B(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_9),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_10),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_12),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_12),
.B(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_12),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_12),
.B(n_194),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_12),
.B(n_205),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_14),
.Y(n_69)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_14),
.Y(n_107)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_14),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_146),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_143),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_124),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_19),
.B(n_124),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_38),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_29),
.C(n_33),
.Y(n_21)
);

XNOR2x2_ASAP7_75t_L g128 ( 
.A(n_22),
.B(n_129),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_25),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_23),
.B(n_25),
.Y(n_131)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_28),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_28),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_29),
.B(n_34),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_56),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_51),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_45),
.Y(n_115)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_55),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_55),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_60)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_63),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_68),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_108),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_88),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_78),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B1(n_86),
.B2(n_87),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_82),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_95),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_123)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.C(n_104),
.Y(n_97)
);

XNOR2x1_ASAP7_75t_SL g110 ( 
.A(n_98),
.B(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_110),
.Y(n_109)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_111),
.C(n_123),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g127 ( 
.A(n_111),
.B(n_123),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_116),
.C(n_119),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_112),
.A2(n_113),
.B1(n_119),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_183),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_119),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_130),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_126),
.B(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_128),
.B(n_130),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.C(n_137),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_131),
.B(n_132),
.Y(n_186)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_135),
.Y(n_161)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_137),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

AO22x1_ASAP7_75t_SL g167 ( 
.A1(n_138),
.A2(n_139),
.B1(n_142),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_142),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_237),
.B(n_242),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_187),
.B(n_236),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_179),
.Y(n_149)
);

NOR2xp67_ASAP7_75t_L g236 ( 
.A(n_150),
.B(n_179),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_165),
.B(n_178),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_152),
.B(n_199),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_158),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_162),
.C(n_164),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_155),
.Y(n_153)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_155),
.Y(n_197)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_158)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_159),
.Y(n_164)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_170),
.A2(n_171),
.B1(n_174),
.B2(n_175),
.Y(n_191)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx4f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_185),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_181),
.B(n_185),
.C(n_239),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_182),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_200),
.B(n_235),
.Y(n_187)
);

NOR2xp67_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_198),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_198),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_192),
.C(n_196),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_190),
.A2(n_191),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_L g234 ( 
.A(n_190),
.B(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_191),
.B(n_215),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_196),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_217),
.B(n_232),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_214),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_202),
.A2(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_208),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_204),
.B1(n_208),
.B2(n_209),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_226),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_225),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_219),
.A2(n_225),
.B(n_227),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_220),
.B(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp33_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_240),
.Y(n_242)
);


endmodule