module real_aes_15501_n_282 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_282);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_282;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_1199;
wire n_951;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_877;
wire n_424;
wire n_802;
wire n_1488;
wire n_337;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_580;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_334;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_769;
wire n_434;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_1457;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_1064;
wire n_540;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_516;
wire n_335;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_1097;
wire n_703;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_0), .A2(n_205), .B1(n_433), .B2(n_1053), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1071 ( .A1(n_0), .A2(n_65), .B1(n_355), .B2(n_1072), .Y(n_1071) );
AOI22xp33_ASAP7_75t_L g1279 ( .A1(n_1), .A2(n_4), .B1(n_1241), .B2(n_1244), .Y(n_1279) );
INVx1_ASAP7_75t_L g572 ( .A(n_2), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_2), .A2(n_102), .B1(n_433), .B2(n_593), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g662 ( .A1(n_3), .A2(n_663), .B(n_666), .C(n_677), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_3), .B(n_315), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1488 ( .A1(n_5), .A2(n_262), .B1(n_574), .B2(n_983), .Y(n_1488) );
INVxp33_ASAP7_75t_SL g1532 ( .A(n_5), .Y(n_1532) );
AOI22xp33_ASAP7_75t_SL g485 ( .A1(n_6), .A2(n_144), .B1(n_366), .B2(n_486), .Y(n_485) );
INVxp67_ASAP7_75t_SL g536 ( .A(n_6), .Y(n_536) );
INVx1_ASAP7_75t_L g1444 ( .A(n_7), .Y(n_1444) );
INVx1_ASAP7_75t_L g1062 ( .A(n_8), .Y(n_1062) );
OAI22xp33_ASAP7_75t_L g1078 ( .A1(n_8), .A2(n_69), .B1(n_496), .B2(n_708), .Y(n_1078) );
AOI22xp33_ASAP7_75t_L g891 ( .A1(n_9), .A2(n_77), .B1(n_695), .B2(n_892), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_9), .A2(n_53), .B1(n_912), .B2(n_913), .Y(n_911) );
INVx1_ASAP7_75t_L g745 ( .A(n_10), .Y(n_745) );
AO22x1_ASAP7_75t_L g784 ( .A1(n_10), .A2(n_142), .B1(n_418), .B2(n_673), .Y(n_784) );
INVx1_ASAP7_75t_L g296 ( .A(n_11), .Y(n_296) );
AND2x2_ASAP7_75t_L g347 ( .A(n_11), .B(n_230), .Y(n_347) );
AND2x2_ASAP7_75t_L g408 ( .A(n_11), .B(n_409), .Y(n_408) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_11), .B(n_306), .Y(n_782) );
INVx1_ASAP7_75t_L g757 ( .A(n_12), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_12), .A2(n_100), .B1(n_423), .B2(n_669), .Y(n_783) );
INVx1_ASAP7_75t_L g1192 ( .A(n_13), .Y(n_1192) );
OAI221xp5_ASAP7_75t_L g1205 ( .A1(n_13), .A2(n_155), .B1(n_627), .B2(n_1206), .C(n_1207), .Y(n_1205) );
INVx2_ASAP7_75t_L g1237 ( .A(n_14), .Y(n_1237) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_14), .B(n_109), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_14), .B(n_1243), .Y(n_1245) );
CKINVDCx5p33_ASAP7_75t_R g1011 ( .A(n_15), .Y(n_1011) );
XNOR2xp5_ASAP7_75t_L g612 ( .A(n_16), .B(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g1017 ( .A(n_17), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g1257 ( .A1(n_18), .A2(n_235), .B1(n_1241), .B2(n_1244), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g1450 ( .A1(n_19), .A2(n_46), .B1(n_381), .B2(n_1451), .Y(n_1450) );
AOI22xp33_ASAP7_75t_L g1460 ( .A1(n_19), .A2(n_279), .B1(n_608), .B2(n_912), .Y(n_1460) );
INVx1_ASAP7_75t_L g598 ( .A(n_20), .Y(n_598) );
AOI22xp33_ASAP7_75t_SL g573 ( .A1(n_21), .A2(n_75), .B1(n_366), .B2(n_574), .Y(n_573) );
AOI221xp5_ASAP7_75t_L g591 ( .A1(n_21), .A2(n_276), .B1(n_426), .B2(n_427), .C(n_515), .Y(n_591) );
INVx1_ASAP7_75t_L g949 ( .A(n_22), .Y(n_949) );
OAI22xp33_ASAP7_75t_L g972 ( .A1(n_22), .A2(n_169), .B1(n_496), .B2(n_973), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g957 ( .A1(n_23), .A2(n_55), .B1(n_524), .B2(n_527), .C(n_958), .Y(n_957) );
INVx1_ASAP7_75t_L g986 ( .A(n_23), .Y(n_986) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_24), .A2(n_153), .B1(n_370), .B2(n_375), .Y(n_369) );
AOI221xp5_ASAP7_75t_L g440 ( .A1(n_24), .A2(n_229), .B1(n_441), .B2(n_445), .C(n_449), .Y(n_440) );
INVx1_ASAP7_75t_L g597 ( .A(n_25), .Y(n_597) );
OAI211xp5_ASAP7_75t_L g678 ( .A1(n_26), .A2(n_679), .B(n_680), .C(n_681), .Y(n_678) );
INVx1_ASAP7_75t_L g721 ( .A(n_26), .Y(n_721) );
INVx1_ASAP7_75t_L g1442 ( .A(n_27), .Y(n_1442) );
OAI221xp5_ASAP7_75t_L g1462 ( .A1(n_27), .A2(n_138), .B1(n_524), .B2(n_1206), .C(n_1463), .Y(n_1462) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_28), .A2(n_97), .B1(n_315), .B2(n_559), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_29), .A2(n_276), .B1(n_366), .B2(n_574), .Y(n_583) );
AOI22xp33_ASAP7_75t_SL g607 ( .A1(n_29), .A2(n_75), .B1(n_439), .B2(n_608), .Y(n_607) );
OAI22xp5_ASAP7_75t_L g1136 ( .A1(n_30), .A2(n_267), .B1(n_1137), .B2(n_1141), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g1175 ( .A1(n_30), .A2(n_267), .B1(n_1176), .B2(n_1179), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g1249 ( .A1(n_31), .A2(n_265), .B1(n_1234), .B2(n_1250), .Y(n_1249) );
AOI22xp33_ASAP7_75t_SL g1199 ( .A1(n_32), .A2(n_91), .B1(n_389), .B2(n_859), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g1217 ( .A1(n_32), .A2(n_161), .B1(n_427), .B2(n_441), .C(n_545), .Y(n_1217) );
NAND2xp5_ASAP7_75t_SL g842 ( .A(n_33), .B(n_422), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_33), .A2(n_157), .B1(n_389), .B2(n_866), .Y(n_865) );
XNOR2xp5_ASAP7_75t_L g1433 ( .A(n_34), .B(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g410 ( .A(n_35), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_36), .A2(n_157), .B1(n_418), .B2(n_595), .Y(n_846) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_36), .A2(n_250), .B1(n_389), .B2(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g1048 ( .A(n_37), .Y(n_1048) );
AOI22xp33_ASAP7_75t_SL g1448 ( .A1(n_38), .A2(n_279), .B1(n_1077), .B2(n_1449), .Y(n_1448) );
AOI221xp5_ASAP7_75t_L g1467 ( .A1(n_38), .A2(n_46), .B1(n_669), .B2(n_671), .C(n_1468), .Y(n_1467) );
AOI22xp33_ASAP7_75t_L g1493 ( .A1(n_39), .A2(n_113), .B1(n_1494), .B2(n_1495), .Y(n_1493) );
INVx1_ASAP7_75t_L g1542 ( .A(n_39), .Y(n_1542) );
AOI22xp5_ASAP7_75t_L g1269 ( .A1(n_40), .A2(n_247), .B1(n_1241), .B2(n_1244), .Y(n_1269) );
AO22x1_ASAP7_75t_L g1254 ( .A1(n_41), .A2(n_60), .B1(n_1234), .B2(n_1238), .Y(n_1254) );
AOI21xp33_ASAP7_75t_L g633 ( .A1(n_42), .A2(n_426), .B(n_449), .Y(n_633) );
INVx1_ASAP7_75t_L g641 ( .A(n_42), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_43), .A2(n_229), .B1(n_370), .B2(n_381), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g429 ( .A1(n_43), .A2(n_153), .B1(n_430), .B2(n_432), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_44), .A2(n_66), .B1(n_595), .B2(n_622), .Y(n_667) );
AOI22xp33_ASAP7_75t_SL g693 ( .A1(n_44), .A2(n_273), .B1(n_366), .B2(n_574), .Y(n_693) );
AOI22xp33_ASAP7_75t_SL g896 ( .A1(n_45), .A2(n_127), .B1(n_897), .B2(n_898), .Y(n_896) );
INVxp67_ASAP7_75t_SL g927 ( .A(n_45), .Y(n_927) );
INVx1_ASAP7_75t_L g322 ( .A(n_47), .Y(n_322) );
INVx1_ASAP7_75t_L g339 ( .A(n_47), .Y(n_339) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_48), .A2(n_124), .B1(n_366), .B2(n_389), .Y(n_388) );
AOI221xp5_ASAP7_75t_L g421 ( .A1(n_48), .A2(n_73), .B1(n_422), .B2(n_425), .C(n_427), .Y(n_421) );
INVx1_ASAP7_75t_L g557 ( .A(n_49), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_50), .A2(n_198), .B1(n_430), .B2(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g642 ( .A(n_50), .Y(n_642) );
INVx1_ASAP7_75t_L g827 ( .A(n_51), .Y(n_827) );
INVxp67_ASAP7_75t_SL g940 ( .A(n_52), .Y(n_940) );
AND4x1_ASAP7_75t_L g989 ( .A(n_52), .B(n_942), .C(n_945), .D(n_970), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_53), .A2(n_133), .B1(n_491), .B2(n_695), .Y(n_893) );
INVx1_ASAP7_75t_L g1445 ( .A(n_54), .Y(n_1445) );
INVx1_ASAP7_75t_L g988 ( .A(n_55), .Y(n_988) );
INVx1_ASAP7_75t_L g289 ( .A(n_56), .Y(n_289) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_57), .A2(n_239), .B1(n_427), .B2(n_618), .C(n_619), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_57), .A2(n_275), .B1(n_355), .B2(n_366), .Y(n_643) );
INVx2_ASAP7_75t_L g325 ( .A(n_58), .Y(n_325) );
INVx1_ASAP7_75t_L g816 ( .A(n_59), .Y(n_816) );
OAI22xp33_ASAP7_75t_L g1508 ( .A1(n_61), .A2(n_228), .B1(n_1509), .B2(n_1510), .Y(n_1508) );
OAI22xp5_ASAP7_75t_L g1523 ( .A1(n_61), .A2(n_228), .B1(n_1524), .B2(n_1526), .Y(n_1523) );
CKINVDCx5p33_ASAP7_75t_R g1437 ( .A(n_62), .Y(n_1437) );
INVx1_ASAP7_75t_L g902 ( .A(n_63), .Y(n_902) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_64), .A2(n_179), .B1(n_1234), .B2(n_1238), .Y(n_1270) );
AOI221xp5_ASAP7_75t_L g1056 ( .A1(n_65), .A2(n_196), .B1(n_427), .B2(n_515), .C(n_1057), .Y(n_1056) );
AOI22xp33_ASAP7_75t_SL g698 ( .A1(n_66), .A2(n_99), .B1(n_366), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g1491 ( .A(n_67), .Y(n_1491) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_68), .A2(n_71), .B1(n_366), .B2(n_368), .Y(n_494) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_68), .A2(n_144), .B1(n_425), .B2(n_513), .C(n_516), .Y(n_512) );
INVx1_ASAP7_75t_L g1061 ( .A(n_69), .Y(n_1061) );
AO221x2_ASAP7_75t_L g1311 ( .A1(n_70), .A2(n_218), .B1(n_1241), .B2(n_1244), .C(n_1312), .Y(n_1311) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_71), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g487 ( .A1(n_72), .A2(n_185), .B1(n_488), .B2(n_491), .Y(n_487) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_72), .A2(n_128), .B1(n_430), .B2(n_432), .Y(n_517) );
AOI22xp33_ASAP7_75t_SL g365 ( .A1(n_73), .A2(n_223), .B1(n_366), .B2(n_368), .Y(n_365) );
INVx1_ASAP7_75t_L g868 ( .A(n_74), .Y(n_868) );
AOI22xp33_ASAP7_75t_SL g1002 ( .A1(n_76), .A2(n_183), .B1(n_389), .B2(n_889), .Y(n_1002) );
AOI22xp33_ASAP7_75t_SL g1035 ( .A1(n_76), .A2(n_241), .B1(n_430), .B2(n_608), .Y(n_1035) );
INVx1_ASAP7_75t_L g924 ( .A(n_77), .Y(n_924) );
INVx1_ASAP7_75t_L g1505 ( .A(n_78), .Y(n_1505) );
AOI21xp33_ASAP7_75t_L g1051 ( .A1(n_79), .A2(n_449), .B(n_619), .Y(n_1051) );
AOI22xp33_ASAP7_75t_L g1073 ( .A1(n_79), .A2(n_171), .B1(n_492), .B2(n_710), .Y(n_1073) );
OAI22xp5_ASAP7_75t_L g1438 ( .A1(n_80), .A2(n_215), .B1(n_461), .B2(n_507), .Y(n_1438) );
OAI211xp5_ASAP7_75t_L g1455 ( .A1(n_80), .A2(n_589), .B(n_1456), .C(n_1461), .Y(n_1455) );
OAI22xp33_ASAP7_75t_L g495 ( .A1(n_81), .A2(n_264), .B1(n_496), .B2(n_502), .Y(n_495) );
INVx1_ASAP7_75t_L g520 ( .A(n_81), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_82), .A2(n_172), .B1(n_381), .B2(n_752), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1216 ( .A1(n_82), .A2(n_90), .B1(n_913), .B2(n_1053), .Y(n_1216) );
OAI22xp5_ASAP7_75t_L g944 ( .A1(n_83), .A2(n_209), .B1(n_461), .B2(n_507), .Y(n_944) );
OAI211xp5_ASAP7_75t_L g946 ( .A1(n_83), .A2(n_510), .B(n_947), .C(n_950), .Y(n_946) );
OAI222xp33_ASAP7_75t_L g768 ( .A1(n_84), .A2(n_206), .B1(n_769), .B2(n_771), .C1(n_773), .C2(n_775), .Y(n_768) );
INVx1_ASAP7_75t_L g788 ( .A(n_84), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g1046 ( .A1(n_85), .A2(n_524), .B(n_1047), .C(n_1049), .Y(n_1046) );
INVx1_ASAP7_75t_L g1069 ( .A(n_85), .Y(n_1069) );
INVx1_ASAP7_75t_L g882 ( .A(n_86), .Y(n_882) );
OAI222xp33_ASAP7_75t_L g916 ( .A1(n_86), .A2(n_123), .B1(n_527), .B2(n_917), .C1(n_918), .C2(n_925), .Y(n_916) );
OAI22xp5_ASAP7_75t_SL g835 ( .A1(n_87), .A2(n_104), .B1(n_836), .B2(n_837), .Y(n_835) );
OAI21xp33_ASAP7_75t_L g848 ( .A1(n_87), .A2(n_708), .B(n_849), .Y(n_848) );
CKINVDCx5p33_ASAP7_75t_R g1094 ( .A(n_88), .Y(n_1094) );
INVx1_ASAP7_75t_L g332 ( .A(n_89), .Y(n_332) );
AOI22xp33_ASAP7_75t_L g1197 ( .A1(n_90), .A2(n_110), .B1(n_381), .B2(n_488), .Y(n_1197) );
INVxp67_ASAP7_75t_SL g1209 ( .A(n_91), .Y(n_1209) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_92), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g956 ( .A1(n_93), .A2(n_271), .B1(n_608), .B2(n_673), .Y(n_956) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_93), .A2(n_114), .B1(n_381), .B2(n_978), .Y(n_980) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_94), .Y(n_291) );
AND2x2_ASAP7_75t_L g1235 ( .A(n_94), .B(n_289), .Y(n_1235) );
AOI22xp33_ASAP7_75t_SL g1003 ( .A1(n_95), .A2(n_281), .B1(n_1004), .B2(n_1006), .Y(n_1003) );
AOI21xp33_ASAP7_75t_L g1032 ( .A1(n_95), .A2(n_606), .B(n_1033), .Y(n_1032) );
CKINVDCx5p33_ASAP7_75t_R g734 ( .A(n_96), .Y(n_734) );
OAI211xp5_ASAP7_75t_SL g1054 ( .A1(n_97), .A2(n_510), .B(n_1055), .C(n_1060), .Y(n_1054) );
CKINVDCx5p33_ASAP7_75t_R g629 ( .A(n_98), .Y(n_629) );
AOI221xp5_ASAP7_75t_SL g674 ( .A1(n_99), .A2(n_273), .B1(n_423), .B2(n_675), .C(n_676), .Y(n_674) );
INVx1_ASAP7_75t_L g753 ( .A(n_100), .Y(n_753) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_101), .Y(n_579) );
INVx1_ASAP7_75t_L g582 ( .A(n_102), .Y(n_582) );
OAI211xp5_ASAP7_75t_L g829 ( .A1(n_103), .A2(n_830), .B(n_831), .C(n_832), .Y(n_829) );
INVxp33_ASAP7_75t_SL g850 ( .A(n_103), .Y(n_850) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_104), .Y(n_872) );
CKINVDCx5p33_ASAP7_75t_R g877 ( .A(n_105), .Y(n_877) );
INVxp67_ASAP7_75t_SL g966 ( .A(n_106), .Y(n_966) );
AOI22xp33_ASAP7_75t_SL g982 ( .A1(n_106), .A2(n_211), .B1(n_983), .B2(n_984), .Y(n_982) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_107), .Y(n_685) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_108), .A2(n_261), .B1(n_502), .B2(n_1019), .Y(n_1018) );
INVx1_ASAP7_75t_L g1027 ( .A(n_108), .Y(n_1027) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_109), .B(n_1237), .Y(n_1236) );
INVx1_ASAP7_75t_L g1243 ( .A(n_109), .Y(n_1243) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_110), .A2(n_172), .B1(n_606), .B2(n_1211), .C(n_1212), .Y(n_1210) );
OAI22xp33_ASAP7_75t_L g1200 ( .A1(n_111), .A2(n_166), .B1(n_502), .B2(n_1019), .Y(n_1200) );
INVx1_ASAP7_75t_L g1220 ( .A(n_111), .Y(n_1220) );
CKINVDCx5p33_ASAP7_75t_R g943 ( .A(n_112), .Y(n_943) );
INVx1_ASAP7_75t_L g1534 ( .A(n_113), .Y(n_1534) );
AOI221xp5_ASAP7_75t_L g967 ( .A1(n_114), .A2(n_222), .B1(n_606), .B2(n_669), .C(n_968), .Y(n_967) );
INVx1_ASAP7_75t_L g567 ( .A(n_115), .Y(n_567) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_115), .A2(n_426), .B(n_606), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g1106 ( .A(n_116), .Y(n_1106) );
INVx2_ASAP7_75t_L g327 ( .A(n_117), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_117), .B(n_325), .Y(n_342) );
INVx1_ASAP7_75t_L g387 ( .A(n_117), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_118), .A2(n_212), .B1(n_1234), .B2(n_1238), .Y(n_1278) );
OAI22xp33_ASAP7_75t_L g1146 ( .A1(n_119), .A2(n_174), .B1(n_1147), .B2(n_1148), .Y(n_1146) );
OAI22xp33_ASAP7_75t_L g1154 ( .A1(n_119), .A2(n_174), .B1(n_1155), .B2(n_1158), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_120), .A2(n_135), .B1(n_679), .B2(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g705 ( .A(n_120), .Y(n_705) );
INVx1_ASAP7_75t_L g763 ( .A(n_121), .Y(n_763) );
NAND2xp33_ASAP7_75t_SL g806 ( .A(n_121), .B(n_423), .Y(n_806) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_122), .A2(n_231), .B1(n_507), .B2(n_559), .Y(n_558) );
OAI211xp5_ASAP7_75t_L g588 ( .A1(n_122), .A2(n_589), .B(n_590), .C(n_596), .Y(n_588) );
INVx1_ASAP7_75t_L g881 ( .A(n_123), .Y(n_881) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_124), .A2(n_223), .B1(n_432), .B2(n_439), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g1095 ( .A(n_125), .Y(n_1095) );
OAI211xp5_ASAP7_75t_SL g1124 ( .A1(n_126), .A2(n_1117), .B(n_1125), .C(n_1128), .Y(n_1124) );
INVx1_ASAP7_75t_L g1174 ( .A(n_126), .Y(n_1174) );
AOI221xp5_ASAP7_75t_L g910 ( .A1(n_127), .A2(n_268), .B1(n_516), .B2(n_543), .C(n_545), .Y(n_910) );
AOI22xp33_ASAP7_75t_SL g493 ( .A1(n_128), .A2(n_243), .B1(n_488), .B2(n_491), .Y(n_493) );
XOR2x2_ASAP7_75t_L g1186 ( .A(n_129), .B(n_1187), .Y(n_1186) );
AOI22xp33_ASAP7_75t_SL g1453 ( .A1(n_130), .A2(n_148), .B1(n_368), .B2(n_1072), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1457 ( .A1(n_130), .A2(n_178), .B1(n_516), .B2(n_952), .C(n_1458), .Y(n_1457) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_131), .Y(n_1102) );
INVx1_ASAP7_75t_L g625 ( .A(n_132), .Y(n_625) );
INVx1_ASAP7_75t_L g920 ( .A(n_133), .Y(n_920) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_134), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1021 ( .A1(n_134), .A2(n_589), .B(n_1022), .C(n_1026), .Y(n_1021) );
INVx1_ASAP7_75t_L g719 ( .A(n_135), .Y(n_719) );
AOI22xp33_ASAP7_75t_SL g1007 ( .A1(n_136), .A2(n_256), .B1(n_1004), .B2(n_1006), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1024 ( .A1(n_136), .A2(n_281), .B1(n_433), .B2(n_1025), .Y(n_1024) );
INVx1_ASAP7_75t_L g1485 ( .A(n_137), .Y(n_1485) );
INVx1_ASAP7_75t_L g1441 ( .A(n_138), .Y(n_1441) );
CKINVDCx16_ASAP7_75t_R g770 ( .A(n_139), .Y(n_770) );
NAND5xp2_ASAP7_75t_L g660 ( .A(n_140), .B(n_661), .C(n_691), .D(n_706), .E(n_716), .Y(n_660) );
INVx1_ASAP7_75t_L g725 ( .A(n_140), .Y(n_725) );
AOI22xp33_ASAP7_75t_SL g634 ( .A1(n_141), .A2(n_275), .B1(n_418), .B2(n_439), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_141), .A2(n_239), .B1(n_366), .B2(n_647), .Y(n_646) );
AOI21xp5_ASAP7_75t_L g764 ( .A1(n_142), .A2(n_702), .B(n_765), .Y(n_764) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_143), .A2(n_168), .B1(n_461), .B2(n_507), .Y(n_506) );
OAI211xp5_ASAP7_75t_SL g509 ( .A1(n_143), .A2(n_510), .B(n_511), .C(n_518), .Y(n_509) );
INVx1_ASAP7_75t_L g810 ( .A(n_145), .Y(n_810) );
AO22x1_ASAP7_75t_L g1255 ( .A1(n_146), .A2(n_233), .B1(n_1241), .B2(n_1244), .Y(n_1255) );
INVx1_ASAP7_75t_L g624 ( .A(n_147), .Y(n_624) );
INVxp67_ASAP7_75t_SL g1466 ( .A(n_148), .Y(n_1466) );
INVx1_ASAP7_75t_L g997 ( .A(n_149), .Y(n_997) );
OAI221xp5_ASAP7_75t_L g1029 ( .A1(n_149), .A2(n_151), .B1(n_528), .B2(n_627), .C(n_1030), .Y(n_1029) );
BUFx3_ASAP7_75t_L g319 ( .A(n_150), .Y(n_319) );
INVx1_ASAP7_75t_L g998 ( .A(n_151), .Y(n_998) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_152), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_154), .A2(n_241), .B1(n_389), .B2(n_897), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g1023 ( .A1(n_154), .A2(n_183), .B1(n_426), .B2(n_427), .C(n_515), .Y(n_1023) );
INVx1_ASAP7_75t_L g1191 ( .A(n_155), .Y(n_1191) );
OAI22xp33_ASAP7_75t_L g1497 ( .A1(n_156), .A2(n_258), .B1(n_298), .B2(n_1498), .Y(n_1497) );
OAI22xp33_ASAP7_75t_L g1514 ( .A1(n_156), .A2(n_258), .B1(n_1515), .B2(n_1517), .Y(n_1514) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_158), .A2(n_173), .B1(n_1241), .B2(n_1244), .Y(n_1240) );
OAI21xp33_ASAP7_75t_L g900 ( .A1(n_159), .A2(n_461), .B(n_901), .Y(n_900) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_160), .Y(n_303) );
AOI22xp33_ASAP7_75t_SL g1194 ( .A1(n_161), .A2(n_237), .B1(n_368), .B2(n_1195), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_162), .A2(n_204), .B1(n_622), .B2(n_673), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_162), .A2(n_197), .B1(n_492), .B2(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g1492 ( .A(n_163), .Y(n_1492) );
CKINVDCx20_ASAP7_75t_R g391 ( .A(n_164), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g1132 ( .A(n_165), .Y(n_1132) );
INVx1_ASAP7_75t_L g1219 ( .A(n_166), .Y(n_1219) );
INVx1_ASAP7_75t_L g1507 ( .A(n_167), .Y(n_1507) );
OAI211xp5_ASAP7_75t_L g1518 ( .A1(n_167), .A2(n_1164), .B(n_1519), .C(n_1521), .Y(n_1518) );
INVx1_ASAP7_75t_L g948 ( .A(n_169), .Y(n_948) );
AOI22xp33_ASAP7_75t_SL g1447 ( .A1(n_170), .A2(n_178), .B1(n_366), .B2(n_898), .Y(n_1447) );
INVx1_ASAP7_75t_L g1465 ( .A(n_170), .Y(n_1465) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_171), .A2(n_254), .B1(n_433), .B2(n_1059), .Y(n_1058) );
INVx1_ASAP7_75t_L g903 ( .A(n_175), .Y(n_903) );
CKINVDCx5p33_ASAP7_75t_R g1091 ( .A(n_176), .Y(n_1091) );
INVx1_ASAP7_75t_L g736 ( .A(n_177), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_177), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g1258 ( .A1(n_180), .A2(n_246), .B1(n_1234), .B2(n_1238), .Y(n_1258) );
XOR2xp5_ASAP7_75t_L g476 ( .A(n_181), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g885 ( .A(n_182), .Y(n_885) );
OAI221xp5_ASAP7_75t_L g626 ( .A1(n_184), .A2(n_240), .B1(n_528), .B2(n_627), .C(n_628), .Y(n_626) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_184), .A2(n_240), .B1(n_393), .B2(n_585), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g542 ( .A1(n_185), .A2(n_243), .B1(n_543), .B2(n_545), .C(n_547), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g845 ( .A1(n_186), .A2(n_426), .B(n_671), .Y(n_845) );
INVx1_ASAP7_75t_L g855 ( .A(n_186), .Y(n_855) );
INVx1_ASAP7_75t_L g1133 ( .A(n_187), .Y(n_1133) );
OAI211xp5_ASAP7_75t_L g1161 ( .A1(n_187), .A2(n_1162), .B(n_1164), .C(n_1166), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g1083 ( .A(n_188), .B(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g715 ( .A(n_189), .Y(n_715) );
CKINVDCx5p33_ASAP7_75t_R g351 ( .A(n_190), .Y(n_351) );
INVxp67_ASAP7_75t_SL g962 ( .A(n_191), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g975 ( .A1(n_191), .A2(n_221), .B1(n_859), .B2(n_976), .Y(n_975) );
INVx1_ASAP7_75t_L g404 ( .A(n_192), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g1202 ( .A(n_193), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1233 ( .A1(n_194), .A2(n_242), .B1(n_1234), .B2(n_1238), .Y(n_1233) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_195), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_196), .A2(n_205), .B1(n_368), .B2(n_1072), .Y(n_1074) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_197), .A2(n_248), .B1(n_423), .B2(n_669), .C(n_671), .Y(n_668) );
INVx1_ASAP7_75t_L g645 ( .A(n_198), .Y(n_645) );
INVx1_ASAP7_75t_L g396 ( .A(n_199), .Y(n_396) );
XOR2x2_ASAP7_75t_L g822 ( .A(n_200), .B(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_201), .A2(n_259), .B1(n_418), .B2(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g857 ( .A(n_201), .Y(n_857) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_202), .Y(n_1050) );
AOI22xp33_ASAP7_75t_SL g1076 ( .A1(n_202), .A2(n_254), .B1(n_372), .B2(n_1077), .Y(n_1076) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_203), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g694 ( .A1(n_204), .A2(n_248), .B1(n_492), .B2(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_R g795 ( .A(n_206), .B(n_796), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_207), .B(n_993), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g1012 ( .A1(n_207), .A2(n_1013), .B1(n_1014), .B2(n_1036), .Y(n_1012) );
INVx1_ASAP7_75t_L g1038 ( .A(n_207), .Y(n_1038) );
AO22x1_ASAP7_75t_L g1288 ( .A1(n_208), .A2(n_236), .B1(n_1234), .B2(n_1289), .Y(n_1288) );
OA22x2_ASAP7_75t_L g1043 ( .A1(n_210), .A2(n_1044), .B1(n_1079), .B2(n_1080), .Y(n_1043) );
CKINVDCx16_ASAP7_75t_R g1079 ( .A(n_210), .Y(n_1079) );
AOI221xp5_ASAP7_75t_L g951 ( .A1(n_211), .A2(n_221), .B1(n_516), .B2(n_952), .C(n_954), .Y(n_951) );
OAI211xp5_ASAP7_75t_L g1499 ( .A1(n_213), .A2(n_1500), .B(n_1503), .C(n_1504), .Y(n_1499) );
INVx1_ASAP7_75t_L g1522 ( .A(n_213), .Y(n_1522) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_214), .A2(n_234), .B1(n_461), .B2(n_507), .Y(n_1203) );
CKINVDCx5p33_ASAP7_75t_R g1089 ( .A(n_216), .Y(n_1089) );
INVx1_ASAP7_75t_L g730 ( .A(n_217), .Y(n_730) );
INVx1_ASAP7_75t_L g481 ( .A(n_219), .Y(n_481) );
OAI221xp5_ASAP7_75t_SL g523 ( .A1(n_219), .A2(n_274), .B1(n_524), .B2(n_527), .C(n_532), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_220), .A2(n_277), .B1(n_507), .B2(n_559), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_222), .A2(n_271), .B1(n_381), .B2(n_978), .Y(n_977) );
AOI22xp33_ASAP7_75t_SL g888 ( .A1(n_224), .A2(n_268), .B1(n_647), .B2(n_889), .Y(n_888) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_224), .Y(n_926) );
INVx1_ASAP7_75t_L g651 ( .A(n_225), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g834 ( .A(n_226), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g1248 ( .A1(n_227), .A2(n_252), .B1(n_1241), .B2(n_1244), .Y(n_1248) );
BUFx3_ASAP7_75t_L g306 ( .A(n_230), .Y(n_306) );
INVx1_ASAP7_75t_L g409 ( .A(n_230), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g1314 ( .A(n_232), .Y(n_1314) );
OAI211xp5_ASAP7_75t_L g1214 ( .A1(n_234), .A2(n_589), .B(n_1215), .C(n_1218), .Y(n_1214) );
INVxp67_ASAP7_75t_SL g1208 ( .A(n_237), .Y(n_1208) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_238), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g1099 ( .A(n_244), .Y(n_1099) );
INVx1_ASAP7_75t_L g331 ( .A(n_245), .Y(n_331) );
INVx1_ASAP7_75t_L g345 ( .A(n_245), .Y(n_345) );
INVx2_ASAP7_75t_L g364 ( .A(n_245), .Y(n_364) );
INVx1_ASAP7_75t_L g747 ( .A(n_249), .Y(n_747) );
AOI22xp33_ASAP7_75t_L g805 ( .A1(n_249), .A2(n_280), .B1(n_622), .B2(n_673), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g839 ( .A(n_250), .B(n_426), .Y(n_839) );
AO22x1_ASAP7_75t_L g1290 ( .A1(n_251), .A2(n_269), .B1(n_1241), .B2(n_1244), .Y(n_1290) );
AOI22xp33_ASAP7_75t_L g1473 ( .A1(n_251), .A2(n_1474), .B1(n_1477), .B2(n_1548), .Y(n_1473) );
XNOR2x1_ASAP7_75t_L g1479 ( .A(n_251), .B(n_1480), .Y(n_1479) );
INVx1_ASAP7_75t_L g475 ( .A(n_253), .Y(n_475) );
INVx1_ASAP7_75t_L g1064 ( .A(n_255), .Y(n_1064) );
INVx1_ASAP7_75t_L g1031 ( .A(n_256), .Y(n_1031) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_257), .A2(n_461), .B(n_470), .Y(n_460) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_259), .Y(n_864) );
OAI22xp33_ASAP7_75t_SL g584 ( .A1(n_260), .A2(n_270), .B1(n_393), .B2(n_585), .Y(n_584) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_260), .A2(n_270), .B1(n_524), .B2(n_528), .C(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g1028 ( .A(n_261), .Y(n_1028) );
INVxp67_ASAP7_75t_SL g1541 ( .A(n_262), .Y(n_1541) );
XNOR2xp5_ASAP7_75t_L g554 ( .A(n_263), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g519 ( .A(n_264), .Y(n_519) );
INVx1_ASAP7_75t_L g930 ( .A(n_265), .Y(n_930) );
INVx1_ASAP7_75t_L g1487 ( .A(n_266), .Y(n_1487) );
CKINVDCx5p33_ASAP7_75t_R g833 ( .A(n_272), .Y(n_833) );
INVx1_ASAP7_75t_L g483 ( .A(n_274), .Y(n_483) );
OAI211xp5_ASAP7_75t_L g615 ( .A1(n_277), .A2(n_589), .B(n_616), .C(n_623), .Y(n_615) );
INVx1_ASAP7_75t_L g844 ( .A(n_278), .Y(n_844) );
INVx1_ASAP7_75t_L g759 ( .A(n_280), .Y(n_759) );
AOI21xp5_ASAP7_75t_L g282 ( .A1(n_283), .A2(n_307), .B(n_1225), .Y(n_282) );
BUFx4f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_292), .Y(n_285) );
NOR2xp33_ASAP7_75t_L g1476 ( .A(n_286), .B(n_295), .Y(n_1476) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_288), .B(n_290), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g1472 ( .A(n_288), .B(n_291), .Y(n_1472) );
INVx1_ASAP7_75t_L g1550 ( .A(n_288), .Y(n_1550) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g1553 ( .A(n_291), .B(n_1550), .Y(n_1553) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_294), .B(n_297), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x4_ASAP7_75t_L g1151 ( .A(n_295), .B(n_1152), .Y(n_1151) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x4_ASAP7_75t_L g428 ( .A(n_296), .B(n_306), .Y(n_428) );
AND2x4_ASAP7_75t_L g450 ( .A(n_296), .B(n_305), .Y(n_450) );
INVx1_ASAP7_75t_L g1147 ( .A(n_297), .Y(n_1147) );
AND2x4_ASAP7_75t_SL g1475 ( .A(n_297), .B(n_1476), .Y(n_1475) );
INVx3_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g298 ( .A(n_299), .B(n_304), .Y(n_298) );
OR2x6_ASAP7_75t_L g1139 ( .A(n_299), .B(n_1140), .Y(n_1139) );
BUFx4f_ASAP7_75t_L g1533 ( .A(n_299), .Y(n_1533) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
BUFx4f_ASAP7_75t_L g535 ( .A(n_300), .Y(n_535) );
INVx3_ASAP7_75t_L g961 ( .A(n_300), .Y(n_961) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx2_ASAP7_75t_L g349 ( .A(n_302), .Y(n_349) );
AND2x2_ASAP7_75t_L g414 ( .A(n_302), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g420 ( .A(n_302), .Y(n_420) );
AND2x2_ASAP7_75t_L g424 ( .A(n_302), .B(n_303), .Y(n_424) );
INVx1_ASAP7_75t_L g465 ( .A(n_302), .Y(n_465) );
NAND2x1_ASAP7_75t_L g604 ( .A(n_302), .B(n_303), .Y(n_604) );
INVx1_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx2_ASAP7_75t_L g415 ( .A(n_303), .Y(n_415) );
AND2x2_ASAP7_75t_L g419 ( .A(n_303), .B(n_420), .Y(n_419) );
BUFx2_ASAP7_75t_L g455 ( .A(n_303), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_303), .B(n_420), .Y(n_540) );
OR2x2_ASAP7_75t_L g804 ( .A(n_303), .B(n_349), .Y(n_804) );
INVxp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g1127 ( .A(n_305), .Y(n_1127) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
BUFx2_ASAP7_75t_L g1131 ( .A(n_306), .Y(n_1131) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_306), .B(n_464), .Y(n_1135) );
OAI22xp33_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_934), .B1(n_935), .B2(n_1224), .Y(n_307) );
INVx1_ASAP7_75t_L g1224 ( .A(n_308), .Y(n_1224) );
AO22x2_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_655), .B1(n_656), .B2(n_933), .Y(n_308) );
INVx1_ASAP7_75t_L g933 ( .A(n_309), .Y(n_933) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_552), .Y(n_309) );
XOR2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_476), .Y(n_310) );
XNOR2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_475), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_401), .Y(n_312) );
AOI221xp5_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_332), .B1(n_333), .B2(n_351), .C(n_352), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx5_ASAP7_75t_L g873 ( .A(n_315), .Y(n_873) );
OR2x6_ASAP7_75t_L g315 ( .A(n_316), .B(n_328), .Y(n_315) );
OR2x2_ASAP7_75t_L g507 ( .A(n_316), .B(n_328), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
INVx8_ASAP7_75t_L g367 ( .A(n_317), .Y(n_367) );
BUFx3_ASAP7_75t_L g765 ( .A(n_317), .Y(n_765) );
BUFx3_ASAP7_75t_L g859 ( .A(n_317), .Y(n_859) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_317), .Y(n_866) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
AND2x4_ASAP7_75t_L g373 ( .A(n_318), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g338 ( .A(n_319), .B(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g356 ( .A(n_319), .B(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
OR2x2_ASAP7_75t_L g499 ( .A(n_319), .B(n_321), .Y(n_499) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVxp67_ASAP7_75t_L g374 ( .A(n_322), .Y(n_374) );
AND2x4_ASAP7_75t_L g358 ( .A(n_323), .B(n_344), .Y(n_358) );
INVx1_ASAP7_75t_L g767 ( .A(n_323), .Y(n_767) );
AND2x6_ASAP7_75t_L g774 ( .A(n_323), .B(n_394), .Y(n_774) );
AND2x2_ASAP7_75t_L g776 ( .A(n_323), .B(n_400), .Y(n_776) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_326), .Y(n_323) );
NAND3x1_ASAP7_75t_L g385 ( .A(n_324), .B(n_386), .C(n_387), .Y(n_385) );
NAND2x1p5_ASAP7_75t_L g702 ( .A(n_324), .B(n_387), .Y(n_702) );
OR2x4_ASAP7_75t_L g1157 ( .A(n_324), .B(n_499), .Y(n_1157) );
INVx1_ASAP7_75t_L g1160 ( .A(n_324), .Y(n_1160) );
AND2x4_ASAP7_75t_L g1165 ( .A(n_324), .B(n_356), .Y(n_1165) );
OR2x6_ASAP7_75t_L g1180 ( .A(n_324), .B(n_571), .Y(n_1180) );
INVx3_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g362 ( .A(n_325), .Y(n_362) );
NAND2xp33_ASAP7_75t_SL g565 ( .A(n_325), .B(n_327), .Y(n_565) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND3x4_ASAP7_75t_L g361 ( .A(n_327), .B(n_362), .C(n_363), .Y(n_361) );
AND2x2_ASAP7_75t_L g754 ( .A(n_327), .B(n_362), .Y(n_754) );
HB1xp67_ASAP7_75t_L g1183 ( .A(n_327), .Y(n_1183) );
INVxp67_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g462 ( .A(n_329), .B(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g713 ( .A(n_329), .Y(n_713) );
OR2x2_ASAP7_75t_L g787 ( .A(n_329), .B(n_463), .Y(n_787) );
INVx1_ASAP7_75t_L g1152 ( .A(n_329), .Y(n_1152) );
BUFx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx2_ASAP7_75t_L g341 ( .A(n_330), .Y(n_341) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_332), .A2(n_417), .B1(n_421), .B2(n_429), .C(n_434), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_333), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_333), .A2(n_557), .B(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_333), .A2(n_651), .B(n_652), .Y(n_650) );
AOI211x1_ASAP7_75t_L g876 ( .A1(n_333), .A2(n_877), .B(n_878), .C(n_900), .Y(n_876) );
AOI21xp33_ASAP7_75t_L g942 ( .A1(n_333), .A2(n_943), .B(n_944), .Y(n_942) );
NAND2xp33_ASAP7_75t_L g1010 ( .A(n_333), .B(n_1011), .Y(n_1010) );
AOI21xp5_ASAP7_75t_L g1063 ( .A1(n_333), .A2(n_1064), .B(n_1065), .Y(n_1063) );
AOI21xp33_ASAP7_75t_SL g1201 ( .A1(n_333), .A2(n_1202), .B(n_1203), .Y(n_1201) );
AOI21xp5_ASAP7_75t_L g1436 ( .A1(n_333), .A2(n_1437), .B(n_1438), .Y(n_1436) );
INVx8_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_343), .Y(n_334) );
INVx1_ASAP7_75t_L g720 ( .A(n_335), .Y(n_720) );
OR2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_340), .Y(n_335) );
BUFx3_ASAP7_75t_L g863 ( .A(n_336), .Y(n_863) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_337), .Y(n_581) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
BUFx2_ASAP7_75t_L g571 ( .A(n_338), .Y(n_571) );
INVx2_ASAP7_75t_L g357 ( .A(n_339), .Y(n_357) );
INVx1_ASAP7_75t_L g469 ( .A(n_339), .Y(n_469) );
OR2x2_ASAP7_75t_L g466 ( .A(n_340), .B(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g473 ( .A(n_340), .Y(n_473) );
INVx1_ASAP7_75t_L g501 ( .A(n_340), .Y(n_501) );
OR2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
OR2x2_ASAP7_75t_L g564 ( .A(n_341), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_SL g800 ( .A(n_341), .B(n_428), .Y(n_800) );
INVx1_ASAP7_75t_L g1122 ( .A(n_341), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1185 ( .A(n_341), .Y(n_1185) );
INVx1_ASAP7_75t_L g741 ( .A(n_342), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_343), .B(n_818), .Y(n_817) );
OR2x2_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g386 ( .A(n_345), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_345), .B(n_408), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
AND2x6_ASAP7_75t_L g434 ( .A(n_347), .B(n_423), .Y(n_434) );
AND2x2_ASAP7_75t_L g453 ( .A(n_347), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_347), .B(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g531 ( .A(n_347), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g792 ( .A(n_347), .B(n_364), .Y(n_792) );
AND2x2_ASAP7_75t_L g407 ( .A(n_348), .B(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g431 ( .A(n_348), .Y(n_431) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_348), .Y(n_595) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_349), .Y(n_684) );
NAND3xp33_ASAP7_75t_SL g352 ( .A(n_353), .B(n_359), .C(n_390), .Y(n_352) );
INVx2_ASAP7_75t_SL g503 ( .A(n_353), .Y(n_503) );
AND5x1_ASAP7_75t_L g823 ( .A(n_353), .B(n_824), .C(n_851), .D(n_867), .E(n_871), .Y(n_823) );
AND4x1_ASAP7_75t_L g970 ( .A(n_353), .B(n_971), .C(n_974), .D(n_985), .Y(n_970) );
NAND4xp75_ASAP7_75t_L g1435 ( .A(n_353), .B(n_1436), .C(n_1439), .D(n_1454), .Y(n_1435) );
INVx3_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_354), .Y(n_561) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_354), .B(n_637), .C(n_649), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g703 ( .A1(n_354), .A2(n_586), .B1(n_682), .B2(n_704), .C(n_705), .Y(n_703) );
INVx3_ASAP7_75t_L g886 ( .A(n_354), .Y(n_886) );
NOR3xp33_ASAP7_75t_L g1066 ( .A(n_354), .B(n_1067), .C(n_1078), .Y(n_1066) );
AND2x4_ASAP7_75t_L g354 ( .A(n_355), .B(n_358), .Y(n_354) );
BUFx2_ASAP7_75t_L g486 ( .A(n_355), .Y(n_486) );
BUFx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx2_ASAP7_75t_L g368 ( .A(n_356), .Y(n_368) );
BUFx3_ASAP7_75t_L g389 ( .A(n_356), .Y(n_389) );
BUFx2_ASAP7_75t_L g574 ( .A(n_356), .Y(n_574) );
INVx2_ASAP7_75t_L g648 ( .A(n_356), .Y(n_648) );
BUFx2_ASAP7_75t_L g976 ( .A(n_356), .Y(n_976) );
BUFx2_ASAP7_75t_L g1495 ( .A(n_356), .Y(n_1495) );
INVx1_ASAP7_75t_L g379 ( .A(n_357), .Y(n_379) );
NAND2x1_ASAP7_75t_L g393 ( .A(n_358), .B(n_394), .Y(n_393) );
AND2x4_ASAP7_75t_L g397 ( .A(n_358), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g482 ( .A(n_358), .B(n_394), .Y(n_482) );
AND2x4_ASAP7_75t_SL g586 ( .A(n_358), .B(n_398), .Y(n_586) );
AND2x4_ASAP7_75t_SL g704 ( .A(n_358), .B(n_394), .Y(n_704) );
AND2x2_ASAP7_75t_L g987 ( .A(n_358), .B(n_394), .Y(n_987) );
AOI33xp33_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_365), .A3(n_369), .B1(n_380), .B2(n_382), .B3(n_388), .Y(n_359) );
AOI33xp33_ASAP7_75t_L g484 ( .A1(n_360), .A2(n_382), .A3(n_485), .B1(n_487), .B2(n_493), .B3(n_494), .Y(n_484) );
AOI33xp33_ASAP7_75t_L g887 ( .A1(n_360), .A2(n_888), .A3(n_891), .B1(n_893), .B2(n_894), .B3(n_896), .Y(n_887) );
AOI33xp33_ASAP7_75t_L g1446 ( .A1(n_360), .A2(n_1009), .A3(n_1447), .B1(n_1448), .B2(n_1450), .B3(n_1453), .Y(n_1446) );
BUFx3_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AOI33xp33_ASAP7_75t_L g692 ( .A1(n_361), .A2(n_693), .A3(n_694), .B1(n_696), .B2(n_698), .B3(n_700), .Y(n_692) );
AOI33xp33_ASAP7_75t_L g974 ( .A1(n_361), .A2(n_975), .A3(n_977), .B1(n_980), .B2(n_981), .B3(n_982), .Y(n_974) );
AOI33xp33_ASAP7_75t_L g1001 ( .A1(n_361), .A2(n_1002), .A3(n_1003), .B1(n_1007), .B2(n_1008), .B3(n_1009), .Y(n_1001) );
AOI33xp33_ASAP7_75t_L g1070 ( .A1(n_361), .A2(n_1071), .A3(n_1073), .B1(n_1074), .B2(n_1075), .B3(n_1076), .Y(n_1070) );
AOI33xp33_ASAP7_75t_L g1193 ( .A1(n_361), .A2(n_1009), .A3(n_1194), .B1(n_1197), .B2(n_1198), .B3(n_1199), .Y(n_1193) );
INVx3_ASAP7_75t_L g1169 ( .A(n_362), .Y(n_1169) );
INVx1_ASAP7_75t_L g551 ( .A(n_363), .Y(n_551) );
OAI31xp33_ASAP7_75t_L g737 ( .A1(n_363), .A2(n_738), .A3(n_742), .B(n_768), .Y(n_737) );
INVx2_ASAP7_75t_SL g1221 ( .A(n_363), .Y(n_1221) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g459 ( .A(n_364), .Y(n_459) );
BUFx2_ASAP7_75t_L g1494 ( .A(n_366), .Y(n_1494) );
INVx8_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_L g472 ( .A(n_367), .Y(n_472) );
INVx3_ASAP7_75t_L g897 ( .A(n_367), .Y(n_897) );
INVx1_ASAP7_75t_L g899 ( .A(n_368), .Y(n_899) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g474 ( .A(n_372), .B(n_473), .Y(n_474) );
INVx2_ASAP7_75t_SL g640 ( .A(n_372), .Y(n_640) );
HB1xp67_ASAP7_75t_L g1449 ( .A(n_372), .Y(n_1449) );
BUFx8_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g490 ( .A(n_373), .Y(n_490) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_373), .Y(n_578) );
BUFx6f_ASAP7_75t_L g752 ( .A(n_373), .Y(n_752) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g892 ( .A(n_376), .Y(n_892) );
INVx5_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g381 ( .A(n_377), .Y(n_381) );
BUFx12f_ASAP7_75t_L g492 ( .A(n_377), .Y(n_492) );
AND2x4_ASAP7_75t_L g819 ( .A(n_377), .B(n_741), .Y(n_819) );
BUFx2_ASAP7_75t_L g1006 ( .A(n_377), .Y(n_1006) );
BUFx3_ASAP7_75t_L g1077 ( .A(n_377), .Y(n_1077) );
AND2x4_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx2_ASAP7_75t_L g395 ( .A(n_378), .Y(n_395) );
NAND2x1p5_ASAP7_75t_L g468 ( .A(n_378), .B(n_469), .Y(n_468) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_378), .Y(n_1170) );
INVx1_ASAP7_75t_L g400 ( .A(n_379), .Y(n_400) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
OAI22xp5_ASAP7_75t_SL g637 ( .A1(n_383), .A2(n_638), .B1(n_639), .B2(n_644), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_384), .Y(n_383) );
INVx2_ASAP7_75t_L g575 ( .A(n_384), .Y(n_575) );
INVx2_ASAP7_75t_L g860 ( .A(n_384), .Y(n_860) );
INVx3_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g895 ( .A(n_385), .Y(n_895) );
AOI22xp33_ASAP7_75t_L g390 ( .A1(n_391), .A2(n_392), .B1(n_396), .B2(n_397), .Y(n_390) );
AOI222xp33_ASAP7_75t_L g435 ( .A1(n_391), .A2(n_396), .B1(n_436), .B2(n_438), .C1(n_440), .C2(n_451), .Y(n_435) );
AOI221x1_ASAP7_75t_L g851 ( .A1(n_392), .A2(n_397), .B1(n_827), .B2(n_833), .C(n_852), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_392), .A2(n_397), .B1(n_997), .B2(n_998), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_392), .A2(n_397), .B1(n_1191), .B2(n_1192), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1440 ( .A1(n_392), .A2(n_397), .B1(n_1441), .B2(n_1442), .Y(n_1440) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx3_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_397), .A2(n_481), .B1(n_482), .B2(n_483), .Y(n_480) );
AO22x1_ASAP7_75t_L g880 ( .A1(n_397), .A2(n_482), .B1(n_881), .B2(n_882), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g985 ( .A1(n_397), .A2(n_986), .B1(n_987), .B2(n_988), .Y(n_985) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_456), .B(n_460), .Y(n_401) );
NAND3xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_416), .C(n_435), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B1(n_410), .B2(n_411), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_404), .A2(n_410), .B1(n_471), .B2(n_474), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_405), .A2(n_519), .B1(n_520), .B2(n_521), .Y(n_518) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_406), .A2(n_412), .B1(n_597), .B2(n_598), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_406), .A2(n_411), .B1(n_948), .B2(n_949), .Y(n_947) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_406), .A2(n_412), .B1(n_1027), .B2(n_1028), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1461 ( .A1(n_406), .A2(n_412), .B1(n_1444), .B2(n_1445), .Y(n_1461) );
BUFx6f_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_407), .A2(n_412), .B1(n_624), .B2(n_625), .Y(n_623) );
AND2x4_ASAP7_75t_L g735 ( .A(n_407), .B(n_713), .Y(n_735) );
INVx1_ASAP7_75t_L g908 ( .A(n_407), .Y(n_908) );
AND2x4_ASAP7_75t_L g412 ( .A(n_408), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g417 ( .A(n_408), .B(n_418), .Y(n_417) );
AND2x4_ASAP7_75t_SL g437 ( .A(n_408), .B(n_423), .Y(n_437) );
AND2x2_ASAP7_75t_L g664 ( .A(n_408), .B(n_665), .Y(n_664) );
BUFx2_ASAP7_75t_L g687 ( .A(n_408), .Y(n_687) );
AND2x2_ASAP7_75t_L g714 ( .A(n_408), .B(n_413), .Y(n_714) );
HB1xp67_ASAP7_75t_L g1140 ( .A(n_409), .Y(n_1140) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_411), .A2(n_907), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1218 ( .A1(n_411), .A2(n_907), .B1(n_1219), .B2(n_1220), .Y(n_1218) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g522 ( .A(n_412), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g906 ( .A1(n_412), .A2(n_902), .B1(n_903), .B2(n_907), .Y(n_906) );
INVx2_ASAP7_75t_L g448 ( .A(n_413), .Y(n_448) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_413), .Y(n_546) );
INVx1_ASAP7_75t_L g620 ( .A(n_413), .Y(n_620) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g426 ( .A(n_414), .Y(n_426) );
INVx2_ASAP7_75t_L g670 ( .A(n_414), .Y(n_670) );
AND2x4_ASAP7_75t_L g1149 ( .A(n_414), .B(n_1140), .Y(n_1149) );
INVx3_ASAP7_75t_L g510 ( .A(n_417), .Y(n_510) );
INVx2_ASAP7_75t_SL g589 ( .A(n_417), .Y(n_589) );
NAND2xp5_ASAP7_75t_R g915 ( .A(n_417), .B(n_885), .Y(n_915) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
BUFx3_ASAP7_75t_L g433 ( .A(n_419), .Y(n_433) );
INVx2_ASAP7_75t_L g609 ( .A(n_419), .Y(n_609) );
BUFx3_ASAP7_75t_L g622 ( .A(n_419), .Y(n_622) );
BUFx3_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx6f_ASAP7_75t_L g515 ( .A(n_423), .Y(n_515) );
BUFx3_ASAP7_75t_L g618 ( .A(n_423), .Y(n_618) );
INVx1_ASAP7_75t_L g953 ( .A(n_423), .Y(n_953) );
AND2x2_ASAP7_75t_L g1126 ( .A(n_423), .B(n_1127), .Y(n_1126) );
BUFx3_ASAP7_75t_L g1211 ( .A(n_423), .Y(n_1211) );
BUFx6f_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g444 ( .A(n_424), .Y(n_444) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g1034 ( .A(n_426), .Y(n_1034) );
HB1xp67_ASAP7_75t_L g1057 ( .A(n_426), .Y(n_1057) );
INVx4_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
INVx1_ASAP7_75t_SL g516 ( .A(n_428), .Y(n_516) );
INVx4_ASAP7_75t_L g676 ( .A(n_428), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g838 ( .A(n_428), .B(n_839), .C(n_840), .D(n_842), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_428), .B(n_1121), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1547 ( .A(n_428), .B(n_1121), .Y(n_1547) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
INVx2_ASAP7_75t_SL g439 ( .A(n_431), .Y(n_439) );
INVx2_ASAP7_75t_L g673 ( .A(n_431), .Y(n_673) );
INVx1_ASAP7_75t_L g841 ( .A(n_431), .Y(n_841) );
INVx2_ASAP7_75t_L g912 ( .A(n_431), .Y(n_912) );
INVx1_ASAP7_75t_L g1053 ( .A(n_431), .Y(n_1053) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_SL g914 ( .A(n_433), .Y(n_914) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_434), .A2(n_512), .B(n_517), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_434), .A2(n_591), .B(n_592), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g616 ( .A1(n_434), .A2(n_617), .B(n_621), .Y(n_616) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_434), .A2(n_910), .B(n_911), .Y(n_909) );
AOI21xp5_ASAP7_75t_L g950 ( .A1(n_434), .A2(n_951), .B(n_956), .Y(n_950) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_434), .A2(n_1023), .B(n_1024), .Y(n_1022) );
AOI21xp5_ASAP7_75t_L g1055 ( .A1(n_434), .A2(n_1056), .B(n_1058), .Y(n_1055) );
AOI21xp5_ASAP7_75t_L g1215 ( .A1(n_434), .A2(n_1216), .B(n_1217), .Y(n_1215) );
AOI21xp5_ASAP7_75t_SL g1456 ( .A1(n_434), .A2(n_1457), .B(n_1460), .Y(n_1456) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_436), .B(n_827), .Y(n_826) );
BUFx3_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g526 ( .A(n_437), .Y(n_526) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
BUFx2_ASAP7_75t_L g544 ( .A(n_444), .Y(n_544) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g1213 ( .A(n_448), .Y(n_1213) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g547 ( .A(n_450), .Y(n_547) );
INVx2_ASAP7_75t_L g606 ( .A(n_450), .Y(n_606) );
INVx3_ASAP7_75t_L g671 ( .A(n_450), .Y(n_671) );
OAI221xp5_ASAP7_75t_L g918 ( .A1(n_450), .A2(n_919), .B1(n_920), .B2(n_921), .C(n_924), .Y(n_918) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g1047 ( .A(n_453), .B(n_1048), .Y(n_1047) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_454), .A2(n_682), .B1(n_683), .B2(n_685), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_454), .A2(n_683), .B1(n_833), .B2(n_834), .Y(n_832) );
BUFx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g530 ( .A(n_455), .Y(n_530) );
INVx1_ASAP7_75t_L g794 ( .A(n_455), .Y(n_794) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_455), .B(n_1131), .Y(n_1130) );
AND2x2_ASAP7_75t_L g1506 ( .A(n_455), .B(n_1131), .Y(n_1506) );
OAI21xp5_ASAP7_75t_L g587 ( .A1(n_456), .A2(n_588), .B(n_599), .Y(n_587) );
OAI21xp5_ASAP7_75t_L g904 ( .A1(n_456), .A2(n_905), .B(n_916), .Y(n_904) );
OAI21xp5_ASAP7_75t_L g1020 ( .A1(n_456), .A2(n_1021), .B(n_1029), .Y(n_1020) );
OAI21xp5_ASAP7_75t_SL g1045 ( .A1(n_456), .A2(n_1046), .B(n_1054), .Y(n_1045) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_458), .B(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g969 ( .A(n_458), .Y(n_969) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
OR2x6_ASAP7_75t_L g701 ( .A(n_459), .B(n_702), .Y(n_701) );
AND2x4_ASAP7_75t_L g781 ( .A(n_459), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g1016 ( .A(n_461), .Y(n_1016) );
AND2x4_ASAP7_75t_L g461 ( .A(n_462), .B(n_466), .Y(n_461) );
AND2x4_ASAP7_75t_L g559 ( .A(n_462), .B(n_466), .Y(n_559) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g717 ( .A(n_466), .Y(n_717) );
INVx3_ASAP7_75t_L g762 ( .A(n_467), .Y(n_762) );
INVx4_ASAP7_75t_L g1520 ( .A(n_467), .Y(n_1520) );
BUFx6f_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
BUFx2_ASAP7_75t_L g749 ( .A(n_468), .Y(n_749) );
BUFx3_ASAP7_75t_L g1101 ( .A(n_468), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_469), .Y(n_1173) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_471), .A2(n_474), .B1(n_597), .B2(n_598), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_471), .A2(n_474), .B1(n_624), .B2(n_625), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_471), .A2(n_474), .B1(n_902), .B2(n_903), .Y(n_901) );
AND2x4_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
AND2x4_ASAP7_75t_L g718 ( .A(n_472), .B(n_473), .Y(n_718) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_472), .A2(n_699), .B1(n_734), .B2(n_770), .Y(n_769) );
INVx2_ASAP7_75t_L g502 ( .A(n_474), .Y(n_502) );
INVx2_ASAP7_75t_L g973 ( .A(n_474), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1443 ( .A1(n_474), .A2(n_718), .B1(n_1444), .B2(n_1445), .Y(n_1443) );
NAND3xp33_ASAP7_75t_L g477 ( .A(n_478), .B(n_504), .C(n_508), .Y(n_477) );
NOR3xp33_ASAP7_75t_L g478 ( .A(n_479), .B(n_495), .C(n_503), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_484), .Y(n_479) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_490), .A2(n_567), .B1(n_568), .B2(n_572), .C(n_573), .Y(n_566) );
INVx3_ASAP7_75t_L g710 ( .A(n_490), .Y(n_710) );
OR2x6_ASAP7_75t_SL g739 ( .A(n_490), .B(n_740), .Y(n_739) );
BUFx2_ASAP7_75t_L g1452 ( .A(n_490), .Y(n_1452) );
BUFx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g869 ( .A(n_496), .B(n_870), .Y(n_869) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_500), .Y(n_496) );
OR2x2_ASAP7_75t_L g1019 ( .A(n_497), .B(n_500), .Y(n_1019) );
INVx2_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx4f_ASAP7_75t_L g744 ( .A(n_499), .Y(n_744) );
OR2x4_ASAP7_75t_L g1178 ( .A(n_499), .B(n_1160), .Y(n_1178) );
INVxp67_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g709 ( .A(n_501), .B(n_710), .Y(n_709) );
NOR3xp33_ASAP7_75t_L g1188 ( .A(n_503), .B(n_1189), .C(n_1200), .Y(n_1188) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_507), .B(n_812), .Y(n_811) );
OAI21xp5_ASAP7_75t_L g508 ( .A1(n_509), .A2(n_523), .B(n_548), .Y(n_508) );
INVx1_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g627 ( .A(n_525), .Y(n_627) );
INVx1_ASAP7_75t_L g917 ( .A(n_525), .Y(n_917) );
INVx4_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g1206 ( .A(n_529), .Y(n_1206) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g686 ( .A(n_531), .Y(n_686) );
OAI221xp5_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_536), .B1(n_537), .B2(n_541), .C(n_542), .Y(n_532) );
OAI22xp5_ASAP7_75t_L g925 ( .A1(n_533), .A2(n_926), .B1(n_927), .B2(n_928), .Y(n_925) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_533), .A2(n_928), .B1(n_1208), .B2(n_1209), .C(n_1210), .Y(n_1207) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx6f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx3_ASAP7_75t_L g679 ( .A(n_535), .Y(n_679) );
INVx4_ASAP7_75t_L g830 ( .A(n_535), .Y(n_830) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx4_ASAP7_75t_L g837 ( .A(n_538), .Y(n_837) );
BUFx6f_ASAP7_75t_L g929 ( .A(n_538), .Y(n_929) );
INVx2_ASAP7_75t_L g965 ( .A(n_538), .Y(n_965) );
INVx8_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g1145 ( .A(n_539), .B(n_1131), .Y(n_1145) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_550), .Y(n_847) );
BUFx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g635 ( .A(n_551), .Y(n_635) );
AOI21x1_ASAP7_75t_L g661 ( .A1(n_551), .A2(n_662), .B(n_690), .Y(n_661) );
HB1xp67_ASAP7_75t_L g1469 ( .A(n_551), .Y(n_1469) );
BUFx3_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AO22x2_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_611), .B1(n_612), .B2(n_654), .Y(n_553) );
INVx1_ASAP7_75t_L g654 ( .A(n_554), .Y(n_654) );
AND4x1_ASAP7_75t_L g555 ( .A(n_556), .B(n_560), .C(n_587), .D(n_610), .Y(n_555) );
NOR3xp33_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .C(n_584), .Y(n_560) );
OAI22xp5_ASAP7_75t_SL g562 ( .A1(n_563), .A2(n_566), .B1(n_575), .B2(n_576), .Y(n_562) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_563), .Y(n_1087) );
BUFx4f_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx8_ASAP7_75t_L g638 ( .A(n_564), .Y(n_638) );
BUFx2_ASAP7_75t_L g853 ( .A(n_564), .Y(n_853) );
OAI221xp5_ASAP7_75t_L g639 ( .A1(n_568), .A2(n_640), .B1(n_641), .B2(n_642), .C(n_643), .Y(n_639) );
INVx3_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g1486 ( .A(n_571), .Y(n_1486) );
OAI221xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_579), .B1(n_580), .B2(n_582), .C(n_583), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx6f_ASAP7_75t_L g695 ( .A(n_578), .Y(n_695) );
BUFx6f_ASAP7_75t_L g697 ( .A(n_578), .Y(n_697) );
INVx2_ASAP7_75t_L g979 ( .A(n_578), .Y(n_979) );
AND2x4_ASAP7_75t_L g1159 ( .A(n_578), .B(n_1160), .Y(n_1159) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_579), .A2(n_601), .B(n_605), .C(n_607), .Y(n_600) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_580), .A2(n_629), .B1(n_640), .B2(n_645), .C(n_646), .Y(n_644) );
CKINVDCx8_ASAP7_75t_R g580 ( .A(n_581), .Y(n_580) );
INVx3_ASAP7_75t_L g746 ( .A(n_581), .Y(n_746) );
INVx3_ASAP7_75t_L g758 ( .A(n_581), .Y(n_758) );
INVx3_ASAP7_75t_L g856 ( .A(n_581), .Y(n_856) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_586), .A2(n_704), .B1(n_1048), .B2(n_1069), .Y(n_1068) );
INVx2_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g1059 ( .A(n_594), .Y(n_1059) );
INVx3_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g1025 ( .A(n_595), .Y(n_1025) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx2_ASAP7_75t_L g680 ( .A(n_602), .Y(n_680) );
INVx2_ASAP7_75t_L g831 ( .A(n_602), .Y(n_831) );
INVx4_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
BUFx4f_ASAP7_75t_L g689 ( .A(n_603), .Y(n_689) );
OR2x6_ASAP7_75t_L g807 ( .A(n_603), .B(n_808), .Y(n_807) );
BUFx4f_ASAP7_75t_L g919 ( .A(n_603), .Y(n_919) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
BUFx3_ASAP7_75t_L g632 ( .A(n_604), .Y(n_632) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g665 ( .A(n_609), .Y(n_665) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND4x1_ASAP7_75t_L g613 ( .A(n_614), .B(n_636), .C(n_650), .D(n_653), .Y(n_613) );
OAI21xp5_ASAP7_75t_L g614 ( .A1(n_615), .A2(n_626), .B(n_635), .Y(n_614) );
INVx2_ASAP7_75t_SL g619 ( .A(n_620), .Y(n_619) );
OAI211xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_630), .B(n_633), .C(n_634), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g843 ( .A1(n_630), .A2(n_844), .B(n_845), .C(n_846), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1114 ( .A1(n_630), .A2(n_836), .B1(n_1094), .B2(n_1099), .Y(n_1114) );
INVx5_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
OR2x2_ASAP7_75t_L g796 ( .A(n_632), .B(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_SL g1117 ( .A(n_632), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1502 ( .A(n_632), .Y(n_1502) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx2_ASAP7_75t_L g699 ( .A(n_648), .Y(n_699) );
INVx1_ASAP7_75t_L g984 ( .A(n_648), .Y(n_984) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AO22x2_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_874), .B1(n_931), .B2(n_932), .Y(n_656) );
INVx1_ASAP7_75t_L g931 ( .A(n_657), .Y(n_931) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_658), .B(n_822), .Y(n_657) );
OAI22xp5_ASAP7_75t_L g658 ( .A1(n_659), .A2(n_729), .B1(n_820), .B2(n_821), .Y(n_658) );
INVx1_ASAP7_75t_L g821 ( .A(n_659), .Y(n_821) );
NAND3xp33_ASAP7_75t_L g659 ( .A(n_660), .B(n_722), .C(n_726), .Y(n_659) );
INVx1_ASAP7_75t_L g723 ( .A(n_661), .Y(n_723) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x4_ASAP7_75t_L g813 ( .A(n_665), .B(n_814), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .B1(n_672), .B2(n_674), .Y(n_666) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g675 ( .A(n_670), .Y(n_675) );
INVx1_ASAP7_75t_L g955 ( .A(n_675), .Y(n_955) );
INVx2_ASAP7_75t_L g1459 ( .A(n_675), .Y(n_1459) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_686), .B1(n_687), .B2(n_688), .Y(n_677) );
INVx2_ASAP7_75t_SL g1111 ( .A(n_679), .Y(n_1111) );
OAI211xp5_ASAP7_75t_L g1030 ( .A1(n_680), .A2(n_1031), .B(n_1032), .C(n_1035), .Y(n_1030) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI222xp33_ASAP7_75t_L g716 ( .A1(n_685), .A2(n_717), .B1(n_718), .B2(n_719), .C1(n_720), .C2(n_721), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g828 ( .A1(n_686), .A2(n_687), .B1(n_829), .B2(n_835), .Y(n_828) );
OAI211xp5_ASAP7_75t_L g1049 ( .A1(n_689), .A2(n_1050), .B(n_1051), .C(n_1052), .Y(n_1049) );
INVx1_ASAP7_75t_L g724 ( .A(n_691), .Y(n_724) );
AND2x2_ASAP7_75t_L g691 ( .A(n_692), .B(n_703), .Y(n_691) );
INVx2_ASAP7_75t_SL g1490 ( .A(n_695), .Y(n_1490) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_SL g1075 ( .A(n_701), .Y(n_1075) );
INVx1_ASAP7_75t_L g728 ( .A(n_706), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_715), .Y(n_706) );
NAND2x1_ASAP7_75t_L g707 ( .A(n_708), .B(n_711), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g1484 ( .A(n_710), .Y(n_1484) );
INVx2_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_712), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
AND2x4_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g727 ( .A(n_716), .Y(n_727) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_717), .A2(n_720), .B1(n_834), .B2(n_850), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g722 ( .A1(n_723), .A2(n_724), .B(n_725), .Y(n_722) );
OAI21xp33_ASAP7_75t_L g726 ( .A1(n_725), .A2(n_727), .B(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g820 ( .A(n_729), .Y(n_820) );
XNOR2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
NOR2x1_ASAP7_75t_L g731 ( .A(n_732), .B(n_777), .Y(n_731) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
INVx3_ASAP7_75t_L g870 ( .A(n_735), .Y(n_870) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_741), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_748), .B1(n_755), .B2(n_760), .C(n_766), .Y(n_742) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_744), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_743) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_744), .Y(n_1090) );
OAI22xp33_ASAP7_75t_L g1104 ( .A1(n_746), .A2(n_1090), .B1(n_1105), .B2(n_1106), .Y(n_1104) );
OAI221xp5_ASAP7_75t_L g748 ( .A1(n_749), .A2(n_750), .B1(n_751), .B2(n_753), .C(n_754), .Y(n_748) );
OR2x6_ASAP7_75t_L g766 ( .A(n_749), .B(n_767), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g801 ( .A1(n_750), .A2(n_802), .B(n_805), .C(n_806), .Y(n_801) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_SL g756 ( .A(n_752), .Y(n_756) );
INVx5_ASAP7_75t_L g862 ( .A(n_752), .Y(n_862) );
INVx2_ASAP7_75t_SL g1005 ( .A(n_752), .Y(n_1005) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B1(n_758), .B2(n_759), .Y(n_755) );
OAI221xp5_ASAP7_75t_L g854 ( .A1(n_756), .A2(n_855), .B1(n_856), .B2(n_857), .C(n_858), .Y(n_854) );
OAI22xp5_ASAP7_75t_L g1093 ( .A1(n_758), .A2(n_979), .B1(n_1094), .B2(n_1095), .Y(n_1093) );
OAI21xp5_ASAP7_75t_SL g760 ( .A1(n_761), .A2(n_763), .B(n_764), .Y(n_760) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g1092 ( .A(n_762), .Y(n_1092) );
BUFx2_ASAP7_75t_L g983 ( .A(n_765), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_770), .A2(n_786), .B1(n_788), .B2(n_789), .Y(n_785) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx4_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVx2_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
NAND3xp33_ASAP7_75t_L g777 ( .A(n_778), .B(n_809), .C(n_815), .Y(n_777) );
NOR3xp33_ASAP7_75t_SL g778 ( .A(n_779), .B(n_795), .C(n_798), .Y(n_778) );
OAI21xp5_ASAP7_75t_SL g779 ( .A1(n_780), .A2(n_784), .B(n_785), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
INVx4_ASAP7_75t_L g1108 ( .A(n_781), .Y(n_1108) );
INVx2_ASAP7_75t_L g1530 ( .A(n_781), .Y(n_1530) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
INVx2_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
NAND2x2_ASAP7_75t_L g790 ( .A(n_791), .B(n_793), .Y(n_790) );
INVx1_ASAP7_75t_L g808 ( .A(n_791), .Y(n_808) );
INVx2_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
INVx2_ASAP7_75t_SL g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g814 ( .A(n_797), .Y(n_814) );
OAI21xp5_ASAP7_75t_L g798 ( .A1(n_799), .A2(n_801), .B(n_807), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx2_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
INVx1_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
BUFx2_ASAP7_75t_L g836 ( .A(n_804), .Y(n_836) );
BUFx2_ASAP7_75t_L g923 ( .A(n_804), .Y(n_923) );
INVx2_ASAP7_75t_L g1540 ( .A(n_804), .Y(n_1540) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_810), .B(n_811), .Y(n_809) );
INVx1_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
AOI21xp5_ASAP7_75t_L g824 ( .A1(n_825), .A2(n_847), .B(n_848), .Y(n_824) );
NAND4xp25_ASAP7_75t_L g825 ( .A(n_826), .B(n_828), .C(n_838), .D(n_843), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_836), .A2(n_1091), .B1(n_1106), .B2(n_1112), .Y(n_1115) );
INVx2_ASAP7_75t_L g1113 ( .A(n_837), .Y(n_1113) );
OAI221xp5_ASAP7_75t_L g861 ( .A1(n_844), .A2(n_862), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_861) );
OAI22xp5_ASAP7_75t_SL g852 ( .A1(n_853), .A2(n_854), .B1(n_860), .B2(n_861), .Y(n_852) );
INVx2_ASAP7_75t_SL g890 ( .A(n_859), .Y(n_890) );
BUFx3_ASAP7_75t_L g1072 ( .A(n_859), .Y(n_1072) );
INVx1_ASAP7_75t_L g1196 ( .A(n_859), .Y(n_1196) );
OAI22xp5_ASAP7_75t_L g1482 ( .A1(n_860), .A2(n_1087), .B1(n_1483), .B2(n_1489), .Y(n_1482) );
INVx8_ASAP7_75t_L g1098 ( .A(n_862), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_873), .B(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g999 ( .A(n_873), .B(n_1000), .Y(n_999) );
INVx2_ASAP7_75t_L g932 ( .A(n_874), .Y(n_932) );
XOR2x2_ASAP7_75t_L g874 ( .A(n_875), .B(n_930), .Y(n_874) );
NAND2xp5_ASAP7_75t_SL g875 ( .A(n_876), .B(n_904), .Y(n_875) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_879), .B(n_887), .Y(n_878) );
NOR2xp33_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .Y(n_879) );
NAND2xp5_ASAP7_75t_SL g883 ( .A(n_884), .B(n_886), .Y(n_883) );
NAND4xp25_ASAP7_75t_SL g995 ( .A(n_886), .B(n_996), .C(n_999), .D(n_1001), .Y(n_995) );
INVx2_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
BUFx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
BUFx2_ASAP7_75t_L g981 ( .A(n_895), .Y(n_981) );
BUFx2_ASAP7_75t_L g1009 ( .A(n_895), .Y(n_1009) );
INVx1_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
NAND3xp33_ASAP7_75t_SL g905 ( .A(n_906), .B(n_909), .C(n_915), .Y(n_905) );
INVx2_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_SL g913 ( .A(n_914), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1537 ( .A1(n_919), .A2(n_1538), .B1(n_1541), .B2(n_1542), .Y(n_1537) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx2_ASAP7_75t_L g1536 ( .A(n_922), .Y(n_1536) );
INVx4_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
OAI22xp33_ASAP7_75t_L g1531 ( .A1(n_928), .A2(n_1532), .B1(n_1533), .B2(n_1534), .Y(n_1531) );
INVx5_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx6_ASAP7_75t_L g1545 ( .A(n_929), .Y(n_1545) );
INVx1_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
XNOR2xp5_ASAP7_75t_L g935 ( .A(n_936), .B(n_1040), .Y(n_935) );
INVx1_ASAP7_75t_L g936 ( .A(n_937), .Y(n_936) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
OAI22x1_ASAP7_75t_L g938 ( .A1(n_939), .A2(n_990), .B1(n_991), .B2(n_1039), .Y(n_938) );
INVx2_ASAP7_75t_L g1039 ( .A(n_939), .Y(n_1039) );
AO21x2_ASAP7_75t_L g939 ( .A1(n_940), .A2(n_941), .B(n_989), .Y(n_939) );
NAND3xp33_ASAP7_75t_SL g941 ( .A(n_942), .B(n_945), .C(n_970), .Y(n_941) );
OAI21xp5_ASAP7_75t_L g945 ( .A1(n_946), .A2(n_957), .B(n_969), .Y(n_945) );
INVx1_ASAP7_75t_L g952 ( .A(n_953), .Y(n_952) );
INVx1_ASAP7_75t_L g968 ( .A(n_953), .Y(n_968) );
INVx1_ASAP7_75t_L g1468 ( .A(n_953), .Y(n_1468) );
INVx1_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g958 ( .A1(n_959), .A2(n_962), .B1(n_963), .B2(n_966), .C(n_967), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g1116 ( .A1(n_959), .A2(n_1095), .B1(n_1102), .B2(n_1117), .Y(n_1116) );
INVx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx2_ASAP7_75t_SL g960 ( .A(n_961), .Y(n_960) );
BUFx6f_ASAP7_75t_L g1464 ( .A(n_961), .Y(n_1464) );
BUFx3_ASAP7_75t_L g1544 ( .A(n_961), .Y(n_1544) );
BUFx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_964), .A2(n_1464), .B1(n_1465), .B2(n_1466), .C(n_1467), .Y(n_1463) );
BUFx6f_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx1_ASAP7_75t_L g971 ( .A(n_972), .Y(n_971) );
INVx1_ASAP7_75t_L g978 ( .A(n_979), .Y(n_978) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
NAND2x1p5_ASAP7_75t_L g991 ( .A(n_992), .B(n_1012), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_994), .B(n_1010), .Y(n_993) );
INVxp67_ASAP7_75t_L g994 ( .A(n_995), .Y(n_994) );
NOR2xp33_ASAP7_75t_SL g1036 ( .A(n_995), .B(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1103 ( .A(n_1009), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_1010), .B(n_1038), .Y(n_1037) );
INVx1_ASAP7_75t_L g1013 ( .A(n_1014), .Y(n_1013) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1020), .Y(n_1014) );
AOI21xp5_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1017), .B(n_1018), .Y(n_1015) );
INVx1_ASAP7_75t_L g1033 ( .A(n_1034), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_1041), .A2(n_1042), .B1(n_1081), .B2(n_1223), .Y(n_1040) );
INVx1_ASAP7_75t_L g1041 ( .A(n_1042), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1044), .Y(n_1080) );
NAND3xp33_ASAP7_75t_L g1044 ( .A(n_1045), .B(n_1063), .C(n_1066), .Y(n_1044) );
NAND2xp5_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1070), .Y(n_1067) );
OAI22xp5_ASAP7_75t_SL g1312 ( .A1(n_1079), .A2(n_1313), .B1(n_1314), .B2(n_1315), .Y(n_1312) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1081), .Y(n_1223) );
AOI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1083), .B1(n_1186), .B2(n_1222), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
NAND3xp33_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1123), .C(n_1153), .Y(n_1084) );
NOR2xp33_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1107), .Y(n_1085) );
OAI33xp33_ASAP7_75t_L g1086 ( .A1(n_1087), .A2(n_1088), .A3(n_1093), .B1(n_1096), .B2(n_1103), .B3(n_1104), .Y(n_1086) );
OAI22xp33_ASAP7_75t_L g1088 ( .A1(n_1089), .A2(n_1090), .B1(n_1091), .B2(n_1092), .Y(n_1088) );
OAI22xp5_ASAP7_75t_L g1109 ( .A1(n_1089), .A2(n_1105), .B1(n_1110), .B2(n_1112), .Y(n_1109) );
OAI22xp5_ASAP7_75t_L g1096 ( .A1(n_1097), .A2(n_1099), .B1(n_1100), .B2(n_1102), .Y(n_1096) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
BUFx6f_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx2_ASAP7_75t_L g1163 ( .A(n_1101), .Y(n_1163) );
OAI33xp33_ASAP7_75t_L g1107 ( .A1(n_1108), .A2(n_1109), .A3(n_1114), .B1(n_1115), .B2(n_1116), .B3(n_1118), .Y(n_1107) );
INVx2_ASAP7_75t_L g1110 ( .A(n_1111), .Y(n_1110) );
INVx2_ASAP7_75t_L g1112 ( .A(n_1113), .Y(n_1112) );
OAI22xp5_ASAP7_75t_L g1535 ( .A1(n_1117), .A2(n_1485), .B1(n_1491), .B2(n_1536), .Y(n_1535) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1119), .Y(n_1118) );
INVx1_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx1_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
OAI31xp33_ASAP7_75t_SL g1123 ( .A1(n_1124), .A2(n_1136), .A3(n_1146), .B(n_1150), .Y(n_1123) );
INVx1_ASAP7_75t_L g1125 ( .A(n_1126), .Y(n_1125) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1126), .Y(n_1503) );
AOI22xp33_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1132), .B1(n_1133), .B2(n_1134), .Y(n_1128) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_1132), .A2(n_1167), .B1(n_1171), .B2(n_1174), .Y(n_1166) );
BUFx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_L g1504 ( .A1(n_1135), .A2(n_1505), .B1(n_1506), .B2(n_1507), .Y(n_1504) );
INVx1_ASAP7_75t_L g1137 ( .A(n_1138), .Y(n_1137) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
BUFx2_ASAP7_75t_L g1509 ( .A(n_1139), .Y(n_1509) );
INVx2_ASAP7_75t_L g1141 ( .A(n_1142), .Y(n_1141) );
INVx2_ASAP7_75t_L g1142 ( .A(n_1143), .Y(n_1142) );
INVx2_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_1145), .Y(n_1144) );
INVx2_ASAP7_75t_L g1511 ( .A(n_1145), .Y(n_1511) );
INVx3_ASAP7_75t_SL g1148 ( .A(n_1149), .Y(n_1148) );
CKINVDCx16_ASAP7_75t_R g1498 ( .A(n_1149), .Y(n_1498) );
BUFx3_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
BUFx2_ASAP7_75t_L g1512 ( .A(n_1151), .Y(n_1512) );
OAI31xp33_ASAP7_75t_SL g1153 ( .A1(n_1154), .A2(n_1161), .A3(n_1175), .B(n_1181), .Y(n_1153) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx2_ASAP7_75t_SL g1516 ( .A(n_1157), .Y(n_1516) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx2_ASAP7_75t_L g1517 ( .A(n_1159), .Y(n_1517) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
CKINVDCx8_ASAP7_75t_R g1164 ( .A(n_1165), .Y(n_1164) );
AOI22xp33_ASAP7_75t_L g1521 ( .A1(n_1167), .A2(n_1171), .B1(n_1505), .B2(n_1522), .Y(n_1521) );
BUFx3_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1170), .Y(n_1168) );
AND2x4_ASAP7_75t_L g1172 ( .A(n_1169), .B(n_1173), .Y(n_1172) );
BUFx6f_ASAP7_75t_L g1171 ( .A(n_1172), .Y(n_1171) );
INVx1_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1177), .Y(n_1526) );
INVx2_ASAP7_75t_SL g1177 ( .A(n_1178), .Y(n_1177) );
BUFx3_ASAP7_75t_L g1179 ( .A(n_1180), .Y(n_1179) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1180), .Y(n_1525) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1184), .Y(n_1181) );
AND2x2_ASAP7_75t_SL g1527 ( .A(n_1182), .B(n_1184), .Y(n_1527) );
INVx1_ASAP7_75t_SL g1182 ( .A(n_1183), .Y(n_1182) );
INVx1_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1186), .Y(n_1222) );
NAND3xp33_ASAP7_75t_L g1187 ( .A(n_1188), .B(n_1201), .C(n_1204), .Y(n_1187) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1193), .Y(n_1189) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1196), .Y(n_1195) );
OAI21xp5_ASAP7_75t_L g1204 ( .A1(n_1205), .A2(n_1214), .B(n_1221), .Y(n_1204) );
BUFx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
OAI221xp5_ASAP7_75t_L g1225 ( .A1(n_1226), .A2(n_1431), .B1(n_1433), .B2(n_1470), .C(n_1473), .Y(n_1225) );
NOR2xp67_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1378), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1342), .Y(n_1227) );
O2A1O1Ixp33_ASAP7_75t_SL g1228 ( .A1(n_1229), .A2(n_1280), .B(n_1309), .C(n_1316), .Y(n_1228) );
O2A1O1Ixp33_ASAP7_75t_L g1229 ( .A1(n_1230), .A2(n_1246), .B(n_1259), .C(n_1275), .Y(n_1229) );
INVx2_ASAP7_75t_L g1262 ( .A(n_1230), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1306 ( .A(n_1230), .B(n_1302), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1230), .B(n_1286), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1345 ( .A(n_1230), .B(n_1346), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1354 ( .A(n_1230), .B(n_1287), .Y(n_1354) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_1230), .A2(n_1262), .B1(n_1412), .B2(n_1414), .C(n_1416), .Y(n_1411) );
INVx2_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1231), .B(n_1277), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g1387 ( .A(n_1231), .B(n_1268), .Y(n_1387) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1284 ( .A(n_1232), .B(n_1285), .Y(n_1284) );
OR2x2_ASAP7_75t_L g1293 ( .A(n_1232), .B(n_1277), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1232), .B(n_1277), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1367 ( .A(n_1232), .B(n_1268), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1392 ( .A(n_1232), .B(n_1268), .Y(n_1392) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1240), .Y(n_1232) );
INVx2_ASAP7_75t_L g1313 ( .A(n_1234), .Y(n_1313) );
AND2x6_ASAP7_75t_L g1234 ( .A(n_1235), .B(n_1236), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1238 ( .A(n_1235), .B(n_1239), .Y(n_1238) );
AND2x4_ASAP7_75t_L g1241 ( .A(n_1235), .B(n_1242), .Y(n_1241) );
AND2x6_ASAP7_75t_L g1244 ( .A(n_1235), .B(n_1245), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1235), .B(n_1239), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1235), .B(n_1239), .Y(n_1289) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1235), .B(n_1242), .Y(n_1432) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1237), .B(n_1243), .Y(n_1242) );
INVxp67_ASAP7_75t_L g1315 ( .A(n_1238), .Y(n_1315) );
HB1xp67_ASAP7_75t_L g1551 ( .A(n_1242), .Y(n_1551) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1246), .Y(n_1349) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_1247), .B(n_1251), .Y(n_1246) );
BUFx2_ASAP7_75t_L g1267 ( .A(n_1247), .Y(n_1267) );
INVx2_ASAP7_75t_L g1301 ( .A(n_1247), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1346 ( .A(n_1247), .B(n_1347), .Y(n_1346) );
AND2x2_ASAP7_75t_L g1356 ( .A(n_1247), .B(n_1272), .Y(n_1356) );
AOI222xp33_ASAP7_75t_L g1416 ( .A1(n_1247), .A2(n_1346), .B1(n_1358), .B2(n_1366), .C1(n_1417), .C2(n_1418), .Y(n_1416) );
AND2x2_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1249), .Y(n_1247) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_1251), .A2(n_1281), .B1(n_1291), .B2(n_1294), .C(n_1296), .Y(n_1280) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1328 ( .A(n_1252), .B(n_1300), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_1252), .B(n_1266), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1415 ( .A(n_1252), .B(n_1302), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1256), .Y(n_1252) );
INVx2_ASAP7_75t_L g1273 ( .A(n_1253), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1347 ( .A(n_1253), .B(n_1274), .Y(n_1347) );
OAI222xp33_ASAP7_75t_L g1405 ( .A1(n_1253), .A2(n_1276), .B1(n_1333), .B2(n_1398), .C1(n_1406), .C2(n_1408), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1430 ( .A(n_1253), .B(n_1267), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1253 ( .A(n_1254), .B(n_1255), .Y(n_1253) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1256), .Y(n_1274) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1256), .B(n_1273), .Y(n_1307) );
AND3x1_ASAP7_75t_L g1324 ( .A(n_1256), .B(n_1273), .C(n_1301), .Y(n_1324) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1256), .B(n_1267), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1256), .B(n_1267), .Y(n_1365) );
NOR2xp33_ASAP7_75t_L g1386 ( .A(n_1256), .B(n_1387), .Y(n_1386) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1256), .B(n_1301), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1256 ( .A(n_1257), .B(n_1258), .Y(n_1256) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1261), .B(n_1263), .Y(n_1260) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1261), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1317 ( .A(n_1261), .B(n_1299), .Y(n_1317) );
INVx2_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
A2O1A1Ixp33_ASAP7_75t_L g1329 ( .A1(n_1262), .A2(n_1310), .B(n_1330), .C(n_1331), .Y(n_1329) );
A2O1A1Ixp33_ASAP7_75t_L g1360 ( .A1(n_1262), .A2(n_1319), .B(n_1361), .C(n_1362), .Y(n_1360) );
NAND2xp5_ASAP7_75t_L g1374 ( .A(n_1262), .B(n_1375), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1262), .B(n_1319), .Y(n_1428) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1264), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1264 ( .A(n_1265), .B(n_1271), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1266), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1266), .B(n_1347), .Y(n_1407) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1268), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1295 ( .A(n_1267), .B(n_1274), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1338 ( .A(n_1267), .B(n_1307), .Y(n_1338) );
OR2x2_ASAP7_75t_L g1339 ( .A(n_1267), .B(n_1273), .Y(n_1339) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1267), .B(n_1273), .Y(n_1361) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1268), .B(n_1287), .Y(n_1297) );
INVx2_ASAP7_75t_L g1302 ( .A(n_1268), .Y(n_1302) );
INVx1_ASAP7_75t_L g1323 ( .A(n_1268), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1268), .B(n_1277), .Y(n_1373) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1268), .B(n_1419), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1429 ( .A(n_1268), .B(n_1430), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1270), .Y(n_1268) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_1271), .A2(n_1291), .B1(n_1369), .B2(n_1373), .C(n_1374), .Y(n_1368) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1272), .B(n_1300), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1272), .B(n_1301), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1273), .B(n_1274), .Y(n_1272) );
AOI321xp33_ASAP7_75t_L g1296 ( .A1(n_1273), .A2(n_1275), .A3(n_1297), .B1(n_1298), .B2(n_1299), .C(n_1303), .Y(n_1296) );
CKINVDCx14_ASAP7_75t_R g1275 ( .A(n_1276), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1276), .B(n_1310), .Y(n_1325) );
INVx3_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1277), .Y(n_1285) );
AND2x2_ASAP7_75t_L g1319 ( .A(n_1277), .B(n_1287), .Y(n_1319) );
OR2x2_ASAP7_75t_L g1331 ( .A(n_1277), .B(n_1286), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1277), .B(n_1367), .Y(n_1366) );
OR2x2_ASAP7_75t_L g1384 ( .A(n_1277), .B(n_1287), .Y(n_1384) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_1277), .B(n_1286), .Y(n_1389) );
AND2x4_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1279), .Y(n_1277) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NOR2xp33_ASAP7_75t_SL g1282 ( .A(n_1283), .B(n_1286), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1284), .B(n_1302), .Y(n_1341) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1284), .B(n_1286), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g1292 ( .A(n_1286), .B(n_1293), .Y(n_1292) );
NAND3xp33_ASAP7_75t_L g1390 ( .A(n_1286), .B(n_1307), .C(n_1391), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1286), .B(n_1377), .Y(n_1422) );
CKINVDCx6p67_ASAP7_75t_R g1286 ( .A(n_1287), .Y(n_1286) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_1287), .B(n_1395), .Y(n_1397) );
NAND2xp5_ASAP7_75t_L g1410 ( .A(n_1287), .B(n_1311), .Y(n_1410) );
OR2x6_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1290), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1308 ( .A(n_1288), .B(n_1290), .Y(n_1308) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1292), .Y(n_1291) );
INVx2_ASAP7_75t_L g1417 ( .A(n_1293), .Y(n_1417) );
OAI332xp33_ASAP7_75t_L g1423 ( .A1(n_1293), .A2(n_1323), .A3(n_1384), .B1(n_1424), .B2(n_1426), .B3(n_1427), .C1(n_1428), .C2(n_1429), .Y(n_1423) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
CKINVDCx14_ASAP7_75t_R g1427 ( .A(n_1297), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1357 ( .A(n_1300), .B(n_1307), .Y(n_1357) );
AND2x2_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1302), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1403 ( .A(n_1301), .B(n_1347), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1301), .B(n_1415), .Y(n_1414) );
NAND2xp5_ASAP7_75t_SL g1424 ( .A(n_1301), .B(n_1425), .Y(n_1424) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_1302), .B(n_1363), .Y(n_1362) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1304), .Y(n_1303) );
NAND3xp33_ASAP7_75t_L g1304 ( .A(n_1305), .B(n_1307), .C(n_1308), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1402 ( .A(n_1305), .B(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1425 ( .A(n_1307), .B(n_1347), .Y(n_1425) );
NOR2xp33_ASAP7_75t_L g1401 ( .A(n_1308), .B(n_1402), .Y(n_1401) );
AOI221xp5_ASAP7_75t_L g1326 ( .A1(n_1309), .A2(n_1327), .B1(n_1329), .B2(n_1332), .C(n_1336), .Y(n_1326) );
A2O1A1Ixp33_ASAP7_75t_L g1379 ( .A1(n_1309), .A2(n_1322), .B(n_1380), .C(n_1383), .Y(n_1379) );
AOI311xp33_ASAP7_75t_L g1393 ( .A1(n_1309), .A2(n_1394), .A3(n_1395), .B(n_1396), .C(n_1401), .Y(n_1393) );
INVx3_ASAP7_75t_L g1309 ( .A(n_1310), .Y(n_1309) );
INVx2_ASAP7_75t_SL g1310 ( .A(n_1311), .Y(n_1310) );
INVx2_ASAP7_75t_SL g1377 ( .A(n_1311), .Y(n_1377) );
OAI221xp5_ASAP7_75t_L g1316 ( .A1(n_1317), .A2(n_1318), .B1(n_1320), .B2(n_1325), .C(n_1326), .Y(n_1316) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1319), .Y(n_1318) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1324), .Y(n_1321) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1322), .Y(n_1352) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1322), .B(n_1372), .Y(n_1376) );
NOR2xp33_ASAP7_75t_L g1399 ( .A(n_1322), .B(n_1363), .Y(n_1399) );
INVx2_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
AND2x2_ASAP7_75t_L g1394 ( .A(n_1323), .B(n_1338), .Y(n_1394) );
NAND2xp5_ASAP7_75t_SL g1408 ( .A(n_1323), .B(n_1334), .Y(n_1408) );
INVx2_ASAP7_75t_L g1335 ( .A(n_1324), .Y(n_1335) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
OAI211xp5_ASAP7_75t_L g1343 ( .A1(n_1331), .A2(n_1344), .B(n_1348), .C(n_1355), .Y(n_1343) );
NOR2xp33_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1335), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AOI21xp33_ASAP7_75t_L g1336 ( .A1(n_1337), .A2(n_1339), .B(n_1340), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1370 ( .A(n_1337), .B(n_1371), .Y(n_1370) );
OAI221xp5_ASAP7_75t_L g1383 ( .A1(n_1337), .A2(n_1384), .B1(n_1385), .B2(n_1388), .C(n_1390), .Y(n_1383) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1338), .Y(n_1337) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
OAI21xp5_ASAP7_75t_SL g1342 ( .A1(n_1343), .A2(n_1368), .B(n_1377), .Y(n_1342) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1351 ( .A(n_1346), .B(n_1352), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1381 ( .A(n_1347), .B(n_1382), .Y(n_1381) );
OAI21xp5_ASAP7_75t_L g1348 ( .A1(n_1349), .A2(n_1350), .B(n_1353), .Y(n_1348) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
O2A1O1Ixp33_ASAP7_75t_L g1355 ( .A1(n_1356), .A2(n_1357), .B(n_1358), .C(n_1359), .Y(n_1355) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1356), .B(n_1413), .Y(n_1412) );
CKINVDCx6p67_ASAP7_75t_R g1395 ( .A(n_1358), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1364), .Y(n_1359) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1366), .Y(n_1364) );
INVx1_ASAP7_75t_L g1426 ( .A(n_1365), .Y(n_1426) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
OAI22xp33_ASAP7_75t_L g1396 ( .A1(n_1371), .A2(n_1397), .B1(n_1398), .B2(n_1400), .Y(n_1396) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
NAND3xp33_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1393), .C(n_1404), .Y(n_1378) );
CKINVDCx5p33_ASAP7_75t_R g1380 ( .A(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1400 ( .A(n_1382), .Y(n_1400) );
INVxp67_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx1_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
AOI221xp5_ASAP7_75t_L g1404 ( .A1(n_1405), .A2(n_1409), .B1(n_1411), .B2(n_1421), .C(n_1423), .Y(n_1404) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
INVx1_ASAP7_75t_L g1419 ( .A(n_1420), .Y(n_1419) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
BUFx2_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
AND3x1_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1443), .C(n_1446), .Y(n_1439) );
INVx2_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
OAI21xp5_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1462), .B(n_1469), .Y(n_1454) );
INVx2_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVxp67_ASAP7_75t_L g1470 ( .A(n_1471), .Y(n_1470) );
BUFx3_ASAP7_75t_L g1471 ( .A(n_1472), .Y(n_1471) );
BUFx4f_ASAP7_75t_L g1474 ( .A(n_1475), .Y(n_1474) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1479), .Y(n_1478) );
NAND4xp75_ASAP7_75t_L g1480 ( .A(n_1481), .B(n_1496), .C(n_1513), .D(n_1528), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
OAI221xp5_ASAP7_75t_L g1483 ( .A1(n_1484), .A2(n_1485), .B1(n_1486), .B2(n_1487), .C(n_1488), .Y(n_1483) );
OAI221xp5_ASAP7_75t_L g1489 ( .A1(n_1486), .A2(n_1490), .B1(n_1491), .B2(n_1492), .C(n_1493), .Y(n_1489) );
OAI22xp5_ASAP7_75t_L g1543 ( .A1(n_1487), .A2(n_1492), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
OAI31xp33_ASAP7_75t_SL g1496 ( .A1(n_1497), .A2(n_1499), .A3(n_1508), .B(n_1512), .Y(n_1496) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1501 ( .A(n_1502), .Y(n_1501) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
OAI31xp33_ASAP7_75t_L g1513 ( .A1(n_1514), .A2(n_1518), .A3(n_1523), .B(n_1527), .Y(n_1513) );
INVx2_ASAP7_75t_SL g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
OA33x2_ASAP7_75t_L g1528 ( .A1(n_1529), .A2(n_1531), .A3(n_1535), .B1(n_1537), .B2(n_1543), .B3(n_1546), .Y(n_1528) );
BUFx6f_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx4_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
BUFx2_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
CKINVDCx5p33_ASAP7_75t_R g1546 ( .A(n_1547), .Y(n_1546) );
HB1xp67_ASAP7_75t_L g1548 ( .A(n_1549), .Y(n_1548) );
OAI21xp5_ASAP7_75t_L g1549 ( .A1(n_1550), .A2(n_1551), .B(n_1552), .Y(n_1549) );
INVx1_ASAP7_75t_L g1552 ( .A(n_1553), .Y(n_1552) );
endmodule