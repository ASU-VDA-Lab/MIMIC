module fake_netlist_5_1067_n_648 (n_137, n_91, n_82, n_122, n_10, n_140, n_24, n_124, n_86, n_136, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_120, n_135, n_30, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_29, n_79, n_131, n_47, n_25, n_53, n_8, n_44, n_40, n_34, n_100, n_62, n_138, n_71, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_12, n_67, n_121, n_36, n_76, n_87, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_11, n_7, n_15, n_48, n_50, n_52, n_88, n_110, n_648);

input n_137;
input n_91;
input n_82;
input n_122;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_120;
input n_135;
input n_30;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_29;
input n_79;
input n_131;
input n_47;
input n_25;
input n_53;
input n_8;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_71;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_11;
input n_7;
input n_15;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_648;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_194;
wire n_316;
wire n_389;
wire n_549;
wire n_418;
wire n_248;
wire n_146;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_619;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_515;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_483;
wire n_544;
wire n_155;
wire n_552;
wire n_547;
wire n_467;
wire n_564;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_590;
wire n_629;
wire n_378;
wire n_551;
wire n_581;
wire n_382;
wire n_554;
wire n_254;
wire n_583;
wire n_302;
wire n_265;
wire n_526;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_621;
wire n_455;
wire n_417;
wire n_612;
wire n_212;
wire n_498;
wire n_516;
wire n_385;
wire n_507;
wire n_497;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_610;
wire n_509;
wire n_568;
wire n_147;
wire n_373;
wire n_307;
wire n_633;
wire n_530;
wire n_150;
wire n_439;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_576;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_492;
wire n_563;
wire n_171;
wire n_153;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_548;
wire n_543;
wire n_260;
wire n_298;
wire n_320;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_519;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_546;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_152;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_308;
wire n_428;
wire n_379;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_297;
wire n_156;
wire n_603;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_157;
wire n_192;
wire n_636;
wire n_600;
wire n_223;
wire n_392;
wire n_158;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_183;
wire n_185;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_169;
wire n_522;
wire n_550;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_555;
wire n_473;
wire n_475;
wire n_422;
wire n_415;
wire n_141;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_584;
wire n_591;
wire n_145;
wire n_521;
wire n_614;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_553;
wire n_311;
wire n_208;
wire n_142;
wire n_214;
wire n_328;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_613;
wire n_241;
wire n_637;
wire n_357;
wire n_598;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_144;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_363;
wire n_413;
wire n_402;
wire n_638;
wire n_197;
wire n_573;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_149;
wire n_477;
wire n_461;
wire n_333;
wire n_571;
wire n_309;
wire n_512;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_151;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_542;
wire n_463;
wire n_488;
wire n_595;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_586;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_627;
wire n_172;
wire n_206;
wire n_217;
wire n_440;
wire n_478;
wire n_545;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_176;
wire n_557;
wire n_182;
wire n_143;
wire n_354;
wire n_575;
wire n_607;
wire n_480;
wire n_647;
wire n_237;
wire n_513;
wire n_425;
wire n_407;
wire n_527;
wire n_180;
wire n_560;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_602;
wire n_574;
wire n_437;
wire n_177;
wire n_453;
wire n_403;
wire n_421;
wire n_623;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_572;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_269;
wire n_529;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_644;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_565;
wire n_426;
wire n_520;
wire n_566;
wire n_409;
wire n_589;
wire n_597;
wire n_500;
wire n_562;
wire n_154;
wire n_148;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_599;
wire n_541;
wire n_391;
wire n_434;
wire n_645;
wire n_539;
wire n_175;
wire n_538;
wire n_262;
wire n_238;
wire n_639;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_360;
wire n_594;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_634;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_626;
wire n_424;
wire n_256;
wire n_305;
wire n_533;
wire n_278;

INVx1_ASAP7_75t_SL g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g142 ( 
.A(n_135),
.Y(n_142)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_SL g144 ( 
.A(n_69),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_103),
.Y(n_145)
);

CKINVDCx5p33_ASAP7_75t_R g146 ( 
.A(n_65),
.Y(n_146)
);

CKINVDCx5p33_ASAP7_75t_R g147 ( 
.A(n_129),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_55),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_60),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_77),
.Y(n_150)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_79),
.Y(n_151)
);

CKINVDCx5p33_ASAP7_75t_R g152 ( 
.A(n_122),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

CKINVDCx5p33_ASAP7_75t_R g154 ( 
.A(n_32),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_62),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_31),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_28),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_38),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_99),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_104),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_90),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_19),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_89),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_52),
.Y(n_166)
);

INVxp33_ASAP7_75t_SL g167 ( 
.A(n_134),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_0),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_1),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_68),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_0),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_14),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_128),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_20),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_25),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_138),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_71),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_43),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_17),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_51),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_16),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_33),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_50),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_118),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_72),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_74),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_46),
.Y(n_193)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_13),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_47),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_131),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_102),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

BUFx5_ASAP7_75t_L g201 ( 
.A(n_49),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_23),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_140),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_75),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_37),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_95),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_56),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_112),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_106),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_64),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_1),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_2),
.Y(n_212)
);

INVx5_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_172),
.B(n_167),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

BUFx12f_ASAP7_75t_L g218 ( 
.A(n_142),
.Y(n_218)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_142),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_169),
.Y(n_220)
);

AND2x4_ASAP7_75t_L g221 ( 
.A(n_145),
.B(n_18),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_155),
.B(n_2),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_3),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_183),
.B(n_3),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_143),
.B(n_4),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_149),
.B(n_4),
.Y(n_228)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_159),
.Y(n_229)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_141),
.B(n_5),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_201),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_182),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_196),
.B(n_5),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_186),
.B(n_6),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_201),
.B(n_6),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_182),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_153),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_160),
.B(n_7),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_182),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_199),
.B(n_7),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_173),
.B(n_164),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_165),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_8),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_201),
.B(n_8),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_166),
.B(n_9),
.Y(n_251)
);

BUFx8_ASAP7_75t_L g252 ( 
.A(n_177),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_181),
.B(n_9),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_185),
.B(n_10),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_188),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_191),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_193),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_237),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_224),
.B(n_147),
.Y(n_259)
);

OAI22xp33_ASAP7_75t_L g260 ( 
.A1(n_214),
.A2(n_178),
.B1(n_209),
.B2(n_208),
.Y(n_260)
);

OAI22xp33_ASAP7_75t_L g261 ( 
.A1(n_211),
.A2(n_200),
.B1(n_207),
.B2(n_206),
.Y(n_261)
);

AND2x4_ASAP7_75t_L g262 ( 
.A(n_221),
.B(n_203),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_222),
.A2(n_210),
.B1(n_205),
.B2(n_204),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_148),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_222),
.A2(n_202),
.B1(n_198),
.B2(n_197),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_247),
.B(n_151),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_236),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_226),
.A2(n_195),
.B1(n_192),
.B2(n_190),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_236),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_226),
.A2(n_163),
.B1(n_184),
.B2(n_180),
.Y(n_270)
);

OAI22xp33_ASAP7_75t_L g271 ( 
.A1(n_225),
.A2(n_189),
.B1(n_179),
.B2(n_176),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_152),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_223),
.A2(n_175),
.B1(n_171),
.B2(n_168),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_223),
.B(n_154),
.Y(n_274)
);

OAI22xp33_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_162),
.B1(n_161),
.B2(n_158),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_246),
.A2(n_156),
.B1(n_157),
.B2(n_12),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_236),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_255),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_278)
);

AND2x2_ASAP7_75t_SL g279 ( 
.A(n_246),
.B(n_11),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g280 ( 
.A(n_255),
.B(n_21),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_218),
.Y(n_281)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_241),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_234),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_234),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_L g285 ( 
.A1(n_249),
.A2(n_15),
.B1(n_22),
.B2(n_24),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_26),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_230),
.B(n_27),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_R g288 ( 
.A1(n_231),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_238),
.A2(n_35),
.B1(n_36),
.B2(n_40),
.Y(n_289)
);

OAI22xp33_ASAP7_75t_L g290 ( 
.A1(n_250),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g291 ( 
.A1(n_227),
.A2(n_240),
.B1(n_228),
.B2(n_218),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_253),
.B(n_45),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_234),
.Y(n_293)
);

BUFx6f_ASAP7_75t_SL g294 ( 
.A(n_221),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_230),
.B(n_48),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_212),
.A2(n_53),
.B1(n_54),
.B2(n_57),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_219),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_221),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_R g299 ( 
.A1(n_244),
.A2(n_63),
.B1(n_66),
.B2(n_67),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_R g300 ( 
.A1(n_220),
.A2(n_78),
.B1(n_80),
.B2(n_81),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_212),
.A2(n_82),
.B1(n_84),
.B2(n_85),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_253),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.Y(n_302)
);

OR2x2_ASAP7_75t_L g303 ( 
.A(n_243),
.B(n_91),
.Y(n_303)
);

AO22x2_ASAP7_75t_L g304 ( 
.A1(n_254),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.Y(n_304)
);

OAI22xp33_ASAP7_75t_SL g305 ( 
.A1(n_243),
.A2(n_96),
.B1(n_97),
.B2(n_98),
.Y(n_305)
);

INVx8_ASAP7_75t_L g306 ( 
.A(n_219),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_220),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_229),
.B(n_107),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_234),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_269),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_277),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_283),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_260),
.B(n_237),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_254),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_258),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_284),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_293),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_303),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

INVxp67_ASAP7_75t_SL g323 ( 
.A(n_262),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_272),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_259),
.B(n_257),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_273),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_268),
.Y(n_327)
);

INVx3_ASAP7_75t_R g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_287),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_294),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

NAND2xp33_ASAP7_75t_R g334 ( 
.A(n_274),
.B(n_257),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_280),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_286),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_263),
.B(n_235),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_302),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_302),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_265),
.B(n_108),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_268),
.B(n_235),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_229),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_261),
.B(n_235),
.Y(n_343)
);

INVxp33_ASAP7_75t_SL g344 ( 
.A(n_270),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_281),
.B(n_257),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_296),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_308),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_301),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_301),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_289),
.Y(n_351)
);

XOR2x2_ASAP7_75t_L g352 ( 
.A(n_276),
.B(n_252),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_282),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_276),
.B(n_248),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_271),
.B(n_248),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_305),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_275),
.B(n_248),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_285),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_307),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_306),
.B(n_229),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_291),
.B(n_229),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_278),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_290),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_288),
.B(n_229),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_299),
.B(n_213),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_300),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_267),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_267),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_260),
.B(n_252),
.Y(n_374)
);

INVx2_ASAP7_75t_SL g375 ( 
.A(n_259),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_325),
.B(n_252),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_323),
.B(n_232),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_323),
.B(n_232),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_329),
.B(n_215),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_375),
.B(n_337),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_318),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_348),
.A2(n_233),
.B(n_239),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_319),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_320),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_314),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_354),
.B(n_233),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g387 ( 
.A(n_314),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_314),
.Y(n_388)
);

HB1xp67_ASAP7_75t_L g389 ( 
.A(n_311),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_239),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_330),
.B(n_217),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_336),
.B(n_217),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_324),
.B(n_217),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_310),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_312),
.Y(n_396)
);

AND2x2_ASAP7_75t_SL g397 ( 
.A(n_338),
.B(n_217),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_313),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_333),
.B(n_217),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_337),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_361),
.B(n_215),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_311),
.B(n_215),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_372),
.Y(n_404)
);

AND2x4_ASAP7_75t_L g405 ( 
.A(n_356),
.B(n_109),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_373),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_321),
.B(n_215),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_368),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_360),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_341),
.B(n_215),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_357),
.Y(n_411)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_339),
.B(n_245),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_346),
.B(n_245),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_347),
.B(n_245),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_357),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_362),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_341),
.B(n_216),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_349),
.B(n_245),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_343),
.B(n_351),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_216),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_355),
.B(n_216),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_353),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_366),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_350),
.A2(n_216),
.B(n_213),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_345),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_344),
.B(n_327),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_358),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_353),
.A2(n_216),
.B(n_213),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_359),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_370),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_245),
.Y(n_432)
);

OR2x2_ASAP7_75t_SL g433 ( 
.A(n_363),
.B(n_242),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g434 ( 
.A(n_316),
.B(n_326),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_331),
.Y(n_435)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_332),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g437 ( 
.A1(n_342),
.A2(n_213),
.B(n_242),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_315),
.B(n_234),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_365),
.B(n_213),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_340),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_377),
.Y(n_441)
);

BUFx8_ASAP7_75t_SL g442 ( 
.A(n_440),
.Y(n_442)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_420),
.B(n_315),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

BUFx8_ASAP7_75t_SL g445 ( 
.A(n_440),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_383),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_399),
.B(n_435),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_395),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_383),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_401),
.B(n_371),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_377),
.B(n_374),
.Y(n_451)
);

AND2x4_ASAP7_75t_L g452 ( 
.A(n_399),
.B(n_364),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_399),
.B(n_374),
.Y(n_453)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

AND2x4_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_436),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_435),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_378),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_404),
.Y(n_458)
);

BUFx8_ASAP7_75t_L g459 ( 
.A(n_435),
.Y(n_459)
);

AND2x4_ASAP7_75t_L g460 ( 
.A(n_436),
.B(n_317),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_110),
.Y(n_461)
);

OR2x2_ASAP7_75t_L g462 ( 
.A(n_416),
.B(n_352),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_436),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g464 ( 
.A(n_416),
.B(n_328),
.Y(n_464)
);

AND2x2_ASAP7_75t_L g465 ( 
.A(n_389),
.B(n_386),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_378),
.B(n_386),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_427),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_431),
.B(n_334),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_434),
.B(n_334),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_411),
.B(n_242),
.Y(n_470)
);

NAND2x1_ASAP7_75t_SL g471 ( 
.A(n_405),
.B(n_113),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_381),
.Y(n_472)
);

AND2x4_ASAP7_75t_L g473 ( 
.A(n_436),
.B(n_115),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_432),
.Y(n_474)
);

INVx6_ASAP7_75t_L g475 ( 
.A(n_432),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_408),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_411),
.B(n_242),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g478 ( 
.A(n_380),
.B(n_242),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_412),
.Y(n_479)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_431),
.B(n_116),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_430),
.Y(n_482)
);

AND2x4_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_119),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_423),
.B(n_120),
.Y(n_484)
);

CKINVDCx6p67_ASAP7_75t_R g485 ( 
.A(n_460),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_465),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_472),
.Y(n_487)
);

INVx4_ASAP7_75t_L g488 ( 
.A(n_454),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_455),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_472),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_455),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_446),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_449),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_459),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_450),
.A2(n_411),
.B1(n_434),
.B2(n_423),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_459),
.Y(n_496)
);

CKINVDCx16_ASAP7_75t_R g497 ( 
.A(n_469),
.Y(n_497)
);

INVx2_ASAP7_75t_SL g498 ( 
.A(n_464),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_482),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_444),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_454),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_441),
.B(n_411),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_454),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_456),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_456),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_456),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_448),
.Y(n_509)
);

BUFx3_ASAP7_75t_L g510 ( 
.A(n_463),
.Y(n_510)
);

INVx4_ASAP7_75t_L g511 ( 
.A(n_463),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_445),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_462),
.Y(n_513)
);

CKINVDCx6p67_ASAP7_75t_R g514 ( 
.A(n_496),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_487),
.Y(n_515)
);

CKINVDCx6p67_ASAP7_75t_R g516 ( 
.A(n_512),
.Y(n_516)
);

OAI22xp33_ASAP7_75t_L g517 ( 
.A1(n_495),
.A2(n_443),
.B1(n_411),
.B2(n_451),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_502),
.A2(n_408),
.B1(n_417),
.B2(n_468),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_492),
.Y(n_519)
);

INVx2_ASAP7_75t_SL g520 ( 
.A(n_498),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_490),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_493),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_486),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_512),
.Y(n_525)
);

BUFx4f_ASAP7_75t_L g526 ( 
.A(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_500),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_502),
.A2(n_408),
.B1(n_417),
.B2(n_466),
.Y(n_528)
);

OAI22xp33_ASAP7_75t_L g529 ( 
.A1(n_497),
.A2(n_408),
.B1(n_441),
.B2(n_457),
.Y(n_529)
);

INVx6_ASAP7_75t_L g530 ( 
.A(n_489),
.Y(n_530)
);

BUFx2_ASAP7_75t_SL g531 ( 
.A(n_503),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_486),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_509),
.A2(n_453),
.B1(n_438),
.B2(n_457),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_485),
.A2(n_479),
.B1(n_409),
.B2(n_474),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g535 ( 
.A1(n_513),
.A2(n_453),
.B1(n_405),
.B2(n_475),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_SL g536 ( 
.A1(n_513),
.A2(n_405),
.B1(n_475),
.B2(n_473),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_489),
.A2(n_382),
.B(n_410),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_494),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_426),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_519),
.Y(n_540)
);

BUFx12f_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_536),
.A2(n_433),
.B1(n_447),
.B2(n_452),
.Y(n_542)
);

AOI22xp33_ASAP7_75t_L g543 ( 
.A1(n_535),
.A2(n_409),
.B1(n_424),
.B2(n_484),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_517),
.A2(n_409),
.B1(n_424),
.B2(n_484),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_532),
.B(n_409),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_SL g546 ( 
.A1(n_531),
.A2(n_461),
.B1(n_473),
.B2(n_397),
.Y(n_546)
);

BUFx6f_ASAP7_75t_SL g547 ( 
.A(n_520),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_515),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_SL g549 ( 
.A1(n_526),
.A2(n_461),
.B1(n_397),
.B2(n_376),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_539),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_517),
.A2(n_424),
.B1(n_483),
.B2(n_480),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_521),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_533),
.A2(n_424),
.B1(n_483),
.B2(n_415),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_527),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_538),
.B(n_525),
.Y(n_556)
);

AOI22xp33_ASAP7_75t_SL g557 ( 
.A1(n_526),
.A2(n_530),
.B1(n_425),
.B2(n_522),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_533),
.A2(n_414),
.B1(n_419),
.B2(n_413),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_529),
.Y(n_559)
);

AOI22xp33_ASAP7_75t_L g560 ( 
.A1(n_534),
.A2(n_529),
.B1(n_415),
.B2(n_419),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_518),
.B(n_414),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_534),
.Y(n_562)
);

OAI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_528),
.A2(n_429),
.B(n_413),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_522),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_530),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_530),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_528),
.A2(n_390),
.B1(n_403),
.B2(n_394),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_518),
.Y(n_568)
);

AND2x2_ASAP7_75t_L g569 ( 
.A(n_550),
.B(n_491),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_SL g570 ( 
.A1(n_561),
.A2(n_537),
.B1(n_429),
.B2(n_481),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_L g571 ( 
.A1(n_546),
.A2(n_514),
.B1(n_516),
.B2(n_476),
.Y(n_571)
);

OAI22xp33_ASAP7_75t_L g572 ( 
.A1(n_563),
.A2(n_402),
.B1(n_458),
.B2(n_477),
.Y(n_572)
);

OAI221xp5_ASAP7_75t_L g573 ( 
.A1(n_549),
.A2(n_471),
.B1(n_398),
.B2(n_396),
.C(n_404),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_562),
.A2(n_394),
.B1(n_406),
.B2(n_398),
.Y(n_574)
);

OAI221xp5_ASAP7_75t_L g575 ( 
.A1(n_558),
.A2(n_396),
.B1(n_406),
.B2(n_478),
.C(n_421),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_541),
.A2(n_390),
.B1(n_403),
.B2(n_400),
.Y(n_576)
);

OAI221xp5_ASAP7_75t_L g577 ( 
.A1(n_543),
.A2(n_422),
.B1(n_418),
.B2(n_392),
.C(n_384),
.Y(n_577)
);

AOI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_561),
.A2(n_428),
.B1(n_470),
.B2(n_510),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_541),
.A2(n_400),
.B1(n_407),
.B2(n_384),
.Y(n_579)
);

OAI22xp33_ASAP7_75t_L g580 ( 
.A1(n_559),
.A2(n_428),
.B1(n_510),
.B2(n_511),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_428),
.B1(n_488),
.B2(n_511),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_407),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_L g583 ( 
.A1(n_560),
.A2(n_488),
.B1(n_505),
.B2(n_507),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g584 ( 
.A1(n_553),
.A2(n_505),
.B1(n_507),
.B2(n_508),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_542),
.A2(n_381),
.B1(n_391),
.B2(n_379),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_551),
.A2(n_385),
.B1(n_393),
.B2(n_388),
.Y(n_586)
);

OAI211xp5_ASAP7_75t_L g587 ( 
.A1(n_557),
.A2(n_437),
.B(n_507),
.C(n_504),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_552),
.B(n_508),
.Y(n_588)
);

OAI221xp5_ASAP7_75t_SL g589 ( 
.A1(n_545),
.A2(n_385),
.B1(n_393),
.B2(n_388),
.C(n_123),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_L g590 ( 
.A1(n_568),
.A2(n_508),
.B1(n_507),
.B2(n_504),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_547),
.A2(n_508),
.B1(n_504),
.B2(n_501),
.Y(n_591)
);

NAND3xp33_ASAP7_75t_L g592 ( 
.A(n_589),
.B(n_548),
.C(n_540),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_569),
.B(n_554),
.Y(n_593)
);

NAND3xp33_ASAP7_75t_L g594 ( 
.A(n_573),
.B(n_548),
.C(n_555),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_582),
.B(n_554),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_588),
.B(n_555),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_564),
.Y(n_597)
);

OAI22xp5_ASAP7_75t_L g598 ( 
.A1(n_571),
.A2(n_547),
.B1(n_568),
.B2(n_565),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_570),
.B(n_578),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_574),
.B(n_564),
.Y(n_600)
);

NOR3xp33_ASAP7_75t_L g601 ( 
.A(n_587),
.B(n_565),
.C(n_556),
.Y(n_601)
);

OAI22xp5_ASAP7_75t_L g602 ( 
.A1(n_579),
.A2(n_576),
.B1(n_575),
.B2(n_547),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_590),
.B(n_565),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_580),
.B(n_566),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_580),
.B(n_566),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_593),
.B(n_585),
.Y(n_606)
);

OR2x2_ASAP7_75t_L g607 ( 
.A(n_596),
.B(n_584),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_601),
.B(n_566),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_595),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_597),
.B(n_591),
.Y(n_610)
);

NOR2x1_ASAP7_75t_L g611 ( 
.A(n_594),
.B(n_577),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_603),
.B(n_566),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_604),
.B(n_566),
.Y(n_613)
);

AND4x1_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_592),
.C(n_599),
.D(n_605),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_609),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_612),
.Y(n_616)
);

XOR2x2_ASAP7_75t_L g617 ( 
.A(n_608),
.B(n_598),
.Y(n_617)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_607),
.B(n_600),
.Y(n_618)
);

NOR2x1_ASAP7_75t_L g619 ( 
.A(n_610),
.B(n_602),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_613),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_615),
.Y(n_621)
);

OR2x6_ASAP7_75t_L g622 ( 
.A(n_619),
.B(n_613),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_618),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_616),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_620),
.Y(n_625)
);

XNOR2x1_ASAP7_75t_L g626 ( 
.A(n_622),
.B(n_617),
.Y(n_626)
);

HB1xp67_ASAP7_75t_L g627 ( 
.A(n_623),
.Y(n_627)
);

OA22x2_ASAP7_75t_L g628 ( 
.A1(n_622),
.A2(n_620),
.B1(n_614),
.B2(n_583),
.Y(n_628)
);

XOR2x2_ASAP7_75t_L g629 ( 
.A(n_625),
.B(n_614),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_621),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_627),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_630),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_630),
.Y(n_633)
);

AOI221xp5_ASAP7_75t_L g634 ( 
.A1(n_631),
.A2(n_621),
.B1(n_626),
.B2(n_624),
.C(n_629),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_631),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_635),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_636),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_637),
.Y(n_638)
);

NAND4xp25_ASAP7_75t_L g639 ( 
.A(n_638),
.B(n_634),
.C(n_633),
.D(n_632),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_639),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_640),
.A2(n_628),
.B1(n_623),
.B2(n_606),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_641),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_642),
.A2(n_581),
.B1(n_504),
.B2(n_501),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_643),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g645 ( 
.A1(n_644),
.A2(n_586),
.B1(n_501),
.B2(n_567),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_645),
.Y(n_646)
);

AOI221xp5_ASAP7_75t_L g647 ( 
.A1(n_646),
.A2(n_387),
.B1(n_439),
.B2(n_130),
.C(n_136),
.Y(n_647)
);

AOI211xp5_ASAP7_75t_L g648 ( 
.A1(n_647),
.A2(n_125),
.B(n_127),
.C(n_137),
.Y(n_648)
);


endmodule