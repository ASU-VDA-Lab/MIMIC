module real_jpeg_23033_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_0),
.B(n_28),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_0),
.B(n_55),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_0),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_0),
.B(n_113),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_0),
.B(n_25),
.Y(n_182)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_2),
.B(n_28),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_32),
.Y(n_31)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_2),
.B(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_4),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_7),
.B(n_35),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_7),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_7),
.B(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_7),
.B(n_73),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_7),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_7),
.B(n_28),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_7),
.B(n_25),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_8),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_8),
.B(n_28),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_32),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g252 ( 
.A(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_8),
.B(n_113),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_8),
.B(n_73),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_8),
.B(n_55),
.Y(n_335)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_10),
.B(n_35),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_10),
.B(n_25),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_10),
.B(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_10),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_10),
.B(n_73),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_10),
.B(n_55),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_10),
.B(n_32),
.Y(n_334)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_12),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_12),
.B(n_113),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_12),
.B(n_73),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_12),
.B(n_55),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_12),
.B(n_32),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_12),
.B(n_28),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_12),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_12),
.B(n_254),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_13),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_13),
.B(n_73),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_13),
.B(n_55),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_13),
.B(n_32),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_13),
.B(n_28),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_13),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_13),
.B(n_254),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_14),
.B(n_55),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_14),
.B(n_32),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_14),
.B(n_73),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_14),
.B(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_14),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_14),
.B(n_28),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_14),
.B(n_25),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_14),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_15),
.B(n_35),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_15),
.B(n_121),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_15),
.B(n_113),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_15),
.B(n_73),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_15),
.B(n_32),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_15),
.B(n_28),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_73),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_16),
.B(n_55),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_16),
.B(n_113),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_16),
.B(n_121),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_16),
.B(n_32),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_16),
.B(n_28),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_16),
.B(n_25),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_16),
.B(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_17),
.Y(n_110)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_17),
.Y(n_122)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_17),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_57),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_44),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_33),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_26),
.C(n_31),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_23),
.A2(n_24),
.B1(n_46),
.B2(n_47),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_27),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_27),
.B1(n_31),
.B2(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_31),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_31),
.B(n_51),
.C(n_53),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_31),
.A2(n_48),
.B1(n_53),
.B2(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_32),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_39),
.Y(n_33)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_38),
.B(n_153),
.Y(n_214)
);

INVx11_ASAP7_75t_L g254 ( 
.A(n_38),
.Y(n_254)
);

INVx8_ASAP7_75t_L g272 ( 
.A(n_38),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_42),
.B(n_267),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_42),
.B(n_299),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_43),
.B(n_277),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_43),
.B(n_250),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_49),
.C(n_50),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_50),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_52),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_SL g69 ( 
.A(n_53),
.B(n_70),
.C(n_72),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_53),
.A2(n_72),
.B1(n_77),
.B2(n_330),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_54),
.B(n_228),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_54),
.B(n_71),
.Y(n_262)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_79),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_58),
.B(n_380),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_69),
.C(n_75),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_59),
.B(n_374),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_60),
.B(n_79),
.Y(n_380)
);

FAx1_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.CI(n_63),
.CON(n_60),
.SN(n_60)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.C(n_67),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_64),
.B(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_65),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_69),
.B(n_75),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_70),
.B(n_355),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g329 ( 
.A1(n_72),
.A2(n_301),
.B1(n_302),
.B2(n_330),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_72),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_SL g359 ( 
.A(n_72),
.B(n_301),
.C(n_328),
.Y(n_359)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_73),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_378),
.C(n_379),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_369),
.C(n_370),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_347),
.C(n_348),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_323),
.C(n_324),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_291),
.C(n_292),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_256),
.C(n_257),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_220),
.C(n_221),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_189),
.C(n_190),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_164),
.C(n_165),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_124),
.C(n_136),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_100),
.C(n_105),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.C(n_98),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_94),
.A2(n_95),
.B1(n_126),
.B2(n_127),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_99),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_101),
.B(n_103),
.C(n_104),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_115),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_106),
.B(n_116),
.C(n_117),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_107),
.B(n_111),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_110),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g250 ( 
.A(n_113),
.Y(n_250)
);

BUFx12f_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_117),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_123),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_118),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_123),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_128),
.C(n_135),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_125),
.B(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_129),
.B1(n_135),
.B2(n_163),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_140)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_134),
.Y(n_277)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_135),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_160),
.C(n_161),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_145),
.C(n_150),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_143),
.C(n_144),
.Y(n_160)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_146),
.B(n_148),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_149),
.Y(n_151)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.C(n_155),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_159),
.B(n_252),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_178),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_179),
.C(n_188),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_174),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_173),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_173),
.C(n_174),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_172),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx24_ASAP7_75t_SL g385 ( 
.A(n_174),
.Y(n_385)
);

FAx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.CI(n_177),
.CON(n_174),
.SN(n_174)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_176),
.C(n_177),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_186),
.B2(n_187),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_182),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_185),
.C(n_187),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_186),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_205),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_194),
.C(n_205),
.Y(n_220)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_196),
.B(n_201),
.C(n_204),
.Y(n_224)
);

BUFx24_ASAP7_75t_SL g382 ( 
.A(n_196),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_198),
.CI(n_199),
.CON(n_196),
.SN(n_196)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_198),
.C(n_199),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_203),
.B2(n_204),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_206),
.B(n_213),
.C(n_218),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_208),
.A2(n_213),
.B1(n_218),
.B2(n_219),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_208),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B(n_212),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_211),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_212),
.B(n_245),
.C(n_246),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_213),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_214),
.B(n_216),
.C(n_217),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_241),
.B2(n_255),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_242),
.C(n_243),
.Y(n_256)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_226),
.C(n_234),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_234),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_229),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_227),
.B(n_230),
.C(n_233),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_228),
.B(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_232),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_240),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_237),
.B1(n_238),
.B2(n_239),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_238),
.Y(n_239)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_247),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_287),
.C(n_288),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_251),
.CI(n_253),
.CON(n_247),
.SN(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_289),
.B2(n_290),
.Y(n_257)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_258),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_259),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_281),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_260),
.B(n_281),
.C(n_289),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_268),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_261),
.B(n_269),
.C(n_270),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_262),
.B(n_264),
.C(n_266),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_280),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_271),
.Y(n_280)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_279),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_275),
.A2(n_276),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_279),
.C(n_280),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_275),
.B(n_298),
.C(n_301),
.Y(n_345)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_282),
.B(n_284),
.C(n_285),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_293),
.B(n_295),
.C(n_322),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_309),
.B2(n_322),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_303),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_297),
.B(n_304),
.C(n_305),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_301),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_305),
.Y(n_381)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_307),
.CI(n_308),
.CON(n_305),
.SN(n_305)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_306),
.B(n_307),
.C(n_308),
.Y(n_332)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_312),
.C(n_313),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_313),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_316),
.B2(n_321),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_317),
.C(n_319),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_316),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_317),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_319),
.B1(n_343),
.B2(n_344),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_344),
.C(n_345),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_346),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_337),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_337),
.C(n_346),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_331),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_332),
.C(n_333),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_333),
.Y(n_331)
);

BUFx24_ASAP7_75t_SL g383 ( 
.A(n_333),
.Y(n_383)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_334),
.B(n_335),
.CI(n_336),
.CON(n_333),
.SN(n_333)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_335),
.C(n_336),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_338),
.B(n_339),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_338),
.B(n_340),
.C(n_341),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_341),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_345),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_343),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_351),
.C(n_361),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_352),
.B1(n_360),
.B2(n_361),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_356),
.B2(n_357),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_353),
.B(n_358),
.C(n_359),
.Y(n_372)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_363),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_364),
.C(n_367),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_364),
.A2(n_365),
.B1(n_366),
.B2(n_367),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_367),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_371),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_370)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_371),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_372),
.B(n_373),
.C(n_377),
.Y(n_378)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_375),
.Y(n_377)
);


endmodule