module real_jpeg_3385_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_1),
.B(n_52),
.Y(n_58)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_50),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_1),
.B(n_27),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_1),
.B(n_25),
.Y(n_133)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_2),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_2),
.B(n_27),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_4),
.B(n_31),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_4),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_4),
.B(n_52),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_4),
.B(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_4),
.B(n_27),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_4),
.B(n_25),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_5),
.B(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_5),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_5),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_5),
.B(n_52),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_8),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_8),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_35),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_8),
.B(n_52),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_8),
.B(n_50),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_9),
.B(n_25),
.Y(n_100)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_25),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_13),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_14),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_SL g98 ( 
.A(n_14),
.B(n_27),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_111),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_109),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_92),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_19),
.B(n_92),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_55),
.Y(n_19)
);

BUFx24_ASAP7_75t_SL g171 ( 
.A(n_20),
.Y(n_171)
);

FAx1_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_37),
.CI(n_41),
.CON(n_20),
.SN(n_20)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_30),
.C(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_22),
.A2(n_23),
.B1(n_107),
.B2(n_108),
.Y(n_106)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_26),
.Y(n_23)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_24),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_28),
.B(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_30),
.B(n_34),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_39),
.B(n_40),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_43),
.B(n_73),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_43),
.B(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_54),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_50),
.Y(n_153)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_75),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_65),
.C(n_69),
.Y(n_56)
);

FAx1_ASAP7_75t_SL g94 ( 
.A(n_57),
.B(n_65),
.CI(n_69),
.CON(n_94),
.SN(n_94)
);

XOR2xp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_59),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_61),
.C(n_62),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_62),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g79 ( 
.A(n_63),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.C(n_68),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_66),
.B(n_68),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_67),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_77),
.B1(n_86),
.B2(n_91),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_81),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_82),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_86),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_88),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_95),
.C(n_106),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_93),
.A2(n_94),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g174 ( 
.A(n_94),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_95),
.B(n_106),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_101),
.C(n_102),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_96),
.B(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g124 ( 
.A(n_102),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_165),
.B(n_170),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_135),
.B(n_164),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_114),
.B(n_126),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_114),
.B(n_126),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_124),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_120),
.B1(n_122),
.B2(n_123),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_118),
.C(n_119),
.Y(n_116)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_117),
.B(n_118),
.CI(n_119),
.CON(n_127),
.SN(n_127)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_120),
.B(n_122),
.C(n_124),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.C(n_134),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_127),
.B(n_161),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_127),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_131),
.B1(n_132),
.B2(n_133),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_158),
.B(n_163),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_148),
.B(n_157),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_138),
.B(n_143),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_143),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_140),
.B(n_141),
.C(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_144),
.B(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_146),
.B1(n_147),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_151),
.B(n_156),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_154),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_159),
.B(n_160),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_166),
.B(n_167),
.Y(n_170)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);


endmodule