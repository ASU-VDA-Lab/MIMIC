module fake_jpeg_27825_n_274 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_274);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_274;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx5_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_6),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_30),
.Y(n_45)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_15),
.Y(n_29)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

OR2x2_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_33),
.B(n_26),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_38),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_42),
.B(n_30),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_32),
.Y(n_61)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_49),
.Y(n_82)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_32),
.B1(n_33),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_57),
.B1(n_28),
.B2(n_44),
.Y(n_77)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_54),
.Y(n_79)
);

NAND2x1_ASAP7_75t_SL g55 ( 
.A(n_47),
.B(n_35),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_27),
.B(n_30),
.C(n_26),
.Y(n_75)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_33),
.B1(n_28),
.B2(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_44),
.A2(n_21),
.B1(n_15),
.B2(n_23),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_45),
.B(n_30),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_64),
.A2(n_66),
.B1(n_35),
.B2(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_51),
.B(n_31),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_71),
.B(n_36),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g73 ( 
.A(n_51),
.B(n_27),
.C(n_47),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_55),
.C(n_31),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g74 ( 
.A1(n_57),
.A2(n_43),
.B1(n_31),
.B2(n_41),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_74),
.A2(n_55),
.B1(n_41),
.B2(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_74),
.Y(n_89)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_60),
.A2(n_29),
.A3(n_36),
.B1(n_34),
.B2(n_28),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_48),
.B1(n_38),
.B2(n_41),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_83),
.A2(n_52),
.B1(n_59),
.B2(n_49),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_86),
.A2(n_92),
.B1(n_95),
.B2(n_98),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_87),
.B(n_81),
.Y(n_120)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVxp33_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_89),
.A2(n_74),
.B1(n_73),
.B2(n_84),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_68),
.A2(n_58),
.B1(n_50),
.B2(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_65),
.Y(n_93)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g124 ( 
.A(n_94),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_83),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_97),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_77),
.A2(n_15),
.B1(n_21),
.B2(n_56),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_65),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_75),
.Y(n_113)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_101),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_82),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_102),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_54),
.B1(n_39),
.B2(n_65),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_103),
.A2(n_70),
.B1(n_69),
.B2(n_82),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_104),
.A2(n_67),
.B(n_81),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_93),
.B(n_80),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_106),
.A2(n_107),
.B(n_111),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_109),
.A2(n_116),
.B1(n_106),
.B2(n_115),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_75),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_113),
.B(n_121),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_85),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_114),
.B(n_120),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_89),
.A2(n_97),
.B1(n_91),
.B2(n_96),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_93),
.B(n_86),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_118),
.A2(n_121),
.B(n_106),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_74),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVxp67_ASAP7_75t_SL g143 ( 
.A(n_122),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_123),
.A2(n_88),
.B1(n_94),
.B2(n_100),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_127),
.A2(n_129),
.B1(n_132),
.B2(n_134),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_119),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_110),
.A2(n_87),
.B1(n_86),
.B2(n_92),
.Y(n_129)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_118),
.A2(n_104),
.B(n_90),
.Y(n_130)
);

OA21x2_ASAP7_75t_L g165 ( 
.A1(n_130),
.A2(n_131),
.B(n_137),
.Y(n_165)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_111),
.A2(n_92),
.B(n_99),
.C(n_95),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_110),
.A2(n_98),
.B1(n_103),
.B2(n_94),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_113),
.B(n_20),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_18),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_88),
.B1(n_72),
.B2(n_102),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_107),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_140),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_145),
.B1(n_140),
.B2(n_117),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_72),
.C(n_101),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_142),
.C(n_106),
.Y(n_155)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_139),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_101),
.C(n_70),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_109),
.A2(n_82),
.B1(n_65),
.B2(n_79),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_79),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_115),
.B(n_18),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_116),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_150),
.B(n_22),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_138),
.B(n_112),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_151),
.B(n_152),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_166),
.B(n_133),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_170),
.C(n_130),
.Y(n_184)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_143),
.Y(n_158)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_129),
.A2(n_132),
.B1(n_148),
.B2(n_135),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_160),
.A2(n_162),
.B1(n_169),
.B2(n_145),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_136),
.A2(n_125),
.B1(n_121),
.B2(n_105),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_125),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_163),
.B(n_144),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_134),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_171),
.Y(n_177)
);

AOI21x1_ASAP7_75t_SL g166 ( 
.A1(n_131),
.A2(n_124),
.B(n_119),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_142),
.B(n_29),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_167),
.B(n_168),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_126),
.B(n_29),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_131),
.A2(n_19),
.B1(n_14),
.B2(n_17),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_146),
.B(n_29),
.C(n_25),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_22),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_141),
.A2(n_10),
.B(n_1),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_172),
.A2(n_13),
.B(n_1),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_179),
.B1(n_165),
.B2(n_19),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_141),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_183),
.Y(n_197)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_178),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_156),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_159),
.A2(n_144),
.B1(n_128),
.B2(n_137),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_180),
.B(n_160),
.Y(n_196)
);

OR2x2_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_193),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_151),
.B(n_130),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_189),
.C(n_191),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_157),
.B(n_127),
.Y(n_185)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_130),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_186),
.B(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_19),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_34),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_188),
.B(n_172),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_168),
.C(n_152),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_25),
.C(n_24),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_13),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_166),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_201),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_161),
.B1(n_158),
.B2(n_159),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_198),
.A2(n_202),
.B1(n_191),
.B2(n_181),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_165),
.C(n_149),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_199),
.B(n_210),
.C(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_203),
.B(n_17),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_174),
.B(n_13),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_205),
.B(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_34),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_17),
.B1(n_14),
.B2(n_2),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_177),
.A2(n_24),
.B1(n_19),
.B2(n_17),
.Y(n_208)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_24),
.Y(n_209)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_175),
.B(n_25),
.C(n_24),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_223),
.B1(n_7),
.B2(n_2),
.Y(n_236)
);

MAJx2_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_7),
.C(n_3),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_211),
.A2(n_187),
.B1(n_190),
.B2(n_189),
.Y(n_216)
);

OR2x2_ASAP7_75t_L g239 ( 
.A(n_216),
.B(n_8),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_175),
.C(n_190),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_218),
.C(n_215),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_194),
.B(n_180),
.C(n_193),
.Y(n_218)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_204),
.Y(n_219)
);

BUFx24_ASAP7_75t_SL g228 ( 
.A(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_222),
.B(n_199),
.Y(n_230)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_196),
.B(n_14),
.CI(n_1),
.CON(n_225),
.SN(n_225)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_195),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_224),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_230),
.B(n_234),
.Y(n_246)
);

NOR2x1_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_204),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_231),
.B(n_235),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_232),
.A2(n_239),
.B(n_5),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_213),
.A2(n_197),
.B(n_198),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_233),
.A2(n_237),
.B(n_225),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_221),
.B(n_201),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_210),
.C(n_2),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_236),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_220),
.A2(n_7),
.B(n_3),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_238),
.B(n_222),
.C(n_212),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_241),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_247),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_231),
.A2(n_212),
.B1(n_3),
.B2(n_4),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_8),
.B1(n_3),
.B2(n_4),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_239),
.B(n_8),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_227),
.A2(n_8),
.B(n_4),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_248),
.A2(n_238),
.B(n_9),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_251),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_228),
.B(n_9),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_11),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_246),
.A2(n_9),
.B(n_10),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_256),
.B(n_11),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_243),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_244),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g267 ( 
.A1(n_260),
.A2(n_258),
.B(n_264),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_253),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_262),
.B(n_263),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_SL g262 ( 
.A1(n_257),
.A2(n_240),
.B(n_245),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_265),
.B(n_254),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_252),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_259),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_270),
.B(n_268),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_271),
.B(n_11),
.C(n_12),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_272),
.B(n_0),
.C(n_12),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_273),
.B(n_12),
.Y(n_274)
);


endmodule