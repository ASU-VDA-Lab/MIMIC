module fake_jpeg_28145_n_37 (n_3, n_2, n_1, n_0, n_4, n_5, n_37);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_37;

wire n_13;
wire n_21;
wire n_33;
wire n_23;
wire n_10;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NOR2xp33_ASAP7_75t_L g6 ( 
.A(n_4),
.B(n_2),
.Y(n_6)
);

INVx8_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_0),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_SL g11 ( 
.A(n_0),
.B(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_13),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_11),
.B(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_11),
.B(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx10_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_17),
.A2(n_8),
.B1(n_12),
.B2(n_9),
.Y(n_22)
);

A2O1A1Ixp33_ASAP7_75t_L g18 ( 
.A1(n_8),
.A2(n_3),
.B(n_4),
.C(n_5),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g25 ( 
.A1(n_18),
.A2(n_19),
.B(n_9),
.Y(n_25)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

AOI21xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_25),
.B(n_18),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_29),
.C(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_13),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

A2O1A1Ixp33_ASAP7_75t_SL g29 ( 
.A1(n_23),
.A2(n_10),
.B(n_0),
.C(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_29),
.Y(n_32)
);

AOI31xp67_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_10),
.A3(n_0),
.B(n_7),
.Y(n_35)
);

AOI322xp5_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_23),
.A3(n_20),
.B1(n_29),
.B2(n_7),
.C1(n_21),
.C2(n_24),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_34),
.A2(n_35),
.B(n_31),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_10),
.B(n_31),
.Y(n_37)
);


endmodule