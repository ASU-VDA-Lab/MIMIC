module fake_ibex_723_n_7788 (n_151, n_85, n_599, n_778, n_822, n_1042, n_507, n_743, n_1060, n_540, n_754, n_395, n_1011, n_84, n_64, n_992, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_1041, n_688, n_130, n_177, n_946, n_707, n_76, n_273, n_309, n_330, n_926, n_9, n_1079, n_1031, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_845, n_947, n_972, n_981, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_956, n_790, n_920, n_452, n_86, n_70, n_664, n_1067, n_255, n_175, n_586, n_773, n_994, n_638, n_398, n_59, n_28, n_125, n_304, n_821, n_191, n_873, n_962, n_593, n_5, n_62, n_71, n_153, n_862, n_545, n_909, n_583, n_887, n_1080, n_957, n_1015, n_678, n_663, n_969, n_194, n_249, n_334, n_634, n_733, n_961, n_991, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_1034, n_371, n_974, n_1036, n_403, n_872, n_423, n_608, n_864, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_930, n_336, n_959, n_258, n_861, n_1018, n_1044, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_1077, n_43, n_216, n_996, n_915, n_911, n_33, n_652, n_781, n_421, n_828, n_738, n_475, n_802, n_166, n_163, n_1045, n_753, n_645, n_500, n_747, n_963, n_542, n_114, n_236, n_900, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_901, n_105, n_187, n_667, n_884, n_1061, n_1, n_154, n_682, n_850, n_182, n_196, n_326, n_327, n_879, n_89, n_1056, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_886, n_840, n_1010, n_561, n_883, n_117, n_417, n_471, n_846, n_739, n_755, n_265, n_853, n_504, n_948, n_158, n_1029, n_859, n_259, n_276, n_339, n_470, n_770, n_965, n_210, n_348, n_220, n_875, n_941, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_876, n_147, n_552, n_251, n_384, n_632, n_989, n_373, n_1051, n_854, n_1008, n_458, n_244, n_73, n_1053, n_343, n_310, n_714, n_1076, n_1032, n_936, n_703, n_426, n_323, n_469, n_829, n_598, n_825, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_939, n_67, n_453, n_591, n_898, n_655, n_333, n_928, n_967, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_1055, n_10, n_673, n_21, n_732, n_798, n_832, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_893, n_590, n_1025, n_465, n_1057, n_1068, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_914, n_120, n_1013, n_982, n_835, n_168, n_526, n_785, n_155, n_824, n_929, n_315, n_441, n_604, n_1024, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_977, n_1075, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_865, n_923, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_907, n_51, n_933, n_1081, n_215, n_279, n_49, n_1037, n_374, n_235, n_464, n_538, n_669, n_838, n_987, n_750, n_1021, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_1052, n_852, n_789, n_880, n_654, n_656, n_1014, n_724, n_437, n_731, n_602, n_904, n_842, n_938, n_355, n_767, n_474, n_878, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_1023, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_944, n_1001, n_156, n_570, n_126, n_623, n_585, n_1030, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_1082, n_222, n_660, n_186, n_524, n_349, n_765, n_849, n_857, n_980, n_454, n_1070, n_1074, n_777, n_1017, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_917, n_185, n_388, n_953, n_625, n_968, n_619, n_536, n_611, n_352, n_290, n_558, n_931, n_666, n_174, n_467, n_427, n_607, n_827, n_157, n_219, n_246, n_31, n_442, n_146, n_1064, n_1071, n_207, n_922, n_438, n_851, n_993, n_1012, n_1028, n_689, n_960, n_1022, n_793, n_167, n_676, n_128, n_937, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_973, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_999, n_1038, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_910, n_1009, n_635, n_979, n_844, n_1066, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_1020, n_847, n_830, n_1062, n_1004, n_473, n_1027, n_445, n_629, n_335, n_413, n_1072, n_82, n_263, n_1069, n_27, n_573, n_353, n_966, n_359, n_826, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_949, n_1007, n_924, n_643, n_137, n_679, n_841, n_772, n_810, n_768, n_839, n_338, n_173, n_696, n_796, n_797, n_837, n_477, n_640, n_954, n_363, n_1006, n_402, n_725, n_180, n_369, n_976, n_596, n_201, n_699, n_14, n_1063, n_351, n_368, n_456, n_834, n_257, n_77, n_998, n_935, n_869, n_925, n_718, n_801, n_918, n_1054, n_44, n_672, n_1039, n_722, n_401, n_1046, n_553, n_554, n_1078, n_1043, n_66, n_735, n_305, n_882, n_942, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_955, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_943, n_1049, n_763, n_745, n_329, n_447, n_940, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_868, n_546, n_199, n_788, n_795, n_1065, n_592, n_986, n_495, n_762, n_410, n_905, n_308, n_975, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_927, n_934, n_658, n_512, n_615, n_950, n_685, n_1026, n_283, n_366, n_397, n_111, n_803, n_894, n_1033, n_692, n_36, n_627, n_990, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_888, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_971, n_101, n_190, n_906, n_138, n_650, n_776, n_409, n_582, n_978, n_818, n_653, n_214, n_238, n_579, n_843, n_899, n_1019, n_1059, n_902, n_332, n_799, n_517, n_211, n_744, n_817, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_881, n_272, n_951, n_511, n_23, n_734, n_468, n_223, n_381, n_1073, n_525, n_815, n_919, n_780, n_535, n_1002, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_863, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_819, n_161, n_237, n_29, n_203, n_268, n_440, n_858, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_952, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_997, n_833, n_217, n_324, n_391, n_831, n_537, n_728, n_78, n_805, n_670, n_820, n_20, n_69, n_892, n_390, n_544, n_891, n_913, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_1016, n_282, n_61, n_680, n_501, n_809, n_752, n_856, n_668, n_779, n_871, n_266, n_42, n_294, n_112, n_958, n_485, n_870, n_46, n_284, n_811, n_1047, n_808, n_80, n_172, n_250, n_945, n_493, n_460, n_609, n_1040, n_476, n_792, n_461, n_575, n_313, n_903, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_1048, n_319, n_195, n_885, n_513, n_212, n_588, n_877, n_693, n_311, n_860, n_661, n_848, n_406, n_606, n_737, n_896, n_97, n_197, n_528, n_181, n_1005, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_836, n_462, n_302, n_450, n_443, n_686, n_985, n_572, n_867, n_983, n_1003, n_644, n_577, n_344, n_393, n_889, n_897, n_436, n_428, n_970, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_816, n_874, n_890, n_912, n_921, n_83, n_32, n_1058, n_107, n_149, n_489, n_677, n_399, n_254, n_908, n_213, n_964, n_424, n_565, n_916, n_823, n_701, n_271, n_995, n_241, n_68, n_503, n_292, n_807, n_984, n_394, n_79, n_1000, n_81, n_35, n_364, n_687, n_895, n_988, n_159, n_202, n_231, n_298, n_587, n_1035, n_760, n_751, n_806, n_932, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_855, n_232, n_380, n_749, n_281, n_866, n_559, n_425, n_1050, n_7788);

input n_151;
input n_85;
input n_599;
input n_778;
input n_822;
input n_1042;
input n_507;
input n_743;
input n_1060;
input n_540;
input n_754;
input n_395;
input n_1011;
input n_84;
input n_64;
input n_992;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_1041;
input n_688;
input n_130;
input n_177;
input n_946;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_926;
input n_9;
input n_1079;
input n_1031;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_845;
input n_947;
input n_972;
input n_981;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_956;
input n_790;
input n_920;
input n_452;
input n_86;
input n_70;
input n_664;
input n_1067;
input n_255;
input n_175;
input n_586;
input n_773;
input n_994;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_821;
input n_191;
input n_873;
input n_962;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_862;
input n_545;
input n_909;
input n_583;
input n_887;
input n_1080;
input n_957;
input n_1015;
input n_678;
input n_663;
input n_969;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_961;
input n_991;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_1034;
input n_371;
input n_974;
input n_1036;
input n_403;
input n_872;
input n_423;
input n_608;
input n_864;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_930;
input n_336;
input n_959;
input n_258;
input n_861;
input n_1018;
input n_1044;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_1077;
input n_43;
input n_216;
input n_996;
input n_915;
input n_911;
input n_33;
input n_652;
input n_781;
input n_421;
input n_828;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_1045;
input n_753;
input n_645;
input n_500;
input n_747;
input n_963;
input n_542;
input n_114;
input n_236;
input n_900;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_901;
input n_105;
input n_187;
input n_667;
input n_884;
input n_1061;
input n_1;
input n_154;
input n_682;
input n_850;
input n_182;
input n_196;
input n_326;
input n_327;
input n_879;
input n_89;
input n_1056;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_886;
input n_840;
input n_1010;
input n_561;
input n_883;
input n_117;
input n_417;
input n_471;
input n_846;
input n_739;
input n_755;
input n_265;
input n_853;
input n_504;
input n_948;
input n_158;
input n_1029;
input n_859;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_965;
input n_210;
input n_348;
input n_220;
input n_875;
input n_941;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_876;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_989;
input n_373;
input n_1051;
input n_854;
input n_1008;
input n_458;
input n_244;
input n_73;
input n_1053;
input n_343;
input n_310;
input n_714;
input n_1076;
input n_1032;
input n_936;
input n_703;
input n_426;
input n_323;
input n_469;
input n_829;
input n_598;
input n_825;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_939;
input n_67;
input n_453;
input n_591;
input n_898;
input n_655;
input n_333;
input n_928;
input n_967;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_1055;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_832;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_893;
input n_590;
input n_1025;
input n_465;
input n_1057;
input n_1068;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_914;
input n_120;
input n_1013;
input n_982;
input n_835;
input n_168;
input n_526;
input n_785;
input n_155;
input n_824;
input n_929;
input n_315;
input n_441;
input n_604;
input n_1024;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_977;
input n_1075;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_865;
input n_923;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_907;
input n_51;
input n_933;
input n_1081;
input n_215;
input n_279;
input n_49;
input n_1037;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_838;
input n_987;
input n_750;
input n_1021;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_1052;
input n_852;
input n_789;
input n_880;
input n_654;
input n_656;
input n_1014;
input n_724;
input n_437;
input n_731;
input n_602;
input n_904;
input n_842;
input n_938;
input n_355;
input n_767;
input n_474;
input n_878;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_1023;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_944;
input n_1001;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_1030;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_1082;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_849;
input n_857;
input n_980;
input n_454;
input n_1070;
input n_1074;
input n_777;
input n_1017;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_917;
input n_185;
input n_388;
input n_953;
input n_625;
input n_968;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_931;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_827;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_1064;
input n_1071;
input n_207;
input n_922;
input n_438;
input n_851;
input n_993;
input n_1012;
input n_1028;
input n_689;
input n_960;
input n_1022;
input n_793;
input n_167;
input n_676;
input n_128;
input n_937;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_973;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_999;
input n_1038;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_910;
input n_1009;
input n_635;
input n_979;
input n_844;
input n_1066;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_1020;
input n_847;
input n_830;
input n_1062;
input n_1004;
input n_473;
input n_1027;
input n_445;
input n_629;
input n_335;
input n_413;
input n_1072;
input n_82;
input n_263;
input n_1069;
input n_27;
input n_573;
input n_353;
input n_966;
input n_359;
input n_826;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_949;
input n_1007;
input n_924;
input n_643;
input n_137;
input n_679;
input n_841;
input n_772;
input n_810;
input n_768;
input n_839;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_837;
input n_477;
input n_640;
input n_954;
input n_363;
input n_1006;
input n_402;
input n_725;
input n_180;
input n_369;
input n_976;
input n_596;
input n_201;
input n_699;
input n_14;
input n_1063;
input n_351;
input n_368;
input n_456;
input n_834;
input n_257;
input n_77;
input n_998;
input n_935;
input n_869;
input n_925;
input n_718;
input n_801;
input n_918;
input n_1054;
input n_44;
input n_672;
input n_1039;
input n_722;
input n_401;
input n_1046;
input n_553;
input n_554;
input n_1078;
input n_1043;
input n_66;
input n_735;
input n_305;
input n_882;
input n_942;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_955;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_943;
input n_1049;
input n_763;
input n_745;
input n_329;
input n_447;
input n_940;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_868;
input n_546;
input n_199;
input n_788;
input n_795;
input n_1065;
input n_592;
input n_986;
input n_495;
input n_762;
input n_410;
input n_905;
input n_308;
input n_975;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_927;
input n_934;
input n_658;
input n_512;
input n_615;
input n_950;
input n_685;
input n_1026;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_894;
input n_1033;
input n_692;
input n_36;
input n_627;
input n_990;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_888;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_971;
input n_101;
input n_190;
input n_906;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_978;
input n_818;
input n_653;
input n_214;
input n_238;
input n_579;
input n_843;
input n_899;
input n_1019;
input n_1059;
input n_902;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_817;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_881;
input n_272;
input n_951;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_1073;
input n_525;
input n_815;
input n_919;
input n_780;
input n_535;
input n_1002;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_863;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_819;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_858;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_952;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_997;
input n_833;
input n_217;
input n_324;
input n_391;
input n_831;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_820;
input n_20;
input n_69;
input n_892;
input n_390;
input n_544;
input n_891;
input n_913;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_1016;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_856;
input n_668;
input n_779;
input n_871;
input n_266;
input n_42;
input n_294;
input n_112;
input n_958;
input n_485;
input n_870;
input n_46;
input n_284;
input n_811;
input n_1047;
input n_808;
input n_80;
input n_172;
input n_250;
input n_945;
input n_493;
input n_460;
input n_609;
input n_1040;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_903;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_1048;
input n_319;
input n_195;
input n_885;
input n_513;
input n_212;
input n_588;
input n_877;
input n_693;
input n_311;
input n_860;
input n_661;
input n_848;
input n_406;
input n_606;
input n_737;
input n_896;
input n_97;
input n_197;
input n_528;
input n_181;
input n_1005;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_836;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_985;
input n_572;
input n_867;
input n_983;
input n_1003;
input n_644;
input n_577;
input n_344;
input n_393;
input n_889;
input n_897;
input n_436;
input n_428;
input n_970;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_816;
input n_874;
input n_890;
input n_912;
input n_921;
input n_83;
input n_32;
input n_1058;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_908;
input n_213;
input n_964;
input n_424;
input n_565;
input n_916;
input n_823;
input n_701;
input n_271;
input n_995;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_984;
input n_394;
input n_79;
input n_1000;
input n_81;
input n_35;
input n_364;
input n_687;
input n_895;
input n_988;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_1035;
input n_760;
input n_751;
input n_806;
input n_932;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_855;
input n_232;
input n_380;
input n_749;
input n_281;
input n_866;
input n_559;
input n_425;
input n_1050;

output n_7788;

wire n_4557;
wire n_6873;
wire n_6210;
wire n_5285;
wire n_6516;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_4983;
wire n_3548;
wire n_5647;
wire n_7170;
wire n_1382;
wire n_2949;
wire n_2840;
wire n_6537;
wire n_3319;
wire n_3915;
wire n_5002;
wire n_5155;
wire n_5130;
wire n_7029;
wire n_4204;
wire n_5899;
wire n_6259;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_3817;
wire n_2038;
wire n_2504;
wire n_7042;
wire n_4607;
wire n_4514;
wire n_3674;
wire n_4249;
wire n_4931;
wire n_1859;
wire n_5827;
wire n_4805;
wire n_1765;
wire n_2392;
wire n_5008;
wire n_6183;
wire n_3280;
wire n_7262;
wire n_7551;
wire n_6616;
wire n_6848;
wire n_4371;
wire n_7766;
wire n_4601;
wire n_6035;
wire n_5858;
wire n_5879;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1782;
wire n_2889;
wire n_6567;
wire n_7063;
wire n_2391;
wire n_4585;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_2396;
wire n_3440;
wire n_4169;
wire n_6744;
wire n_7707;
wire n_3570;
wire n_5760;
wire n_4875;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2506;
wire n_7589;
wire n_6229;
wire n_7643;
wire n_3598;
wire n_1752;
wire n_4172;
wire n_6639;
wire n_1730;
wire n_5243;
wire n_3479;
wire n_5587;
wire n_3751;
wire n_3262;
wire n_4673;
wire n_3537;
wire n_5667;
wire n_2343;
wire n_5615;
wire n_1480;
wire n_7147;
wire n_6327;
wire n_1463;
wire n_1823;
wire n_4781;
wire n_6256;
wire n_4423;
wire n_5517;
wire n_1766;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_7067;
wire n_5962;
wire n_3347;
wire n_3395;
wire n_4808;
wire n_6658;
wire n_4507;
wire n_3577;
wire n_2995;
wire n_6842;
wire n_4526;
wire n_6286;
wire n_3472;
wire n_7485;
wire n_5922;
wire n_1981;
wire n_7636;
wire n_3976;
wire n_4348;
wire n_5931;
wire n_7450;
wire n_7492;
wire n_6760;
wire n_7396;
wire n_3807;
wire n_2998;
wire n_3845;
wire n_7082;
wire n_2163;
wire n_4450;
wire n_4467;
wire n_6159;
wire n_6517;
wire n_7313;
wire n_7305;
wire n_4801;
wire n_6005;
wire n_3639;
wire n_5809;
wire n_7332;
wire n_1664;
wire n_4144;
wire n_3298;
wire n_1427;
wire n_4447;
wire n_4955;
wire n_3208;
wire n_5588;
wire n_4569;
wire n_5404;
wire n_3671;
wire n_7673;
wire n_1778;
wire n_7151;
wire n_2839;
wire n_7013;
wire n_4998;
wire n_1698;
wire n_1496;
wire n_2333;
wire n_2705;
wire n_5505;
wire n_1214;
wire n_1274;
wire n_1595;
wire n_6530;
wire n_4510;
wire n_5658;
wire n_4567;
wire n_7672;
wire n_5151;
wire n_2362;
wire n_5478;
wire n_2822;
wire n_1306;
wire n_5994;
wire n_1493;
wire n_2597;
wire n_2774;
wire n_7776;
wire n_6602;
wire n_7753;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_5037;
wire n_5878;
wire n_5716;
wire n_1960;
wire n_6562;
wire n_7397;
wire n_7324;
wire n_3979;
wire n_3714;
wire n_6534;
wire n_6629;
wire n_7105;
wire n_2844;
wire n_6192;
wire n_3565;
wire n_7560;
wire n_5304;
wire n_3883;
wire n_5866;
wire n_5941;
wire n_3943;
wire n_4563;
wire n_1309;
wire n_5882;
wire n_1316;
wire n_1562;
wire n_6102;
wire n_7187;
wire n_4854;
wire n_6732;
wire n_3769;
wire n_6456;
wire n_1445;
wire n_6026;
wire n_2147;
wire n_5591;
wire n_6083;
wire n_7229;
wire n_2253;
wire n_4479;
wire n_5381;
wire n_3858;
wire n_4173;
wire n_6674;
wire n_6486;
wire n_5261;
wire n_5895;
wire n_7099;
wire n_5944;
wire n_6328;
wire n_5673;
wire n_7251;
wire n_7189;
wire n_4422;
wire n_5743;
wire n_6868;
wire n_1865;
wire n_5033;
wire n_6491;
wire n_4842;
wire n_4786;
wire n_1170;
wire n_3842;
wire n_2980;
wire n_7706;
wire n_6219;
wire n_5075;
wire n_1322;
wire n_4457;
wire n_4060;
wire n_6241;
wire n_7507;
wire n_1305;
wire n_2088;
wire n_6724;
wire n_1248;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_7097;
wire n_3780;
wire n_5571;
wire n_1653;
wire n_1375;
wire n_6254;
wire n_1118;
wire n_6066;
wire n_7241;
wire n_1881;
wire n_3798;
wire n_4809;
wire n_5241;
wire n_3060;
wire n_5129;
wire n_4124;
wire n_4499;
wire n_1350;
wire n_3627;
wire n_5191;
wire n_7264;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_2412;
wire n_2783;
wire n_5259;
wire n_3293;
wire n_7372;
wire n_2550;
wire n_5913;
wire n_6302;
wire n_6580;
wire n_7607;
wire n_5266;
wire n_3381;
wire n_2750;
wire n_1650;
wire n_1453;
wire n_5580;
wire n_1108;
wire n_6078;
wire n_7521;
wire n_1423;
wire n_3836;
wire n_1239;
wire n_4714;
wire n_5660;
wire n_5955;
wire n_1209;
wire n_5419;
wire n_3732;
wire n_6070;
wire n_6926;
wire n_3295;
wire n_3199;
wire n_1616;
wire n_6625;
wire n_7628;
wire n_2389;
wire n_5612;
wire n_6408;
wire n_6638;
wire n_7358;
wire n_2107;
wire n_3435;
wire n_4828;
wire n_4480;
wire n_1613;
wire n_3874;
wire n_6878;
wire n_2782;
wire n_4258;
wire n_1549;
wire n_4290;
wire n_1531;
wire n_2919;
wire n_6019;
wire n_4577;
wire n_7316;
wire n_1424;
wire n_2625;
wire n_2444;
wire n_3652;
wire n_4913;
wire n_2199;
wire n_1610;
wire n_4398;
wire n_7207;
wire n_1298;
wire n_1844;
wire n_6485;
wire n_4055;
wire n_3194;
wire n_4692;
wire n_7112;
wire n_7083;
wire n_5987;
wire n_6421;
wire n_6009;
wire n_2431;
wire n_2084;
wire n_1243;
wire n_7026;
wire n_3572;
wire n_6114;
wire n_6996;
wire n_1121;
wire n_4823;
wire n_7366;
wire n_5195;
wire n_7657;
wire n_5541;
wire n_7033;
wire n_6081;
wire n_3951;
wire n_4927;
wire n_3355;
wire n_2019;
wire n_1407;
wire n_4680;
wire n_1821;
wire n_7103;
wire n_5609;
wire n_5904;
wire n_4757;
wire n_5254;
wire n_6334;
wire n_3698;
wire n_2731;
wire n_4451;
wire n_5423;
wire n_4653;
wire n_3466;
wire n_3370;
wire n_6606;
wire n_1504;
wire n_6864;
wire n_1781;
wire n_4331;
wire n_7733;
wire n_2028;
wire n_3678;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_5732;
wire n_5141;
wire n_1293;
wire n_7711;
wire n_3968;
wire n_4825;
wire n_6178;
wire n_3950;
wire n_5252;
wire n_6209;
wire n_7445;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_4623;
wire n_4523;
wire n_4411;
wire n_3811;
wire n_6941;
wire n_1271;
wire n_6011;
wire n_7667;
wire n_3416;
wire n_6824;
wire n_3147;
wire n_3983;
wire n_3628;
wire n_2425;
wire n_2800;
wire n_7140;
wire n_4225;
wire n_7169;
wire n_5238;
wire n_6533;
wire n_3859;
wire n_6540;
wire n_4489;
wire n_6912;
wire n_3455;
wire n_6940;
wire n_1591;
wire n_7048;
wire n_2289;
wire n_2841;
wire n_4271;
wire n_7303;
wire n_1409;
wire n_2744;
wire n_3524;
wire n_6085;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_4404;
wire n_1521;
wire n_5502;
wire n_3054;
wire n_2456;
wire n_2924;
wire n_5288;
wire n_2264;
wire n_1987;
wire n_7192;
wire n_5749;
wire n_1129;
wire n_1244;
wire n_7639;
wire n_3365;
wire n_4974;
wire n_6802;
wire n_4725;
wire n_6691;
wire n_6431;
wire n_1932;
wire n_3775;
wire n_6196;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_7394;
wire n_4658;
wire n_2655;
wire n_3487;
wire n_1715;
wire n_6377;
wire n_3300;
wire n_5920;
wire n_5969;
wire n_1713;
wire n_3621;
wire n_2036;
wire n_1255;
wire n_6855;
wire n_2740;
wire n_2622;
wire n_4250;
wire n_7003;
wire n_1218;
wire n_4572;
wire n_5705;
wire n_4374;
wire n_6146;
wire n_7161;
wire n_3708;
wire n_2626;
wire n_1446;
wire n_7723;
wire n_7748;
wire n_6958;
wire n_3218;
wire n_2880;
wire n_5887;
wire n_5948;
wire n_7226;
wire n_2423;
wire n_3849;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_4469;
wire n_2580;
wire n_3529;
wire n_3222;
wire n_6711;
wire n_6124;
wire n_3352;
wire n_4180;
wire n_2964;
wire n_4062;
wire n_1498;
wire n_7356;
wire n_5199;
wire n_7377;
wire n_1207;
wire n_1735;
wire n_3813;
wire n_1825;
wire n_4232;
wire n_7360;
wire n_7315;
wire n_4199;
wire n_6061;
wire n_5099;
wire n_1210;
wire n_7081;
wire n_6136;
wire n_7559;
wire n_4033;
wire n_2522;
wire n_4608;
wire n_7446;
wire n_1201;
wire n_5859;
wire n_7224;
wire n_1246;
wire n_5258;
wire n_4231;
wire n_7541;
wire n_6187;
wire n_1724;
wire n_2838;
wire n_1540;
wire n_3243;
wire n_7583;
wire n_3214;
wire n_1890;
wire n_3128;
wire n_4073;
wire n_6402;
wire n_2549;
wire n_4325;
wire n_7131;
wire n_2440;
wire n_4113;
wire n_7777;
wire n_1440;
wire n_4646;
wire n_7155;
wire n_6305;
wire n_1751;
wire n_2146;
wire n_2341;
wire n_1737;
wire n_4819;
wire n_4261;
wire n_4884;
wire n_1083;
wire n_3205;
wire n_4490;
wire n_2358;
wire n_6971;
wire n_7553;
wire n_6128;
wire n_2361;
wire n_6804;
wire n_4128;
wire n_5213;
wire n_6469;
wire n_5354;
wire n_2062;
wire n_7700;
wire n_3932;
wire n_2339;
wire n_7338;
wire n_1963;
wire n_1418;
wire n_1137;
wire n_2552;
wire n_7221;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_3345;
wire n_6714;
wire n_4114;
wire n_6983;
wire n_1776;
wire n_6113;
wire n_3544;
wire n_5049;
wire n_1279;
wire n_6857;
wire n_4209;
wire n_3692;
wire n_5163;
wire n_1408;
wire n_5707;
wire n_3913;
wire n_3535;
wire n_6859;
wire n_2287;
wire n_3597;
wire n_4190;
wire n_7101;
wire n_2954;
wire n_6379;
wire n_6911;
wire n_6766;
wire n_2046;
wire n_6454;
wire n_4443;
wire n_4151;
wire n_4625;
wire n_4170;
wire n_7692;
wire n_7173;
wire n_4424;
wire n_6570;
wire n_1465;
wire n_6071;
wire n_4674;
wire n_6893;
wire n_6450;
wire n_1232;
wire n_2715;
wire n_6270;
wire n_4679;
wire n_6065;
wire n_7530;
wire n_1345;
wire n_4456;
wire n_5574;
wire n_1590;
wire n_7729;
wire n_7349;
wire n_2133;
wire n_3553;
wire n_5081;
wire n_6850;
wire n_6332;
wire n_6345;
wire n_1471;
wire n_5385;
wire n_3441;
wire n_4559;
wire n_5336;
wire n_2551;
wire n_4641;
wire n_4064;
wire n_5668;
wire n_4110;
wire n_4379;
wire n_3397;
wire n_5310;
wire n_4145;
wire n_6507;
wire n_1627;
wire n_3880;
wire n_7749;
wire n_5192;
wire n_4664;
wire n_3829;
wire n_7690;
wire n_1864;
wire n_6827;
wire n_5206;
wire n_2010;
wire n_2733;
wire n_6120;
wire n_7068;
wire n_3796;
wire n_5719;
wire n_6544;
wire n_5157;
wire n_1836;
wire n_6384;
wire n_4753;
wire n_1420;
wire n_2651;
wire n_1699;
wire n_6699;
wire n_4894;
wire n_5892;
wire n_5216;
wire n_6901;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3954;
wire n_3978;
wire n_4321;
wire n_5375;
wire n_2418;
wire n_1087;
wire n_1599;
wire n_3070;
wire n_3477;
wire n_1575;
wire n_6773;
wire n_4416;
wire n_7430;
wire n_5998;
wire n_4024;
wire n_5521;
wire n_3975;
wire n_3164;
wire n_6314;
wire n_1448;
wire n_3034;
wire n_6765;
wire n_7703;
wire n_6605;
wire n_5433;
wire n_2628;
wire n_4361;
wire n_1705;
wire n_4237;
wire n_2263;
wire n_3495;
wire n_3169;
wire n_6349;
wire n_3759;
wire n_4777;
wire n_7391;
wire n_4800;
wire n_3629;
wire n_5573;
wire n_7695;
wire n_5620;
wire n_4117;
wire n_6527;
wire n_7283;
wire n_2884;
wire n_3383;
wire n_7148;
wire n_3687;
wire n_6626;
wire n_4154;
wire n_3459;
wire n_6105;
wire n_6704;
wire n_2691;
wire n_2243;
wire n_3092;
wire n_7592;
wire n_5330;
wire n_4385;
wire n_2759;
wire n_3434;
wire n_7254;
wire n_2654;
wire n_7199;
wire n_5729;
wire n_2975;
wire n_2503;
wire n_4072;
wire n_1512;
wire n_4908;
wire n_3885;
wire n_7509;
wire n_1426;
wire n_2365;
wire n_6528;
wire n_2245;
wire n_3877;
wire n_6939;
wire n_5083;
wire n_3260;
wire n_6463;
wire n_2776;
wire n_6727;
wire n_2630;
wire n_6348;
wire n_1967;
wire n_1095;
wire n_6883;
wire n_5801;
wire n_3834;
wire n_5579;
wire n_1378;
wire n_7457;
wire n_3257;
wire n_2459;
wire n_6652;
wire n_2439;
wire n_7619;
wire n_7760;
wire n_1430;
wire n_5365;
wire n_2450;
wire n_6459;
wire n_4195;
wire n_1475;
wire n_3337;
wire n_5263;
wire n_6950;
wire n_4851;
wire n_4963;
wire n_1122;
wire n_3387;
wire n_7327;
wire n_6126;
wire n_4495;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_2728;
wire n_4685;
wire n_6915;
wire n_6115;
wire n_3428;
wire n_5959;
wire n_6282;
wire n_2427;
wire n_5017;
wire n_1127;
wire n_5938;
wire n_7025;
wire n_1845;
wire n_3835;
wire n_7645;
wire n_3723;
wire n_3389;
wire n_5292;
wire n_2422;
wire n_6277;
wire n_5190;
wire n_1679;
wire n_2342;
wire n_5926;
wire n_2755;
wire n_6531;
wire n_2301;
wire n_6922;
wire n_1578;
wire n_2712;
wire n_5316;
wire n_4314;
wire n_6731;
wire n_6502;
wire n_2788;
wire n_2089;
wire n_7090;
wire n_1857;
wire n_7587;
wire n_7574;
wire n_1997;
wire n_7174;
wire n_3314;
wire n_5135;
wire n_1349;
wire n_7250;
wire n_3891;
wire n_4704;
wire n_1777;
wire n_3409;
wire n_6646;
wire n_1546;
wire n_6394;
wire n_4003;
wire n_4775;
wire n_3420;
wire n_5840;
wire n_4192;
wire n_4633;
wire n_1950;
wire n_6439;
wire n_6084;
wire n_4593;
wire n_3914;
wire n_3289;
wire n_6902;
wire n_1834;
wire n_3372;
wire n_7641;
wire n_4121;
wire n_2862;
wire n_3850;
wire n_4488;
wire n_3405;
wire n_6837;
wire n_1657;
wire n_1741;
wire n_4264;
wire n_4183;
wire n_4118;
wire n_4302;
wire n_2138;
wire n_4916;
wire n_6767;
wire n_7102;
wire n_4858;
wire n_6733;
wire n_1914;
wire n_3833;
wire n_5833;
wire n_6723;
wire n_3339;
wire n_7177;
wire n_6900;
wire n_3673;
wire n_5792;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_3556;
wire n_5617;
wire n_1340;
wire n_2562;
wire n_6191;
wire n_3269;
wire n_7539;
wire n_5491;
wire n_2223;
wire n_5024;
wire n_3876;
wire n_4971;
wire n_1267;
wire n_2683;
wire n_3432;
wire n_5696;
wire n_1816;
wire n_7233;
wire n_4645;
wire n_4619;
wire n_2318;
wire n_2141;
wire n_1422;
wire n_6044;
wire n_4339;
wire n_5493;
wire n_4085;
wire n_3190;
wire n_3878;
wire n_4661;
wire n_2947;
wire n_4080;
wire n_5406;
wire n_1754;
wire n_3686;
wire n_6595;
wire n_7742;
wire n_2679;
wire n_4028;
wire n_5704;
wire n_7031;
wire n_1517;
wire n_5973;
wire n_7012;
wire n_7238;
wire n_3670;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_4289;
wire n_7030;
wire n_7110;
wire n_5555;
wire n_1895;
wire n_1860;
wire n_5727;
wire n_6856;
wire n_5770;
wire n_1763;
wire n_6976;
wire n_3912;
wire n_5169;
wire n_1607;
wire n_6682;
wire n_2959;
wire n_2380;
wire n_2420;
wire n_3265;
wire n_2221;
wire n_1774;
wire n_5274;
wire n_7517;
wire n_2516;
wire n_2031;
wire n_7121;
wire n_1348;
wire n_7317;
wire n_1191;
wire n_4099;
wire n_7190;
wire n_3899;
wire n_6153;
wire n_4729;
wire n_5957;
wire n_7429;
wire n_1617;
wire n_2639;
wire n_5323;
wire n_6777;
wire n_3099;
wire n_6412;
wire n_4745;
wire n_4057;
wire n_7390;
wire n_2410;
wire n_7145;
wire n_3206;
wire n_2633;
wire n_2049;
wire n_6245;
wire n_2113;
wire n_7787;
wire n_1690;
wire n_6553;
wire n_4466;
wire n_4132;
wire n_3361;
wire n_6543;
wire n_5566;
wire n_7561;
wire n_7529;
wire n_6185;
wire n_6706;
wire n_5342;
wire n_6884;
wire n_4603;
wire n_1135;
wire n_4300;
wire n_3277;
wire n_7533;
wire n_2758;
wire n_5787;
wire n_6745;
wire n_7210;
wire n_4417;
wire n_5967;
wire n_1550;
wire n_1169;
wire n_6224;
wire n_1938;
wire n_3452;
wire n_7563;
wire n_4022;
wire n_5843;
wire n_2194;
wire n_6072;
wire n_4320;
wire n_1173;
wire n_2736;
wire n_2845;
wire n_3886;
wire n_7191;
wire n_1901;
wire n_5332;
wire n_6073;
wire n_3096;
wire n_6097;
wire n_2059;
wire n_1278;
wire n_5553;
wire n_4730;
wire n_5763;
wire n_4616;
wire n_4760;
wire n_1710;
wire n_3021;
wire n_6881;
wire n_1603;
wire n_5864;
wire n_5227;
wire n_7136;
wire n_3404;
wire n_2072;
wire n_2963;
wire n_1489;
wire n_1993;
wire n_4859;
wire n_7213;
wire n_1455;
wire n_2182;
wire n_3115;
wire n_5352;
wire n_4583;
wire n_7034;
wire n_1502;
wire n_4923;
wire n_3920;
wire n_5370;
wire n_4082;
wire n_3273;
wire n_4367;
wire n_4282;
wire n_5600;
wire n_4475;
wire n_2286;
wire n_2563;
wire n_4893;
wire n_6990;
wire n_3650;
wire n_6948;
wire n_5014;
wire n_3513;
wire n_2677;
wire n_2531;
wire n_6591;
wire n_4029;
wire n_3212;
wire n_1321;
wire n_1779;
wire n_2489;
wire n_6816;
wire n_7512;
wire n_2950;
wire n_2272;
wire n_3574;
wire n_2608;
wire n_6712;
wire n_5824;
wire n_6280;
wire n_7682;
wire n_5472;
wire n_5950;
wire n_3739;
wire n_2825;
wire n_7098;
wire n_4338;
wire n_5546;
wire n_6222;
wire n_5972;
wire n_4985;
wire n_2742;
wire n_3604;
wire n_1740;
wire n_3540;
wire n_2680;
wire n_1343;
wire n_1371;
wire n_4198;
wire n_5924;
wire n_4529;
wire n_2861;
wire n_2976;
wire n_6656;
wire n_7323;
wire n_2366;
wire n_6318;
wire n_6200;
wire n_7149;
wire n_7219;
wire n_4919;
wire n_7320;
wire n_7175;
wire n_4111;
wire n_4200;
wire n_1659;
wire n_4575;
wire n_4847;
wire n_4803;
wire n_1878;
wire n_1374;
wire n_7357;
wire n_2851;
wire n_2973;
wire n_3651;
wire n_6637;
wire n_4666;
wire n_5752;
wire n_1242;
wire n_2810;
wire n_1119;
wire n_3027;
wire n_4189;
wire n_4076;
wire n_5233;
wire n_3438;
wire n_4835;
wire n_3464;
wire n_4390;
wire n_5977;
wire n_4722;
wire n_1530;
wire n_3215;
wire n_5968;
wire n_2871;
wire n_2764;
wire n_5713;
wire n_3648;
wire n_3234;
wire n_6577;
wire n_4058;
wire n_6268;
wire n_5403;
wire n_7593;
wire n_4611;
wire n_5527;
wire n_2714;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_5831;
wire n_1459;
wire n_4032;
wire n_6032;
wire n_2232;
wire n_4541;
wire n_4530;
wire n_1570;
wire n_5048;
wire n_5671;
wire n_6129;
wire n_1303;
wire n_1994;
wire n_7449;
wire n_6058;
wire n_1526;
wire n_4268;
wire n_2367;
wire n_3236;
wire n_1961;
wire n_3013;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_3256;
wire n_3126;
wire n_5834;
wire n_1257;
wire n_6641;
wire n_2864;
wire n_1632;
wire n_3104;
wire n_5951;
wire n_4895;
wire n_5480;
wire n_7663;
wire n_3354;
wire n_4069;
wire n_5289;
wire n_3373;
wire n_7218;
wire n_6863;
wire n_2784;
wire n_4140;
wire n_1909;
wire n_7292;
wire n_4125;
wire n_2495;
wire n_4531;
wire n_6556;
wire n_4789;
wire n_4778;
wire n_2703;
wire n_6152;
wire n_7582;
wire n_2574;
wire n_7659;
wire n_7142;
wire n_5492;
wire n_1887;
wire n_6106;
wire n_7428;
wire n_3504;
wire n_3511;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_3101;
wire n_6805;
wire n_5260;
wire n_6416;
wire n_7602;
wire n_5069;
wire n_2364;
wire n_7133;
wire n_2641;
wire n_7306;
wire n_7202;
wire n_6771;
wire n_4751;
wire n_7730;
wire n_5930;
wire n_5309;
wire n_6695;
wire n_3774;
wire n_2494;
wire n_3863;
wire n_5782;
wire n_2228;
wire n_4474;
wire n_5646;
wire n_7691;
wire n_1518;
wire n_4350;
wire n_5327;
wire n_4478;
wire n_2872;
wire n_2411;
wire n_3539;
wire n_2266;
wire n_4473;
wire n_6673;
wire n_7138;
wire n_7370;
wire n_3761;
wire n_2830;
wire n_4675;
wire n_3083;
wire n_6978;
wire n_7626;
wire n_5927;
wire n_3844;
wire n_4049;
wire n_2044;
wire n_2091;
wire n_4945;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_5019;
wire n_4891;
wire n_6910;
wire n_2394;
wire n_1572;
wire n_7236;
wire n_1245;
wire n_4867;
wire n_7387;
wire n_2929;
wire n_6346;
wire n_4911;
wire n_5414;
wire n_1329;
wire n_2409;
wire n_6403;
wire n_2405;
wire n_2601;
wire n_4405;
wire n_3118;
wire n_6172;
wire n_7122;
wire n_3742;
wire n_6004;
wire n_3532;
wire n_6347;
wire n_6482;
wire n_7698;
wire n_5280;
wire n_5466;
wire n_5469;
wire n_7024;
wire n_6925;
wire n_6483;
wire n_4686;
wire n_7466;
wire n_6358;
wire n_4682;
wire n_5750;
wire n_5305;
wire n_2914;
wire n_1833;
wire n_6598;
wire n_6800;
wire n_7410;
wire n_5186;
wire n_7257;
wire n_1986;
wire n_2882;
wire n_4301;
wire n_2493;
wire n_6499;
wire n_6944;
wire n_6215;
wire n_2115;
wire n_2013;
wire n_1556;
wire n_3547;
wire n_4898;
wire n_6980;
wire n_3700;
wire n_5180;
wire n_6594;
wire n_6233;
wire n_4733;
wire n_5368;
wire n_6338;
wire n_5757;
wire n_3947;
wire n_4684;
wire n_3663;
wire n_2129;
wire n_3230;
wire n_6621;
wire n_7282;
wire n_2532;
wire n_3782;
wire n_1720;
wire n_3831;
wire n_2293;
wire n_7495;
wire n_7334;
wire n_3068;
wire n_3071;
wire n_3919;
wire n_3683;
wire n_6053;
wire n_2734;
wire n_1166;
wire n_7346;
wire n_5267;
wire n_7649;
wire n_6020;
wire n_2310;
wire n_2674;
wire n_1284;
wire n_7532;
wire n_7740;
wire n_6432;
wire n_6426;
wire n_2689;
wire n_1992;
wire n_4493;
wire n_4797;
wire n_5397;
wire n_4962;
wire n_2596;
wire n_1488;
wire n_7401;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_3606;
wire n_5232;
wire n_7245;
wire n_1866;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_6946;
wire n_5890;
wire n_4644;
wire n_4412;
wire n_6068;
wire n_5802;
wire n_4266;
wire n_5815;
wire n_5605;
wire n_6897;
wire n_3124;
wire n_2982;
wire n_2634;
wire n_5384;
wire n_6550;
wire n_3015;
wire n_3321;
wire n_3081;
wire n_4639;
wire n_2291;
wire n_5664;
wire n_4102;
wire n_3612;
wire n_2172;
wire n_1728;
wire n_5863;
wire n_1230;
wire n_7075;
wire n_7710;
wire n_3622;
wire n_5276;
wire n_3857;
wire n_6847;
wire n_6042;
wire n_2357;
wire n_5197;
wire n_4354;
wire n_5320;
wire n_2937;
wire n_3728;
wire n_5087;
wire n_5265;
wire n_4401;
wire n_4727;
wire n_7367;
wire n_6265;
wire n_4296;
wire n_5312;
wire n_5534;
wire n_2967;
wire n_6737;
wire n_3005;
wire n_4627;
wire n_6936;
wire n_5107;
wire n_6780;
wire n_4309;
wire n_4027;
wire n_7132;
wire n_7486;
wire n_6758;
wire n_2056;
wire n_2054;
wire n_2226;
wire n_1402;
wire n_3267;
wire n_3008;
wire n_6452;
wire n_2802;
wire n_4728;
wire n_7419;
wire n_2279;
wire n_1536;
wire n_1719;
wire n_5281;
wire n_4046;
wire n_7201;
wire n_2961;
wire n_6458;
wire n_3689;
wire n_4631;
wire n_3283;
wire n_7555;
wire n_1736;
wire n_6176;
wire n_7265;
wire n_7232;
wire n_2907;
wire n_1948;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_6092;
wire n_7023;
wire n_3675;
wire n_7227;
wire n_2378;
wire n_2749;
wire n_3658;
wire n_4901;
wire n_3133;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_5025;
wire n_4539;
wire n_1205;
wire n_5575;
wire n_2969;
wire n_6052;
wire n_5753;
wire n_3550;
wire n_5401;
wire n_7642;
wire n_5509;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_6468;
wire n_1414;
wire n_5506;
wire n_6063;
wire n_7273;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_3275;
wire n_2645;
wire n_7623;
wire n_5417;
wire n_1714;
wire n_1958;
wire n_1611;
wire n_7774;
wire n_5015;
wire n_5372;
wire n_1675;
wire n_6909;
wire n_1551;
wire n_1533;
wire n_3792;
wire n_2515;
wire n_3089;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3988;
wire n_3406;
wire n_3758;
wire n_6418;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_3662;
wire n_6344;
wire n_1354;
wire n_3329;
wire n_1277;
wire n_5995;
wire n_3233;
wire n_3193;
wire n_2582;
wire n_7070;
wire n_5253;
wire n_3789;
wire n_6308;
wire n_2174;
wire n_6989;
wire n_2510;
wire n_7634;
wire n_2435;
wire n_3934;
wire n_2583;
wire n_1678;
wire n_4606;
wire n_1287;
wire n_1525;
wire n_6662;
wire n_6461;
wire n_7046;
wire n_1150;
wire n_1674;
wire n_6304;
wire n_3980;
wire n_2912;
wire n_2710;
wire n_6617;
wire n_2970;
wire n_1393;
wire n_4691;
wire n_5937;
wire n_2978;
wire n_5291;
wire n_3502;
wire n_5460;
wire n_3935;
wire n_5379;
wire n_1854;
wire n_1084;
wire n_2804;
wire n_5390;
wire n_5691;
wire n_4926;
wire n_5043;
wire n_6549;
wire n_7194;
wire n_4688;
wire n_5097;
wire n_5675;
wire n_3144;
wire n_4234;
wire n_4146;
wire n_2835;
wire n_4656;
wire n_4932;
wire n_6179;
wire n_1930;
wire n_5577;
wire n_1234;
wire n_4881;
wire n_7527;
wire n_7290;
wire n_3755;
wire n_1469;
wire n_4632;
wire n_7146;
wire n_3255;
wire n_1652;
wire n_2183;
wire n_6607;
wire n_1883;
wire n_2037;
wire n_4550;
wire n_6960;
wire n_1226;
wire n_7253;
wire n_4651;
wire n_1873;
wire n_1619;
wire n_2682;
wire n_1666;
wire n_3605;
wire n_5181;
wire n_3105;
wire n_3146;
wire n_4892;
wire n_4343;
wire n_7615;
wire n_3931;
wire n_5745;
wire n_7434;
wire n_4421;
wire n_2322;
wire n_7477;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_7452;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_5893;
wire n_3843;
wire n_2847;
wire n_4399;
wire n_1308;
wire n_5067;
wire n_6823;
wire n_3904;
wire n_4378;
wire n_6455;
wire n_3729;
wire n_5637;
wire n_3484;
wire n_7414;
wire n_2485;
wire n_5614;
wire n_4477;
wire n_5177;
wire n_5643;
wire n_2179;
wire n_6725;
wire n_4654;
wire n_3984;
wire n_4233;
wire n_4765;
wire n_7475;
wire n_7775;
wire n_7184;
wire n_3086;
wire n_2475;
wire n_3721;
wire n_5695;
wire n_3726;
wire n_6914;
wire n_5438;
wire n_4277;
wire n_4431;
wire n_7152;
wire n_4771;
wire n_4652;
wire n_4970;
wire n_6927;
wire n_5179;
wire n_3804;
wire n_1908;
wire n_6457;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_4285;
wire n_4928;
wire n_3251;
wire n_6916;
wire n_6973;
wire n_2921;
wire n_3724;
wire n_3192;
wire n_3753;
wire n_5683;
wire n_3566;
wire n_7554;
wire n_6564;
wire n_2820;
wire n_2311;
wire n_5701;
wire n_4403;
wire n_3242;
wire n_6566;
wire n_7114;
wire n_1654;
wire n_6428;
wire n_5774;
wire n_3330;
wire n_2707;
wire n_4746;
wire n_7354;
wire n_4382;
wire n_4002;
wire n_3631;
wire n_6808;
wire n_7609;
wire n_7037;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_4545;
wire n_2336;
wire n_3987;
wire n_7709;
wire n_3969;
wire n_4437;
wire n_6747;
wire n_7335;
wire n_3856;
wire n_6496;
wire n_1155;
wire n_5394;
wire n_1292;
wire n_5462;
wire n_2432;
wire n_3043;
wire n_2273;
wire n_5428;
wire n_4491;
wire n_4672;
wire n_5001;
wire n_2421;
wire n_3237;
wire n_6095;
wire n_6787;
wire n_1970;
wire n_3946;
wire n_7183;
wire n_2953;
wire n_3949;
wire n_3507;
wire n_6150;
wire n_3926;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_2436;
wire n_1663;
wire n_6784;
wire n_4267;
wire n_5933;
wire n_4723;
wire n_7433;
wire n_2269;
wire n_6741;
wire n_2472;
wire n_2846;
wire n_3699;
wire n_4312;
wire n_5874;
wire n_5104;
wire n_2249;
wire n_3022;
wire n_4014;
wire n_3766;
wire n_3707;
wire n_7669;
wire n_4217;
wire n_3973;
wire n_5964;
wire n_5551;
wire n_5319;
wire n_4769;
wire n_4724;
wire n_2260;
wire n_5543;
wire n_4721;
wire n_2663;
wire n_3882;
wire n_6807;
wire n_2595;
wire n_5723;
wire n_5621;
wire n_6795;
wire n_7437;
wire n_6898;
wire n_5386;
wire n_4433;
wire n_5133;
wire n_5056;
wire n_6785;
wire n_7384;
wire n_7588;
wire n_6738;
wire n_3030;
wire n_5631;
wire n_6818;
wire n_5983;
wire n_7516;
wire n_5796;
wire n_4503;
wire n_6232;
wire n_3917;
wire n_3679;
wire n_7393;
wire n_4517;
wire n_6021;
wire n_4511;
wire n_3221;
wire n_3210;
wire n_6966;
wire n_1672;
wire n_4171;
wire n_3764;
wire n_5405;
wire n_6389;
wire n_3795;
wire n_6055;
wire n_4788;
wire n_4754;
wire n_1817;
wire n_5848;
wire n_5221;
wire n_1301;
wire n_5997;
wire n_4166;
wire n_2242;
wire n_4845;
wire n_1561;
wire n_5122;
wire n_2247;
wire n_3177;
wire n_3399;
wire n_5439;
wire n_6899;
wire n_4850;
wire n_1869;
wire n_7614;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_3676;
wire n_1753;
wire n_6351;
wire n_7503;
wire n_4610;
wire n_6441;
wire n_5854;
wire n_6754;
wire n_4067;
wire n_6822;
wire n_6796;
wire n_6849;
wire n_6836;
wire n_4997;
wire n_5906;
wire n_7355;
wire n_6755;
wire n_7608;
wire n_4393;
wire n_5205;
wire n_3777;
wire n_7084;
wire n_5916;
wire n_7685;
wire n_5993;
wire n_4553;
wire n_5240;
wire n_3961;
wire n_1520;
wire n_7515;
wire n_2509;
wire n_5714;
wire n_4283;
wire n_4174;
wire n_4870;
wire n_2399;
wire n_1370;
wire n_1708;
wire n_3038;
wire n_7483;
wire n_6476;
wire n_5828;
wire n_7648;
wire n_6276;
wire n_5907;
wire n_5284;
wire n_4804;
wire n_3716;
wire n_1649;
wire n_3450;
wire n_6669;
wire n_5357;
wire n_6717;
wire n_4994;
wire n_4518;
wire n_4732;
wire n_1936;
wire n_1717;
wire n_6040;
wire n_2257;
wire n_4856;
wire n_5088;
wire n_5250;
wire n_1467;
wire n_6388;
wire n_3217;
wire n_2511;
wire n_5461;
wire n_6298;
wire n_6988;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2661;
wire n_4079;
wire n_7256;
wire n_3573;
wire n_7652;
wire n_3563;
wire n_4993;
wire n_3510;
wire n_7172;
wire n_4248;
wire n_2334;
wire n_2350;
wire n_5958;
wire n_5619;
wire n_7117;
wire n_1709;
wire n_6655;
wire n_6541;
wire n_2649;
wire n_3607;
wire n_4476;
wire n_6460;
wire n_3241;
wire n_2746;
wire n_5471;
wire n_2256;
wire n_5210;
wire n_2445;
wire n_1980;
wire n_6790;
wire n_3583;
wire n_4987;
wire n_3832;
wire n_4649;
wire n_3508;
wire n_6295;
wire n_1862;
wire n_4693;
wire n_3415;
wire n_2355;
wire n_4992;
wire n_1543;
wire n_3386;
wire n_4568;
wire n_4359;
wire n_3814;
wire n_1441;
wire n_4573;
wire n_4105;
wire n_4206;
wire n_5273;
wire n_7722;
wire n_4177;
wire n_1888;
wire n_6497;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_5877;
wire n_6535;
wire n_5457;
wire n_5482;
wire n_4700;
wire n_2828;
wire n_1964;
wire n_6090;
wire n_3720;
wire n_1196;
wire n_6840;
wire n_1182;
wire n_4074;
wire n_5237;
wire n_5360;
wire n_3633;
wire n_1731;
wire n_5596;
wire n_2879;
wire n_3514;
wire n_3091;
wire n_5625;
wire n_4037;
wire n_4582;
wire n_5539;
wire n_3426;
wire n_7287;
wire n_4308;
wire n_2288;
wire n_3075;
wire n_1671;
wire n_6748;
wire n_3448;
wire n_3788;
wire n_6164;
wire n_6211;
wire n_2076;
wire n_3733;
wire n_1831;
wire n_4853;
wire n_6676;
wire n_6117;
wire n_6563;
wire n_1312;
wire n_5844;
wire n_6470;
wire n_7301;
wire n_6448;
wire n_3684;
wire n_6667;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_6018;
wire n_6094;
wire n_3970;
wire n_3291;
wire n_2454;
wire n_4008;
wire n_4973;
wire n_7786;
wire n_2829;
wire n_4966;
wire n_2968;
wire n_4494;
wire n_3473;
wire n_5362;
wire n_6236;
wire n_6208;
wire n_5294;
wire n_6197;
wire n_3263;
wire n_4501;
wire n_7156;
wire n_1772;
wire n_2858;
wire n_7780;
wire n_1283;
wire n_6552;
wire n_1421;
wire n_4922;
wire n_6237;
wire n_5089;
wire n_2573;
wire n_1793;
wire n_2424;
wire n_6993;
wire n_2390;
wire n_7544;
wire n_7203;
wire n_4402;
wire n_2793;
wire n_4813;
wire n_6653;
wire n_3098;
wire n_7732;
wire n_6449;
wire n_1711;
wire n_3069;
wire n_5465;
wire n_3107;
wire n_5488;
wire n_4134;
wire n_4131;
wire n_6539;
wire n_4330;
wire n_5832;
wire n_2176;
wire n_2805;
wire n_5165;
wire n_2319;
wire n_5678;
wire n_7658;
wire n_3757;
wire n_5811;
wire n_1933;
wire n_7408;
wire n_7605;
wire n_1842;
wire n_3364;
wire n_3429;
wire n_3306;
wire n_5234;
wire n_3787;
wire n_5140;
wire n_3445;
wire n_2080;
wire n_5655;
wire n_5514;
wire n_2554;
wire n_6130;
wire n_1676;
wire n_7476;
wire n_7624;
wire n_5020;
wire n_5225;
wire n_1136;
wire n_1918;
wire n_3642;
wire n_2461;
wire n_1229;
wire n_1490;
wire n_1179;
wire n_4818;
wire n_7566;
wire n_4462;
wire n_1153;
wire n_6560;
wire n_7307;
wire n_2787;
wire n_4540;
wire n_6987;
wire n_4187;
wire n_7684;
wire n_1273;
wire n_3821;
wire n_2930;
wire n_2616;
wire n_4979;
wire n_7409;
wire n_7087;
wire n_3503;
wire n_2441;
wire n_7280;
wire n_7680;
wire n_4063;
wire n_4362;
wire n_5318;
wire n_3312;
wire n_1848;
wire n_4009;
wire n_7107;
wire n_2650;
wire n_2888;
wire n_3614;
wire n_5946;
wire n_6131;
wire n_3394;
wire n_6207;
wire n_6984;
wire n_5942;
wire n_2530;
wire n_2792;
wire n_2372;
wire n_4191;
wire n_4965;
wire n_1522;
wire n_2523;
wire n_6701;
wire n_6326;
wire n_3488;
wire n_6365;
wire n_7288;
wire n_7248;
wire n_2832;
wire n_4991;
wire n_4525;
wire n_4011;
wire n_3526;
wire n_5242;
wire n_2142;
wire n_6519;
wire n_3703;
wire n_5116;
wire n_6635;
wire n_6907;
wire n_4554;
wire n_1260;
wire n_7038;
wire n_4097;
wire n_4861;
wire n_3239;
wire n_6155;
wire n_5953;
wire n_2600;
wire n_3952;
wire n_1171;
wire n_1126;
wire n_6151;
wire n_6074;
wire n_4596;
wire n_2434;
wire n_3578;
wire n_4734;
wire n_5947;
wire n_6661;
wire n_6730;
wire n_4492;
wire n_3470;
wire n_1738;
wire n_6370;
wire n_1729;
wire n_5563;
wire n_2094;
wire n_1479;
wire n_2306;
wire n_7153;
wire n_5194;
wire n_7230;
wire n_4579;
wire n_5628;
wire n_6994;
wire n_2568;
wire n_2629;
wire n_3587;
wire n_4936;
wire n_2097;
wire n_2109;
wire n_2648;
wire n_6262;
wire n_2398;
wire n_7572;
wire n_1593;
wire n_7308;
wire n_1775;
wire n_6889;
wire n_6361;
wire n_6803;
wire n_7481;
wire n_2570;
wire n_4025;
wire n_6751;
wire n_2184;
wire n_3948;
wire n_2842;
wire n_1400;
wire n_7403;
wire n_2469;
wire n_6024;
wire n_3074;
wire n_4640;
wire n_5790;
wire n_6523;
wire n_5746;
wire n_5883;
wire n_7369;
wire n_5630;
wire n_3136;
wire n_3108;
wire n_6696;
wire n_2395;
wire n_7089;
wire n_6062;
wire n_4059;
wire n_7258;
wire n_4130;
wire n_2752;
wire n_2124;
wire n_3991;
wire n_3974;
wire n_4642;
wire n_3625;
wire n_1746;
wire n_2716;
wire n_2212;
wire n_6943;
wire n_4878;
wire n_1832;
wire n_1128;
wire n_2376;
wire n_3398;
wire n_3718;
wire n_6252;
wire n_7080;
wire n_7718;
wire n_5193;
wire n_2170;
wire n_6407;
wire n_4904;
wire n_1785;
wire n_3999;
wire n_1405;
wire n_4087;
wire n_7002;
wire n_5153;
wire n_6235;
wire n_5369;
wire n_7745;
wire n_6726;
wire n_7689;
wire n_3238;
wire n_6740;
wire n_4318;
wire n_3731;
wire n_3555;
wire n_3254;
wire n_5007;
wire n_4717;
wire n_4052;
wire n_6447;
wire n_6799;
wire n_2463;
wire n_6932;
wire n_6434;
wire n_2478;
wire n_3178;
wire n_4245;
wire n_7008;
wire n_3378;
wire n_5689;
wire n_3350;
wire n_6391;
wire n_5399;
wire n_4873;
wire n_6630;
wire n_6631;
wire n_3936;
wire n_1560;
wire n_5513;
wire n_3166;
wire n_3953;
wire n_3385;
wire n_1265;
wire n_2488;
wire n_2042;
wire n_5891;
wire n_1925;
wire n_6489;
wire n_7049;
wire n_1251;
wire n_6657;
wire n_3090;
wire n_1247;
wire n_5030;
wire n_3816;
wire n_5098;
wire n_5755;
wire n_4636;
wire n_7062;
wire n_7493;
wire n_5408;
wire n_4256;
wire n_1185;
wire n_3575;
wire n_6716;
wire n_6797;
wire n_2765;
wire n_4278;
wire n_6165;
wire n_6263;
wire n_6481;
wire n_4609;
wire n_5148;
wire n_7215;
wire n_7340;
wire n_4822;
wire n_6694;
wire n_2936;
wire n_7154;
wire n_2985;
wire n_3106;
wire n_6597;
wire n_4030;
wire n_4276;
wire n_6238;
wire n_4612;
wire n_1148;
wire n_1667;
wire n_6272;
wire n_5454;
wire n_3902;
wire n_1707;
wire n_4203;
wire n_5650;
wire n_2055;
wire n_4866;
wire n_2385;
wire n_6965;
wire n_3864;
wire n_3026;
wire n_3294;
wire n_4831;
wire n_5656;
wire n_1143;
wire n_6647;
wire n_7279;
wire n_7499;
wire n_2584;
wire n_4381;
wire n_5183;
wire n_7771;
wire n_2442;
wire n_5072;
wire n_4441;
wire n_2000;
wire n_4083;
wire n_2696;
wire n_4960;
wire n_5146;
wire n_6846;
wire n_5131;
wire n_1894;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_4228;
wire n_4699;
wire n_5803;
wire n_1331;
wire n_1223;
wire n_5754;
wire n_1739;
wire n_3130;
wire n_1353;
wire n_7052;
wire n_5018;
wire n_2386;
wire n_7662;
wire n_3324;
wire n_3073;
wire n_2029;
wire n_4254;
wire n_4536;
wire n_7728;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_6931;
wire n_4924;
wire n_2238;
wire n_6398;
wire n_6700;
wire n_5786;
wire n_4138;
wire n_3100;
wire n_1727;
wire n_6366;
wire n_6853;
wire n_1294;
wire n_1351;
wire n_6679;
wire n_5035;
wire n_5425;
wire n_1380;
wire n_6036;
wire n_3336;
wire n_6104;
wire n_1291;
wire n_5742;
wire n_5901;
wire n_3763;
wire n_7158;
wire n_4284;
wire n_5943;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_6253;
wire n_7299;
wire n_1830;
wire n_6770;
wire n_3476;
wire n_3990;
wire n_2011;
wire n_4044;
wire n_5499;
wire n_7095;
wire n_7464;
wire n_1662;
wire n_7426;
wire n_3443;
wire n_5143;
wire n_3029;
wire n_4135;
wire n_7076;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_5302;
wire n_1660;
wire n_5640;
wire n_4000;
wire n_5841;
wire n_5011;
wire n_2556;
wire n_1537;
wire n_3908;
wire n_3696;
wire n_2902;
wire n_6242;
wire n_6660;
wire n_3608;
wire n_4269;
wire n_4016;
wire n_4915;
wire n_4286;
wire n_3048;
wire n_6414;
wire n_7666;
wire n_1962;
wire n_5296;
wire n_7246;
wire n_5159;
wire n_1952;
wire n_1624;
wire n_4795;
wire n_1598;
wire n_2952;
wire n_7459;
wire n_2250;
wire n_1491;
wire n_3778;
wire n_7570;
wire n_2075;
wire n_4816;
wire n_6951;
wire n_3335;
wire n_4846;
wire n_3669;
wire n_1899;
wire n_4001;
wire n_6029;
wire n_2892;
wire n_3356;
wire n_4377;
wire n_3220;
wire n_3422;
wire n_5798;
wire n_2309;
wire n_2274;
wire n_6278;
wire n_6949;
wire n_5096;
wire n_6480;
wire n_7380;
wire n_6443;
wire n_3712;
wire n_5805;
wire n_5171;
wire n_2143;
wire n_4637;
wire n_4976;
wire n_4021;
wire n_5351;
wire n_2739;
wire n_2528;
wire n_7167;
wire n_7537;
wire n_2548;
wire n_3216;
wire n_6157;
wire n_6453;
wire n_3061;
wire n_3717;
wire n_3424;
wire n_3745;
wire n_3245;
wire n_6693;
wire n_4855;
wire n_5851;
wire n_4643;
wire n_5217;
wire n_6030;
wire n_4736;
wire n_2817;
wire n_1790;
wire n_4202;
wire n_3196;
wire n_5767;
wire n_4287;
wire n_2809;
wire n_6615;
wire n_3921;
wire n_3480;
wire n_7455;
wire n_1494;
wire n_2060;
wire n_2214;
wire n_7755;
wire n_1726;
wire n_5751;
wire n_6819;
wire n_1241;
wire n_5929;
wire n_2589;
wire n_5928;
wire n_1231;
wire n_1208;
wire n_1604;
wire n_4947;
wire n_3506;
wire n_1976;
wire n_1337;
wire n_2984;
wire n_4890;
wire n_4538;
wire n_4023;
wire n_3031;
wire n_4920;
wire n_5869;
wire n_5862;
wire n_1238;
wire n_3959;
wire n_6937;
wire n_4288;
wire n_7629;
wire n_2452;
wire n_6274;
wire n_2144;
wire n_4763;
wire n_7725;
wire n_2592;
wire n_2251;
wire n_5201;
wire n_1644;
wire n_4586;
wire n_6190;
wire n_3860;
wire n_5353;
wire n_1871;
wire n_3044;
wire n_2868;
wire n_3493;
wire n_2818;
wire n_7474;
wire n_3486;
wire n_2426;
wire n_1403;
wire n_2181;
wire n_4034;
wire n_3253;
wire n_5444;
wire n_1149;
wire n_6860;
wire n_7739;
wire n_4905;
wire n_6100;
wire n_1457;
wire n_3172;
wire n_6833;
wire n_2159;
wire n_6865;
wire n_2700;
wire n_1222;
wire n_1630;
wire n_1959;
wire n_1198;
wire n_7135;
wire n_6794;
wire n_3637;
wire n_7216;
wire n_3393;
wire n_5772;
wire n_1261;
wire n_5520;
wire n_3327;
wire n_1114;
wire n_7487;
wire n_5277;
wire n_5900;
wire n_7421;
wire n_7694;
wire n_3647;
wire n_6240;
wire n_3928;
wire n_3619;
wire n_4043;
wire n_1846;
wire n_1573;
wire n_7399;
wire n_1956;
wire n_7186;
wire n_5569;
wire n_5779;
wire n_4270;
wire n_2983;
wire n_4273;
wire n_7580;
wire n_7632;
wire n_6498;
wire n_6720;
wire n_1669;
wire n_7562;
wire n_6247;
wire n_5109;
wire n_1885;
wire n_1989;
wire n_5837;
wire n_5402;
wire n_1801;
wire n_3740;
wire n_3001;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_2576;
wire n_6854;
wire n_4344;
wire n_1342;
wire n_6574;
wire n_2756;
wire n_7197;
wire n_7015;
wire n_7747;
wire n_1175;
wire n_4408;
wire n_6832;
wire n_5473;
wire n_1221;
wire n_3875;
wire n_5113;
wire n_7066;
wire n_4341;
wire n_4759;
wire n_7688;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_6779;
wire n_2567;
wire n_5645;
wire n_7044;
wire n_1085;
wire n_2981;
wire n_2222;
wire n_4439;
wire n_5102;
wire n_6258;
wire n_7329;
wire n_6139;
wire n_5167;
wire n_7756;
wire n_4565;
wire n_5562;
wire n_7713;
wire n_1451;
wire n_7438;
wire n_4663;
wire n_2471;
wire n_5666;
wire n_1288;
wire n_1275;
wire n_4519;
wire n_2757;
wire n_1622;
wire n_3121;
wire n_2121;
wire n_6887;
wire n_4515;
wire n_1893;
wire n_5639;
wire n_5607;
wire n_7735;
wire n_2278;
wire n_6769;
wire n_6903;
wire n_2433;
wire n_7255;
wire n_2798;
wire n_3425;
wire n_1771;
wire n_3308;
wire n_6169;
wire n_1507;
wire n_5914;
wire n_1206;
wire n_3576;
wire n_5275;
wire n_3109;
wire n_4838;
wire n_2553;
wire n_4524;
wire n_2218;
wire n_6861;
wire n_2130;
wire n_4862;
wire n_7270;
wire n_5114;
wire n_7071;
wire n_7773;
wire n_6697;
wire n_4260;
wire n_4628;
wire n_4696;
wire n_1097;
wire n_3122;
wire n_3012;
wire n_6826;
wire n_5005;
wire n_5004;
wire n_7768;
wire n_3368;
wire n_3586;
wire n_2381;
wire n_2313;
wire n_7235;
wire n_4597;
wire n_1812;
wire n_5090;
wire n_4574;
wire n_7129;
wire n_4242;
wire n_7243;
wire n_4949;
wire n_4748;
wire n_4959;
wire n_1747;
wire n_7342;
wire n_3400;
wire n_2508;
wire n_4243;
wire n_2540;
wire n_7547;
wire n_3820;
wire n_5395;
wire n_6494;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_2316;
wire n_5489;
wire n_5649;
wire n_7581;
wire n_1995;
wire n_4677;
wire n_1631;
wire n_7310;
wire n_2911;
wire n_1828;
wire n_6972;
wire n_1389;
wire n_6380;
wire n_7200;
wire n_7751;
wire n_5791;
wire n_1798;
wire n_5559;
wire n_6703;
wire n_7116;
wire n_4562;
wire n_1584;
wire n_7540;
wire n_7720;
wire n_5009;
wire n_6034;
wire n_1438;
wire n_1973;
wire n_2156;
wire n_6719;
wire n_6526;
wire n_4986;
wire n_4453;
wire n_1366;
wire n_7208;
wire n_1187;
wire n_3173;
wire n_6212;
wire n_4281;
wire n_4332;
wire n_7337;
wire n_3433;
wire n_3998;
wire n_1686;
wire n_4464;
wire n_3017;
wire n_4605;
wire n_4737;
wire n_6111;
wire n_2542;
wire n_2843;
wire n_3305;
wire n_1635;
wire n_7055;
wire n_5295;
wire n_6427;
wire n_4310;
wire n_3752;
wire n_7073;
wire n_2637;
wire n_7417;
wire n_7159;
wire n_5047;
wire n_5504;
wire n_7494;
wire n_7784;
wire n_5076;
wire n_3543;
wire n_5693;
wire n_3655;
wire n_7314;
wire n_3791;
wire n_6904;
wire n_6778;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_7294;
wire n_6520;
wire n_4906;
wire n_4257;
wire n_7016;
wire n_5712;
wire n_4516;
wire n_2913;
wire n_5028;
wire n_2254;
wire n_1381;
wire n_1597;
wire n_1486;
wire n_6444;
wire n_7422;
wire n_5622;
wire n_4196;
wire n_5255;
wire n_2371;
wire n_6362;
wire n_3898;
wire n_6749;
wire n_3366;
wire n_3453;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_6648;
wire n_2408;
wire n_6985;
wire n_4961;
wire n_6330;
wire n_5013;
wire n_2140;
wire n_6622;
wire n_2134;
wire n_2483;
wire n_2466;
wire n_3661;
wire n_5348;
wire n_6405;
wire n_2048;
wire n_2760;
wire n_1299;
wire n_2942;
wire n_4420;
wire n_4964;
wire n_5251;
wire n_5036;
wire n_3665;
wire n_2079;
wire n_4807;
wire n_4886;
wire n_6488;
wire n_7783;
wire n_4342;
wire n_5554;
wire n_2671;
wire n_3296;
wire n_5919;
wire n_5978;
wire n_6220;
wire n_1390;
wire n_2775;
wire n_7178;
wire n_7330;
wire n_3223;
wire n_2005;
wire n_7764;
wire n_1116;
wire n_7704;
wire n_2811;
wire n_1758;
wire n_7388;
wire n_2848;
wire n_6087;
wire n_1784;
wire n_3200;
wire n_1213;
wire n_3483;
wire n_5702;
wire n_3207;
wire n_5450;
wire n_7697;
wire n_5806;
wire n_1180;
wire n_4657;
wire n_3869;
wire n_3852;
wire n_1220;
wire n_5071;
wire n_5308;
wire n_5982;
wire n_6692;
wire n_7079;
wire n_6590;
wire n_7536;
wire n_3036;
wire n_7209;
wire n_5012;
wire n_5376;
wire n_6501;
wire n_5778;
wire n_4207;
wire n_1760;
wire n_5208;
wire n_6396;
wire n_2173;
wire n_2824;
wire n_7467;
wire n_4038;
wire n_5503;
wire n_7206;
wire n_4793;
wire n_4472;
wire n_2588;
wire n_6702;
wire n_3046;
wire n_7505;
wire n_6551;
wire n_1142;
wire n_1385;
wire n_4395;
wire n_4274;
wire n_5644;
wire n_7501;
wire n_6368;
wire n_2533;
wire n_1500;
wire n_2706;
wire n_1868;
wire n_2303;
wire n_7490;
wire n_4532;
wire n_5235;
wire n_5062;
wire n_6309;
wire n_3332;
wire n_5161;
wire n_4413;
wire n_4743;
wire n_2403;
wire n_5016;
wire n_2702;
wire n_3922;
wire n_7051;
wire n_7278;
wire n_2791;
wire n_1450;
wire n_7416;
wire n_2092;
wire n_6248;
wire n_5996;
wire n_3189;
wire n_7611;
wire n_2797;
wire n_7600;
wire n_1089;
wire n_4275;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_7447;
wire n_2996;
wire n_2836;
wire n_1404;
wire n_3582;
wire n_4830;
wire n_7520;
wire n_4442;
wire n_7702;
wire n_5700;
wire n_7274;
wire n_2168;
wire n_1442;
wire n_7668;
wire n_4689;
wire n_2886;
wire n_5699;
wire n_6287;
wire n_6022;
wire n_1968;
wire n_6579;
wire n_6820;
wire n_4018;
wire n_2609;
wire n_6633;
wire n_4613;
wire n_5940;
wire n_6614;
wire n_1483;
wire n_1703;
wire n_7591;
wire n_1953;
wire n_3715;
wire n_6952;
wire n_7617;
wire n_3261;
wire n_5324;
wire n_7534;
wire n_6547;
wire n_7065;
wire n_5421;
wire n_3861;
wire n_5175;
wire n_3161;
wire n_3313;
wire n_1807;
wire n_1310;
wire n_3198;
wire n_5820;
wire n_3463;
wire n_2559;
wire n_6589;
wire n_6995;
wire n_4188;
wire n_2619;
wire n_2726;
wire n_2917;
wire n_5340;
wire n_3738;
wire n_1640;
wire n_5694;
wire n_5022;
wire n_7461;
wire n_1145;
wire n_2307;
wire n_3546;
wire n_1511;
wire n_1651;
wire n_6297;
wire n_5245;
wire n_7326;
wire n_5651;
wire n_3944;
wire n_3595;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1696;
wire n_6367;
wire n_7761;
wire n_6198;
wire n_1355;
wire n_5364;
wire n_5459;
wire n_4534;
wire n_3635;
wire n_7423;
wire n_3270;
wire n_5168;
wire n_7443;
wire n_4590;
wire n_4602;
wire n_5329;
wire n_5510;
wire n_7746;
wire n_6251;
wire n_1335;
wire n_3213;
wire n_4394;
wire n_1900;
wire n_6583;
wire n_3418;
wire n_2614;
wire n_5581;
wire n_7556;
wire n_1091;
wire n_1780;
wire n_3865;
wire n_2769;
wire n_4220;
wire n_6879;
wire n_5812;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_4742;
wire n_2100;
wire n_4948;
wire n_3903;
wire n_3895;
wire n_1194;
wire n_3851;
wire n_4508;
wire n_4934;
wire n_7104;
wire n_7631;
wire n_3482;
wire n_2282;
wire n_3654;
wire n_4939;
wire n_4213;
wire n_2430;
wire n_2673;
wire n_2926;
wire n_1534;
wire n_5711;
wire n_3268;
wire n_4703;
wire n_1655;
wire n_3494;
wire n_7106;
wire n_3615;
wire n_7693;
wire n_7198;
wire n_7656;
wire n_7381;
wire n_5970;
wire n_3363;
wire n_7731;
wire n_1186;
wire n_3180;
wire n_5570;
wire n_1743;
wire n_7182;
wire n_6310;
wire n_6852;
wire n_1506;
wire n_5061;
wire n_2594;
wire n_1474;
wire n_3150;
wire n_5550;
wire n_4773;
wire n_3853;
wire n_6961;
wire n_2512;
wire n_4449;
wire n_5219;
wire n_6618;
wire n_7670;
wire n_2607;
wire n_4615;
wire n_3911;
wire n_7126;
wire n_5132;
wire n_4883;
wire n_6249;
wire n_3559;
wire n_6956;
wire n_5184;
wire n_6440;
wire n_7564;
wire n_5747;
wire n_6575;
wire n_5821;
wire n_4943;
wire n_2498;
wire n_7524;
wire n_4630;
wire n_3812;
wire n_6584;
wire n_6689;
wire n_2017;
wire n_1227;
wire n_5326;
wire n_3750;
wire n_5909;
wire n_6050;
wire n_3838;
wire n_5868;
wire n_1954;
wire n_4749;
wire n_1125;
wire n_6643;
wire n_2687;
wire n_3456;
wire n_6569;
wire n_6814;
wire n_3132;
wire n_5618;
wire n_6596;
wire n_7176;
wire n_4159;
wire n_7056;
wire n_4372;
wire n_5528;
wire n_4731;
wire n_4004;
wire n_1134;
wire n_1684;
wire n_7594;
wire n_4353;
wire n_5593;
wire n_3334;
wire n_3819;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_5740;
wire n_1233;
wire n_5108;
wire n_3653;
wire n_4360;
wire n_6123;
wire n_4897;
wire n_2139;
wire n_3693;
wire n_5477;
wire n_5934;
wire n_5218;
wire n_1138;
wire n_2943;
wire n_5272;
wire n_1096;
wire n_7535;
wire n_3135;
wire n_4239;
wire n_3175;
wire n_6273;
wire n_7368;
wire n_5464;
wire n_6895;
wire n_6548;
wire n_7627;
wire n_6420;
wire n_6474;
wire n_1268;
wire n_3187;
wire n_3830;
wire n_2724;
wire n_6890;
wire n_5688;
wire n_6141;
wire n_1829;
wire n_1338;
wire n_6234;
wire n_1327;
wire n_5204;
wire n_6789;
wire n_5400;
wire n_3407;
wire n_3315;
wire n_4470;
wire n_4690;
wire n_3982;
wire n_6311;
wire n_6867;
wire n_2565;
wire n_4201;
wire n_6634;
wire n_6288;
wire n_1636;
wire n_1687;
wire n_5303;
wire n_4584;
wire n_3184;
wire n_6290;
wire n_5804;
wire n_6764;
wire n_4155;
wire n_3890;
wire n_5519;
wire n_5023;
wire n_2032;
wire n_3392;
wire n_4802;
wire n_6935;
wire n_1258;
wire n_2208;
wire n_1344;
wire n_5971;
wire n_2198;
wire n_1929;
wire n_5095;
wire n_1680;
wire n_1195;
wire n_5902;
wire n_4304;
wire n_4975;
wire n_4821;
wire n_4160;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_4910;
wire n_5064;
wire n_6478;
wire n_7382;
wire n_3641;
wire n_5203;
wire n_5065;
wire n_4887;
wire n_5436;
wire n_7579;
wire n_3996;
wire n_7130;
wire n_6942;
wire n_6056;
wire n_7647;
wire n_2873;
wire n_1576;
wire n_6772;
wire n_6466;
wire n_3049;
wire n_4015;
wire n_4211;
wire n_4119;
wire n_3620;
wire n_2558;
wire n_2347;
wire n_3884;
wire n_3103;
wire n_3770;
wire n_4591;
wire n_2527;
wire n_5314;
wire n_7469;
wire n_5044;
wire n_1509;
wire n_2944;
wire n_1648;
wire n_4349;
wire n_1886;
wire n_6228;
wire n_1841;
wire n_6955;
wire n_5886;
wire n_2685;
wire n_5344;
wire n_1313;
wire n_4223;
wire n_2090;
wire n_5173;
wire n_5585;
wire n_3722;
wire n_5981;
wire n_3802;
wire n_5343;
wire n_5783;
wire n_2215;
wire n_1449;
wire n_1723;
wire n_3129;
wire n_5515;
wire n_4806;
wire n_2116;
wire n_5784;
wire n_5337;
wire n_3592;
wire n_5545;
wire n_1645;
wire n_3186;
wire n_6393;
wire n_7654;
wire n_6375;
wire n_7762;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_5209;
wire n_1269;
wire n_2773;
wire n_2906;
wire n_3097;
wire n_5495;
wire n_7427;
wire n_6908;
wire n_3910;
wire n_4238;
wire n_1466;
wire n_3667;
wire n_6424;
wire n_7506;
wire n_3822;
wire n_1276;
wire n_6874;
wire n_1637;
wire n_2900;
wire n_5799;
wire n_6296;
wire n_3765;
wire n_2216;
wire n_5888;
wire n_6736;
wire n_4259;
wire n_1620;
wire n_7376;
wire n_5196;
wire n_5086;
wire n_7018;
wire n_6025;
wire n_6168;
wire n_7498;
wire n_3518;
wire n_5885;
wire n_2022;
wire n_7134;
wire n_3967;
wire n_2373;
wire n_7456;
wire n_1853;
wire n_2275;
wire n_5398;
wire n_5434;
wire n_5797;
wire n_2899;
wire n_5830;
wire n_5896;
wire n_3351;
wire n_7480;
wire n_2008;
wire n_5052;
wire n_2859;
wire n_5952;
wire n_6003;
wire n_2564;
wire n_5110;
wire n_7348;
wire n_5918;
wire n_4799;
wire n_1356;
wire n_2591;
wire n_3965;
wire n_1969;
wire n_5808;
wire n_6119;
wire n_1296;
wire n_4444;
wire n_4676;
wire n_5212;
wire n_6525;
wire n_1764;
wire n_7383;
wire n_1250;
wire n_1190;
wire n_5733;
wire n_4598;
wire n_3259;
wire n_7053;
wire n_7660;
wire n_5483;
wire n_6713;
wire n_6919;
wire n_4533;
wire n_4078;
wire n_1794;
wire n_7557;
wire n_3779;
wire n_3203;
wire n_7240;
wire n_7468;
wire n_3923;
wire n_4392;
wire n_3808;
wire n_6750;
wire n_4455;
wire n_3093;
wire n_2664;
wire n_1434;
wire n_4129;
wire n_5278;
wire n_2114;
wire n_6204;
wire n_1609;
wire n_5522;
wire n_3530;
wire n_6981;
wire n_1132;
wire n_5584;
wire n_4548;
wire n_6675;
wire n_1803;
wire n_5264;
wire n_6321;
wire n_1281;
wire n_4535;
wire n_1447;
wire n_2150;
wire n_6337;
wire n_4999;
wire n_5328;
wire n_7604;
wire n_2660;
wire n_5447;
wire n_5029;
wire n_5127;
wire n_5006;
wire n_5679;
wire n_4604;
wire n_7585;
wire n_6828;
wire n_5123;
wire n_6160;
wire n_7043;
wire n_3467;
wire n_6156;
wire n_4240;
wire n_7074;
wire n_7119;
wire n_7596;
wire n_2219;
wire n_6116;
wire n_4522;
wire n_1387;
wire n_3371;
wire n_4713;
wire n_1368;
wire n_1154;
wire n_6267;
wire n_2539;
wire n_6875;
wire n_1701;
wire n_5236;
wire n_7567;
wire n_6678;
wire n_5239;
wire n_5307;
wire n_2387;
wire n_3375;
wire n_2397;
wire n_3317;
wire n_3963;
wire n_6870;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_6561;
wire n_6715;
wire n_2529;
wire n_4103;
wire n_4126;
wire n_4710;
wire n_5576;
wire n_3282;
wire n_5144;
wire n_2708;
wire n_5164;
wire n_6557;
wire n_2748;
wire n_5359;
wire n_7386;
wire n_6503;
wire n_5925;
wire n_2224;
wire n_5526;
wire n_5810;
wire n_2233;
wire n_2499;
wire n_6333;
wire n_5172;
wire n_3888;
wire n_4549;
wire n_3309;
wire n_5126;
wire n_1924;
wire n_3024;
wire n_7701;
wire n_4767;
wire n_7007;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_7027;
wire n_5999;
wire n_5147;
wire n_7616;
wire n_5407;
wire n_7432;
wire n_1553;
wire n_3542;
wire n_5536;
wire n_1090;
wire n_6002;
wire n_3374;
wire n_3704;
wire n_7661;
wire n_2786;
wire n_1905;
wire n_4355;
wire n_2958;
wire n_7009;
wire n_6140;
wire n_5903;
wire n_7263;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_4834;
wire n_6336;
wire n_3660;
wire n_2718;
wire n_4712;
wire n_5849;
wire n_7772;
wire n_6663;
wire n_1795;
wire n_7610;
wire n_3634;
wire n_4096;
wire n_6844;
wire n_2101;
wire n_5378;
wire n_1152;
wire n_3626;
wire n_2599;
wire n_6999;
wire n_4571;
wire n_7214;
wire n_6982;
wire n_5389;
wire n_6166;
wire n_3171;
wire n_6170;
wire n_1733;
wire n_6257;
wire n_7613;
wire n_3986;
wire n_2853;
wire n_1552;
wire n_6620;
wire n_4930;
wire n_5345;
wire n_2217;
wire n_3594;
wire n_2866;
wire n_5138;
wire n_3153;
wire n_6202;
wire n_1189;
wire n_4995;
wire n_6529;
wire n_4039;
wire n_4253;
wire n_4681;
wire n_2623;
wire n_6843;
wire n_3232;
wire n_5228;
wire n_2178;
wire n_1181;
wire n_3815;
wire n_4375;
wire n_5629;
wire n_5945;
wire n_4205;
wire n_6161;
wire n_3790;
wire n_6147;
wire n_2404;
wire n_5601;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_1203;
wire n_6554;
wire n_3640;
wire n_6877;
wire n_2821;
wire n_6892;
wire n_4768;
wire n_6133;
wire n_6109;
wire n_6585;
wire n_5985;
wire n_7162;
wire n_5435;
wire n_5665;
wire n_3299;
wire n_4070;
wire n_4558;
wire n_6436;
wire n_3065;
wire n_2375;
wire n_2572;
wire n_1656;
wire n_2063;
wire n_3082;
wire n_5709;
wire n_4504;
wire n_5176;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_4864;
wire n_3855;
wire n_3357;
wire n_4485;
wire n_1510;
wire n_5003;
wire n_2852;
wire n_2132;
wire n_5567;
wire n_1236;
wire n_3412;
wire n_5765;
wire n_1712;
wire n_6409;
wire n_4537;
wire n_5771;
wire n_5271;
wire n_1184;
wire n_2585;
wire n_7510;
wire n_2220;
wire n_4005;
wire n_1364;
wire n_3183;
wire n_4323;
wire n_5068;
wire n_4184;
wire n_2468;
wire n_5078;
wire n_7268;
wire n_3248;
wire n_2606;
wire n_5980;
wire n_7465;
wire n_4337;
wire n_4826;
wire n_7398;
wire n_2152;
wire n_5073;
wire n_5420;
wire n_6386;
wire n_5599;
wire n_4952;
wire n_3785;
wire n_3525;
wire n_5508;
wire n_2779;
wire n_1117;
wire n_2547;
wire n_6473;
wire n_1748;
wire n_7304;
wire n_7036;
wire n_2935;
wire n_5084;
wire n_6651;
wire n_7462;
wire n_2490;
wire n_3127;
wire n_7171;
wire n_3496;
wire n_3568;
wire n_5789;
wire n_4876;
wire n_5322;
wire n_6490;
wire n_3841;
wire n_4626;
wire n_1334;
wire n_7678;
wire n_7597;
wire n_3879;
wire n_6558;
wire n_2402;
wire n_1200;
wire n_2379;
wire n_2300;
wire n_1120;
wire n_6500;
wire n_5590;
wire n_5638;
wire n_4747;
wire n_5152;
wire n_3341;
wire n_4347;
wire n_1852;
wire n_3868;
wire n_4791;
wire n_5497;
wire n_2481;
wire n_4409;
wire n_5361;
wire n_7293;
wire n_1264;
wire n_6752;
wire n_2808;
wire n_5010;
wire n_6363;
wire n_3396;
wire n_6007;
wire n_2102;
wire n_7568;
wire n_3492;
wire n_3558;
wire n_2751;
wire n_1548;
wire n_4824;
wire n_5117;
wire n_2977;
wire n_1682;
wire n_6142;
wire n_3599;
wire n_7363;
wire n_6244;
wire n_1896;
wire n_1704;
wire n_2234;
wire n_6369;
wire n_6518;
wire n_5050;
wire n_5608;
wire n_5610;
wire n_4152;
wire n_6698;
wire n_1352;
wire n_5125;
wire n_2328;
wire n_6977;
wire n_6578;
wire n_4587;
wire n_6118;
wire n_6429;
wire n_6158;
wire n_2332;
wire n_7511;
wire n_7028;
wire n_1628;
wire n_6810;
wire n_1773;
wire n_7237;
wire n_3580;
wire n_2369;
wire n_5474;
wire n_3584;
wire n_4500;
wire n_5845;
wire n_1115;
wire n_1395;
wire n_7039;
wire n_4660;
wire n_2823;
wire n_3274;
wire n_2613;
wire n_6049;
wire n_2419;
wire n_6671;
wire n_6791;
wire n_5794;
wire n_5299;
wire n_2807;
wire n_4047;
wire n_5905;
wire n_4157;
wire n_3956;
wire n_1431;
wire n_5202;
wire n_6967;
wire n_5170;
wire n_5724;
wire n_6610;
wire n_7442;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_6108;
wire n_2241;
wire n_7618;
wire n_6768;
wire n_2458;
wire n_7489;
wire n_7144;
wire n_3401;
wire n_3032;
wire n_7362;
wire n_5042;
wire n_1750;
wire n_2833;
wire n_3179;
wire n_6382;
wire n_5662;
wire n_1563;
wire n_4051;
wire n_3123;
wire n_6576;
wire n_1875;
wire n_6947;
wire n_1615;
wire n_3719;
wire n_5334;
wire n_5595;
wire n_6938;
wire n_7765;
wire n_6260;
wire n_5244;
wire n_7453;
wire n_2635;
wire n_4077;
wire n_3897;
wire n_3475;
wire n_2077;
wire n_2520;
wire n_2193;
wire n_4010;
wire n_4942;
wire n_4255;
wire n_5692;
wire n_2908;
wire n_4561;
wire n_6906;
wire n_4957;
wire n_2053;
wire n_1580;
wire n_5728;
wire n_7758;
wire n_2200;
wire n_2304;
wire n_4683;
wire n_6148;
wire n_6404;
wire n_1439;
wire n_2352;
wire n_4839;
wire n_2185;
wire n_7124;
wire n_2476;
wire n_1266;
wire n_4814;
wire n_2781;
wire n_6217;
wire n_6324;
wire n_6918;
wire n_2460;
wire n_4694;
wire n_3600;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_2308;
wire n_3498;
wire n_4520;
wire n_1428;
wire n_4026;
wire n_7143;
wire n_2903;
wire n_3659;
wire n_5795;
wire n_4496;
wire n_6048;
wire n_1528;
wire n_3840;
wire n_5889;
wire n_5856;
wire n_7606;
wire n_3481;
wire n_4719;
wire n_4100;
wire n_3517;
wire n_5722;
wire n_2464;
wire n_1413;
wire n_6834;
wire n_5498;
wire n_2925;
wire n_2270;
wire n_5034;
wire n_5725;
wire n_6812;
wire n_1706;
wire n_1592;
wire n_6110;
wire n_1461;
wire n_2695;
wire n_6300;
wire n_5657;
wire n_3656;
wire n_3137;
wire n_3116;
wire n_4426;
wire n_5282;
wire n_5511;
wire n_7123;
wire n_2414;
wire n_5736;
wire n_5642;
wire n_6624;
wire n_3316;
wire n_2465;
wire n_3925;
wire n_4089;
wire n_1683;
wire n_7072;
wire n_4175;
wire n_4458;
wire n_7488;
wire n_6001;
wire n_3955;
wire n_3158;
wire n_3657;
wire n_5776;
wire n_5826;
wire n_6687;
wire n_2684;
wire n_1104;
wire n_2205;
wire n_2875;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_5932;
wire n_4185;
wire n_2064;
wire n_3088;
wire n_1497;
wire n_2002;
wire n_7734;
wire n_6088;
wire n_6762;
wire n_4815;
wire n_2545;
wire n_2050;
wire n_3695;
wire n_6239;
wire n_2500;
wire n_6992;
wire n_7109;
wire n_1917;
wire n_1444;
wire n_6091;
wire n_4316;
wire n_5453;
wire n_3328;
wire n_2763;
wire n_7644;
wire n_5136;
wire n_6352;
wire n_2761;
wire n_4020;
wire n_5494;
wire n_6101;
wire n_1920;
wire n_4306;
wire n_6319;
wire n_2997;
wire n_3735;
wire n_2127;
wire n_6188;
wire n_5718;
wire n_5634;
wire n_3028;
wire n_3228;
wire n_5079;
wire n_3706;
wire n_6395;
wire n_1432;
wire n_3322;
wire n_7325;
wire n_1174;
wire n_6037;
wire n_4512;
wire n_4483;
wire n_3499;
wire n_3552;
wire n_4164;
wire n_1286;
wire n_6759;
wire n_3784;
wire n_4142;
wire n_6206;
wire n_7137;
wire n_4621;
wire n_7526;
wire n_3016;
wire n_7699;
wire n_1629;
wire n_5706;
wire n_7350;
wire n_2694;
wire n_6177;
wire n_3609;
wire n_3447;
wire n_3771;
wire n_4678;
wire n_2647;
wire n_1850;
wire n_1670;
wire n_4123;
wire n_7311;
wire n_7458;
wire n_2317;
wire n_1384;
wire n_1612;
wire n_5496;
wire n_1099;
wire n_3113;
wire n_4305;
wire n_2909;
wire n_4007;
wire n_3960;
wire n_7244;
wire n_1524;
wire n_7681;
wire n_4707;
wire n_4429;
wire n_1991;
wire n_2566;
wire n_7339;
wire n_2210;
wire n_5606;
wire n_6322;
wire n_1225;
wire n_7247;
wire n_2346;
wire n_4695;
wire n_7331;
wire n_7128;
wire n_2180;
wire n_3376;
wire n_6313;
wire n_5989;
wire n_2617;
wire n_5870;
wire n_7284;
wire n_4163;
wire n_7321;
wire n_2831;
wire n_6504;
wire n_2865;
wire n_1625;
wire n_4638;
wire n_5530;
wire n_4498;
wire n_2240;
wire n_7309;
wire n_1797;
wire n_4750;
wire n_3993;
wire n_7163;
wire n_2120;
wire n_1289;
wire n_1557;
wire n_1567;
wire n_2007;
wire n_2004;
wire n_5424;
wire n_5230;
wire n_2086;
wire n_6886;
wire n_4832;
wire n_5229;
wire n_7054;
wire n_3666;
wire n_6374;
wire n_1839;
wire n_5160;
wire n_2330;
wire n_1587;
wire n_2555;
wire n_6356;
wire n_6640;
wire n_5313;
wire n_2108;
wire n_6462;
wire n_5333;
wire n_5207;
wire n_2535;
wire n_6959;
wire n_5158;
wire n_2945;
wire n_5154;
wire n_3057;
wire n_7413;
wire n_4319;
wire n_3760;
wire n_5721;
wire n_7185;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_5654;
wire n_2196;
wire n_5860;
wire n_1538;
wire n_3773;
wire n_6710;
wire n_5884;
wire n_2604;
wire n_3462;
wire n_4373;
wire n_6945;
wire n_2351;
wire n_2437;
wire n_1889;
wire n_6776;
wire n_1124;
wire n_5839;
wire n_2688;
wire n_4990;
wire n_7336;
wire n_3302;
wire n_1673;
wire n_5058;
wire n_2085;
wire n_3304;
wire n_1725;
wire n_6231;
wire n_2149;
wire n_7630;
wire n_2001;
wire n_1800;
wire n_3746;
wire n_6905;
wire n_7737;
wire n_7120;
wire n_3645;
wire n_5823;
wire n_4262;
wire n_4019;
wire n_2735;
wire n_6401;
wire n_2035;
wire n_4436;
wire n_4697;
wire n_1906;
wire n_1647;
wire n_4357;
wire n_7374;
wire n_6521;
wire n_4849;
wire n_5101;
wire n_5532;
wire n_4366;
wire n_6582;
wire n_7491;
wire n_6964;
wire n_4139;
wire n_1270;
wire n_5297;
wire n_4340;
wire n_1476;
wire n_7001;
wire n_2027;
wire n_5611;
wire n_2012;
wire n_3512;
wire n_4720;
wire n_3892;
wire n_7111;
wire n_6623;
wire n_1880;
wire n_6225;
wire n_7519;
wire n_1642;
wire n_5744;
wire n_6798;
wire n_2447;
wire n_3358;
wire n_5538;
wire n_2894;
wire n_5249;
wire n_5669;
wire n_2587;
wire n_1605;
wire n_6134;
wire n_2099;
wire n_1202;
wire n_5793;
wire n_3410;
wire n_4900;
wire n_6493;
wire n_6364;
wire n_5715;
wire n_6665;
wire n_7538;
wire n_3408;
wire n_3182;
wire n_1879;
wire n_4941;
wire n_1311;
wire n_5966;
wire n_2299;
wire n_2078;
wire n_6284;
wire n_3709;
wire n_3011;
wire n_5383;
wire n_6649;
wire n_5775;
wire n_2315;
wire n_3623;
wire n_6230;
wire n_5558;
wire n_7165;
wire n_2157;
wire n_6546;
wire n_3446;
wire n_5547;
wire n_5572;
wire n_5659;
wire n_5223;
wire n_6555;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_6010;
wire n_3058;
wire n_4334;
wire n_6331;
wire n_6888;
wire n_2211;
wire n_6047;
wire n_5708;
wire n_7599;
wire n_6532;
wire n_5817;
wire n_3384;
wire n_4698;
wire n_6677;
wire n_2225;
wire n_1411;
wire n_5867;
wire n_7389;
wire n_1501;
wire n_7418;
wire n_5636;
wire n_5106;
wire n_5800;
wire n_7375;
wire n_7671;
wire n_7096;
wire n_5257;
wire n_7719;
wire n_7281;
wire n_7300;
wire n_4397;
wire n_6920;
wire n_3611;
wire n_4186;
wire n_2093;
wire n_2675;
wire n_5371;
wire n_6524;
wire n_6781;
wire n_4229;
wire n_4294;
wire n_7085;
wire n_1919;
wire n_4351;
wire n_6811;
wire n_6226;
wire n_2893;
wire n_6281;
wire n_2009;
wire n_6514;
wire n_5731;
wire n_4162;
wire n_1416;
wire n_3465;
wire n_7683;
wire n_1515;
wire n_6921;
wire n_4127;
wire n_4620;
wire n_1314;
wire n_3059;
wire n_3085;
wire n_2867;
wire n_2229;
wire n_4770;
wire n_7212;
wire n_7285;
wire n_7676;
wire n_3871;
wire n_2388;
wire n_6685;
wire n_7590;
wire n_3112;
wire n_5623;
wire n_5921;
wire n_6082;
wire n_3413;
wire n_4580;
wire n_7032;
wire n_2624;
wire n_1813;
wire n_4581;
wire n_4618;
wire n_7125;
wire n_5178;
wire n_6609;
wire n_5853;
wire n_7160;
wire n_7100;
wire n_1105;
wire n_5898;
wire n_5198;
wire n_2898;
wire n_5437;
wire n_6627;
wire n_2519;
wire n_2231;
wire n_2816;
wire n_2803;
wire n_3402;
wire n_5053;
wire n_1256;
wire n_4670;
wire n_7319;
wire n_6162;
wire n_7638;
wire n_5592;
wire n_5484;
wire n_6650;
wire n_5418;
wire n_4982;
wire n_6079;
wire n_6013;
wire n_5432;
wire n_1769;
wire n_7635;
wire n_5270;
wire n_1372;
wire n_1847;
wire n_5166;
wire n_5358;
wire n_3805;
wire n_2406;
wire n_4017;
wire n_7504;
wire n_1586;
wire n_3497;
wire n_6722;
wire n_5156;
wire n_6592;
wire n_3382;
wire n_4236;
wire n_4313;
wire n_5548;
wire n_5687;
wire n_3561;
wire n_2543;
wire n_6512;
wire n_2992;
wire n_1541;
wire n_6008;
wire n_6522;
wire n_4907;
wire n_4659;
wire n_2128;
wire n_1697;
wire n_1872;
wire n_5822;
wire n_2690;
wire n_3942;
wire n_2020;
wire n_5758;
wire n_1939;
wire n_7767;
wire n_5366;
wire n_4053;
wire n_5392;
wire n_4279;
wire n_3937;
wire n_6400;
wire n_7371;
wire n_3303;
wire n_5115;
wire n_5046;
wire n_7361;
wire n_5139;
wire n_4555;
wire n_5829;
wire n_5686;
wire n_7440;
wire n_5735;
wire n_3549;
wire n_1481;
wire n_6613;
wire n_1928;
wire n_4235;
wire n_3972;
wire n_5674;
wire n_2314;
wire n_2126;
wire n_3403;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_1361;
wire n_5039;
wire n_6538;
wire n_1693;
wire n_2081;
wire n_5341;
wire n_2993;
wire n_7010;
wire n_5032;
wire n_3018;
wire n_4820;
wire n_2449;
wire n_2131;
wire n_7289;
wire n_2526;
wire n_4794;
wire n_1302;
wire n_5041;
wire n_6505;
wire n_3989;
wire n_6581;
wire n_5565;
wire n_7004;
wire n_7021;
wire n_6350;
wire n_4752;
wire n_4546;
wire n_7234;
wire n_3918;
wire n_6378;
wire n_3191;
wire n_3051;
wire n_6975;
wire n_7266;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_4415;
wire n_2487;
wire n_3343;
wire n_3163;
wire n_6243;
wire n_3786;
wire n_4061;
wire n_4432;
wire n_6484;
wire n_1912;
wire n_4552;
wire n_3143;
wire n_1876;
wire n_7754;
wire n_6573;
wire n_6786;
wire n_6774;
wire n_6419;
wire n_4790;
wire n_1811;
wire n_1285;
wire n_5448;
wire n_4263;
wire n_3725;
wire n_5974;
wire n_5852;
wire n_6143;
wire n_6851;
wire n_1529;
wire n_1824;
wire n_3522;
wire n_4528;
wire n_4888;
wire n_4502;
wire n_5085;
wire n_7211;
wire n_4335;
wire n_7141;
wire n_3444;
wire n_4218;
wire n_4705;
wire n_6112;
wire n_6138;
wire n_3009;
wire n_4471;
wire n_1141;
wire n_3297;
wire n_6729;
wire n_7150;
wire n_6882;
wire n_1168;
wire n_5500;
wire n_7378;
wire n_6045;
wire n_5293;
wire n_6203;
wire n_7470;
wire n_3000;
wire n_2305;
wire n_1192;
wire n_1290;
wire n_2514;
wire n_4386;
wire n_6568;
wire n_4547;
wire n_7633;
wire n_4836;
wire n_5458;
wire n_3545;
wire n_1101;
wire n_4193;
wire n_5670;
wire n_7420;
wire n_1336;
wire n_6433;
wire n_6023;
wire n_1358;
wire n_3318;
wire n_5684;
wire n_1397;
wire n_1359;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_4984;
wire n_1532;
wire n_5624;
wire n_3430;
wire n_1685;
wire n_7558;
wire n_5325;
wire n_2801;
wire n_3225;
wire n_3067;
wire n_6189;
wire n_6167;
wire n_5059;
wire n_1462;
wire n_5825;
wire n_3823;
wire n_4718;
wire n_3185;
wire n_2326;
wire n_5586;
wire n_6998;
wire n_1398;
wire n_5222;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_4634;
wire n_6335;
wire n_5741;
wire n_1692;
wire n_5875;
wire n_6721;
wire n_4796;
wire n_6312;
wire n_4560;
wire n_1240;
wire n_3285;
wire n_5045;
wire n_7640;
wire n_1814;
wire n_4882;
wire n_1808;
wire n_2768;
wire n_1658;
wire n_6611;
wire n_7484;
wire n_5038;
wire n_5769;
wire n_3837;
wire n_7708;
wire n_4841;
wire n_6213;
wire n_3076;
wire n_6264;
wire n_4954;
wire n_4635;
wire n_4521;
wire n_5703;
wire n_3893;
wire n_4272;
wire n_2148;
wire n_2104;
wire n_2653;
wire n_2855;
wire n_6301;
wire n_2618;
wire n_7598;
wire n_4448;
wire n_3359;
wire n_5501;
wire n_6216;
wire n_2331;
wire n_1600;
wire n_7271;
wire n_5894;
wire n_4701;
wire n_5248;
wire n_5872;
wire n_4088;
wire n_2136;
wire n_7322;
wire n_7549;
wire n_7022;
wire n_5443;
wire n_6193;
wire n_1913;
wire n_6885;
wire n_7217;
wire n_7166;
wire n_3056;
wire n_4208;
wire n_5363;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_6806;
wire n_4865;
wire n_2066;
wire n_7584;
wire n_1974;
wire n_1158;
wire n_6588;
wire n_4589;
wire n_3924;
wire n_6933;
wire n_1915;
wire n_2534;
wire n_5908;
wire n_4972;
wire n_5597;
wire n_4617;
wire n_3311;
wire n_1160;
wire n_4094;
wire n_4772;
wire n_4857;
wire n_7297;
wire n_7664;
wire n_3613;
wire n_1383;
wire n_7546;
wire n_2057;
wire n_7179;
wire n_5984;
wire n_6385;
wire n_7415;
wire n_5533;
wire n_1822;
wire n_6051;
wire n_1804;
wire n_1581;
wire n_7057;
wire n_5387;
wire n_4776;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_2246;
wire n_2738;
wire n_6793;
wire n_1851;
wire n_1755;
wire n_5589;
wire n_6746;
wire n_4702;
wire n_1341;
wire n_7411;
wire n_4486;
wire n_4946;
wire n_2202;
wire n_5380;
wire n_2262;
wire n_5134;
wire n_1333;
wire n_4506;
wire n_7108;
wire n_7736;
wire n_3157;
wire n_4669;
wire n_4226;
wire n_4153;
wire n_7220;
wire n_6015;
wire n_4329;
wire n_6435;
wire n_4877;
wire n_3442;
wire n_2327;
wire n_4780;
wire n_6411;
wire n_4327;
wire n_5954;
wire n_5412;
wire n_2656;
wire n_6323;
wire n_4168;
wire n_2258;
wire n_4396;
wire n_2039;
wire n_5174;
wire n_4465;
wire n_6174;
wire n_7223;
wire n_2544;
wire n_7261;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_3266;
wire n_7092;
wire n_5468;
wire n_1843;
wire n_2030;
wire n_4576;
wire n_6728;
wire n_4075;
wire n_5429;
wire n_3593;
wire n_6586;
wire n_2536;
wire n_1399;
wire n_3685;
wire n_5269;
wire n_4833;
wire n_1903;
wire n_1849;
wire n_7275;
wire n_3768;
wire n_4224;
wire n_7272;
wire n_4868;
wire n_5124;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_7436;
wire n_3181;
wire n_7249;
wire n_3644;
wire n_5287;
wire n_4387;
wire n_5865;
wire n_2368;
wire n_6437;
wire n_4896;
wire n_1157;
wire n_7168;
wire n_2065;
wire n_2901;
wire n_5583;
wire n_3818;
wire n_4368;
wire n_1295;
wire n_1983;
wire n_4798;
wire n_2201;
wire n_1582;
wire n_7712;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3610;
wire n_5416;
wire n_7743;
wire n_2569;
wire n_7705;
wire n_1998;
wire n_1596;
wire n_3077;
wire n_7091;
wire n_1100;
wire n_4158;
wire n_4687;
wire n_4756;
wire n_4095;
wire n_2177;
wire n_2123;
wire n_4364;
wire n_3019;
wire n_2235;
wire n_5373;
wire n_4967;
wire n_6067;
wire n_6858;
wire n_7679;
wire n_5377;
wire n_2290;
wire n_6479;
wire n_7228;
wire n_3272;
wire n_7353;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_5350;
wire n_6279;
wire n_6841;
wire n_4668;
wire n_7696;
wire n_2383;
wire n_5632;
wire n_2640;
wire n_7687;
wire n_1492;
wire n_6425;
wire n_1478;
wire n_6896;
wire n_1796;
wire n_3569;
wire n_2374;
wire n_1614;
wire n_4648;
wire n_2598;
wire n_1722;
wire n_5290;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_4785;
wire n_5120;
wire n_2230;
wire n_5535;
wire n_3033;
wire n_2151;
wire n_5382;
wire n_6354;
wire n_4912;
wire n_6320;
wire n_1971;
wire n_5759;
wire n_2479;
wire n_4914;
wire n_6954;
wire n_2359;
wire n_2360;
wire n_4902;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_6612;
wire n_6376;
wire n_2571;
wire n_7000;
wire n_5479;
wire n_6006;
wire n_5598;
wire n_7040;
wire n_6132;
wire n_7196;
wire n_2799;
wire n_7655;
wire n_4708;
wire n_4592;
wire n_1307;
wire n_5578;
wire n_2644;
wire n_4445;
wire n_3211;
wire n_1840;
wire n_2837;
wire n_6872;
wire n_6089;
wire n_5211;
wire n_7205;
wire n_1668;
wire n_7260;
wire n_7500;
wire n_5861;
wire n_7086;
wire n_6417;
wire n_1681;
wire n_4031;
wire n_7569;
wire n_4120;
wire n_3533;
wire n_3896;
wire n_2192;
wire n_7763;
wire n_4578;
wire n_3323;
wire n_1937;
wire n_3839;
wire n_3509;
wire n_1749;
wire n_2918;
wire n_3353;
wire n_5092;
wire n_1945;
wire n_5182;
wire n_5430;
wire n_2638;
wire n_3939;
wire n_7577;
wire n_4874;
wire n_1228;
wire n_7047;
wire n_7412;
wire n_4840;
wire n_7717;
wire n_2354;
wire n_5956;
wire n_6027;
wire n_6477;
wire n_4311;
wire n_5766;
wire n_6269;
wire n_1133;
wire n_1926;
wire n_2363;
wire n_2814;
wire n_5094;
wire n_6275;
wire n_3264;
wire n_3204;
wire n_6390;
wire n_2003;
wire n_3727;
wire n_2621;
wire n_2922;
wire n_6306;
wire n_3881;
wire n_1910;
wire n_5446;
wire n_1606;
wire n_5315;
wire n_3711;
wire n_7077;
wire n_2164;
wire n_7565;
wire n_1618;
wire n_3748;
wire n_4389;
wire n_3668;
wire n_3197;
wire n_1955;
wire n_4556;
wire n_2413;
wire n_3148;
wire n_4779;
wire n_6122;
wire n_1253;
wire n_1484;
wire n_2686;
wire n_4214;
wire n_4430;
wire n_3151;
wire n_3977;
wire n_3125;
wire n_2812;
wire n_4889;
wire n_4221;
wire n_1638;
wire n_6831;
wire n_6175;
wire n_5279;
wire n_6506;
wire n_6690;
wire n_4650;
wire n_6968;
wire n_6415;
wire n_2280;
wire n_7576;
wire n_4428;
wire n_4784;
wire n_2393;
wire n_4766;
wire n_7523;
wire n_3809;
wire n_1999;
wire n_3810;
wire n_5103;
wire n_5835;
wire n_4968;
wire n_1215;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_5311;
wire n_2283;
wire n_2806;
wire n_6184;
wire n_2813;
wire n_5268;
wire n_4295;
wire n_1716;
wire n_1412;
wire n_6285;
wire n_5773;
wire n_3310;
wire n_4182;
wire n_7750;
wire n_1401;
wire n_2951;
wire n_5451;
wire n_7578;
wire n_5452;
wire n_2145;
wire n_2122;
wire n_6644;
wire n_1588;
wire n_2579;
wire n_6688;
wire n_7402;
wire n_2876;
wire n_6670;
wire n_7473;
wire n_3301;
wire n_2370;
wire n_5321;
wire n_5215;
wire n_4600;
wire n_2025;
wire n_3451;
wire n_1219;
wire n_6680;
wire n_4513;
wire n_5635;
wire n_1252;
wire n_2730;
wire n_1927;
wire n_5356;
wire n_4735;
wire n_2767;
wire n_4667;
wire n_5150;
wire n_2826;
wire n_2112;
wire n_6180;
wire n_5613;
wire n_7405;
wire n_6137;
wire n_2762;
wire n_4774;
wire n_4711;
wire n_3023;
wire n_7343;
wire n_3224;
wire n_7721;
wire n_4481;
wire n_3762;
wire n_6410;
wire n_5063;
wire n_4671;
wire n_6046;
wire n_1326;
wire n_4981;
wire n_1799;
wire n_7252;
wire n_1689;
wire n_1304;
wire n_6465;
wire n_5653;
wire n_2541;
wire n_4879;
wire n_2987;
wire n_5788;
wire n_1702;
wire n_3916;
wire n_3630;
wire n_1558;
wire n_2722;
wire n_5057;
wire n_3618;
wire n_2727;
wire n_6991;
wire n_5560;
wire n_2719;
wire n_2213;
wire n_5476;
wire n_3521;
wire n_6121;
wire n_2723;
wire n_6077;
wire n_4054;
wire n_1569;
wire n_6000;
wire n_6205;
wire n_4012;
wire n_5582;
wire n_6705;
wire n_3567;
wire n_7601;
wire n_4352;
wire n_1988;
wire n_5935;
wire n_6201;
wire n_2401;
wire n_1787;
wire n_3094;
wire n_2166;
wire n_2451;
wire n_4665;
wire n_2631;
wire n_1867;
wire n_5697;
wire n_4252;
wire n_4505;
wire n_4219;
wire n_5119;
wire n_2292;
wire n_7451;
wire n_6471;
wire n_3560;
wire n_5813;
wire n_1742;
wire n_1818;
wire n_5100;
wire n_3847;
wire n_2203;
wire n_5427;
wire n_4909;
wire n_2693;
wire n_1159;
wire n_2281;
wire n_3202;
wire n_7603;
wire n_7575;
wire n_7188;
wire n_6913;
wire n_5467;
wire n_2646;
wire n_7525;
wire n_5346;
wire n_3887;
wire n_3800;
wire n_7528;
wire n_7113;
wire n_4435;
wire n_1235;
wire n_6355;
wire n_4755;
wire n_6329;
wire n_3827;
wire n_6145;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_5633;
wire n_7637;
wire n_1835;
wire n_2697;
wire n_3531;
wire n_2470;
wire n_5726;
wire n_2890;
wire n_6734;
wire n_4400;
wire n_1519;
wire n_1425;
wire n_4812;
wire n_5415;
wire n_2069;
wire n_2602;
wire n_4090;
wire n_5445;
wire n_6446;
wire n_4996;
wire n_4136;
wire n_5040;
wire n_7471;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_5031;
wire n_1360;
wire n_5814;
wire n_5374;
wire n_2070;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3039;
wire n_7296;
wire n_3900;
wire n_3478;
wire n_3701;
wire n_2766;
wire n_3756;
wire n_3754;
wire n_4156;
wire n_6057;
wire n_5818;
wire n_7781;
wire n_2416;
wire n_2962;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_6221;
wire n_5876;
wire n_5529;
wire n_3006;
wire n_3348;
wire n_4758;
wire n_2236;
wire n_5317;
wire n_3957;
wire n_2377;
wire n_2577;
wire n_3165;
wire n_4419;
wire n_2795;
wire n_7741;
wire n_5490;
wire n_3520;
wire n_2632;
wire n_4406;
wire n_7727;
wire n_6825;
wire n_5897;
wire n_5331;
wire n_6107;
wire n_6743;
wire n_1106;
wire n_4655;
wire n_6080;
wire n_1634;
wire n_5556;
wire n_1452;
wire n_4953;
wire n_7345;
wire n_7472;
wire n_6339;
wire n_4570;
wire n_5391;
wire n_5431;
wire n_3966;
wire n_4293;
wire n_6371;
wire n_6014;
wire n_1577;
wire n_1700;
wire n_4122;
wire n_4542;
wire n_5021;
wire n_2819;
wire n_5456;
wire n_5523;
wire n_1985;
wire n_1140;
wire n_4740;
wire n_3007;
wire n_1487;
wire n_6373;
wire n_1237;
wire n_4230;
wire n_7157;
wire n_1109;
wire n_2741;
wire n_4333;
wire n_7674;
wire n_5231;
wire n_6809;
wire n_5512;
wire n_6406;
wire n_3436;
wire n_6223;
wire n_4460;
wire n_2312;
wire n_2946;
wire n_4040;
wire n_7622;
wire n_7115;
wire n_1884;
wire n_6632;
wire n_2717;
wire n_1589;
wire n_5720;
wire n_7286;
wire n_4527;
wire n_2877;
wire n_5881;
wire n_1996;
wire n_5857;
wire n_5256;
wire n_3964;
wire n_3110;
wire n_5717;
wire n_1677;
wire n_4384;
wire n_2297;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_1792;
wire n_6654;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_4762;
wire n_5561;
wire n_1877;
wire n_6871;
wire n_1477;
wire n_3155;
wire n_4938;
wire n_5487;
wire n_4407;
wire n_5961;
wire n_5077;
wire n_6672;
wire n_5214;
wire n_1249;
wire n_3468;
wire n_7344;
wire n_2006;
wire n_7714;
wire n_1990;
wire n_5413;
wire n_3680;
wire n_6227;
wire n_7612;
wire n_3624;
wire n_6098;
wire n_4989;
wire n_7744;
wire n_2467;
wire n_5066;
wire n_4292;
wire n_6953;
wire n_7779;
wire n_3145;
wire n_5682;
wire n_6891;
wire n_2662;
wire n_3872;
wire n_5602;
wire n_3801;
wire n_2883;
wire n_1178;
wire n_6163;
wire n_1464;
wire n_1566;
wire n_7127;
wire n_6565;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_6601;
wire n_2277;
wire n_1982;
wire n_2252;
wire n_1695;
wire n_3331;
wire n_2999;
wire n_2910;
wire n_4414;
wire n_6979;
wire n_2294;
wire n_2295;
wire n_4977;
wire n_4706;
wire n_1602;
wire n_2965;
wire n_6076;
wire n_7650;
wire n_5347;
wire n_2382;
wire n_2557;
wire n_2505;
wire n_7050;
wire n_3554;
wire n_7431;
wire n_6199;
wire n_3730;
wire n_4307;
wire n_4356;
wire n_6930;
wire n_1935;
wire n_7770;
wire n_5568;
wire n_3367;
wire n_1146;
wire n_2785;
wire n_7118;
wire n_7259;
wire n_5060;
wire n_4929;
wire n_5121;
wire n_1608;
wire n_3776;
wire n_4951;
wire n_5756;
wire n_5162;
wire n_5224;
wire n_2160;
wire n_2699;
wire n_2991;
wire n_6513;
wire n_6214;
wire n_1436;
wire n_6821;
wire n_4137;
wire n_1485;
wire n_7448;
wire n_2239;
wire n_6289;
wire n_3826;
wire n_4365;
wire n_1979;
wire n_3781;
wire n_6775;
wire n_4215;
wire n_4315;
wire n_6559;
wire n_2971;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_7518;
wire n_3797;
wire n_6683;
wire n_3281;
wire n_3505;
wire n_4427;
wire n_4564;
wire n_2934;
wire n_6815;
wire n_6430;
wire n_4042;
wire n_5663;
wire n_2525;
wire n_5552;
wire n_4624;
wire n_6043;
wire n_4317;
wire n_3087;
wire n_7726;
wire n_4925;
wire n_2197;
wire n_7069;
wire n_1470;
wire n_2098;
wire n_1761;
wire n_4041;
wire n_5672;
wire n_7478;
wire n_4958;
wire n_5051;
wire n_4297;
wire n_5367;
wire n_5339;
wire n_4709;
wire n_3379;
wire n_4425;
wire n_3390;
wire n_5000;
wire n_1806;
wire n_1539;
wire n_2711;
wire n_3646;
wire n_7011;
wire n_2209;
wire n_3020;
wire n_3142;
wire n_2612;
wire n_5226;
wire n_2095;
wire n_2486;
wire n_5855;
wire n_5819;
wire n_2521;
wire n_5388;
wire n_1574;
wire n_6608;
wire n_7686;
wire n_6186;
wire n_4764;
wire n_4899;
wire n_6283;
wire n_6445;
wire n_7716;
wire n_4141;
wire n_4614;
wire n_2979;
wire n_4739;
wire n_1300;
wire n_4035;
wire n_4291;
wire n_6372;
wire n_3419;
wire n_4935;
wire n_4880;
wire n_7759;
wire n_3167;
wire n_5188;
wire n_2986;
wire n_4969;
wire n_7675;
wire n_2400;
wire n_6467;
wire n_6144;
wire n_5681;
wire n_2507;
wire n_3682;
wire n_3131;
wire n_1495;
wire n_6291;
wire n_1357;
wire n_6593;
wire n_7482;
wire n_4566;
wire n_5262;
wire n_2794;
wire n_6542;
wire n_3672;
wire n_2496;
wire n_4918;
wire n_2974;
wire n_6763;
wire n_6782;
wire n_7621;
wire n_5604;
wire n_3449;
wire n_2923;
wire n_2990;
wire n_1339;
wire n_1544;
wire n_4933;
wire n_4872;
wire n_5910;
wire n_1315;
wire n_4647;
wire n_7552;
wire n_6839;
wire n_2340;
wire n_6125;
wire n_2117;
wire n_5990;
wire n_1328;
wire n_4837;
wire n_6218;
wire n_3638;
wire n_2106;
wire n_5880;
wire n_5685;
wire n_7164;
wire n_6619;
wire n_6515;
wire n_6060;
wire n_1263;
wire n_4940;
wire n_4176;
wire n_4454;
wire n_7017;
wire n_7454;
wire n_6664;
wire n_5992;
wire n_5105;
wire n_6761;
wire n_5807;
wire n_3772;
wire n_7769;
wire n_2948;
wire n_4322;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_5449;
wire n_3867;
wire n_4956;
wire n_2045;
wire n_1535;
wire n_4227;
wire n_6599;
wire n_2190;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_3929;
wire n_6974;
wire n_1898;
wire n_1254;
wire n_7312;
wire n_6894;
wire n_2524;
wire n_3927;
wire n_7045;
wire n_1941;
wire n_5338;
wire n_5070;
wire n_3564;
wire n_3095;
wire n_1783;
wire n_5842;
wire n_3279;
wire n_1815;
wire n_3344;
wire n_6173;
wire n_4133;
wire n_6093;
wire n_3985;
wire n_7277;
wire n_6099;
wire n_5939;
wire n_7502;
wire n_5481;
wire n_5187;
wire n_5762;
wire n_3252;
wire n_1162;
wire n_2578;
wire n_5486;
wire n_5426;
wire n_2745;
wire n_2110;
wire n_6031;
wire n_6064;
wire n_6997;
wire n_3747;
wire n_1323;
wire n_6753;
wire n_5846;
wire n_6033;
wire n_3710;
wire n_1429;
wire n_6316;
wire n_3209;
wire n_2026;
wire n_5537;
wire n_3588;
wire n_7778;
wire n_5220;
wire n_6341;
wire n_2103;
wire n_4497;
wire n_4388;
wire n_7359;
wire n_3632;
wire n_5200;
wire n_7225;
wire n_1874;
wire n_7651;
wire n_4116;
wire n_3377;
wire n_5816;
wire n_1601;
wire n_3414;
wire n_2933;
wire n_7020;
wire n_3828;
wire n_1367;
wire n_3240;
wire n_2895;
wire n_1458;
wire n_1694;
wire n_7392;
wire n_2271;
wire n_2356;
wire n_5676;
wire n_5463;
wire n_2261;
wire n_4066;
wire n_2994;
wire n_4980;
wire n_2105;
wire n_2187;
wire n_5780;
wire n_2642;
wire n_6924;
wire n_5485;
wire n_5737;
wire n_6876;
wire n_7424;
wire n_1643;
wire n_1789;
wire n_7625;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_3589;
wire n_6571;
wire n_1112;
wire n_2384;
wire n_6962;
wire n_1376;
wire n_1858;
wire n_3523;
wire n_2815;
wire n_2446;
wire n_3388;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_6039;
wire n_5355;
wire n_4048;
wire n_7059;
wire n_4084;
wire n_5149;
wire n_1527;
wire n_3174;
wire n_4848;
wire n_6970;
wire n_5185;
wire n_6829;
wire n_2849;
wire n_6509;
wire n_6642;
wire n_5847;
wire n_5091;
wire n_5936;
wire n_1177;
wire n_3292;
wire n_6442;
wire n_7522;
wire n_6636;
wire n_3940;
wire n_6475;
wire n_2502;
wire n_5396;
wire n_4860;
wire n_4438;
wire n_5300;
wire n_6830;
wire n_3290;
wire n_7365;
wire n_3585;
wire n_7094;
wire n_2878;
wire n_1810;
wire n_7439;
wire n_6342;
wire n_3047;
wire n_2610;
wire n_5917;
wire n_7035;
wire n_5306;
wire n_3427;
wire n_1188;
wire n_3431;
wire n_2024;
wire n_3783;
wire n_1503;
wire n_1942;
wire n_4326;
wire n_3141;
wire n_6838;
wire n_2698;
wire n_6869;
wire n_3930;
wire n_4149;
wire n_5518;
wire n_5531;
wire n_1259;
wire n_4101;
wire n_6735;
wire n_4792;
wire n_2916;
wire n_3736;
wire n_2611;
wire n_6012;
wire n_6866;
wire n_4383;
wire n_7395;
wire n_2709;
wire n_5074;
wire n_6492;
wire n_7005;
wire n_2244;
wire n_6387;
wire n_3664;
wire n_1456;
wire n_3907;
wire n_5246;
wire n_2665;
wire n_5544;
wire n_6742;
wire n_3063;
wire n_4543;
wire n_6969;
wire n_2881;
wire n_3862;
wire n_2018;
wire n_3134;
wire n_5652;
wire n_7180;
wire n_5409;
wire n_2581;
wire n_6271;
wire n_5540;
wire n_2237;
wire n_2268;
wire n_2320;
wire n_6929;
wire n_2255;
wire n_1820;
wire n_6986;
wire n_3906;
wire n_3474;
wire n_1946;
wire n_3111;
wire n_4212;
wire n_7752;
wire n_6709;
wire n_4827;
wire n_1639;
wire n_2154;
wire n_6149;
wire n_3162;
wire n_4599;
wire n_2732;
wire n_3004;
wire n_3333;
wire n_4509;
wire n_3705;
wire n_4783;
wire n_3276;
wire n_2956;
wire n_1415;
wire n_3743;
wire n_7724;
wire n_4068;
wire n_7385;
wire n_2153;
wire n_5777;
wire n_2891;
wire n_2457;
wire n_3825;
wire n_6545;
wire n_4434;
wire n_2737;
wire n_5557;
wire n_1406;
wire n_3591;
wire n_6054;
wire n_2137;
wire n_7444;
wire n_6756;
wire n_5442;
wire n_1473;
wire n_3140;
wire n_2125;
wire n_1176;
wire n_7620;
wire n_3848;
wire n_1897;
wire n_2477;
wire n_4622;
wire n_5549;
wire n_3139;
wire n_4715;
wire n_7441;
wire n_6250;
wire n_6718;
wire n_4222;
wire n_5730;
wire n_2206;
wire n_3734;
wire n_7078;
wire n_3538;
wire n_4716;
wire n_4588;
wire n_2265;
wire n_5054;
wire n_5349;
wire n_7093;
wire n_1167;
wire n_7333;
wire n_3231;
wire n_6423;
wire n_6659;
wire n_3138;
wire n_6303;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_3349;
wire n_7508;
wire n_4988;
wire n_5128;
wire n_3454;
wire n_6668;
wire n_6299;
wire n_4143;
wire n_5027;
wire n_4410;
wire n_5026;
wire n_5189;
wire n_1718;
wire n_3229;
wire n_6757;
wire n_2546;
wire n_4741;
wire n_6383;
wire n_5516;
wire n_1139;
wire n_2345;
wire n_1324;
wire n_4440;
wire n_7496;
wire n_3649;
wire n_1838;
wire n_6880;
wire n_3824;
wire n_7425;
wire n_3439;
wire n_5525;
wire n_1513;
wire n_5836;
wire n_5677;
wire n_6182;
wire n_6510;
wire n_1788;
wire n_5764;
wire n_2348;
wire n_6171;
wire n_2417;
wire n_7550;
wire n_2043;
wire n_3601;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_7715;
wire n_5768;
wire n_6353;
wire n_7302;
wire n_6472;
wire n_2248;
wire n_3500;
wire n_2850;
wire n_3962;
wire n_6360;
wire n_3846;
wire n_4328;
wire n_7548;
wire n_5142;
wire n_1433;
wire n_6934;
wire n_5082;
wire n_1907;
wire n_6686;
wire n_7019;
wire n_3994;
wire n_5911;
wire n_5118;
wire n_2135;
wire n_5781;
wire n_5739;
wire n_7595;
wire n_1088;
wire n_7088;
wire n_6666;
wire n_6075;
wire n_1102;
wire n_5145;
wire n_7542;
wire n_4487;
wire n_7204;
wire n_7014;
wire n_1165;
wire n_6708;
wire n_5111;
wire n_4148;
wire n_3066;
wire n_6135;
wire n_2869;
wire n_6422;
wire n_4829;
wire n_2455;
wire n_2874;
wire n_4937;
wire n_7665;
wire n_4463;
wire n_2284;
wire n_1931;
wire n_7341;
wire n_7407;
wire n_6266;
wire n_5748;
wire n_1809;
wire n_7757;
wire n_3491;
wire n_4844;
wire n_3271;
wire n_5734;
wire n_2667;
wire n_7514;
wire n_6317;
wire n_7646;
wire n_7653;
wire n_6059;
wire n_5247;
wire n_1565;
wire n_2325;
wire n_6041;
wire n_3346;
wire n_5411;
wire n_5422;
wire n_3391;
wire n_6801;
wire n_1547;
wire n_1542;
wire n_5991;
wire n_1362;
wire n_6343;
wire n_4178;
wire n_4324;
wire n_7193;
wire n_3288;
wire n_2518;
wire n_6069;
wire n_3045;
wire n_3014;
wire n_5475;
wire n_6511;
wire n_1951;
wire n_1330;
wire n_5850;
wire n_6307;
wire n_7373;
wire n_5440;
wire n_1940;
wire n_3767;
wire n_1212;
wire n_1199;
wire n_4852;
wire n_1978;
wire n_1767;
wire n_1443;
wire n_5641;
wire n_1861;
wire n_1564;
wire n_7291;
wire n_2593;
wire n_1623;
wire n_6413;
wire n_6603;
wire n_1131;
wire n_6707;
wire n_3120;
wire n_1554;
wire n_4843;
wire n_7239;
wire n_6255;
wire n_4761;
wire n_6294;
wire n_2021;
wire n_6835;
wire n_7406;
wire n_2713;
wire n_2938;
wire n_3227;
wire n_3342;
wire n_5441;
wire n_2939;
wire n_6587;
wire n_6792;
wire n_4036;
wire n_1147;
wire n_5055;
wire n_4380;
wire n_2790;
wire n_2034;
wire n_3102;
wire n_4345;
wire n_6487;
wire n_1892;
wire n_5761;
wire n_6195;
wire n_2061;
wire n_6038;
wire n_1373;
wire n_7677;
wire n_3866;
wire n_3803;
wire n_2083;
wire n_2119;
wire n_5976;
wire n_7513;
wire n_2207;
wire n_4210;
wire n_7782;
wire n_3485;
wire n_4810;
wire n_3149;
wire n_5871;
wire n_2827;
wire n_5680;
wire n_3278;
wire n_2701;
wire n_6928;
wire n_2337;
wire n_4045;
wire n_4871;
wire n_2513;
wire n_1369;
wire n_1297;
wire n_1734;
wire n_4461;
wire n_2323;
wire n_7242;
wire n_6086;
wire n_5915;
wire n_5524;
wire n_7573;
wire n_5112;
wire n_3042;
wire n_5542;
wire n_5627;
wire n_2561;
wire n_5785;
wire n_2491;
wire n_6438;
wire n_5298;
wire n_7181;
wire n_1161;
wire n_1103;
wire n_6739;
wire n_4363;
wire n_5564;
wire n_5603;
wire n_3551;
wire n_3992;
wire n_4147;
wire n_6451;
wire n_4811;
wire n_6495;
wire n_5093;
wire n_5710;
wire n_3176;
wire n_2429;
wire n_3326;
wire n_5986;
wire n_3581;
wire n_3423;
wire n_1646;
wire n_4161;
wire n_5137;
wire n_1759;
wire n_2096;
wire n_5912;
wire n_2296;
wire n_7139;
wire n_6194;
wire n_1911;
wire n_7586;
wire n_6381;
wire n_7404;
wire n_2870;
wire n_6862;
wire n_4869;
wire n_6397;
wire n_4013;
wire n_1211;
wire n_4482;
wire n_3794;
wire n_6628;
wire n_5283;
wire n_1419;
wire n_7328;
wire n_6783;
wire n_4738;
wire n_7231;
wire n_6604;
wire n_1193;
wire n_2928;
wire n_3380;
wire n_3557;
wire n_7435;
wire n_2227;
wire n_2652;
wire n_3596;
wire n_7058;
wire n_5286;
wire n_2627;
wire n_1827;
wire n_3369;
wire n_5626;
wire n_4086;
wire n_5410;
wire n_4112;
wire n_2501;
wire n_2051;
wire n_1805;
wire n_3737;
wire n_1183;
wire n_7041;
wire n_3160;
wire n_4744;
wire n_1204;
wire n_1151;
wire n_3286;
wire n_1092;
wire n_6788;
wire n_2668;
wire n_6684;
wire n_1386;
wire n_2931;
wire n_7364;
wire n_2492;
wire n_5960;
wire n_3636;
wire n_4787;
wire n_4885;
wire n_2927;
wire n_4459;
wire n_7738;
wire n_1516;
wire n_4551;
wire n_4484;
wire n_5988;
wire n_1499;
wire n_5838;
wire n_2155;
wire n_3938;
wire n_6103;
wire n_7006;
wire n_6016;
wire n_3114;
wire n_3905;
wire n_6817;
wire n_1661;
wire n_6261;
wire n_7276;
wire n_1965;
wire n_5616;
wire n_1757;
wire n_7571;
wire n_7269;
wire n_6399;
wire n_4726;
wire n_3617;
wire n_3602;
wire n_4298;
wire n_6181;
wire n_3053;
wire n_5965;
wire n_3894;
wire n_6645;
wire n_2407;
wire n_6845;
wire n_2267;
wire n_2302;
wire n_2082;
wire n_2560;
wire n_2453;
wire n_6572;
wire n_4544;
wire n_7531;
wire n_7222;
wire n_4595;
wire n_4418;
wire n_2770;
wire n_7463;
wire n_2704;
wire n_6246;
wire n_1762;
wire n_7347;
wire n_4944;
wire n_7060;
wire n_4468;
wire n_5923;
wire n_6357;
wire n_6508;
wire n_6536;
wire n_3421;
wire n_7064;
wire n_4950;
wire n_3247;
wire n_1454;
wire n_4108;
wire n_6917;
wire n_7545;
wire n_4594;
wire n_6359;
wire n_5949;
wire n_7479;
wire n_1325;
wire n_2754;
wire n_4629;
wire n_4903;
wire n_3041;
wire n_7400;
wire n_4194;
wire n_3713;
wire n_2692;
wire n_5738;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_2324;
wire n_6096;
wire n_4921;
wire n_1111;
wire n_1819;
wire n_4863;
wire n_6813;
wire n_2670;
wire n_7379;
wire n_1745;
wire n_7318;
wire n_7352;
wire n_3941;
wire n_3516;
wire n_3933;
wire n_7295;
wire n_3562;
wire n_1916;
wire n_3873;
wire n_7785;
wire n_7267;
wire n_2073;
wire n_4093;
wire n_1947;
wire n_2165;
wire n_2016;
wire n_3793;
wire n_5080;
wire n_7497;
wire n_5975;
wire n_1791;
wire n_5301;
wire n_6464;
wire n_1113;
wire n_6963;
wire n_4817;
wire n_1468;
wire n_4917;
wire n_6017;
wire n_5507;
wire n_1164;
wire n_6340;
wire n_7543;
wire n_3749;
wire n_5470;
wire n_6315;
wire n_6923;
wire n_3691;
wire n_4452;
wire n_3501;
wire n_2538;
wire n_1559;
wire n_4446;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_6392;
wire n_4280;
wire n_2285;
wire n_5979;
wire n_1934;
wire n_2040;
wire n_3246;
wire n_2186;
wire n_5648;
wire n_1665;
wire n_5335;
wire n_5594;
wire n_3417;
wire n_2725;
wire n_6681;
wire n_1482;
wire n_4782;
wire n_5393;
wire n_5661;
wire n_4978;
wire n_6292;
wire n_5690;
wire n_2349;
wire n_1902;
wire n_2474;
wire n_6154;
wire n_7460;
wire n_5963;
wire n_6293;
wire n_1417;
wire n_5455;
wire n_7061;
wire n_7351;
wire n_3536;
wire n_1346;
wire n_5873;
wire n_2834;
wire n_6127;
wire n_1123;
wire n_1272;
wire n_7298;
wire n_2497;
wire n_7195;
wire n_3040;
wire n_6028;
wire n_6325;
wire n_1410;
wire n_6600;
wire n_3528;
wire n_3677;
wire n_2657;
wire n_6957;
wire n_2743;
wire n_5698;
wire n_4662;
wire n_2658;

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_1048),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_195),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_578),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_996),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_1039),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_47),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_121),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_417),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_183),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_459),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_446),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_570),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_1021),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_799),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_495),
.Y(n_1097)
);

BUFx6f_ASAP7_75t_L g1098 ( 
.A(n_48),
.Y(n_1098)
);

BUFx10_ASAP7_75t_L g1099 ( 
.A(n_646),
.Y(n_1099)
);

CKINVDCx20_ASAP7_75t_R g1100 ( 
.A(n_757),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1077),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_136),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_454),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_622),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_33),
.Y(n_1105)
);

CKINVDCx20_ASAP7_75t_R g1106 ( 
.A(n_621),
.Y(n_1106)
);

CKINVDCx5p33_ASAP7_75t_R g1107 ( 
.A(n_846),
.Y(n_1107)
);

CKINVDCx5p33_ASAP7_75t_R g1108 ( 
.A(n_344),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_1018),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_910),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_1041),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_307),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_177),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_963),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_739),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_252),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_990),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_964),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_147),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1035),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_985),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_260),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_959),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_174),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_111),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_138),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_155),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_734),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_473),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_776),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_62),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_326),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1058),
.Y(n_1133)
);

INVx2_ASAP7_75t_SL g1134 ( 
.A(n_773),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_723),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_171),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1064),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_739),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_612),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_805),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_1000),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_877),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_238),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_387),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_203),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_866),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_287),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_399),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_704),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_974),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_806),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_855),
.Y(n_1152)
);

INVxp67_ASAP7_75t_SL g1153 ( 
.A(n_489),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_686),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_510),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_987),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_90),
.Y(n_1157)
);

CKINVDCx5p33_ASAP7_75t_R g1158 ( 
.A(n_65),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1010),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_1030),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_936),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_982),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_73),
.Y(n_1163)
);

INVx1_ASAP7_75t_SL g1164 ( 
.A(n_218),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_547),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1026),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_269),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_193),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_778),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1008),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1043),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_418),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_1007),
.Y(n_1173)
);

CKINVDCx20_ASAP7_75t_R g1174 ( 
.A(n_430),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1036),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_886),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_841),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_1044),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_633),
.Y(n_1179)
);

INVxp67_ASAP7_75t_L g1180 ( 
.A(n_463),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_916),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_615),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_651),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_1061),
.Y(n_1184)
);

INVx1_ASAP7_75t_SL g1185 ( 
.A(n_1005),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_426),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_544),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_949),
.Y(n_1188)
);

CKINVDCx16_ASAP7_75t_R g1189 ( 
.A(n_447),
.Y(n_1189)
);

BUFx6f_ASAP7_75t_L g1190 ( 
.A(n_349),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_37),
.Y(n_1191)
);

BUFx5_ASAP7_75t_L g1192 ( 
.A(n_966),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_108),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_986),
.Y(n_1194)
);

INVx1_ASAP7_75t_SL g1195 ( 
.A(n_793),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_515),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_162),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_123),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_868),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_503),
.Y(n_1200)
);

BUFx3_ASAP7_75t_L g1201 ( 
.A(n_123),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_413),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_902),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1042),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_63),
.Y(n_1205)
);

CKINVDCx20_ASAP7_75t_R g1206 ( 
.A(n_1073),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_377),
.Y(n_1207)
);

BUFx8_ASAP7_75t_SL g1208 ( 
.A(n_261),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_933),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_241),
.Y(n_1210)
);

CKINVDCx5p33_ASAP7_75t_R g1211 ( 
.A(n_17),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_303),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_714),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_250),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_969),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_243),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_279),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_575),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_12),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_815),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_849),
.Y(n_1221)
);

CKINVDCx16_ASAP7_75t_R g1222 ( 
.A(n_1032),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_585),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_389),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_179),
.Y(n_1225)
);

BUFx6f_ASAP7_75t_L g1226 ( 
.A(n_630),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_751),
.Y(n_1227)
);

BUFx10_ASAP7_75t_L g1228 ( 
.A(n_154),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_421),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_45),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_345),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_495),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_791),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_95),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_228),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_313),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_674),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_637),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_505),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_884),
.Y(n_1240)
);

CKINVDCx16_ASAP7_75t_R g1241 ( 
.A(n_151),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_372),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_718),
.Y(n_1243)
);

INVx1_ASAP7_75t_SL g1244 ( 
.A(n_1001),
.Y(n_1244)
);

CKINVDCx5p33_ASAP7_75t_R g1245 ( 
.A(n_709),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_852),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_216),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_981),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_566),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_976),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_308),
.Y(n_1251)
);

CKINVDCx5p33_ASAP7_75t_R g1252 ( 
.A(n_30),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_355),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_778),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_807),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_962),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_1040),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_456),
.Y(n_1258)
);

BUFx3_ASAP7_75t_L g1259 ( 
.A(n_1049),
.Y(n_1259)
);

CKINVDCx5p33_ASAP7_75t_R g1260 ( 
.A(n_1012),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_61),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_979),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_514),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_492),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_742),
.Y(n_1265)
);

CKINVDCx5p33_ASAP7_75t_R g1266 ( 
.A(n_426),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_110),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_232),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1057),
.Y(n_1269)
);

CKINVDCx16_ASAP7_75t_R g1270 ( 
.A(n_105),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_139),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1064),
.Y(n_1272)
);

CKINVDCx5p33_ASAP7_75t_R g1273 ( 
.A(n_630),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_312),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_529),
.Y(n_1275)
);

INVx2_ASAP7_75t_SL g1276 ( 
.A(n_358),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_264),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_585),
.Y(n_1278)
);

CKINVDCx5p33_ASAP7_75t_R g1279 ( 
.A(n_531),
.Y(n_1279)
);

CKINVDCx5p33_ASAP7_75t_R g1280 ( 
.A(n_556),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_637),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_734),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_385),
.Y(n_1283)
);

INVx1_ASAP7_75t_SL g1284 ( 
.A(n_745),
.Y(n_1284)
);

CKINVDCx5p33_ASAP7_75t_R g1285 ( 
.A(n_1020),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_964),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_77),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_516),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_230),
.Y(n_1289)
);

BUFx2_ASAP7_75t_L g1290 ( 
.A(n_492),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1030),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_821),
.Y(n_1292)
);

CKINVDCx5p33_ASAP7_75t_R g1293 ( 
.A(n_995),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_519),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_353),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_184),
.Y(n_1296)
);

HB1xp67_ASAP7_75t_L g1297 ( 
.A(n_526),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_186),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_707),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_584),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_178),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1002),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_241),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_77),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_229),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_1064),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_357),
.Y(n_1307)
);

INVx1_ASAP7_75t_SL g1308 ( 
.A(n_566),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_663),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_606),
.Y(n_1310)
);

INVx4_ASAP7_75t_R g1311 ( 
.A(n_964),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_418),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_715),
.Y(n_1313)
);

CKINVDCx5p33_ASAP7_75t_R g1314 ( 
.A(n_448),
.Y(n_1314)
);

CKINVDCx5p33_ASAP7_75t_R g1315 ( 
.A(n_968),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_749),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_889),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_1038),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_957),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_898),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1034),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1033),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_332),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_456),
.Y(n_1324)
);

CKINVDCx5p33_ASAP7_75t_R g1325 ( 
.A(n_545),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_620),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_253),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_639),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_247),
.Y(n_1329)
);

CKINVDCx14_ASAP7_75t_R g1330 ( 
.A(n_435),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_298),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_999),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1035),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_980),
.Y(n_1334)
);

INVx1_ASAP7_75t_SL g1335 ( 
.A(n_711),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_333),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_648),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_224),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_78),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_626),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_128),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_953),
.Y(n_1342)
);

CKINVDCx5p33_ASAP7_75t_R g1343 ( 
.A(n_185),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_381),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1027),
.Y(n_1345)
);

CKINVDCx16_ASAP7_75t_R g1346 ( 
.A(n_906),
.Y(n_1346)
);

INVxp67_ASAP7_75t_L g1347 ( 
.A(n_455),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_71),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1062),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_349),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_373),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_1009),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_148),
.Y(n_1353)
);

INVxp67_ASAP7_75t_SL g1354 ( 
.A(n_117),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_411),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_617),
.Y(n_1356)
);

CKINVDCx5p33_ASAP7_75t_R g1357 ( 
.A(n_254),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_783),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_577),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_1012),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_983),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_823),
.Y(n_1362)
);

BUFx6f_ASAP7_75t_L g1363 ( 
.A(n_1014),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_398),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_575),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1061),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_752),
.Y(n_1367)
);

CKINVDCx5p33_ASAP7_75t_R g1368 ( 
.A(n_1024),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_443),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_956),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_998),
.Y(n_1371)
);

CKINVDCx5p33_ASAP7_75t_R g1372 ( 
.A(n_109),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_965),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_751),
.Y(n_1374)
);

CKINVDCx5p33_ASAP7_75t_R g1375 ( 
.A(n_956),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_20),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1029),
.Y(n_1377)
);

CKINVDCx14_ASAP7_75t_R g1378 ( 
.A(n_902),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_588),
.Y(n_1379)
);

BUFx5_ASAP7_75t_L g1380 ( 
.A(n_613),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_191),
.Y(n_1381)
);

HB1xp67_ASAP7_75t_L g1382 ( 
.A(n_325),
.Y(n_1382)
);

INVx1_ASAP7_75t_SL g1383 ( 
.A(n_1016),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_625),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_389),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1011),
.Y(n_1386)
);

CKINVDCx5p33_ASAP7_75t_R g1387 ( 
.A(n_749),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_250),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_65),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_514),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_130),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1031),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_967),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_203),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_229),
.Y(n_1395)
);

CKINVDCx5p33_ASAP7_75t_R g1396 ( 
.A(n_361),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_807),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1028),
.Y(n_1398)
);

INVx1_ASAP7_75t_SL g1399 ( 
.A(n_65),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1037),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_688),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_769),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_824),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_799),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_402),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_836),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_221),
.Y(n_1407)
);

BUFx2_ASAP7_75t_L g1408 ( 
.A(n_978),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_887),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_720),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_747),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_681),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_593),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_985),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_863),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_248),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_276),
.Y(n_1417)
);

CKINVDCx5p33_ASAP7_75t_R g1418 ( 
.A(n_416),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_657),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_820),
.Y(n_1420)
);

CKINVDCx5p33_ASAP7_75t_R g1421 ( 
.A(n_780),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_210),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_943),
.Y(n_1423)
);

CKINVDCx16_ASAP7_75t_R g1424 ( 
.A(n_512),
.Y(n_1424)
);

CKINVDCx20_ASAP7_75t_R g1425 ( 
.A(n_690),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_595),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_360),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_359),
.Y(n_1428)
);

BUFx3_ASAP7_75t_L g1429 ( 
.A(n_31),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_518),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_316),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_728),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_897),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_669),
.Y(n_1434)
);

CKINVDCx5p33_ASAP7_75t_R g1435 ( 
.A(n_614),
.Y(n_1435)
);

CKINVDCx5p33_ASAP7_75t_R g1436 ( 
.A(n_1003),
.Y(n_1436)
);

CKINVDCx5p33_ASAP7_75t_R g1437 ( 
.A(n_1056),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_604),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_533),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_617),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1071),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_663),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_882),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_643),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_220),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1013),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1060),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1035),
.Y(n_1448)
);

CKINVDCx20_ASAP7_75t_R g1449 ( 
.A(n_888),
.Y(n_1449)
);

CKINVDCx20_ASAP7_75t_R g1450 ( 
.A(n_289),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_357),
.Y(n_1451)
);

CKINVDCx5p33_ASAP7_75t_R g1452 ( 
.A(n_909),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_383),
.Y(n_1453)
);

CKINVDCx20_ASAP7_75t_R g1454 ( 
.A(n_975),
.Y(n_1454)
);

CKINVDCx20_ASAP7_75t_R g1455 ( 
.A(n_659),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_438),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_545),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_303),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_434),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1053),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_483),
.Y(n_1461)
);

INVx1_ASAP7_75t_SL g1462 ( 
.A(n_887),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_377),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1043),
.Y(n_1464)
);

BUFx10_ASAP7_75t_L g1465 ( 
.A(n_109),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_886),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_283),
.Y(n_1467)
);

CKINVDCx20_ASAP7_75t_R g1468 ( 
.A(n_415),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_373),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1023),
.Y(n_1470)
);

CKINVDCx5p33_ASAP7_75t_R g1471 ( 
.A(n_925),
.Y(n_1471)
);

CKINVDCx14_ASAP7_75t_R g1472 ( 
.A(n_302),
.Y(n_1472)
);

BUFx3_ASAP7_75t_L g1473 ( 
.A(n_654),
.Y(n_1473)
);

INVx1_ASAP7_75t_SL g1474 ( 
.A(n_249),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_57),
.Y(n_1475)
);

BUFx3_ASAP7_75t_L g1476 ( 
.A(n_613),
.Y(n_1476)
);

INVxp67_ASAP7_75t_SL g1477 ( 
.A(n_719),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_661),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_787),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_634),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_148),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1022),
.Y(n_1482)
);

CKINVDCx5p33_ASAP7_75t_R g1483 ( 
.A(n_246),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_85),
.Y(n_1484)
);

CKINVDCx5p33_ASAP7_75t_R g1485 ( 
.A(n_43),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_934),
.Y(n_1486)
);

CKINVDCx5p33_ASAP7_75t_R g1487 ( 
.A(n_942),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_304),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_439),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_989),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_901),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_84),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_876),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_544),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_961),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_970),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1044),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_821),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_146),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_476),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1004),
.Y(n_1501)
);

CKINVDCx5p33_ASAP7_75t_R g1502 ( 
.A(n_792),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_320),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_412),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_275),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_424),
.Y(n_1506)
);

CKINVDCx20_ASAP7_75t_R g1507 ( 
.A(n_485),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_684),
.Y(n_1508)
);

CKINVDCx5p33_ASAP7_75t_R g1509 ( 
.A(n_963),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_971),
.Y(n_1510)
);

INVx3_ASAP7_75t_L g1511 ( 
.A(n_1009),
.Y(n_1511)
);

CKINVDCx5p33_ASAP7_75t_R g1512 ( 
.A(n_993),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_358),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_836),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_772),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1025),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_54),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_756),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1006),
.Y(n_1519)
);

CKINVDCx5p33_ASAP7_75t_R g1520 ( 
.A(n_503),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_459),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_633),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_276),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_339),
.Y(n_1524)
);

CKINVDCx5p33_ASAP7_75t_R g1525 ( 
.A(n_39),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_603),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_88),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_810),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_635),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_853),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_787),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_297),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_366),
.Y(n_1533)
);

CKINVDCx20_ASAP7_75t_R g1534 ( 
.A(n_404),
.Y(n_1534)
);

BUFx5_ASAP7_75t_L g1535 ( 
.A(n_612),
.Y(n_1535)
);

BUFx3_ASAP7_75t_L g1536 ( 
.A(n_803),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_971),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1043),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_480),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_309),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_277),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_270),
.Y(n_1542)
);

BUFx6f_ASAP7_75t_L g1543 ( 
.A(n_267),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_390),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_695),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_663),
.Y(n_1546)
);

CKINVDCx20_ASAP7_75t_R g1547 ( 
.A(n_96),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_890),
.Y(n_1548)
);

INVx1_ASAP7_75t_SL g1549 ( 
.A(n_112),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_755),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_571),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_151),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_74),
.Y(n_1553)
);

CKINVDCx16_ASAP7_75t_R g1554 ( 
.A(n_947),
.Y(n_1554)
);

CKINVDCx5p33_ASAP7_75t_R g1555 ( 
.A(n_251),
.Y(n_1555)
);

INVx1_ASAP7_75t_SL g1556 ( 
.A(n_557),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_958),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_994),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_988),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_976),
.Y(n_1560)
);

CKINVDCx20_ASAP7_75t_R g1561 ( 
.A(n_253),
.Y(n_1561)
);

BUFx3_ASAP7_75t_L g1562 ( 
.A(n_389),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_991),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_73),
.Y(n_1564)
);

CKINVDCx5p33_ASAP7_75t_R g1565 ( 
.A(n_508),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_665),
.Y(n_1566)
);

INVx2_ASAP7_75t_SL g1567 ( 
.A(n_1015),
.Y(n_1567)
);

CKINVDCx5p33_ASAP7_75t_R g1568 ( 
.A(n_197),
.Y(n_1568)
);

CKINVDCx5p33_ASAP7_75t_R g1569 ( 
.A(n_834),
.Y(n_1569)
);

CKINVDCx5p33_ASAP7_75t_R g1570 ( 
.A(n_158),
.Y(n_1570)
);

CKINVDCx5p33_ASAP7_75t_R g1571 ( 
.A(n_511),
.Y(n_1571)
);

CKINVDCx20_ASAP7_75t_R g1572 ( 
.A(n_536),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_709),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_993),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_614),
.Y(n_1575)
);

CKINVDCx20_ASAP7_75t_R g1576 ( 
.A(n_873),
.Y(n_1576)
);

CKINVDCx5p33_ASAP7_75t_R g1577 ( 
.A(n_385),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_938),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_304),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1048),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_463),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_144),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_384),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_311),
.Y(n_1584)
);

CKINVDCx5p33_ASAP7_75t_R g1585 ( 
.A(n_650),
.Y(n_1585)
);

CKINVDCx5p33_ASAP7_75t_R g1586 ( 
.A(n_149),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_893),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_217),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_812),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_70),
.Y(n_1590)
);

INVx4_ASAP7_75t_R g1591 ( 
.A(n_883),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_648),
.Y(n_1592)
);

CKINVDCx20_ASAP7_75t_R g1593 ( 
.A(n_451),
.Y(n_1593)
);

CKINVDCx5p33_ASAP7_75t_R g1594 ( 
.A(n_557),
.Y(n_1594)
);

CKINVDCx5p33_ASAP7_75t_R g1595 ( 
.A(n_42),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_595),
.Y(n_1596)
);

CKINVDCx5p33_ASAP7_75t_R g1597 ( 
.A(n_784),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_643),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1046),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_302),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_977),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_917),
.Y(n_1602)
);

BUFx6f_ASAP7_75t_L g1603 ( 
.A(n_133),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_984),
.Y(n_1604)
);

CKINVDCx5p33_ASAP7_75t_R g1605 ( 
.A(n_266),
.Y(n_1605)
);

CKINVDCx20_ASAP7_75t_R g1606 ( 
.A(n_545),
.Y(n_1606)
);

CKINVDCx5p33_ASAP7_75t_R g1607 ( 
.A(n_697),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_312),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_997),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_24),
.Y(n_1610)
);

CKINVDCx5p33_ASAP7_75t_R g1611 ( 
.A(n_598),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1005),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_660),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_822),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_443),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_259),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_849),
.Y(n_1617)
);

CKINVDCx20_ASAP7_75t_R g1618 ( 
.A(n_227),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1019),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1001),
.Y(n_1620)
);

BUFx2_ASAP7_75t_L g1621 ( 
.A(n_325),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_546),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_23),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1068),
.Y(n_1624)
);

CKINVDCx5p33_ASAP7_75t_R g1625 ( 
.A(n_669),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_768),
.Y(n_1626)
);

INVx3_ASAP7_75t_L g1627 ( 
.A(n_287),
.Y(n_1627)
);

CKINVDCx5p33_ASAP7_75t_R g1628 ( 
.A(n_579),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_603),
.Y(n_1629)
);

CKINVDCx5p33_ASAP7_75t_R g1630 ( 
.A(n_911),
.Y(n_1630)
);

CKINVDCx20_ASAP7_75t_R g1631 ( 
.A(n_976),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_454),
.Y(n_1632)
);

CKINVDCx5p33_ASAP7_75t_R g1633 ( 
.A(n_447),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_320),
.Y(n_1634)
);

BUFx3_ASAP7_75t_L g1635 ( 
.A(n_944),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_868),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_917),
.Y(n_1637)
);

BUFx10_ASAP7_75t_L g1638 ( 
.A(n_297),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_967),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_166),
.Y(n_1640)
);

CKINVDCx5p33_ASAP7_75t_R g1641 ( 
.A(n_869),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_944),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_772),
.Y(n_1643)
);

CKINVDCx5p33_ASAP7_75t_R g1644 ( 
.A(n_235),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_574),
.Y(n_1645)
);

BUFx10_ASAP7_75t_L g1646 ( 
.A(n_650),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_732),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1027),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_524),
.Y(n_1649)
);

INVx1_ASAP7_75t_SL g1650 ( 
.A(n_953),
.Y(n_1650)
);

CKINVDCx5p33_ASAP7_75t_R g1651 ( 
.A(n_1046),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_345),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_307),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_533),
.Y(n_1654)
);

CKINVDCx5p33_ASAP7_75t_R g1655 ( 
.A(n_143),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_98),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_687),
.Y(n_1657)
);

CKINVDCx5p33_ASAP7_75t_R g1658 ( 
.A(n_770),
.Y(n_1658)
);

CKINVDCx5p33_ASAP7_75t_R g1659 ( 
.A(n_293),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_328),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_193),
.Y(n_1661)
);

CKINVDCx5p33_ASAP7_75t_R g1662 ( 
.A(n_411),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_340),
.Y(n_1663)
);

CKINVDCx5p33_ASAP7_75t_R g1664 ( 
.A(n_622),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_419),
.Y(n_1665)
);

CKINVDCx5p33_ASAP7_75t_R g1666 ( 
.A(n_836),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_52),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_596),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_660),
.Y(n_1669)
);

CKINVDCx5p33_ASAP7_75t_R g1670 ( 
.A(n_270),
.Y(n_1670)
);

CKINVDCx20_ASAP7_75t_R g1671 ( 
.A(n_445),
.Y(n_1671)
);

INVx1_ASAP7_75t_SL g1672 ( 
.A(n_1010),
.Y(n_1672)
);

CKINVDCx5p33_ASAP7_75t_R g1673 ( 
.A(n_21),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_311),
.Y(n_1674)
);

BUFx2_ASAP7_75t_L g1675 ( 
.A(n_747),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_234),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_119),
.Y(n_1677)
);

CKINVDCx5p33_ASAP7_75t_R g1678 ( 
.A(n_1050),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_972),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_362),
.Y(n_1680)
);

BUFx8_ASAP7_75t_SL g1681 ( 
.A(n_95),
.Y(n_1681)
);

CKINVDCx5p33_ASAP7_75t_R g1682 ( 
.A(n_17),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_164),
.Y(n_1683)
);

CKINVDCx20_ASAP7_75t_R g1684 ( 
.A(n_6),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_37),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_842),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_774),
.Y(n_1687)
);

CKINVDCx5p33_ASAP7_75t_R g1688 ( 
.A(n_182),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_683),
.Y(n_1689)
);

CKINVDCx5p33_ASAP7_75t_R g1690 ( 
.A(n_316),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_145),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_513),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_755),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_853),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_960),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_526),
.Y(n_1696)
);

CKINVDCx5p33_ASAP7_75t_R g1697 ( 
.A(n_499),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_865),
.Y(n_1698)
);

CKINVDCx20_ASAP7_75t_R g1699 ( 
.A(n_506),
.Y(n_1699)
);

INVx1_ASAP7_75t_SL g1700 ( 
.A(n_252),
.Y(n_1700)
);

INVx2_ASAP7_75t_SL g1701 ( 
.A(n_426),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_973),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_305),
.Y(n_1703)
);

CKINVDCx5p33_ASAP7_75t_R g1704 ( 
.A(n_992),
.Y(n_1704)
);

CKINVDCx5p33_ASAP7_75t_R g1705 ( 
.A(n_27),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_571),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1029),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_270),
.Y(n_1708)
);

BUFx5_ASAP7_75t_L g1709 ( 
.A(n_33),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_336),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_177),
.Y(n_1711)
);

CKINVDCx5p33_ASAP7_75t_R g1712 ( 
.A(n_785),
.Y(n_1712)
);

HB1xp67_ASAP7_75t_L g1713 ( 
.A(n_113),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_534),
.Y(n_1714)
);

BUFx5_ASAP7_75t_L g1715 ( 
.A(n_606),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_560),
.Y(n_1716)
);

CKINVDCx5p33_ASAP7_75t_R g1717 ( 
.A(n_1026),
.Y(n_1717)
);

CKINVDCx5p33_ASAP7_75t_R g1718 ( 
.A(n_83),
.Y(n_1718)
);

CKINVDCx20_ASAP7_75t_R g1719 ( 
.A(n_141),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_44),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_215),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1017),
.Y(n_1722)
);

CKINVDCx5p33_ASAP7_75t_R g1723 ( 
.A(n_1025),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_900),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_705),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_375),
.Y(n_1726)
);

INVx2_ASAP7_75t_SL g1727 ( 
.A(n_30),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1114),
.B(n_0),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1610),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1685),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1720),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1727),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1097),
.Y(n_1733)
);

INVx1_ASAP7_75t_L g1734 ( 
.A(n_1134),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1330),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1149),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1276),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1323),
.Y(n_1738)
);

CKINVDCx16_ASAP7_75t_R g1739 ( 
.A(n_1189),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1330),
.Y(n_1740)
);

CKINVDCx14_ASAP7_75t_R g1741 ( 
.A(n_1378),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1208),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1429),
.Y(n_1743)
);

CKINVDCx5p33_ASAP7_75t_R g1744 ( 
.A(n_1378),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1446),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1475),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1506),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1567),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1472),
.Y(n_1749)
);

BUFx3_ASAP7_75t_L g1750 ( 
.A(n_1709),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1701),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1116),
.Y(n_1752)
);

CKINVDCx16_ASAP7_75t_R g1753 ( 
.A(n_1222),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1472),
.Y(n_1754)
);

CKINVDCx5p33_ASAP7_75t_R g1755 ( 
.A(n_1208),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1197),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1290),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1709),
.Y(n_1758)
);

CKINVDCx20_ASAP7_75t_R g1759 ( 
.A(n_1681),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1322),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1408),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1592),
.Y(n_1762)
);

CKINVDCx5p33_ASAP7_75t_R g1763 ( 
.A(n_1681),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1621),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1709),
.Y(n_1765)
);

CKINVDCx5p33_ASAP7_75t_R g1766 ( 
.A(n_1105),
.Y(n_1766)
);

CKINVDCx5p33_ASAP7_75t_R g1767 ( 
.A(n_1211),
.Y(n_1767)
);

CKINVDCx5p33_ASAP7_75t_R g1768 ( 
.A(n_1219),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1098),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1675),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1145),
.Y(n_1771)
);

CKINVDCx14_ASAP7_75t_R g1772 ( 
.A(n_1099),
.Y(n_1772)
);

CKINVDCx5p33_ASAP7_75t_R g1773 ( 
.A(n_1252),
.Y(n_1773)
);

INVxp67_ASAP7_75t_L g1774 ( 
.A(n_1429),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1145),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1416),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1416),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1376),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1511),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1511),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1485),
.B(n_0),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1627),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1709),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1297),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1627),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1683),
.Y(n_1786)
);

BUFx6f_ASAP7_75t_L g1787 ( 
.A(n_1098),
.Y(n_1787)
);

INVx3_ASAP7_75t_L g1788 ( 
.A(n_1099),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1683),
.Y(n_1789)
);

BUFx3_ASAP7_75t_L g1790 ( 
.A(n_1709),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1382),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1684),
.Y(n_1792)
);

BUFx10_ASAP7_75t_L g1793 ( 
.A(n_1525),
.Y(n_1793)
);

CKINVDCx20_ASAP7_75t_R g1794 ( 
.A(n_1106),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1494),
.Y(n_1795)
);

CKINVDCx20_ASAP7_75t_R g1796 ( 
.A(n_1106),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1713),
.Y(n_1797)
);

BUFx6f_ASAP7_75t_L g1798 ( 
.A(n_1098),
.Y(n_1798)
);

INVxp67_ASAP7_75t_SL g1799 ( 
.A(n_1191),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1709),
.Y(n_1800)
);

CKINVDCx5p33_ASAP7_75t_R g1801 ( 
.A(n_1595),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1709),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1089),
.Y(n_1803)
);

CKINVDCx5p33_ASAP7_75t_R g1804 ( 
.A(n_1623),
.Y(n_1804)
);

CKINVDCx20_ASAP7_75t_R g1805 ( 
.A(n_1100),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1090),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1095),
.Y(n_1807)
);

INVxp67_ASAP7_75t_SL g1808 ( 
.A(n_1191),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1101),
.Y(n_1809)
);

CKINVDCx5p33_ASAP7_75t_R g1810 ( 
.A(n_1673),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1117),
.Y(n_1811)
);

CKINVDCx5p33_ASAP7_75t_R g1812 ( 
.A(n_1682),
.Y(n_1812)
);

INVxp67_ASAP7_75t_SL g1813 ( 
.A(n_1172),
.Y(n_1813)
);

BUFx3_ASAP7_75t_L g1814 ( 
.A(n_1192),
.Y(n_1814)
);

CKINVDCx16_ASAP7_75t_R g1815 ( 
.A(n_1241),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1118),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1130),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1705),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1131),
.Y(n_1819)
);

BUFx3_ASAP7_75t_L g1820 ( 
.A(n_1192),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1133),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1192),
.Y(n_1822)
);

CKINVDCx5p33_ASAP7_75t_R g1823 ( 
.A(n_1270),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1137),
.Y(n_1824)
);

CKINVDCx20_ASAP7_75t_R g1825 ( 
.A(n_1100),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1346),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1138),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1143),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1144),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1146),
.Y(n_1830)
);

CKINVDCx5p33_ASAP7_75t_R g1831 ( 
.A(n_1424),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1162),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1433),
.Y(n_1833)
);

CKINVDCx5p33_ASAP7_75t_R g1834 ( 
.A(n_1554),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1165),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1083),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1168),
.Y(n_1837)
);

INVxp67_ASAP7_75t_L g1838 ( 
.A(n_1172),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1192),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1170),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1156),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1175),
.Y(n_1842)
);

CKINVDCx5p33_ASAP7_75t_R g1843 ( 
.A(n_1085),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1176),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1179),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1187),
.Y(n_1846)
);

CKINVDCx5p33_ASAP7_75t_R g1847 ( 
.A(n_1086),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1192),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1204),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1209),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1180),
.Y(n_1851)
);

BUFx2_ASAP7_75t_L g1852 ( 
.A(n_1201),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1213),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1216),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1201),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1347),
.Y(n_1856)
);

BUFx2_ASAP7_75t_L g1857 ( 
.A(n_1224),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1217),
.Y(n_1858)
);

CKINVDCx5p33_ASAP7_75t_R g1859 ( 
.A(n_1087),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1220),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1221),
.Y(n_1861)
);

CKINVDCx5p33_ASAP7_75t_R g1862 ( 
.A(n_1088),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1091),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1225),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1772),
.Y(n_1865)
);

CKINVDCx20_ASAP7_75t_R g1866 ( 
.A(n_1792),
.Y(n_1866)
);

CKINVDCx5p33_ASAP7_75t_R g1867 ( 
.A(n_1766),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1743),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1767),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1768),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1743),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1774),
.Y(n_1872)
);

INVxp67_ASAP7_75t_SL g1873 ( 
.A(n_1774),
.Y(n_1873)
);

CKINVDCx20_ASAP7_75t_R g1874 ( 
.A(n_1794),
.Y(n_1874)
);

INVx2_ASAP7_75t_L g1875 ( 
.A(n_1814),
.Y(n_1875)
);

CKINVDCx20_ASAP7_75t_R g1876 ( 
.A(n_1796),
.Y(n_1876)
);

HB1xp67_ASAP7_75t_L g1877 ( 
.A(n_1773),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1778),
.Y(n_1878)
);

CKINVDCx16_ASAP7_75t_R g1879 ( 
.A(n_1733),
.Y(n_1879)
);

CKINVDCx5p33_ASAP7_75t_R g1880 ( 
.A(n_1801),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1852),
.Y(n_1881)
);

CKINVDCx16_ASAP7_75t_R g1882 ( 
.A(n_1739),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1857),
.Y(n_1883)
);

CKINVDCx5p33_ASAP7_75t_R g1884 ( 
.A(n_1804),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1838),
.Y(n_1885)
);

CKINVDCx5p33_ASAP7_75t_R g1886 ( 
.A(n_1810),
.Y(n_1886)
);

INVxp33_ASAP7_75t_SL g1887 ( 
.A(n_1812),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

BUFx2_ASAP7_75t_L g1889 ( 
.A(n_1818),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1793),
.Y(n_1890)
);

CKINVDCx20_ASAP7_75t_R g1891 ( 
.A(n_1805),
.Y(n_1891)
);

INVxp33_ASAP7_75t_SL g1892 ( 
.A(n_1735),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1855),
.Y(n_1893)
);

CKINVDCx5p33_ASAP7_75t_R g1894 ( 
.A(n_1793),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1755),
.Y(n_1895)
);

CKINVDCx5p33_ASAP7_75t_R g1896 ( 
.A(n_1763),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1855),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1799),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1808),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1732),
.Y(n_1900)
);

INVxp67_ASAP7_75t_SL g1901 ( 
.A(n_1784),
.Y(n_1901)
);

INVx2_ASAP7_75t_L g1902 ( 
.A(n_1820),
.Y(n_1902)
);

HB1xp67_ASAP7_75t_L g1903 ( 
.A(n_1741),
.Y(n_1903)
);

INVx3_ASAP7_75t_L g1904 ( 
.A(n_1788),
.Y(n_1904)
);

CKINVDCx5p33_ASAP7_75t_R g1905 ( 
.A(n_1753),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1813),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1734),
.Y(n_1907)
);

CKINVDCx5p33_ASAP7_75t_R g1908 ( 
.A(n_1815),
.Y(n_1908)
);

CKINVDCx20_ASAP7_75t_R g1909 ( 
.A(n_1825),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1736),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1737),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1788),
.B(n_1092),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1750),
.Y(n_1913)
);

CKINVDCx5p33_ASAP7_75t_R g1914 ( 
.A(n_1742),
.Y(n_1914)
);

CKINVDCx5p33_ASAP7_75t_R g1915 ( 
.A(n_1759),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1738),
.Y(n_1916)
);

CKINVDCx20_ASAP7_75t_R g1917 ( 
.A(n_1841),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1823),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1745),
.Y(n_1919)
);

CKINVDCx20_ASAP7_75t_R g1920 ( 
.A(n_1826),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1746),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1747),
.Y(n_1922)
);

CKINVDCx20_ASAP7_75t_R g1923 ( 
.A(n_1831),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1748),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1751),
.Y(n_1925)
);

CKINVDCx20_ASAP7_75t_R g1926 ( 
.A(n_1833),
.Y(n_1926)
);

CKINVDCx5p33_ASAP7_75t_R g1927 ( 
.A(n_1836),
.Y(n_1927)
);

CKINVDCx5p33_ASAP7_75t_R g1928 ( 
.A(n_1843),
.Y(n_1928)
);

CKINVDCx20_ASAP7_75t_R g1929 ( 
.A(n_1834),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1771),
.Y(n_1930)
);

CKINVDCx20_ASAP7_75t_R g1931 ( 
.A(n_1847),
.Y(n_1931)
);

INVxp67_ASAP7_75t_L g1932 ( 
.A(n_1851),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1775),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1776),
.Y(n_1934)
);

CKINVDCx20_ASAP7_75t_R g1935 ( 
.A(n_1859),
.Y(n_1935)
);

NOR2xp67_ASAP7_75t_L g1936 ( 
.A(n_1856),
.B(n_1224),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1777),
.Y(n_1937)
);

HB1xp67_ASAP7_75t_L g1938 ( 
.A(n_1862),
.Y(n_1938)
);

CKINVDCx20_ASAP7_75t_R g1939 ( 
.A(n_1863),
.Y(n_1939)
);

INVxp67_ASAP7_75t_SL g1940 ( 
.A(n_1781),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1779),
.Y(n_1941)
);

CKINVDCx5p33_ASAP7_75t_R g1942 ( 
.A(n_1740),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1744),
.Y(n_1943)
);

INVxp67_ASAP7_75t_SL g1944 ( 
.A(n_1781),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1780),
.Y(n_1945)
);

CKINVDCx20_ASAP7_75t_R g1946 ( 
.A(n_1749),
.Y(n_1946)
);

CKINVDCx5p33_ASAP7_75t_R g1947 ( 
.A(n_1754),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1790),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1752),
.B(n_1094),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1782),
.Y(n_1950)
);

CKINVDCx5p33_ASAP7_75t_R g1951 ( 
.A(n_1791),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1785),
.Y(n_1952)
);

CKINVDCx5p33_ASAP7_75t_R g1953 ( 
.A(n_1795),
.Y(n_1953)
);

CKINVDCx20_ASAP7_75t_R g1954 ( 
.A(n_1728),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1786),
.Y(n_1955)
);

CKINVDCx5p33_ASAP7_75t_R g1956 ( 
.A(n_1797),
.Y(n_1956)
);

CKINVDCx5p33_ASAP7_75t_R g1957 ( 
.A(n_1756),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1789),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1729),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1730),
.Y(n_1960)
);

CKINVDCx5p33_ASAP7_75t_R g1961 ( 
.A(n_1757),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1760),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1731),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1803),
.Y(n_1964)
);

CKINVDCx20_ASAP7_75t_R g1965 ( 
.A(n_1761),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1758),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1762),
.B(n_1096),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1806),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1764),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1807),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1809),
.Y(n_1971)
);

CKINVDCx5p33_ASAP7_75t_R g1972 ( 
.A(n_1770),
.Y(n_1972)
);

CKINVDCx20_ASAP7_75t_R g1973 ( 
.A(n_1811),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1816),
.Y(n_1974)
);

CKINVDCx5p33_ASAP7_75t_R g1975 ( 
.A(n_1817),
.Y(n_1975)
);

CKINVDCx16_ASAP7_75t_R g1976 ( 
.A(n_1819),
.Y(n_1976)
);

INVx2_ASAP7_75t_L g1977 ( 
.A(n_1765),
.Y(n_1977)
);

CKINVDCx20_ASAP7_75t_R g1978 ( 
.A(n_1821),
.Y(n_1978)
);

CKINVDCx20_ASAP7_75t_R g1979 ( 
.A(n_1824),
.Y(n_1979)
);

CKINVDCx16_ASAP7_75t_R g1980 ( 
.A(n_1827),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1828),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1829),
.Y(n_1982)
);

CKINVDCx5p33_ASAP7_75t_R g1983 ( 
.A(n_1830),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1832),
.Y(n_1984)
);

CKINVDCx20_ASAP7_75t_R g1985 ( 
.A(n_1835),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1837),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1840),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1842),
.Y(n_1988)
);

INVxp67_ASAP7_75t_SL g1989 ( 
.A(n_1844),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1845),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1846),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1849),
.Y(n_1992)
);

NOR2xp33_ASAP7_75t_L g1993 ( 
.A(n_1850),
.B(n_1102),
.Y(n_1993)
);

BUFx6f_ASAP7_75t_SL g1994 ( 
.A(n_1853),
.Y(n_1994)
);

CKINVDCx20_ASAP7_75t_R g1995 ( 
.A(n_1854),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1858),
.Y(n_1996)
);

INVx1_ASAP7_75t_L g1997 ( 
.A(n_1860),
.Y(n_1997)
);

NOR2xp67_ASAP7_75t_L g1998 ( 
.A(n_1861),
.B(n_1259),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1864),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1800),
.B(n_1103),
.Y(n_2000)
);

CKINVDCx20_ASAP7_75t_R g2001 ( 
.A(n_1802),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1783),
.Y(n_2002)
);

HB1xp67_ASAP7_75t_L g2003 ( 
.A(n_1822),
.Y(n_2003)
);

CKINVDCx5p33_ASAP7_75t_R g2004 ( 
.A(n_1839),
.Y(n_2004)
);

CKINVDCx5p33_ASAP7_75t_R g2005 ( 
.A(n_1848),
.Y(n_2005)
);

NOR2xp33_ASAP7_75t_R g2006 ( 
.A(n_1769),
.B(n_1104),
.Y(n_2006)
);

CKINVDCx20_ASAP7_75t_R g2007 ( 
.A(n_1798),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1798),
.B(n_1107),
.Y(n_2008)
);

INVx3_ASAP7_75t_L g2009 ( 
.A(n_1769),
.Y(n_2009)
);

INVxp33_ASAP7_75t_SL g2010 ( 
.A(n_1769),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1787),
.Y(n_2011)
);

CKINVDCx14_ASAP7_75t_R g2012 ( 
.A(n_1787),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1787),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1798),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1743),
.Y(n_2015)
);

NOR2xp67_ASAP7_75t_L g2016 ( 
.A(n_1788),
.B(n_1259),
.Y(n_2016)
);

INVxp67_ASAP7_75t_SL g2017 ( 
.A(n_1743),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1743),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1743),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1743),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1743),
.Y(n_2021)
);

CKINVDCx20_ASAP7_75t_R g2022 ( 
.A(n_1792),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1772),
.Y(n_2023)
);

NOR2xp67_ASAP7_75t_L g2024 ( 
.A(n_1788),
.B(n_1272),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1814),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1743),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1743),
.Y(n_2027)
);

CKINVDCx5p33_ASAP7_75t_R g2028 ( 
.A(n_1772),
.Y(n_2028)
);

CKINVDCx5p33_ASAP7_75t_R g2029 ( 
.A(n_1772),
.Y(n_2029)
);

CKINVDCx5p33_ASAP7_75t_R g2030 ( 
.A(n_1772),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1743),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1743),
.Y(n_2032)
);

NOR2xp67_ASAP7_75t_L g2033 ( 
.A(n_1788),
.B(n_1272),
.Y(n_2033)
);

NOR2xp33_ASAP7_75t_L g2034 ( 
.A(n_1788),
.B(n_1108),
.Y(n_2034)
);

HB1xp67_ASAP7_75t_L g2035 ( 
.A(n_1772),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1743),
.Y(n_2036)
);

INVxp67_ASAP7_75t_SL g2037 ( 
.A(n_1743),
.Y(n_2037)
);

CKINVDCx20_ASAP7_75t_R g2038 ( 
.A(n_1792),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1772),
.Y(n_2039)
);

CKINVDCx20_ASAP7_75t_R g2040 ( 
.A(n_1792),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1743),
.Y(n_2041)
);

CKINVDCx5p33_ASAP7_75t_R g2042 ( 
.A(n_1772),
.Y(n_2042)
);

CKINVDCx16_ASAP7_75t_R g2043 ( 
.A(n_1772),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1743),
.Y(n_2044)
);

CKINVDCx5p33_ASAP7_75t_R g2045 ( 
.A(n_1772),
.Y(n_2045)
);

INVxp67_ASAP7_75t_SL g2046 ( 
.A(n_1743),
.Y(n_2046)
);

INVxp67_ASAP7_75t_SL g2047 ( 
.A(n_1743),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1743),
.Y(n_2048)
);

CKINVDCx5p33_ASAP7_75t_R g2049 ( 
.A(n_1772),
.Y(n_2049)
);

CKINVDCx20_ASAP7_75t_R g2050 ( 
.A(n_1792),
.Y(n_2050)
);

CKINVDCx5p33_ASAP7_75t_R g2051 ( 
.A(n_1772),
.Y(n_2051)
);

CKINVDCx16_ASAP7_75t_R g2052 ( 
.A(n_1772),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1743),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1772),
.Y(n_2054)
);

CKINVDCx5p33_ASAP7_75t_R g2055 ( 
.A(n_1772),
.Y(n_2055)
);

CKINVDCx20_ASAP7_75t_R g2056 ( 
.A(n_1792),
.Y(n_2056)
);

CKINVDCx20_ASAP7_75t_R g2057 ( 
.A(n_1792),
.Y(n_2057)
);

CKINVDCx5p33_ASAP7_75t_R g2058 ( 
.A(n_1772),
.Y(n_2058)
);

CKINVDCx16_ASAP7_75t_R g2059 ( 
.A(n_1772),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1743),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1772),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1743),
.Y(n_2062)
);

CKINVDCx5p33_ASAP7_75t_R g2063 ( 
.A(n_1772),
.Y(n_2063)
);

CKINVDCx5p33_ASAP7_75t_R g2064 ( 
.A(n_1772),
.Y(n_2064)
);

CKINVDCx5p33_ASAP7_75t_R g2065 ( 
.A(n_1772),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_1743),
.Y(n_2066)
);

CKINVDCx16_ASAP7_75t_R g2067 ( 
.A(n_1772),
.Y(n_2067)
);

INVx2_ASAP7_75t_L g2068 ( 
.A(n_1814),
.Y(n_2068)
);

CKINVDCx5p33_ASAP7_75t_R g2069 ( 
.A(n_1772),
.Y(n_2069)
);

BUFx2_ASAP7_75t_SL g2070 ( 
.A(n_1793),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1743),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1743),
.Y(n_2072)
);

NOR2xp33_ASAP7_75t_L g2073 ( 
.A(n_1788),
.B(n_1109),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1772),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1743),
.Y(n_2075)
);

CKINVDCx20_ASAP7_75t_R g2076 ( 
.A(n_1792),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1814),
.Y(n_2077)
);

CKINVDCx20_ASAP7_75t_R g2078 ( 
.A(n_1792),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1743),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_R g2080 ( 
.A(n_1772),
.B(n_1110),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1743),
.Y(n_2081)
);

CKINVDCx5p33_ASAP7_75t_R g2082 ( 
.A(n_1772),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1743),
.Y(n_2083)
);

CKINVDCx20_ASAP7_75t_R g2084 ( 
.A(n_1792),
.Y(n_2084)
);

CKINVDCx20_ASAP7_75t_R g2085 ( 
.A(n_1792),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1743),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1743),
.Y(n_2087)
);

INVxp67_ASAP7_75t_L g2088 ( 
.A(n_1784),
.Y(n_2088)
);

CKINVDCx5p33_ASAP7_75t_R g2089 ( 
.A(n_1772),
.Y(n_2089)
);

INVxp33_ASAP7_75t_L g2090 ( 
.A(n_1784),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1743),
.Y(n_2091)
);

HB1xp67_ASAP7_75t_L g2092 ( 
.A(n_1772),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1940),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1940),
.Y(n_2094)
);

CKINVDCx5p33_ASAP7_75t_R g2095 ( 
.A(n_2080),
.Y(n_2095)
);

BUFx3_ASAP7_75t_L g2096 ( 
.A(n_2007),
.Y(n_2096)
);

CKINVDCx5p33_ASAP7_75t_R g2097 ( 
.A(n_2043),
.Y(n_2097)
);

NOR2xp67_ASAP7_75t_L g2098 ( 
.A(n_2035),
.B(n_0),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1944),
.Y(n_2099)
);

AND2x2_ASAP7_75t_L g2100 ( 
.A(n_2090),
.B(n_1901),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_1901),
.B(n_1099),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1904),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1944),
.Y(n_2103)
);

INVx1_ASAP7_75t_L g2104 ( 
.A(n_1963),
.Y(n_2104)
);

OA21x2_ASAP7_75t_L g2105 ( 
.A1(n_2000),
.A2(n_1977),
.B(n_1966),
.Y(n_2105)
);

INVx5_ASAP7_75t_L g2106 ( 
.A(n_1904),
.Y(n_2106)
);

OR2x2_ASAP7_75t_L g2107 ( 
.A(n_2088),
.B(n_1164),
.Y(n_2107)
);

HB1xp67_ASAP7_75t_L g2108 ( 
.A(n_1976),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_1930),
.Y(n_2109)
);

INVx2_ASAP7_75t_L g2110 ( 
.A(n_1933),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1963),
.Y(n_2111)
);

BUFx2_ASAP7_75t_L g2112 ( 
.A(n_1973),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_1873),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1934),
.Y(n_2114)
);

INVx2_ASAP7_75t_L g2115 ( 
.A(n_1937),
.Y(n_2115)
);

NOR2xp33_ASAP7_75t_R g2116 ( 
.A(n_1865),
.B(n_1155),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_1932),
.B(n_1228),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1873),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2017),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2017),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2037),
.B(n_1192),
.Y(n_2121)
);

INVx6_ASAP7_75t_L g2122 ( 
.A(n_2052),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2037),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_2047),
.Y(n_2124)
);

NAND2xp5_ASAP7_75t_L g2125 ( 
.A(n_2047),
.B(n_1192),
.Y(n_2125)
);

NOR2xp33_ASAP7_75t_L g2126 ( 
.A(n_1912),
.B(n_1112),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_2046),
.B(n_1380),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_1971),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1941),
.Y(n_2129)
);

AND2x4_ASAP7_75t_L g2130 ( 
.A(n_2054),
.B(n_1155),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1971),
.Y(n_2131)
);

INVx2_ASAP7_75t_L g2132 ( 
.A(n_1945),
.Y(n_2132)
);

CKINVDCx5p33_ASAP7_75t_R g2133 ( 
.A(n_2059),
.Y(n_2133)
);

CKINVDCx20_ASAP7_75t_R g2134 ( 
.A(n_1866),
.Y(n_2134)
);

CKINVDCx20_ASAP7_75t_R g2135 ( 
.A(n_2022),
.Y(n_2135)
);

CKINVDCx5p33_ASAP7_75t_R g2136 ( 
.A(n_2067),
.Y(n_2136)
);

AND2x4_ASAP7_75t_L g2137 ( 
.A(n_2092),
.B(n_1156),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1989),
.Y(n_2138)
);

INVxp67_ASAP7_75t_L g2139 ( 
.A(n_1889),
.Y(n_2139)
);

CKINVDCx20_ASAP7_75t_R g2140 ( 
.A(n_2038),
.Y(n_2140)
);

INVx1_ASAP7_75t_L g2141 ( 
.A(n_1989),
.Y(n_2141)
);

INVx2_ASAP7_75t_L g2142 ( 
.A(n_1950),
.Y(n_2142)
);

NOR2xp33_ASAP7_75t_L g2143 ( 
.A(n_1906),
.B(n_1113),
.Y(n_2143)
);

INVx2_ASAP7_75t_SL g2144 ( 
.A(n_1975),
.Y(n_2144)
);

CKINVDCx20_ASAP7_75t_R g2145 ( 
.A(n_2040),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_1900),
.Y(n_2146)
);

INVx3_ASAP7_75t_L g2147 ( 
.A(n_1994),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_1898),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2091),
.B(n_1380),
.Y(n_2149)
);

CKINVDCx20_ASAP7_75t_R g2150 ( 
.A(n_2050),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1980),
.B(n_1228),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_1952),
.Y(n_2152)
);

CKINVDCx5p33_ASAP7_75t_R g2153 ( 
.A(n_2070),
.Y(n_2153)
);

INVx2_ASAP7_75t_L g2154 ( 
.A(n_1955),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1958),
.Y(n_2155)
);

OA21x2_ASAP7_75t_L g2156 ( 
.A1(n_2002),
.A2(n_1960),
.B(n_1959),
.Y(n_2156)
);

AOI22xp5_ASAP7_75t_L g2157 ( 
.A1(n_1983),
.A2(n_1119),
.B1(n_1121),
.B2(n_1115),
.Y(n_2157)
);

CKINVDCx20_ASAP7_75t_R g2158 ( 
.A(n_2056),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1899),
.Y(n_2159)
);

CKINVDCx16_ASAP7_75t_R g2160 ( 
.A(n_1879),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2003),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_1974),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_1964),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_1994),
.Y(n_2164)
);

AND2x6_ASAP7_75t_L g2165 ( 
.A(n_1969),
.B(n_1473),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2034),
.B(n_1122),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1907),
.Y(n_2167)
);

OA21x2_ASAP7_75t_L g2168 ( 
.A1(n_1968),
.A2(n_1981),
.B(n_1970),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1982),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_1910),
.Y(n_2170)
);

AND2x2_ASAP7_75t_L g2171 ( 
.A(n_1951),
.B(n_1228),
.Y(n_2171)
);

OA21x2_ASAP7_75t_L g2172 ( 
.A1(n_1984),
.A2(n_1987),
.B(n_1986),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_1868),
.B(n_1380),
.Y(n_2173)
);

INVx2_ASAP7_75t_L g2174 ( 
.A(n_1988),
.Y(n_2174)
);

INVx3_ASAP7_75t_L g2175 ( 
.A(n_1911),
.Y(n_2175)
);

INVx2_ASAP7_75t_L g2176 ( 
.A(n_1990),
.Y(n_2176)
);

CKINVDCx5p33_ASAP7_75t_R g2177 ( 
.A(n_2057),
.Y(n_2177)
);

HB1xp67_ASAP7_75t_L g2178 ( 
.A(n_1978),
.Y(n_2178)
);

HB1xp67_ASAP7_75t_L g2179 ( 
.A(n_1979),
.Y(n_2179)
);

BUFx2_ASAP7_75t_L g2180 ( 
.A(n_1985),
.Y(n_2180)
);

INVx2_ASAP7_75t_L g2181 ( 
.A(n_1991),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1916),
.Y(n_2182)
);

CKINVDCx20_ASAP7_75t_R g2183 ( 
.A(n_2076),
.Y(n_2183)
);

CKINVDCx5p33_ASAP7_75t_R g2184 ( 
.A(n_2078),
.Y(n_2184)
);

INVx5_ASAP7_75t_L g2185 ( 
.A(n_2009),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1919),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1921),
.Y(n_2187)
);

AND2x4_ASAP7_75t_L g2188 ( 
.A(n_2023),
.B(n_1174),
.Y(n_2188)
);

CKINVDCx20_ASAP7_75t_R g2189 ( 
.A(n_2084),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1922),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_1924),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1925),
.Y(n_2192)
);

BUFx6f_ASAP7_75t_L g2193 ( 
.A(n_2028),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1998),
.Y(n_2194)
);

INVx2_ASAP7_75t_L g2195 ( 
.A(n_1992),
.Y(n_2195)
);

AND2x4_ASAP7_75t_L g2196 ( 
.A(n_2029),
.B(n_1174),
.Y(n_2196)
);

HB1xp67_ASAP7_75t_L g2197 ( 
.A(n_1995),
.Y(n_2197)
);

INVx2_ASAP7_75t_L g2198 ( 
.A(n_1996),
.Y(n_2198)
);

CKINVDCx20_ASAP7_75t_R g2199 ( 
.A(n_2085),
.Y(n_2199)
);

INVxp67_ASAP7_75t_L g2200 ( 
.A(n_1869),
.Y(n_2200)
);

INVx3_ASAP7_75t_L g2201 ( 
.A(n_1890),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_1953),
.B(n_1465),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_1894),
.Y(n_2203)
);

AND2x4_ASAP7_75t_L g2204 ( 
.A(n_2030),
.B(n_1450),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2016),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_L g2206 ( 
.A(n_1871),
.B(n_1380),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1872),
.B(n_2015),
.Y(n_2207)
);

AND2x4_ASAP7_75t_L g2208 ( 
.A(n_2039),
.B(n_1450),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2018),
.B(n_2019),
.Y(n_2209)
);

INVx2_ASAP7_75t_L g2210 ( 
.A(n_1997),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2024),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2033),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_2042),
.Y(n_2213)
);

AOI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_1956),
.A2(n_1124),
.B1(n_1125),
.B2(n_1123),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_2045),
.Y(n_2215)
);

XNOR2xp5_ASAP7_75t_L g2216 ( 
.A(n_1874),
.B(n_1454),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_2073),
.B(n_1885),
.Y(n_2217)
);

HB1xp67_ASAP7_75t_L g2218 ( 
.A(n_1954),
.Y(n_2218)
);

INVx2_ASAP7_75t_L g2219 ( 
.A(n_1999),
.Y(n_2219)
);

AND2x2_ASAP7_75t_L g2220 ( 
.A(n_1877),
.B(n_1465),
.Y(n_2220)
);

INVx6_ASAP7_75t_L g2221 ( 
.A(n_1882),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_2020),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1887),
.Y(n_2223)
);

NAND2xp33_ASAP7_75t_L g2224 ( 
.A(n_2049),
.B(n_2051),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2021),
.Y(n_2225)
);

AND2x4_ASAP7_75t_L g2226 ( 
.A(n_2055),
.B(n_2058),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_2026),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2027),
.Y(n_2228)
);

BUFx6f_ASAP7_75t_L g2229 ( 
.A(n_2089),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2031),
.Y(n_2230)
);

BUFx8_ASAP7_75t_L g2231 ( 
.A(n_1881),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2032),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_2036),
.Y(n_2233)
);

CKINVDCx16_ASAP7_75t_R g2234 ( 
.A(n_1931),
.Y(n_2234)
);

HB1xp67_ASAP7_75t_L g2235 ( 
.A(n_1867),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2041),
.Y(n_2236)
);

NAND2xp5_ASAP7_75t_L g2237 ( 
.A(n_2087),
.B(n_1380),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2044),
.Y(n_2238)
);

INVx2_ASAP7_75t_L g2239 ( 
.A(n_2048),
.Y(n_2239)
);

AND2x4_ASAP7_75t_L g2240 ( 
.A(n_2061),
.B(n_1454),
.Y(n_2240)
);

CKINVDCx11_ASAP7_75t_R g2241 ( 
.A(n_1876),
.Y(n_2241)
);

OAI22x1_ASAP7_75t_L g2242 ( 
.A1(n_1905),
.A2(n_1468),
.B1(n_1507),
.B2(n_1455),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2053),
.Y(n_2243)
);

AND2x4_ASAP7_75t_L g2244 ( 
.A(n_1936),
.B(n_1153),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2060),
.Y(n_2245)
);

NOR2xp33_ASAP7_75t_L g2246 ( 
.A(n_1888),
.B(n_1126),
.Y(n_2246)
);

CKINVDCx5p33_ASAP7_75t_R g2247 ( 
.A(n_2063),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_2064),
.B(n_1455),
.Y(n_2248)
);

INVx4_ASAP7_75t_L g2249 ( 
.A(n_2065),
.Y(n_2249)
);

BUFx6f_ASAP7_75t_L g2250 ( 
.A(n_2069),
.Y(n_2250)
);

CKINVDCx5p33_ASAP7_75t_R g2251 ( 
.A(n_2074),
.Y(n_2251)
);

OA21x2_ASAP7_75t_L g2252 ( 
.A1(n_1913),
.A2(n_1236),
.B(n_1233),
.Y(n_2252)
);

CKINVDCx5p33_ASAP7_75t_R g2253 ( 
.A(n_2082),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2062),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2086),
.B(n_1380),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1893),
.B(n_1897),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1870),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2083),
.B(n_2066),
.Y(n_2258)
);

OAI22xp5_ASAP7_75t_SL g2259 ( 
.A1(n_1891),
.A2(n_1507),
.B1(n_1522),
.B2(n_1468),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2071),
.Y(n_2260)
);

BUFx6f_ASAP7_75t_L g2261 ( 
.A(n_1878),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_L g2262 ( 
.A(n_2072),
.B(n_1380),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2081),
.B(n_1535),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2075),
.Y(n_2264)
);

BUFx6f_ASAP7_75t_L g2265 ( 
.A(n_1880),
.Y(n_2265)
);

NOR2xp33_ASAP7_75t_L g2266 ( 
.A(n_1883),
.B(n_1127),
.Y(n_2266)
);

CKINVDCx5p33_ASAP7_75t_R g2267 ( 
.A(n_1935),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2079),
.B(n_1354),
.Y(n_2268)
);

INVx6_ASAP7_75t_L g2269 ( 
.A(n_1892),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2008),
.Y(n_2270)
);

INVx4_ASAP7_75t_L g2271 ( 
.A(n_1884),
.Y(n_2271)
);

AND2x4_ASAP7_75t_L g2272 ( 
.A(n_1938),
.B(n_1477),
.Y(n_2272)
);

BUFx6f_ASAP7_75t_L g2273 ( 
.A(n_1886),
.Y(n_2273)
);

AOI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_1957),
.A2(n_1129),
.B1(n_1132),
.B2(n_1128),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2004),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1993),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_SL g2277 ( 
.A1(n_1909),
.A2(n_1528),
.B1(n_1534),
.B2(n_1522),
.Y(n_2277)
);

AND2x4_ASAP7_75t_L g2278 ( 
.A(n_1903),
.B(n_1473),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2005),
.Y(n_2279)
);

NAND2xp5_ASAP7_75t_L g2280 ( 
.A(n_1949),
.B(n_1535),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_1967),
.Y(n_2281)
);

AOI22xp5_ASAP7_75t_L g2282 ( 
.A1(n_1961),
.A2(n_1136),
.B1(n_1139),
.B2(n_1135),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_1962),
.A2(n_1141),
.B1(n_1142),
.B2(n_1140),
.Y(n_2283)
);

AND2x4_ASAP7_75t_L g2284 ( 
.A(n_2001),
.B(n_1476),
.Y(n_2284)
);

INVx4_ASAP7_75t_L g2285 ( 
.A(n_1927),
.Y(n_2285)
);

INVx2_ASAP7_75t_L g2286 ( 
.A(n_2011),
.Y(n_2286)
);

INVx3_ASAP7_75t_L g2287 ( 
.A(n_1928),
.Y(n_2287)
);

HB1xp67_ASAP7_75t_L g2288 ( 
.A(n_1908),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1942),
.Y(n_2289)
);

INVx2_ASAP7_75t_L g2290 ( 
.A(n_2009),
.Y(n_2290)
);

BUFx6f_ASAP7_75t_L g2291 ( 
.A(n_1943),
.Y(n_2291)
);

INVx2_ASAP7_75t_L g2292 ( 
.A(n_2013),
.Y(n_2292)
);

INVx5_ASAP7_75t_L g2293 ( 
.A(n_1875),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_SL g2294 ( 
.A1(n_1917),
.A2(n_1534),
.B1(n_1538),
.B2(n_1528),
.Y(n_2294)
);

INVx1_ASAP7_75t_L g2295 ( 
.A(n_1972),
.Y(n_2295)
);

INVx1_ASAP7_75t_L g2296 ( 
.A(n_2006),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_L g2297 ( 
.A(n_1948),
.B(n_1535),
.Y(n_2297)
);

AND2x2_ASAP7_75t_L g2298 ( 
.A(n_1947),
.B(n_1465),
.Y(n_2298)
);

INVx2_ASAP7_75t_SL g2299 ( 
.A(n_1939),
.Y(n_2299)
);

AOI22xp5_ASAP7_75t_L g2300 ( 
.A1(n_1965),
.A2(n_1148),
.B1(n_1151),
.B2(n_1147),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_1902),
.B(n_1523),
.Y(n_2301)
);

INVxp67_ASAP7_75t_L g2302 ( 
.A(n_1895),
.Y(n_2302)
);

BUFx3_ASAP7_75t_L g2303 ( 
.A(n_1896),
.Y(n_2303)
);

AND2x4_ASAP7_75t_L g2304 ( 
.A(n_1946),
.B(n_1476),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2012),
.Y(n_2305)
);

CKINVDCx5p33_ASAP7_75t_R g2306 ( 
.A(n_1914),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_2014),
.Y(n_2307)
);

NAND2xp5_ASAP7_75t_SL g2308 ( 
.A(n_2025),
.B(n_1523),
.Y(n_2308)
);

BUFx3_ASAP7_75t_L g2309 ( 
.A(n_1918),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_2010),
.Y(n_2310)
);

NAND2x1p5_ASAP7_75t_L g2311 ( 
.A(n_1920),
.B(n_1482),
.Y(n_2311)
);

CKINVDCx5p33_ASAP7_75t_R g2312 ( 
.A(n_1915),
.Y(n_2312)
);

INVx2_ASAP7_75t_L g2313 ( 
.A(n_2068),
.Y(n_2313)
);

NAND2xp5_ASAP7_75t_L g2314 ( 
.A(n_2077),
.B(n_1535),
.Y(n_2314)
);

HB1xp67_ASAP7_75t_L g2315 ( 
.A(n_1923),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1926),
.B(n_1152),
.Y(n_2316)
);

AND2x2_ASAP7_75t_L g2317 ( 
.A(n_1929),
.B(n_1523),
.Y(n_2317)
);

AND2x6_ASAP7_75t_L g2318 ( 
.A(n_1906),
.B(n_1482),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_1940),
.Y(n_2319)
);

INVx2_ASAP7_75t_L g2320 ( 
.A(n_1904),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1940),
.Y(n_2321)
);

INVx2_ASAP7_75t_L g2322 ( 
.A(n_1904),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_1901),
.Y(n_2323)
);

INVx2_ASAP7_75t_L g2324 ( 
.A(n_1904),
.Y(n_2324)
);

BUFx6f_ASAP7_75t_L g2325 ( 
.A(n_1865),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1940),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_2007),
.Y(n_2327)
);

BUFx6f_ASAP7_75t_L g2328 ( 
.A(n_1865),
.Y(n_2328)
);

NAND2xp5_ASAP7_75t_SL g2329 ( 
.A(n_1975),
.B(n_1638),
.Y(n_2329)
);

INVx1_ASAP7_75t_L g2330 ( 
.A(n_1940),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1940),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1940),
.Y(n_2332)
);

NAND2xp5_ASAP7_75t_L g2333 ( 
.A(n_1940),
.B(n_1535),
.Y(n_2333)
);

OA21x2_ASAP7_75t_L g2334 ( 
.A1(n_2000),
.A2(n_1243),
.B(n_1239),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1940),
.Y(n_2335)
);

BUFx2_ASAP7_75t_L g2336 ( 
.A(n_1940),
.Y(n_2336)
);

AND2x2_ASAP7_75t_L g2337 ( 
.A(n_2090),
.B(n_1638),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2090),
.B(n_1638),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_1904),
.Y(n_2339)
);

NAND2xp5_ASAP7_75t_L g2340 ( 
.A(n_1940),
.B(n_1535),
.Y(n_2340)
);

INVx3_ASAP7_75t_L g2341 ( 
.A(n_1904),
.Y(n_2341)
);

BUFx12f_ASAP7_75t_L g2342 ( 
.A(n_1905),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2080),
.Y(n_2343)
);

CKINVDCx16_ASAP7_75t_R g2344 ( 
.A(n_2043),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_1940),
.B(n_1536),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_1940),
.B(n_1535),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_1940),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2348)
);

INVx3_ASAP7_75t_L g2349 ( 
.A(n_1904),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_1904),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1940),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_1940),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2353)
);

AND2x4_ASAP7_75t_L g2354 ( 
.A(n_2035),
.B(n_1538),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_1904),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_1940),
.Y(n_2356)
);

NAND2xp5_ASAP7_75t_L g2357 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_1940),
.Y(n_2358)
);

AND2x2_ASAP7_75t_SL g2359 ( 
.A(n_2043),
.B(n_1311),
.Y(n_2359)
);

INVx1_ASAP7_75t_L g2360 ( 
.A(n_1940),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1940),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_1940),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_2035),
.B(n_1547),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_1904),
.Y(n_2364)
);

AND2x6_ASAP7_75t_L g2365 ( 
.A(n_1906),
.B(n_1536),
.Y(n_2365)
);

AOI22xp5_ASAP7_75t_L g2366 ( 
.A1(n_1940),
.A2(n_1157),
.B1(n_1158),
.B2(n_1154),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1940),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_1904),
.Y(n_2369)
);

BUFx6f_ASAP7_75t_L g2370 ( 
.A(n_1865),
.Y(n_2370)
);

CKINVDCx16_ASAP7_75t_R g2371 ( 
.A(n_2043),
.Y(n_2371)
);

NOR2xp33_ASAP7_75t_R g2372 ( 
.A(n_1865),
.B(n_1547),
.Y(n_2372)
);

AOI22x1_ASAP7_75t_SL g2373 ( 
.A1(n_1866),
.A2(n_1561),
.B1(n_1572),
.B2(n_1560),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_1940),
.Y(n_2374)
);

BUFx8_ASAP7_75t_L g2375 ( 
.A(n_1994),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_1940),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_1904),
.Y(n_2377)
);

AND2x4_ASAP7_75t_L g2378 ( 
.A(n_2035),
.B(n_1560),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1865),
.Y(n_2379)
);

CKINVDCx5p33_ASAP7_75t_R g2380 ( 
.A(n_2080),
.Y(n_2380)
);

AND2x2_ASAP7_75t_L g2381 ( 
.A(n_2090),
.B(n_1646),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_1865),
.Y(n_2382)
);

HB1xp67_ASAP7_75t_L g2383 ( 
.A(n_1976),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_SL g2385 ( 
.A(n_1887),
.B(n_1561),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_1940),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_1940),
.Y(n_2387)
);

BUFx6f_ASAP7_75t_L g2388 ( 
.A(n_1865),
.Y(n_2388)
);

OAI22xp5_ASAP7_75t_SL g2389 ( 
.A1(n_1866),
.A2(n_1576),
.B1(n_1578),
.B2(n_1572),
.Y(n_2389)
);

AND2x2_ASAP7_75t_L g2390 ( 
.A(n_2090),
.B(n_1646),
.Y(n_2390)
);

INVx2_ASAP7_75t_L g2391 ( 
.A(n_1904),
.Y(n_2391)
);

AOI22xp5_ASAP7_75t_L g2392 ( 
.A1(n_1940),
.A2(n_1160),
.B1(n_1161),
.B2(n_1159),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_SL g2393 ( 
.A(n_1975),
.B(n_1646),
.Y(n_2393)
);

AOI22xp5_ASAP7_75t_L g2394 ( 
.A1(n_1940),
.A2(n_1166),
.B1(n_1167),
.B2(n_1163),
.Y(n_2394)
);

BUFx3_ASAP7_75t_L g2395 ( 
.A(n_2007),
.Y(n_2395)
);

NOR2xp67_ASAP7_75t_L g2396 ( 
.A(n_2035),
.B(n_0),
.Y(n_2396)
);

AND2x2_ASAP7_75t_SL g2397 ( 
.A(n_2043),
.B(n_1591),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_1904),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_L g2399 ( 
.A(n_1940),
.B(n_1715),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_R g2400 ( 
.A(n_1865),
.B(n_1576),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2090),
.B(n_1169),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1940),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2336),
.Y(n_2403)
);

BUFx6f_ASAP7_75t_L g2404 ( 
.A(n_2336),
.Y(n_2404)
);

INVx2_ASAP7_75t_L g2405 ( 
.A(n_2156),
.Y(n_2405)
);

BUFx2_ASAP7_75t_L g2406 ( 
.A(n_2108),
.Y(n_2406)
);

OR2x2_ASAP7_75t_L g2407 ( 
.A(n_2107),
.B(n_1185),
.Y(n_2407)
);

INVx2_ASAP7_75t_L g2408 ( 
.A(n_2156),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2093),
.Y(n_2409)
);

NAND2xp5_ASAP7_75t_L g2410 ( 
.A(n_2345),
.B(n_1171),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2094),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2099),
.Y(n_2412)
);

CKINVDCx16_ASAP7_75t_R g2413 ( 
.A(n_2385),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_L g2414 ( 
.A(n_2345),
.B(n_1173),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2103),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2319),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2321),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2326),
.Y(n_2418)
);

BUFx4f_ASAP7_75t_L g2419 ( 
.A(n_2122),
.Y(n_2419)
);

NOR2xp33_ASAP7_75t_L g2420 ( 
.A(n_2100),
.B(n_1206),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2330),
.Y(n_2421)
);

AND2x2_ASAP7_75t_L g2422 ( 
.A(n_2401),
.B(n_1578),
.Y(n_2422)
);

AOI22xp5_ASAP7_75t_L g2423 ( 
.A1(n_2323),
.A2(n_1593),
.B1(n_1606),
.B2(n_1587),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2331),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2332),
.Y(n_2425)
);

INVx2_ASAP7_75t_L g2426 ( 
.A(n_2335),
.Y(n_2426)
);

INVxp33_ASAP7_75t_SL g2427 ( 
.A(n_2223),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2347),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_L g2429 ( 
.A(n_2351),
.B(n_1177),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2352),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2356),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2358),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_SL g2433 ( 
.A(n_2360),
.B(n_1178),
.Y(n_2433)
);

CKINVDCx5p33_ASAP7_75t_R g2434 ( 
.A(n_2241),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2361),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2362),
.Y(n_2436)
);

OAI22xp33_ASAP7_75t_L g2437 ( 
.A1(n_2383),
.A2(n_1593),
.B1(n_1606),
.B2(n_1587),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_2368),
.B(n_2374),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2376),
.Y(n_2439)
);

INVx2_ASAP7_75t_L g2440 ( 
.A(n_2386),
.Y(n_2440)
);

INVx2_ASAP7_75t_L g2441 ( 
.A(n_2387),
.Y(n_2441)
);

INVx2_ASAP7_75t_L g2442 ( 
.A(n_2402),
.Y(n_2442)
);

INVx2_ASAP7_75t_L g2443 ( 
.A(n_2163),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_SL g2444 ( 
.A(n_2101),
.B(n_2144),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2168),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2169),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2168),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2174),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2176),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2172),
.Y(n_2450)
);

INVx2_ASAP7_75t_SL g2451 ( 
.A(n_2151),
.Y(n_2451)
);

AND2x2_ASAP7_75t_L g2452 ( 
.A(n_2337),
.B(n_1618),
.Y(n_2452)
);

CKINVDCx5p33_ASAP7_75t_R g2453 ( 
.A(n_2342),
.Y(n_2453)
);

INVx8_ASAP7_75t_L g2454 ( 
.A(n_2165),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2218),
.B(n_1195),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2181),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_2106),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2172),
.Y(n_2458)
);

NOR2xp33_ASAP7_75t_L g2459 ( 
.A(n_2117),
.B(n_1242),
.Y(n_2459)
);

NAND3xp33_ASAP7_75t_L g2460 ( 
.A(n_2316),
.B(n_1182),
.C(n_1181),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2195),
.Y(n_2461)
);

CKINVDCx5p33_ASAP7_75t_R g2462 ( 
.A(n_2116),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2198),
.Y(n_2463)
);

INVx2_ASAP7_75t_L g2464 ( 
.A(n_2210),
.Y(n_2464)
);

INVx8_ASAP7_75t_L g2465 ( 
.A(n_2165),
.Y(n_2465)
);

INVx3_ASAP7_75t_L g2466 ( 
.A(n_2106),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2148),
.Y(n_2467)
);

INVx1_ASAP7_75t_L g2468 ( 
.A(n_2159),
.Y(n_2468)
);

INVx2_ASAP7_75t_L g2469 ( 
.A(n_2219),
.Y(n_2469)
);

AND2x2_ASAP7_75t_L g2470 ( 
.A(n_2338),
.B(n_1618),
.Y(n_2470)
);

NOR2xp33_ASAP7_75t_L g2471 ( 
.A(n_2200),
.B(n_1294),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2102),
.Y(n_2472)
);

INVxp33_ASAP7_75t_SL g2473 ( 
.A(n_2216),
.Y(n_2473)
);

AND2x2_ASAP7_75t_L g2474 ( 
.A(n_2381),
.B(n_1620),
.Y(n_2474)
);

INVx2_ASAP7_75t_L g2475 ( 
.A(n_2320),
.Y(n_2475)
);

BUFx6f_ASAP7_75t_L g2476 ( 
.A(n_2252),
.Y(n_2476)
);

CKINVDCx5p33_ASAP7_75t_R g2477 ( 
.A(n_2372),
.Y(n_2477)
);

NOR2x1_ASAP7_75t_L g2478 ( 
.A(n_2271),
.B(n_1620),
.Y(n_2478)
);

AND2x2_ASAP7_75t_L g2479 ( 
.A(n_2390),
.B(n_1631),
.Y(n_2479)
);

INVx1_ASAP7_75t_L g2480 ( 
.A(n_2161),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_SL g2481 ( 
.A(n_2171),
.B(n_1183),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2322),
.Y(n_2482)
);

BUFx6f_ASAP7_75t_L g2483 ( 
.A(n_2252),
.Y(n_2483)
);

CKINVDCx6p67_ASAP7_75t_R g2484 ( 
.A(n_2309),
.Y(n_2484)
);

AO21x2_ASAP7_75t_L g2485 ( 
.A1(n_2280),
.A2(n_1249),
.B(n_1247),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2139),
.B(n_1631),
.Y(n_2486)
);

INVx2_ASAP7_75t_L g2487 ( 
.A(n_2324),
.Y(n_2487)
);

NAND2xp5_ASAP7_75t_L g2488 ( 
.A(n_2104),
.B(n_1184),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2111),
.B(n_1186),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2339),
.Y(n_2490)
);

INVx4_ASAP7_75t_L g2491 ( 
.A(n_2153),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2128),
.B(n_1188),
.Y(n_2492)
);

NOR2xp33_ASAP7_75t_L g2493 ( 
.A(n_2202),
.B(n_2220),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_2350),
.Y(n_2494)
);

INVx2_ASAP7_75t_L g2495 ( 
.A(n_2355),
.Y(n_2495)
);

INVx2_ASAP7_75t_L g2496 ( 
.A(n_2364),
.Y(n_2496)
);

NAND2xp5_ASAP7_75t_SL g2497 ( 
.A(n_2281),
.B(n_1193),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2131),
.B(n_1194),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2369),
.Y(n_2499)
);

INVx2_ASAP7_75t_L g2500 ( 
.A(n_2377),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2391),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2284),
.B(n_1671),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2333),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2398),
.Y(n_2504)
);

INVx2_ASAP7_75t_L g2505 ( 
.A(n_2313),
.Y(n_2505)
);

INVx2_ASAP7_75t_SL g2506 ( 
.A(n_2221),
.Y(n_2506)
);

NOR2xp33_ASAP7_75t_L g2507 ( 
.A(n_2295),
.B(n_1321),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2340),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2175),
.Y(n_2509)
);

INVx3_ASAP7_75t_L g2510 ( 
.A(n_2106),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2138),
.B(n_1196),
.Y(n_2511)
);

INVx2_ASAP7_75t_L g2512 ( 
.A(n_2105),
.Y(n_2512)
);

INVx2_ASAP7_75t_L g2513 ( 
.A(n_2105),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2346),
.Y(n_2514)
);

NAND2xp5_ASAP7_75t_SL g2515 ( 
.A(n_2284),
.B(n_1198),
.Y(n_2515)
);

AOI21x1_ASAP7_75t_L g2516 ( 
.A1(n_2297),
.A2(n_1251),
.B(n_1250),
.Y(n_2516)
);

INVx2_ASAP7_75t_L g2517 ( 
.A(n_2109),
.Y(n_2517)
);

INVx2_ASAP7_75t_L g2518 ( 
.A(n_2110),
.Y(n_2518)
);

BUFx3_ASAP7_75t_L g2519 ( 
.A(n_2122),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2348),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2353),
.Y(n_2521)
);

INVx2_ASAP7_75t_L g2522 ( 
.A(n_2114),
.Y(n_2522)
);

INVxp67_ASAP7_75t_SL g2523 ( 
.A(n_2096),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_SL g2524 ( 
.A(n_2366),
.B(n_1199),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2272),
.B(n_1671),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2115),
.Y(n_2526)
);

NOR2x1p5_ASAP7_75t_L g2527 ( 
.A(n_2285),
.B(n_1200),
.Y(n_2527)
);

INVxp33_ASAP7_75t_SL g2528 ( 
.A(n_2216),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2357),
.Y(n_2529)
);

INVx2_ASAP7_75t_L g2530 ( 
.A(n_2129),
.Y(n_2530)
);

INVx2_ASAP7_75t_SL g2531 ( 
.A(n_2221),
.Y(n_2531)
);

INVx2_ASAP7_75t_L g2532 ( 
.A(n_2132),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2142),
.Y(n_2533)
);

INVx1_ASAP7_75t_SL g2534 ( 
.A(n_2112),
.Y(n_2534)
);

AO21x2_ASAP7_75t_L g2535 ( 
.A1(n_2314),
.A2(n_1264),
.B(n_1263),
.Y(n_2535)
);

INVx1_ASAP7_75t_SL g2536 ( 
.A(n_2112),
.Y(n_2536)
);

INVx2_ASAP7_75t_L g2537 ( 
.A(n_2152),
.Y(n_2537)
);

NOR2xp33_ASAP7_75t_L g2538 ( 
.A(n_2298),
.B(n_1367),
.Y(n_2538)
);

INVx2_ASAP7_75t_L g2539 ( 
.A(n_2154),
.Y(n_2539)
);

NOR3xp33_ASAP7_75t_L g2540 ( 
.A(n_2389),
.B(n_1284),
.C(n_1244),
.Y(n_2540)
);

NAND2xp33_ASAP7_75t_L g2541 ( 
.A(n_2318),
.B(n_1715),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2392),
.B(n_1202),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_SL g2543 ( 
.A(n_2394),
.B(n_1203),
.Y(n_2543)
);

NAND2xp5_ASAP7_75t_L g2544 ( 
.A(n_2141),
.B(n_1205),
.Y(n_2544)
);

INVx1_ASAP7_75t_SL g2545 ( 
.A(n_2180),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2155),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2146),
.Y(n_2547)
);

HB1xp67_ASAP7_75t_L g2548 ( 
.A(n_2162),
.Y(n_2548)
);

BUFx2_ASAP7_75t_L g2549 ( 
.A(n_2400),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2367),
.Y(n_2550)
);

NAND2xp5_ASAP7_75t_SL g2551 ( 
.A(n_2276),
.B(n_1210),
.Y(n_2551)
);

NOR2xp33_ASAP7_75t_L g2552 ( 
.A(n_2275),
.B(n_1373),
.Y(n_2552)
);

INVx2_ASAP7_75t_L g2553 ( 
.A(n_2167),
.Y(n_2553)
);

INVx2_ASAP7_75t_SL g2554 ( 
.A(n_2327),
.Y(n_2554)
);

INVx2_ASAP7_75t_SL g2555 ( 
.A(n_2395),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2384),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2334),
.Y(n_2557)
);

INVx2_ASAP7_75t_L g2558 ( 
.A(n_2170),
.Y(n_2558)
);

INVxp33_ASAP7_75t_L g2559 ( 
.A(n_2178),
.Y(n_2559)
);

OR2x6_ASAP7_75t_L g2560 ( 
.A(n_2269),
.B(n_1562),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_L g2561 ( 
.A(n_2113),
.B(n_1212),
.Y(n_2561)
);

INVx2_ASAP7_75t_SL g2562 ( 
.A(n_2165),
.Y(n_2562)
);

INVx2_ASAP7_75t_L g2563 ( 
.A(n_2182),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2399),
.Y(n_2564)
);

INVx8_ASAP7_75t_L g2565 ( 
.A(n_2318),
.Y(n_2565)
);

INVx2_ASAP7_75t_L g2566 ( 
.A(n_2186),
.Y(n_2566)
);

INVx3_ASAP7_75t_L g2567 ( 
.A(n_2293),
.Y(n_2567)
);

AND2x2_ASAP7_75t_L g2568 ( 
.A(n_2272),
.B(n_1391),
.Y(n_2568)
);

INVx8_ASAP7_75t_L g2569 ( 
.A(n_2318),
.Y(n_2569)
);

NAND3xp33_ASAP7_75t_L g2570 ( 
.A(n_2266),
.B(n_1215),
.C(n_1214),
.Y(n_2570)
);

INVx2_ASAP7_75t_SL g2571 ( 
.A(n_2269),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2187),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2190),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2191),
.Y(n_2574)
);

INVx4_ASAP7_75t_L g2575 ( 
.A(n_2257),
.Y(n_2575)
);

INVx2_ASAP7_75t_L g2576 ( 
.A(n_2192),
.Y(n_2576)
);

INVx2_ASAP7_75t_L g2577 ( 
.A(n_2334),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2341),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_SL g2579 ( 
.A(n_2279),
.B(n_1218),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2375),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_SL g2581 ( 
.A(n_2157),
.B(n_1229),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2149),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2349),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2173),
.Y(n_2584)
);

INVx8_ASAP7_75t_L g2585 ( 
.A(n_2365),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_SL g2586 ( 
.A(n_2214),
.B(n_1230),
.Y(n_2586)
);

NAND2xp5_ASAP7_75t_L g2587 ( 
.A(n_2118),
.B(n_2119),
.Y(n_2587)
);

BUFx6f_ASAP7_75t_L g2588 ( 
.A(n_2365),
.Y(n_2588)
);

INVx2_ASAP7_75t_L g2589 ( 
.A(n_2227),
.Y(n_2589)
);

CKINVDCx20_ASAP7_75t_R g2590 ( 
.A(n_2234),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2206),
.Y(n_2591)
);

NAND3xp33_ASAP7_75t_L g2592 ( 
.A(n_2166),
.B(n_1232),
.C(n_1231),
.Y(n_2592)
);

AND2x2_ASAP7_75t_L g2593 ( 
.A(n_2317),
.B(n_1398),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2233),
.Y(n_2594)
);

NOR2xp33_ASAP7_75t_L g2595 ( 
.A(n_2329),
.B(n_1400),
.Y(n_2595)
);

INVx2_ASAP7_75t_L g2596 ( 
.A(n_2239),
.Y(n_2596)
);

INVx2_ASAP7_75t_L g2597 ( 
.A(n_2243),
.Y(n_2597)
);

INVx3_ASAP7_75t_L g2598 ( 
.A(n_2293),
.Y(n_2598)
);

NOR2xp33_ASAP7_75t_L g2599 ( 
.A(n_2393),
.B(n_1425),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2120),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2237),
.Y(n_2601)
);

INVx2_ASAP7_75t_L g2602 ( 
.A(n_2123),
.Y(n_2602)
);

INVx2_ASAP7_75t_L g2603 ( 
.A(n_2124),
.Y(n_2603)
);

INVx2_ASAP7_75t_L g2604 ( 
.A(n_2222),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2225),
.Y(n_2605)
);

BUFx10_ASAP7_75t_L g2606 ( 
.A(n_2226),
.Y(n_2606)
);

INVx1_ASAP7_75t_L g2607 ( 
.A(n_2255),
.Y(n_2607)
);

INVx4_ASAP7_75t_L g2608 ( 
.A(n_2257),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2228),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2230),
.Y(n_2610)
);

BUFx3_ASAP7_75t_L g2611 ( 
.A(n_2193),
.Y(n_2611)
);

BUFx3_ASAP7_75t_L g2612 ( 
.A(n_2193),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_L g2613 ( 
.A(n_2126),
.B(n_1234),
.Y(n_2613)
);

AND2x2_ASAP7_75t_L g2614 ( 
.A(n_2300),
.B(n_1449),
.Y(n_2614)
);

NAND2xp5_ASAP7_75t_SL g2615 ( 
.A(n_2274),
.B(n_1235),
.Y(n_2615)
);

NOR2xp33_ASAP7_75t_L g2616 ( 
.A(n_2268),
.B(n_1699),
.Y(n_2616)
);

INVx3_ASAP7_75t_L g2617 ( 
.A(n_2293),
.Y(n_2617)
);

INVx2_ASAP7_75t_L g2618 ( 
.A(n_2232),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2262),
.Y(n_2619)
);

NAND2xp33_ASAP7_75t_L g2620 ( 
.A(n_2365),
.B(n_1237),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2263),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2236),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_SL g2623 ( 
.A(n_2282),
.B(n_1238),
.Y(n_2623)
);

INVx3_ASAP7_75t_L g2624 ( 
.A(n_2238),
.Y(n_2624)
);

INVxp33_ASAP7_75t_L g2625 ( 
.A(n_2179),
.Y(n_2625)
);

OAI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2235),
.A2(n_1719),
.B1(n_1706),
.B2(n_1245),
.Y(n_2626)
);

INVx5_ASAP7_75t_L g2627 ( 
.A(n_2147),
.Y(n_2627)
);

INVx2_ASAP7_75t_L g2628 ( 
.A(n_2245),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2283),
.B(n_1240),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2254),
.Y(n_2630)
);

NOR2xp33_ASAP7_75t_SL g2631 ( 
.A(n_2302),
.B(n_1248),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_L g2632 ( 
.A(n_2217),
.B(n_1253),
.Y(n_2632)
);

BUFx4f_ASAP7_75t_L g2633 ( 
.A(n_2229),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2121),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2311),
.B(n_1254),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2125),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2127),
.Y(n_2637)
);

INVx2_ASAP7_75t_L g2638 ( 
.A(n_2260),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2264),
.Y(n_2639)
);

INVx3_ASAP7_75t_L g2640 ( 
.A(n_2286),
.Y(n_2640)
);

INVx2_ASAP7_75t_L g2641 ( 
.A(n_2194),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2207),
.Y(n_2642)
);

INVx1_ASAP7_75t_L g2643 ( 
.A(n_2209),
.Y(n_2643)
);

INVx3_ASAP7_75t_L g2644 ( 
.A(n_2205),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2258),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2211),
.Y(n_2646)
);

INVx2_ASAP7_75t_SL g2647 ( 
.A(n_2278),
.Y(n_2647)
);

AND3x2_ASAP7_75t_L g2648 ( 
.A(n_2180),
.B(n_1286),
.C(n_1269),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2212),
.Y(n_2649)
);

BUFx10_ASAP7_75t_L g2650 ( 
.A(n_2261),
.Y(n_2650)
);

NAND2xp5_ASAP7_75t_SL g2651 ( 
.A(n_2278),
.B(n_1255),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2256),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2270),
.Y(n_2653)
);

BUFx6f_ASAP7_75t_L g2654 ( 
.A(n_2185),
.Y(n_2654)
);

INVx2_ASAP7_75t_L g2655 ( 
.A(n_2292),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2307),
.Y(n_2656)
);

BUFx10_ASAP7_75t_L g2657 ( 
.A(n_2261),
.Y(n_2657)
);

OR2x6_ASAP7_75t_L g2658 ( 
.A(n_2265),
.B(n_1562),
.Y(n_2658)
);

INVx8_ASAP7_75t_L g2659 ( 
.A(n_2265),
.Y(n_2659)
);

NAND2xp5_ASAP7_75t_SL g2660 ( 
.A(n_2098),
.B(n_1256),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2268),
.Y(n_2661)
);

AND2x6_ASAP7_75t_L g2662 ( 
.A(n_2164),
.B(n_1635),
.Y(n_2662)
);

NOR2xp33_ASAP7_75t_L g2663 ( 
.A(n_2305),
.B(n_1257),
.Y(n_2663)
);

INVx2_ASAP7_75t_L g2664 ( 
.A(n_2290),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2143),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2244),
.Y(n_2666)
);

INVx2_ASAP7_75t_L g2667 ( 
.A(n_2244),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2185),
.Y(n_2668)
);

INVx5_ASAP7_75t_L g2669 ( 
.A(n_2273),
.Y(n_2669)
);

NAND2xp5_ASAP7_75t_L g2670 ( 
.A(n_2246),
.B(n_1258),
.Y(n_2670)
);

CKINVDCx11_ASAP7_75t_R g2671 ( 
.A(n_2134),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2301),
.Y(n_2672)
);

INVx2_ASAP7_75t_L g2673 ( 
.A(n_2185),
.Y(n_2673)
);

INVx2_ASAP7_75t_L g2674 ( 
.A(n_2308),
.Y(n_2674)
);

CKINVDCx6p67_ASAP7_75t_R g2675 ( 
.A(n_2344),
.Y(n_2675)
);

INVx2_ASAP7_75t_L g2676 ( 
.A(n_2310),
.Y(n_2676)
);

INVx2_ASAP7_75t_SL g2677 ( 
.A(n_2304),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2203),
.B(n_1260),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2296),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2304),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2359),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2397),
.Y(n_2682)
);

NAND2xp5_ASAP7_75t_L g2683 ( 
.A(n_2396),
.B(n_1261),
.Y(n_2683)
);

INVx3_ASAP7_75t_L g2684 ( 
.A(n_2249),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2287),
.B(n_1262),
.Y(n_2685)
);

INVx2_ASAP7_75t_L g2686 ( 
.A(n_2201),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2197),
.Y(n_2687)
);

INVx2_ASAP7_75t_L g2688 ( 
.A(n_2213),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2215),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_SL g2690 ( 
.A(n_2273),
.B(n_2289),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2130),
.Y(n_2691)
);

INVx2_ASAP7_75t_L g2692 ( 
.A(n_2289),
.Y(n_2692)
);

CKINVDCx5p33_ASAP7_75t_R g2693 ( 
.A(n_2267),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_SL g2694 ( 
.A(n_2291),
.B(n_1265),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2137),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2354),
.B(n_1266),
.Y(n_2696)
);

CKINVDCx6p67_ASAP7_75t_R g2697 ( 
.A(n_2371),
.Y(n_2697)
);

HB1xp67_ASAP7_75t_L g2698 ( 
.A(n_2259),
.Y(n_2698)
);

INVx2_ASAP7_75t_L g2699 ( 
.A(n_2291),
.Y(n_2699)
);

INVx2_ASAP7_75t_L g2700 ( 
.A(n_2231),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2229),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2363),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2378),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2242),
.Y(n_2704)
);

OR2x2_ASAP7_75t_L g2705 ( 
.A(n_2277),
.B(n_1308),
.Y(n_2705)
);

BUFx8_ASAP7_75t_SL g2706 ( 
.A(n_2135),
.Y(n_2706)
);

INVx2_ASAP7_75t_L g2707 ( 
.A(n_2250),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2250),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2325),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_SL g2710 ( 
.A(n_2095),
.B(n_1267),
.Y(n_2710)
);

INVx2_ASAP7_75t_L g2711 ( 
.A(n_2325),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2328),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_SL g2713 ( 
.A(n_2343),
.B(n_1268),
.Y(n_2713)
);

INVx2_ASAP7_75t_L g2714 ( 
.A(n_2328),
.Y(n_2714)
);

INVx1_ASAP7_75t_L g2715 ( 
.A(n_2303),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2370),
.Y(n_2716)
);

INVx2_ASAP7_75t_L g2717 ( 
.A(n_2370),
.Y(n_2717)
);

INVx2_ASAP7_75t_L g2718 ( 
.A(n_2379),
.Y(n_2718)
);

BUFx3_ASAP7_75t_L g2719 ( 
.A(n_2379),
.Y(n_2719)
);

INVx2_ASAP7_75t_L g2720 ( 
.A(n_2382),
.Y(n_2720)
);

HB1xp67_ASAP7_75t_L g2721 ( 
.A(n_2294),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2288),
.Y(n_2722)
);

NAND2xp5_ASAP7_75t_SL g2723 ( 
.A(n_2380),
.B(n_1271),
.Y(n_2723)
);

INVx1_ASAP7_75t_L g2724 ( 
.A(n_2382),
.Y(n_2724)
);

INVx3_ASAP7_75t_L g2725 ( 
.A(n_2388),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2388),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2188),
.Y(n_2727)
);

CKINVDCx5p33_ASAP7_75t_R g2728 ( 
.A(n_2160),
.Y(n_2728)
);

CKINVDCx5p33_ASAP7_75t_R g2729 ( 
.A(n_2140),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2196),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2204),
.Y(n_2731)
);

BUFx3_ASAP7_75t_L g2732 ( 
.A(n_2097),
.Y(n_2732)
);

INVx2_ASAP7_75t_L g2733 ( 
.A(n_2208),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2240),
.B(n_1273),
.Y(n_2734)
);

CKINVDCx6p67_ASAP7_75t_R g2735 ( 
.A(n_2145),
.Y(n_2735)
);

INVx2_ASAP7_75t_L g2736 ( 
.A(n_2248),
.Y(n_2736)
);

NAND2xp5_ASAP7_75t_L g2737 ( 
.A(n_2247),
.B(n_1274),
.Y(n_2737)
);

INVx3_ASAP7_75t_L g2738 ( 
.A(n_2251),
.Y(n_2738)
);

INVx2_ASAP7_75t_L g2739 ( 
.A(n_2133),
.Y(n_2739)
);

INVx1_ASAP7_75t_L g2740 ( 
.A(n_2315),
.Y(n_2740)
);

AND2x2_ASAP7_75t_L g2741 ( 
.A(n_2299),
.B(n_1275),
.Y(n_2741)
);

CKINVDCx5p33_ASAP7_75t_R g2742 ( 
.A(n_2150),
.Y(n_2742)
);

AO22x2_ASAP7_75t_L g2743 ( 
.A1(n_2373),
.A2(n_1383),
.B1(n_1394),
.B2(n_1335),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2224),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2136),
.Y(n_2745)
);

NAND3xp33_ASAP7_75t_L g2746 ( 
.A(n_2253),
.B(n_1280),
.C(n_1279),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2306),
.Y(n_2747)
);

INVx2_ASAP7_75t_L g2748 ( 
.A(n_2312),
.Y(n_2748)
);

INVx1_ASAP7_75t_L g2749 ( 
.A(n_2177),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2184),
.Y(n_2750)
);

INVx5_ASAP7_75t_L g2751 ( 
.A(n_2158),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_SL g2752 ( 
.A(n_2183),
.B(n_1281),
.Y(n_2752)
);

HB1xp67_ASAP7_75t_L g2753 ( 
.A(n_2189),
.Y(n_2753)
);

INVxp33_ASAP7_75t_L g2754 ( 
.A(n_2199),
.Y(n_2754)
);

NAND2xp33_ASAP7_75t_SL g2755 ( 
.A(n_2336),
.B(n_1282),
.Y(n_2755)
);

AOI21x1_ASAP7_75t_L g2756 ( 
.A1(n_2297),
.A2(n_1291),
.B(n_1287),
.Y(n_2756)
);

INVx2_ASAP7_75t_L g2757 ( 
.A(n_2336),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2336),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2336),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2336),
.Y(n_2760)
);

NAND3xp33_ASAP7_75t_L g2761 ( 
.A(n_2316),
.B(n_1285),
.C(n_1283),
.Y(n_2761)
);

INVx3_ASAP7_75t_L g2762 ( 
.A(n_2345),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2336),
.Y(n_2763)
);

INVx1_ASAP7_75t_SL g2764 ( 
.A(n_2107),
.Y(n_2764)
);

NAND3xp33_ASAP7_75t_L g2765 ( 
.A(n_2316),
.B(n_1289),
.C(n_1288),
.Y(n_2765)
);

INVx2_ASAP7_75t_SL g2766 ( 
.A(n_2108),
.Y(n_2766)
);

INVx2_ASAP7_75t_L g2767 ( 
.A(n_2336),
.Y(n_2767)
);

CKINVDCx5p33_ASAP7_75t_R g2768 ( 
.A(n_2241),
.Y(n_2768)
);

CKINVDCx5p33_ASAP7_75t_R g2769 ( 
.A(n_2241),
.Y(n_2769)
);

INVx11_ASAP7_75t_L g2770 ( 
.A(n_2375),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2336),
.B(n_1292),
.Y(n_2771)
);

INVx2_ASAP7_75t_L g2772 ( 
.A(n_2336),
.Y(n_2772)
);

INVx2_ASAP7_75t_L g2773 ( 
.A(n_2336),
.Y(n_2773)
);

OR2x2_ASAP7_75t_L g2774 ( 
.A(n_2107),
.B(n_1399),
.Y(n_2774)
);

BUFx3_ASAP7_75t_L g2775 ( 
.A(n_2122),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2336),
.Y(n_2776)
);

BUFx2_ASAP7_75t_L g2777 ( 
.A(n_2108),
.Y(n_2777)
);

NAND2xp5_ASAP7_75t_SL g2778 ( 
.A(n_2336),
.B(n_1293),
.Y(n_2778)
);

INVx2_ASAP7_75t_L g2779 ( 
.A(n_2336),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2336),
.B(n_1296),
.Y(n_2780)
);

INVx1_ASAP7_75t_L g2781 ( 
.A(n_2336),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2336),
.Y(n_2782)
);

INVx2_ASAP7_75t_L g2783 ( 
.A(n_2336),
.Y(n_2783)
);

INVx2_ASAP7_75t_SL g2784 ( 
.A(n_2108),
.Y(n_2784)
);

INVx2_ASAP7_75t_L g2785 ( 
.A(n_2336),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2336),
.B(n_1298),
.Y(n_2786)
);

INVx2_ASAP7_75t_SL g2787 ( 
.A(n_2108),
.Y(n_2787)
);

INVx2_ASAP7_75t_L g2788 ( 
.A(n_2336),
.Y(n_2788)
);

NOR2xp33_ASAP7_75t_L g2789 ( 
.A(n_2100),
.B(n_1300),
.Y(n_2789)
);

BUFx6f_ASAP7_75t_SL g2790 ( 
.A(n_2309),
.Y(n_2790)
);

INVx1_ASAP7_75t_L g2791 ( 
.A(n_2336),
.Y(n_2791)
);

AND3x2_ASAP7_75t_L g2792 ( 
.A(n_2385),
.B(n_1299),
.C(n_1295),
.Y(n_2792)
);

CKINVDCx5p33_ASAP7_75t_R g2793 ( 
.A(n_2241),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2336),
.B(n_1301),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2336),
.Y(n_2795)
);

NAND2xp5_ASAP7_75t_SL g2796 ( 
.A(n_2336),
.B(n_1302),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2336),
.Y(n_2797)
);

NAND3x1_ASAP7_75t_L g2798 ( 
.A(n_2540),
.B(n_1313),
.C(n_1304),
.Y(n_2798)
);

CKINVDCx5p33_ASAP7_75t_R g2799 ( 
.A(n_2706),
.Y(n_2799)
);

INVx3_ASAP7_75t_L g2800 ( 
.A(n_2404),
.Y(n_2800)
);

NOR2xp33_ASAP7_75t_L g2801 ( 
.A(n_2459),
.B(n_1303),
.Y(n_2801)
);

INVx1_ASAP7_75t_L g2802 ( 
.A(n_2573),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2631),
.B(n_1305),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2764),
.B(n_1462),
.Y(n_2804)
);

NAND2xp5_ASAP7_75t_L g2805 ( 
.A(n_2642),
.B(n_1306),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2405),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2573),
.Y(n_2807)
);

CKINVDCx5p33_ASAP7_75t_R g2808 ( 
.A(n_2671),
.Y(n_2808)
);

INVx2_ASAP7_75t_L g2809 ( 
.A(n_2408),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2574),
.Y(n_2810)
);

BUFx6f_ASAP7_75t_L g2811 ( 
.A(n_2404),
.Y(n_2811)
);

BUFx6f_ASAP7_75t_L g2812 ( 
.A(n_2404),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2642),
.B(n_1307),
.Y(n_2813)
);

INVx4_ASAP7_75t_L g2814 ( 
.A(n_2659),
.Y(n_2814)
);

INVx4_ASAP7_75t_L g2815 ( 
.A(n_2659),
.Y(n_2815)
);

INVx3_ASAP7_75t_L g2816 ( 
.A(n_2654),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2574),
.Y(n_2817)
);

INVx4_ASAP7_75t_SL g2818 ( 
.A(n_2580),
.Y(n_2818)
);

BUFx3_ASAP7_75t_L g2819 ( 
.A(n_2669),
.Y(n_2819)
);

INVx2_ASAP7_75t_L g2820 ( 
.A(n_2557),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2409),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2409),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2407),
.B(n_2774),
.Y(n_2823)
);

INVx2_ASAP7_75t_L g2824 ( 
.A(n_2557),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2411),
.Y(n_2825)
);

CKINVDCx5p33_ASAP7_75t_R g2826 ( 
.A(n_2770),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2411),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_L g2828 ( 
.A(n_2643),
.B(n_1310),
.Y(n_2828)
);

INVx5_ASAP7_75t_L g2829 ( 
.A(n_2560),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2412),
.Y(n_2830)
);

INVx1_ASAP7_75t_L g2831 ( 
.A(n_2412),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2415),
.Y(n_2832)
);

NAND3xp33_ASAP7_75t_L g2833 ( 
.A(n_2678),
.B(n_1314),
.C(n_1312),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2476),
.Y(n_2834)
);

BUFx3_ASAP7_75t_L g2835 ( 
.A(n_2669),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_SL g2836 ( 
.A(n_2755),
.B(n_2413),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2415),
.Y(n_2837)
);

OR2x2_ASAP7_75t_SL g2838 ( 
.A(n_2698),
.B(n_1316),
.Y(n_2838)
);

INVx1_ASAP7_75t_L g2839 ( 
.A(n_2416),
.Y(n_2839)
);

NAND2xp5_ASAP7_75t_SL g2840 ( 
.A(n_2643),
.B(n_1315),
.Y(n_2840)
);

OAI22xp5_ASAP7_75t_SL g2841 ( 
.A1(n_2473),
.A2(n_1319),
.B1(n_1320),
.B2(n_1317),
.Y(n_2841)
);

NOR2x1p5_ASAP7_75t_L g2842 ( 
.A(n_2735),
.B(n_1325),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2654),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2416),
.Y(n_2844)
);

BUFx2_ASAP7_75t_L g2845 ( 
.A(n_2560),
.Y(n_2845)
);

BUFx2_ASAP7_75t_L g2846 ( 
.A(n_2406),
.Y(n_2846)
);

INVx2_ASAP7_75t_L g2847 ( 
.A(n_2557),
.Y(n_2847)
);

INVx4_ASAP7_75t_L g2848 ( 
.A(n_2669),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2480),
.Y(n_2849)
);

AND2x2_ASAP7_75t_SL g2850 ( 
.A(n_2620),
.B(n_1084),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2639),
.Y(n_2851)
);

AOI22xp5_ASAP7_75t_L g2852 ( 
.A1(n_2471),
.A2(n_1336),
.B1(n_1337),
.B2(n_1328),
.Y(n_2852)
);

AND2x2_ASAP7_75t_L g2853 ( 
.A(n_2645),
.B(n_1339),
.Y(n_2853)
);

INVx1_ASAP7_75t_SL g2854 ( 
.A(n_2777),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2417),
.Y(n_2855)
);

INVxp67_ASAP7_75t_SL g2856 ( 
.A(n_2437),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2639),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2418),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2421),
.Y(n_2859)
);

INVx1_ASAP7_75t_SL g2860 ( 
.A(n_2658),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2645),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2467),
.Y(n_2862)
);

INVx1_ASAP7_75t_L g2863 ( 
.A(n_2468),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2547),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_SL g2865 ( 
.A(n_2766),
.B(n_1340),
.Y(n_2865)
);

BUFx6f_ASAP7_75t_L g2866 ( 
.A(n_2476),
.Y(n_2866)
);

BUFx10_ASAP7_75t_L g2867 ( 
.A(n_2658),
.Y(n_2867)
);

INVxp67_ASAP7_75t_SL g2868 ( 
.A(n_2476),
.Y(n_2868)
);

AND2x2_ASAP7_75t_L g2869 ( 
.A(n_2422),
.B(n_2525),
.Y(n_2869)
);

AND2x6_ASAP7_75t_L g2870 ( 
.A(n_2588),
.B(n_1635),
.Y(n_2870)
);

AND2x6_ASAP7_75t_L g2871 ( 
.A(n_2588),
.B(n_1692),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2553),
.Y(n_2872)
);

INVx2_ASAP7_75t_L g2873 ( 
.A(n_2424),
.Y(n_2873)
);

NAND2xp5_ASAP7_75t_L g2874 ( 
.A(n_2403),
.B(n_2760),
.Y(n_2874)
);

BUFx2_ASAP7_75t_L g2875 ( 
.A(n_2784),
.Y(n_2875)
);

INVx1_ASAP7_75t_SL g2876 ( 
.A(n_2534),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2434),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2650),
.Y(n_2878)
);

INVx1_ASAP7_75t_L g2879 ( 
.A(n_2558),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2403),
.B(n_1342),
.Y(n_2880)
);

AND2x6_ASAP7_75t_L g2881 ( 
.A(n_2588),
.B(n_1692),
.Y(n_2881)
);

CKINVDCx5p33_ASAP7_75t_R g2882 ( 
.A(n_2768),
.Y(n_2882)
);

NOR2xp33_ASAP7_75t_L g2883 ( 
.A(n_2538),
.B(n_1343),
.Y(n_2883)
);

INVx1_ASAP7_75t_L g2884 ( 
.A(n_2563),
.Y(n_2884)
);

AND2x2_ASAP7_75t_SL g2885 ( 
.A(n_2633),
.B(n_1084),
.Y(n_2885)
);

NOR2xp33_ASAP7_75t_L g2886 ( 
.A(n_2451),
.B(n_1344),
.Y(n_2886)
);

INVx6_ASAP7_75t_L g2887 ( 
.A(n_2650),
.Y(n_2887)
);

BUFx4f_ASAP7_75t_L g2888 ( 
.A(n_2675),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2657),
.Y(n_2889)
);

NAND2xp5_ASAP7_75t_SL g2890 ( 
.A(n_2787),
.B(n_1348),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2566),
.Y(n_2891)
);

NAND2x1p5_ASAP7_75t_L g2892 ( 
.A(n_2633),
.B(n_1474),
.Y(n_2892)
);

AOI22xp5_ASAP7_75t_L g2893 ( 
.A1(n_2626),
.A2(n_1352),
.B1(n_1353),
.B2(n_1349),
.Y(n_2893)
);

AND2x4_ASAP7_75t_L g2894 ( 
.A(n_2744),
.B(n_1324),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2572),
.Y(n_2895)
);

AND2x4_ASAP7_75t_L g2896 ( 
.A(n_2653),
.B(n_1326),
.Y(n_2896)
);

AND2x2_ASAP7_75t_L g2897 ( 
.A(n_2486),
.B(n_1355),
.Y(n_2897)
);

HB1xp67_ASAP7_75t_L g2898 ( 
.A(n_2536),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2576),
.Y(n_2899)
);

AND2x2_ASAP7_75t_L g2900 ( 
.A(n_2452),
.B(n_1356),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2425),
.Y(n_2901)
);

INVxp33_ASAP7_75t_L g2902 ( 
.A(n_2753),
.Y(n_2902)
);

INVx1_ASAP7_75t_L g2903 ( 
.A(n_2604),
.Y(n_2903)
);

INVx4_ASAP7_75t_L g2904 ( 
.A(n_2565),
.Y(n_2904)
);

BUFx3_ASAP7_75t_L g2905 ( 
.A(n_2657),
.Y(n_2905)
);

INVx6_ASAP7_75t_L g2906 ( 
.A(n_2575),
.Y(n_2906)
);

INVx2_ASAP7_75t_L g2907 ( 
.A(n_2426),
.Y(n_2907)
);

CKINVDCx5p33_ASAP7_75t_R g2908 ( 
.A(n_2769),
.Y(n_2908)
);

AOI22xp33_ASAP7_75t_L g2909 ( 
.A1(n_2420),
.A2(n_1358),
.B1(n_1359),
.B2(n_1357),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2605),
.Y(n_2910)
);

INVx2_ASAP7_75t_L g2911 ( 
.A(n_2430),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_SL g2912 ( 
.A(n_2685),
.B(n_1360),
.Y(n_2912)
);

INVx2_ASAP7_75t_L g2913 ( 
.A(n_2432),
.Y(n_2913)
);

AND2x4_ASAP7_75t_L g2914 ( 
.A(n_2760),
.B(n_1327),
.Y(n_2914)
);

AND2x4_ASAP7_75t_L g2915 ( 
.A(n_2776),
.B(n_1329),
.Y(n_2915)
);

NAND2xp5_ASAP7_75t_SL g2916 ( 
.A(n_2757),
.B(n_1364),
.Y(n_2916)
);

AND2x6_ASAP7_75t_L g2917 ( 
.A(n_2577),
.B(n_1098),
.Y(n_2917)
);

OR2x2_ASAP7_75t_L g2918 ( 
.A(n_2423),
.B(n_1532),
.Y(n_2918)
);

NAND2xp5_ASAP7_75t_L g2919 ( 
.A(n_2776),
.B(n_1365),
.Y(n_2919)
);

INVx2_ASAP7_75t_L g2920 ( 
.A(n_2439),
.Y(n_2920)
);

BUFx3_ASAP7_75t_L g2921 ( 
.A(n_2519),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2781),
.B(n_1366),
.Y(n_2922)
);

INVxp67_ASAP7_75t_SL g2923 ( 
.A(n_2483),
.Y(n_2923)
);

INVx2_ASAP7_75t_L g2924 ( 
.A(n_2440),
.Y(n_2924)
);

NAND2x1p5_ASAP7_75t_L g2925 ( 
.A(n_2575),
.B(n_1549),
.Y(n_2925)
);

NOR2xp33_ASAP7_75t_L g2926 ( 
.A(n_2493),
.B(n_1368),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2781),
.B(n_2791),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2470),
.B(n_1370),
.Y(n_2928)
);

INVxp33_ASAP7_75t_L g2929 ( 
.A(n_2455),
.Y(n_2929)
);

AND2x4_ASAP7_75t_L g2930 ( 
.A(n_2791),
.B(n_1333),
.Y(n_2930)
);

BUFx6f_ASAP7_75t_L g2931 ( 
.A(n_2483),
.Y(n_2931)
);

NOR3xp33_ASAP7_75t_L g2932 ( 
.A(n_2460),
.B(n_1632),
.C(n_1556),
.Y(n_2932)
);

BUFx6f_ASAP7_75t_SL g2933 ( 
.A(n_2732),
.Y(n_2933)
);

BUFx6f_ASAP7_75t_L g2934 ( 
.A(n_2483),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2428),
.Y(n_2935)
);

NAND2xp5_ASAP7_75t_L g2936 ( 
.A(n_2797),
.B(n_2652),
.Y(n_2936)
);

INVx2_ASAP7_75t_L g2937 ( 
.A(n_2441),
.Y(n_2937)
);

AO22x2_ASAP7_75t_L g2938 ( 
.A1(n_2512),
.A2(n_1672),
.B1(n_1700),
.B2(n_1650),
.Y(n_2938)
);

INVx1_ASAP7_75t_L g2939 ( 
.A(n_2428),
.Y(n_2939)
);

AND2x2_ASAP7_75t_L g2940 ( 
.A(n_2474),
.B(n_2479),
.Y(n_2940)
);

NOR2xp33_ASAP7_75t_L g2941 ( 
.A(n_2593),
.B(n_2559),
.Y(n_2941)
);

CKINVDCx5p33_ASAP7_75t_R g2942 ( 
.A(n_2793),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2431),
.Y(n_2943)
);

AND2x2_ASAP7_75t_L g2944 ( 
.A(n_2614),
.B(n_1372),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_L g2945 ( 
.A(n_2625),
.B(n_1374),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2609),
.Y(n_2946)
);

BUFx6f_ASAP7_75t_L g2947 ( 
.A(n_2654),
.Y(n_2947)
);

INVxp67_ASAP7_75t_L g2948 ( 
.A(n_2548),
.Y(n_2948)
);

AOI22xp33_ASAP7_75t_L g2949 ( 
.A1(n_2721),
.A2(n_1381),
.B1(n_1386),
.B2(n_1375),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2610),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2797),
.B(n_1387),
.Y(n_2951)
);

AND2x6_ASAP7_75t_L g2952 ( 
.A(n_2503),
.B(n_1111),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2618),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2568),
.B(n_1388),
.Y(n_2954)
);

BUFx6f_ASAP7_75t_L g2955 ( 
.A(n_2513),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2652),
.B(n_1389),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2622),
.Y(n_2957)
);

NOR2xp33_ASAP7_75t_L g2958 ( 
.A(n_2616),
.B(n_1390),
.Y(n_2958)
);

AND2x6_ASAP7_75t_L g2959 ( 
.A(n_2503),
.B(n_1111),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2628),
.Y(n_2960)
);

INVx1_ASAP7_75t_L g2961 ( 
.A(n_2630),
.Y(n_2961)
);

INVx3_ASAP7_75t_L g2962 ( 
.A(n_2457),
.Y(n_2962)
);

BUFx6f_ASAP7_75t_L g2963 ( 
.A(n_2565),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2442),
.Y(n_2964)
);

BUFx6f_ASAP7_75t_L g2965 ( 
.A(n_2569),
.Y(n_2965)
);

AND2x4_ASAP7_75t_L g2966 ( 
.A(n_2638),
.B(n_1334),
.Y(n_2966)
);

NOR2xp33_ASAP7_75t_L g2967 ( 
.A(n_2545),
.B(n_1392),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_SL g2968 ( 
.A(n_2758),
.B(n_1393),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2431),
.Y(n_2969)
);

BUFx2_ASAP7_75t_L g2970 ( 
.A(n_2729),
.Y(n_2970)
);

CKINVDCx5p33_ASAP7_75t_R g2971 ( 
.A(n_2697),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2759),
.B(n_1396),
.Y(n_2972)
);

INVx1_ASAP7_75t_L g2973 ( 
.A(n_2435),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2624),
.Y(n_2974)
);

AND2x4_ASAP7_75t_L g2975 ( 
.A(n_2684),
.B(n_1341),
.Y(n_2975)
);

INVx2_ASAP7_75t_L g2976 ( 
.A(n_2624),
.Y(n_2976)
);

BUFx6f_ASAP7_75t_L g2977 ( 
.A(n_2569),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2435),
.Y(n_2978)
);

INVx1_ASAP7_75t_L g2979 ( 
.A(n_2436),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2763),
.B(n_2767),
.Y(n_2980)
);

AND2x2_ASAP7_75t_SL g2981 ( 
.A(n_2549),
.B(n_1093),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2436),
.Y(n_2982)
);

NAND2x1p5_ASAP7_75t_L g2983 ( 
.A(n_2608),
.B(n_1111),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2600),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2602),
.Y(n_2985)
);

BUFx2_ASAP7_75t_L g2986 ( 
.A(n_2742),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2603),
.Y(n_2987)
);

AND2x4_ASAP7_75t_L g2988 ( 
.A(n_2684),
.B(n_2491),
.Y(n_2988)
);

BUFx6f_ASAP7_75t_L g2989 ( 
.A(n_2585),
.Y(n_2989)
);

BUFx3_ASAP7_75t_L g2990 ( 
.A(n_2775),
.Y(n_2990)
);

BUFx6f_ASAP7_75t_L g2991 ( 
.A(n_2585),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_2453),
.Y(n_2992)
);

AND2x6_ASAP7_75t_L g2993 ( 
.A(n_2508),
.B(n_2514),
.Y(n_2993)
);

INVx5_ASAP7_75t_L g2994 ( 
.A(n_2608),
.Y(n_2994)
);

NOR2xp33_ASAP7_75t_L g2995 ( 
.A(n_2507),
.B(n_1397),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2454),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2589),
.Y(n_2997)
);

INVx3_ASAP7_75t_L g2998 ( 
.A(n_2457),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2594),
.Y(n_2999)
);

NAND2xp33_ASAP7_75t_L g3000 ( 
.A(n_2662),
.B(n_1401),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2438),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2596),
.Y(n_3002)
);

BUFx6f_ASAP7_75t_L g3003 ( 
.A(n_2454),
.Y(n_3003)
);

AND2x6_ASAP7_75t_L g3004 ( 
.A(n_2508),
.B(n_2514),
.Y(n_3004)
);

INVx2_ASAP7_75t_SL g3005 ( 
.A(n_2419),
.Y(n_3005)
);

INVx4_ASAP7_75t_L g3006 ( 
.A(n_2465),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2772),
.B(n_1402),
.Y(n_3007)
);

BUFx10_ASAP7_75t_L g3008 ( 
.A(n_2790),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_L g3009 ( 
.A(n_2465),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2587),
.Y(n_3010)
);

CKINVDCx5p33_ASAP7_75t_R g3011 ( 
.A(n_2427),
.Y(n_3011)
);

INVx2_ASAP7_75t_SL g3012 ( 
.A(n_2419),
.Y(n_3012)
);

CKINVDCx5p33_ASAP7_75t_R g3013 ( 
.A(n_2728),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2773),
.B(n_2779),
.Y(n_3014)
);

INVx2_ASAP7_75t_SL g3015 ( 
.A(n_2751),
.Y(n_3015)
);

NOR2xp33_ASAP7_75t_L g3016 ( 
.A(n_2552),
.B(n_1404),
.Y(n_3016)
);

HB1xp67_ASAP7_75t_L g3017 ( 
.A(n_2611),
.Y(n_3017)
);

OR2x6_ASAP7_75t_L g3018 ( 
.A(n_2700),
.B(n_1093),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_SL g3019 ( 
.A(n_2782),
.B(n_1405),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2520),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2520),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2783),
.B(n_1410),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_SL g3023 ( 
.A(n_2785),
.B(n_1414),
.Y(n_3023)
);

NOR2xp33_ASAP7_75t_L g3024 ( 
.A(n_2444),
.B(n_1415),
.Y(n_3024)
);

INVx3_ASAP7_75t_L g3025 ( 
.A(n_2466),
.Y(n_3025)
);

INVx5_ASAP7_75t_L g3026 ( 
.A(n_2662),
.Y(n_3026)
);

AND2x2_ASAP7_75t_L g3027 ( 
.A(n_2502),
.B(n_1417),
.Y(n_3027)
);

NOR2xp33_ASAP7_75t_L g3028 ( 
.A(n_2703),
.B(n_1418),
.Y(n_3028)
);

BUFx3_ASAP7_75t_L g3029 ( 
.A(n_2612),
.Y(n_3029)
);

NOR2xp33_ASAP7_75t_L g3030 ( 
.A(n_2515),
.B(n_1419),
.Y(n_3030)
);

INVx1_ASAP7_75t_SL g3031 ( 
.A(n_2635),
.Y(n_3031)
);

CKINVDCx5p33_ASAP7_75t_R g3032 ( 
.A(n_2590),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2788),
.B(n_1420),
.Y(n_3033)
);

INVxp67_ASAP7_75t_L g3034 ( 
.A(n_2741),
.Y(n_3034)
);

AOI22xp33_ASAP7_75t_L g3035 ( 
.A1(n_2687),
.A2(n_1423),
.B1(n_1426),
.B2(n_1421),
.Y(n_3035)
);

INVx3_ASAP7_75t_L g3036 ( 
.A(n_2466),
.Y(n_3036)
);

INVx2_ASAP7_75t_SL g3037 ( 
.A(n_2751),
.Y(n_3037)
);

INVx4_ASAP7_75t_L g3038 ( 
.A(n_2792),
.Y(n_3038)
);

NAND2xp5_ASAP7_75t_L g3039 ( 
.A(n_2795),
.B(n_1430),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2665),
.B(n_1431),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_L g3041 ( 
.A(n_2677),
.B(n_1432),
.Y(n_3041)
);

CKINVDCx11_ASAP7_75t_R g3042 ( 
.A(n_2484),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2521),
.Y(n_3043)
);

INVx5_ASAP7_75t_L g3044 ( 
.A(n_2662),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2521),
.Y(n_3045)
);

NOR2xp33_ASAP7_75t_L g3046 ( 
.A(n_2727),
.B(n_1434),
.Y(n_3046)
);

INVx5_ASAP7_75t_L g3047 ( 
.A(n_2662),
.Y(n_3047)
);

NAND2xp5_ASAP7_75t_SL g3048 ( 
.A(n_2491),
.B(n_1435),
.Y(n_3048)
);

BUFx4f_ASAP7_75t_L g3049 ( 
.A(n_2738),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2529),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2597),
.Y(n_3051)
);

AND3x2_ASAP7_75t_L g3052 ( 
.A(n_2595),
.B(n_1350),
.C(n_1345),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2771),
.B(n_1436),
.Y(n_3053)
);

INVx3_ASAP7_75t_L g3054 ( 
.A(n_2510),
.Y(n_3054)
);

AND2x2_ASAP7_75t_SL g3055 ( 
.A(n_2705),
.B(n_1120),
.Y(n_3055)
);

AND2x2_ASAP7_75t_L g3056 ( 
.A(n_2789),
.B(n_1437),
.Y(n_3056)
);

AND2x4_ASAP7_75t_L g3057 ( 
.A(n_2527),
.B(n_1351),
.Y(n_3057)
);

INVxp33_ASAP7_75t_L g3058 ( 
.A(n_2696),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2780),
.B(n_1438),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2529),
.Y(n_3060)
);

BUFx6f_ASAP7_75t_L g3061 ( 
.A(n_2510),
.Y(n_3061)
);

BUFx6f_ASAP7_75t_L g3062 ( 
.A(n_2567),
.Y(n_3062)
);

INVx2_ASAP7_75t_L g3063 ( 
.A(n_2443),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2550),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2550),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2556),
.Y(n_3066)
);

AO22x2_ASAP7_75t_L g3067 ( 
.A1(n_2704),
.A2(n_1371),
.B1(n_1385),
.B2(n_1369),
.Y(n_3067)
);

INVx4_ASAP7_75t_SL g3068 ( 
.A(n_2790),
.Y(n_3068)
);

INVx5_ASAP7_75t_L g3069 ( 
.A(n_2725),
.Y(n_3069)
);

NAND2xp5_ASAP7_75t_SL g3070 ( 
.A(n_2786),
.B(n_2794),
.Y(n_3070)
);

NAND2xp5_ASAP7_75t_SL g3071 ( 
.A(n_2556),
.B(n_1439),
.Y(n_3071)
);

NAND2xp5_ASAP7_75t_L g3072 ( 
.A(n_2665),
.B(n_2762),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2762),
.B(n_1443),
.Y(n_3073)
);

NAND2xp5_ASAP7_75t_SL g3074 ( 
.A(n_2564),
.B(n_1445),
.Y(n_3074)
);

INVx5_ASAP7_75t_L g3075 ( 
.A(n_2725),
.Y(n_3075)
);

INVx3_ASAP7_75t_L g3076 ( 
.A(n_2509),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2564),
.Y(n_3077)
);

INVx1_ASAP7_75t_SL g3078 ( 
.A(n_2719),
.Y(n_3078)
);

INVx1_ASAP7_75t_L g3079 ( 
.A(n_2446),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2448),
.Y(n_3080)
);

AND2x6_ASAP7_75t_L g3081 ( 
.A(n_2634),
.B(n_2636),
.Y(n_3081)
);

NAND2xp5_ASAP7_75t_L g3082 ( 
.A(n_2666),
.B(n_1447),
.Y(n_3082)
);

AND2x2_ASAP7_75t_L g3083 ( 
.A(n_2661),
.B(n_1451),
.Y(n_3083)
);

BUFx2_ASAP7_75t_L g3084 ( 
.A(n_2693),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2478),
.B(n_1452),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2449),
.Y(n_3086)
);

BUFx10_ASAP7_75t_L g3087 ( 
.A(n_2571),
.Y(n_3087)
);

INVx1_ASAP7_75t_L g3088 ( 
.A(n_2456),
.Y(n_3088)
);

INVx5_ASAP7_75t_L g3089 ( 
.A(n_2606),
.Y(n_3089)
);

NOR2xp33_ASAP7_75t_L g3090 ( 
.A(n_2730),
.B(n_1453),
.Y(n_3090)
);

INVx1_ASAP7_75t_L g3091 ( 
.A(n_2461),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2666),
.B(n_1457),
.Y(n_3092)
);

INVx1_ASAP7_75t_L g3093 ( 
.A(n_2463),
.Y(n_3093)
);

INVx4_ASAP7_75t_SL g3094 ( 
.A(n_2554),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2632),
.B(n_2429),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2464),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2469),
.Y(n_3097)
);

INVx4_ASAP7_75t_L g3098 ( 
.A(n_2606),
.Y(n_3098)
);

BUFx3_ASAP7_75t_L g3099 ( 
.A(n_2751),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2488),
.B(n_1458),
.Y(n_3100)
);

BUFx10_ASAP7_75t_L g3101 ( 
.A(n_2648),
.Y(n_3101)
);

INVx8_ASAP7_75t_L g3102 ( 
.A(n_2627),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2731),
.B(n_1459),
.Y(n_3103)
);

NAND2xp5_ASAP7_75t_L g3104 ( 
.A(n_2489),
.B(n_1460),
.Y(n_3104)
);

BUFx3_ASAP7_75t_L g3105 ( 
.A(n_2506),
.Y(n_3105)
);

BUFx2_ASAP7_75t_L g3106 ( 
.A(n_2722),
.Y(n_3106)
);

INVx1_ASAP7_75t_L g3107 ( 
.A(n_2517),
.Y(n_3107)
);

INVx2_ASAP7_75t_L g3108 ( 
.A(n_2518),
.Y(n_3108)
);

INVx1_ASAP7_75t_L g3109 ( 
.A(n_2522),
.Y(n_3109)
);

INVx1_ASAP7_75t_L g3110 ( 
.A(n_2526),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2530),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2492),
.B(n_1463),
.Y(n_3112)
);

INVx4_ASAP7_75t_L g3113 ( 
.A(n_2738),
.Y(n_3113)
);

AND2x2_ASAP7_75t_L g3114 ( 
.A(n_2647),
.B(n_1464),
.Y(n_3114)
);

OR2x2_ASAP7_75t_L g3115 ( 
.A(n_2410),
.B(n_1469),
.Y(n_3115)
);

INVx1_ASAP7_75t_L g3116 ( 
.A(n_2532),
.Y(n_3116)
);

INVx1_ASAP7_75t_L g3117 ( 
.A(n_2533),
.Y(n_3117)
);

INVx2_ASAP7_75t_SL g3118 ( 
.A(n_2627),
.Y(n_3118)
);

BUFx10_ASAP7_75t_L g3119 ( 
.A(n_2531),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2537),
.Y(n_3120)
);

BUFx10_ASAP7_75t_L g3121 ( 
.A(n_2555),
.Y(n_3121)
);

INVx2_ASAP7_75t_L g3122 ( 
.A(n_2539),
.Y(n_3122)
);

INVx2_ASAP7_75t_L g3123 ( 
.A(n_2546),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2599),
.B(n_1471),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2567),
.Y(n_3125)
);

OR2x6_ASAP7_75t_L g3126 ( 
.A(n_2739),
.B(n_1714),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2445),
.Y(n_3127)
);

AND2x6_ASAP7_75t_L g3128 ( 
.A(n_2634),
.B(n_1111),
.Y(n_3128)
);

HB1xp67_ASAP7_75t_L g3129 ( 
.A(n_2687),
.Y(n_3129)
);

AND2x4_ASAP7_75t_L g3130 ( 
.A(n_2672),
.B(n_1395),
.Y(n_3130)
);

AND2x4_ASAP7_75t_L g3131 ( 
.A(n_2672),
.B(n_1406),
.Y(n_3131)
);

NAND2xp5_ASAP7_75t_L g3132 ( 
.A(n_2498),
.B(n_1479),
.Y(n_3132)
);

INVx3_ASAP7_75t_L g3133 ( 
.A(n_2598),
.Y(n_3133)
);

BUFx4f_ASAP7_75t_L g3134 ( 
.A(n_2747),
.Y(n_3134)
);

BUFx2_ASAP7_75t_L g3135 ( 
.A(n_2523),
.Y(n_3135)
);

INVx1_ASAP7_75t_L g3136 ( 
.A(n_2667),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2445),
.Y(n_3137)
);

INVx1_ASAP7_75t_L g3138 ( 
.A(n_2676),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_L g3139 ( 
.A(n_2511),
.B(n_1481),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2680),
.B(n_1483),
.Y(n_3140)
);

AND2x4_ASAP7_75t_L g3141 ( 
.A(n_2692),
.B(n_2699),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2544),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2447),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2447),
.Y(n_3144)
);

INVx3_ASAP7_75t_L g3145 ( 
.A(n_2598),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2561),
.B(n_1484),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2450),
.Y(n_3147)
);

INVxp67_ASAP7_75t_SL g3148 ( 
.A(n_2450),
.Y(n_3148)
);

CKINVDCx11_ASAP7_75t_R g3149 ( 
.A(n_2745),
.Y(n_3149)
);

INVx4_ASAP7_75t_L g3150 ( 
.A(n_2627),
.Y(n_3150)
);

INVx3_ASAP7_75t_L g3151 ( 
.A(n_2617),
.Y(n_3151)
);

INVx2_ASAP7_75t_L g3152 ( 
.A(n_2458),
.Y(n_3152)
);

INVx4_ASAP7_75t_L g3153 ( 
.A(n_2462),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2458),
.Y(n_3154)
);

AND2x4_ASAP7_75t_L g3155 ( 
.A(n_2674),
.B(n_2701),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2505),
.Y(n_3156)
);

BUFx6f_ASAP7_75t_L g3157 ( 
.A(n_2617),
.Y(n_3157)
);

NOR2x1p5_ASAP7_75t_L g3158 ( 
.A(n_2477),
.B(n_1487),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2414),
.B(n_2691),
.Y(n_3159)
);

INVxp33_ASAP7_75t_L g3160 ( 
.A(n_2754),
.Y(n_3160)
);

AOI22xp33_ASAP7_75t_L g3161 ( 
.A1(n_2691),
.A2(n_1491),
.B1(n_1492),
.B2(n_1489),
.Y(n_3161)
);

BUFx6f_ASAP7_75t_L g3162 ( 
.A(n_2668),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_2695),
.B(n_1493),
.Y(n_3163)
);

NAND3xp33_ASAP7_75t_L g3164 ( 
.A(n_2592),
.B(n_1498),
.C(n_1495),
.Y(n_3164)
);

INVx2_ASAP7_75t_L g3165 ( 
.A(n_2655),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2695),
.B(n_1502),
.Y(n_3166)
);

INVx2_ASAP7_75t_L g3167 ( 
.A(n_2656),
.Y(n_3167)
);

NOR2xp33_ASAP7_75t_SL g3168 ( 
.A(n_2528),
.B(n_1503),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2613),
.B(n_1508),
.Y(n_3169)
);

BUFx2_ASAP7_75t_L g3170 ( 
.A(n_2748),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_SL g3171 ( 
.A(n_2746),
.B(n_1509),
.Y(n_3171)
);

BUFx6f_ASAP7_75t_L g3172 ( 
.A(n_2673),
.Y(n_3172)
);

OR2x6_ASAP7_75t_L g3173 ( 
.A(n_2747),
.B(n_1714),
.Y(n_3173)
);

BUFx3_ASAP7_75t_L g3174 ( 
.A(n_2707),
.Y(n_3174)
);

OR2x2_ASAP7_75t_L g3175 ( 
.A(n_2733),
.B(n_1510),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2640),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_2516),
.Y(n_3177)
);

NOR2xp33_ASAP7_75t_R g3178 ( 
.A(n_2749),
.B(n_1512),
.Y(n_3178)
);

INVx1_ASAP7_75t_L g3179 ( 
.A(n_2640),
.Y(n_3179)
);

OR2x6_ASAP7_75t_L g3180 ( 
.A(n_2736),
.B(n_1120),
.Y(n_3180)
);

BUFx3_ASAP7_75t_L g3181 ( 
.A(n_2708),
.Y(n_3181)
);

NOR2xp33_ASAP7_75t_L g3182 ( 
.A(n_2481),
.B(n_1513),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2756),
.Y(n_3183)
);

NOR2xp33_ASAP7_75t_L g3184 ( 
.A(n_2702),
.B(n_1515),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2636),
.Y(n_3185)
);

HB1xp67_ASAP7_75t_L g3186 ( 
.A(n_2740),
.Y(n_3186)
);

OAI22xp5_ASAP7_75t_L g3187 ( 
.A1(n_2637),
.A2(n_2582),
.B1(n_2591),
.B2(n_2584),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2582),
.Y(n_3188)
);

AND2x6_ASAP7_75t_L g3189 ( 
.A(n_2637),
.B(n_2584),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_2734),
.B(n_1518),
.Y(n_3190)
);

NAND3xp33_ASAP7_75t_L g3191 ( 
.A(n_2761),
.B(n_1723),
.C(n_1524),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_2591),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2702),
.B(n_1520),
.Y(n_3193)
);

INVx2_ASAP7_75t_L g3194 ( 
.A(n_2641),
.Y(n_3194)
);

BUFx3_ASAP7_75t_L g3195 ( 
.A(n_2709),
.Y(n_3195)
);

AO22x2_ASAP7_75t_L g3196 ( 
.A1(n_2562),
.A2(n_1409),
.B1(n_1411),
.B2(n_1407),
.Y(n_3196)
);

AOI22xp33_ASAP7_75t_L g3197 ( 
.A1(n_2778),
.A2(n_1533),
.B1(n_1537),
.B2(n_1531),
.Y(n_3197)
);

BUFx10_ASAP7_75t_L g3198 ( 
.A(n_2715),
.Y(n_3198)
);

INVxp67_ASAP7_75t_SL g3199 ( 
.A(n_2541),
.Y(n_3199)
);

CKINVDCx20_ASAP7_75t_R g3200 ( 
.A(n_2752),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_SL g3201 ( 
.A(n_2737),
.B(n_1544),
.Y(n_3201)
);

INVx2_ASAP7_75t_L g3202 ( 
.A(n_2646),
.Y(n_3202)
);

AND2x2_ASAP7_75t_L g3203 ( 
.A(n_2796),
.B(n_1546),
.Y(n_3203)
);

BUFx3_ASAP7_75t_L g3204 ( 
.A(n_2711),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_2601),
.Y(n_3205)
);

NAND2xp5_ASAP7_75t_L g3206 ( 
.A(n_2670),
.B(n_2433),
.Y(n_3206)
);

BUFx6f_ASAP7_75t_L g3207 ( 
.A(n_2578),
.Y(n_3207)
);

AND2x2_ASAP7_75t_L g3208 ( 
.A(n_2663),
.B(n_1548),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_2524),
.B(n_1550),
.Y(n_3209)
);

INVx5_ASAP7_75t_L g3210 ( 
.A(n_2712),
.Y(n_3210)
);

OR2x6_ASAP7_75t_L g3211 ( 
.A(n_2749),
.B(n_1207),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_2686),
.B(n_1551),
.Y(n_3212)
);

INVxp33_ASAP7_75t_L g3213 ( 
.A(n_2750),
.Y(n_3213)
);

INVx1_ASAP7_75t_L g3214 ( 
.A(n_2646),
.Y(n_3214)
);

INVx1_ASAP7_75t_L g3215 ( 
.A(n_2649),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2583),
.Y(n_3216)
);

AND2x2_ASAP7_75t_SL g3217 ( 
.A(n_2750),
.B(n_1207),
.Y(n_3217)
);

INVx1_ASAP7_75t_L g3218 ( 
.A(n_2649),
.Y(n_3218)
);

INVx4_ASAP7_75t_L g3219 ( 
.A(n_2714),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2679),
.Y(n_3220)
);

AND2x4_ASAP7_75t_L g3221 ( 
.A(n_2716),
.B(n_1412),
.Y(n_3221)
);

INVx2_ASAP7_75t_L g3222 ( 
.A(n_2472),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_SL g3223 ( 
.A(n_2765),
.B(n_1553),
.Y(n_3223)
);

OR2x6_ASAP7_75t_L g3224 ( 
.A(n_2690),
.B(n_2743),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_2683),
.B(n_1555),
.Y(n_3225)
);

AND2x4_ASAP7_75t_L g3226 ( 
.A(n_2717),
.B(n_1413),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_2743),
.B(n_1564),
.Y(n_3227)
);

INVx2_ASAP7_75t_L g3228 ( 
.A(n_2475),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2482),
.Y(n_3229)
);

AOI22xp5_ASAP7_75t_L g3230 ( 
.A1(n_2542),
.A2(n_1568),
.B1(n_1569),
.B2(n_1565),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_SL g3231 ( 
.A(n_2688),
.B(n_1570),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_2651),
.B(n_1571),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_2681),
.B(n_1573),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_SL g3234 ( 
.A(n_2689),
.B(n_1574),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2487),
.Y(n_3235)
);

AND2x6_ASAP7_75t_L g3236 ( 
.A(n_2601),
.B(n_1150),
.Y(n_3236)
);

BUFx2_ASAP7_75t_L g3237 ( 
.A(n_2724),
.Y(n_3237)
);

INVx1_ASAP7_75t_L g3238 ( 
.A(n_2490),
.Y(n_3238)
);

NOR2xp33_ASAP7_75t_L g3239 ( 
.A(n_2581),
.B(n_1575),
.Y(n_3239)
);

BUFx10_ASAP7_75t_L g3240 ( 
.A(n_2726),
.Y(n_3240)
);

INVx1_ASAP7_75t_SL g3241 ( 
.A(n_2718),
.Y(n_3241)
);

INVx4_ASAP7_75t_L g3242 ( 
.A(n_2720),
.Y(n_3242)
);

INVx4_ASAP7_75t_L g3243 ( 
.A(n_2494),
.Y(n_3243)
);

HB1xp67_ASAP7_75t_L g3244 ( 
.A(n_2535),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2495),
.Y(n_3245)
);

INVx4_ASAP7_75t_L g3246 ( 
.A(n_2496),
.Y(n_3246)
);

INVx2_ASAP7_75t_SL g3247 ( 
.A(n_2694),
.Y(n_3247)
);

INVx4_ASAP7_75t_L g3248 ( 
.A(n_2499),
.Y(n_3248)
);

INVx1_ASAP7_75t_L g3249 ( 
.A(n_2500),
.Y(n_3249)
);

AND2x2_ASAP7_75t_SL g3250 ( 
.A(n_2682),
.B(n_1223),
.Y(n_3250)
);

INVx2_ASAP7_75t_L g3251 ( 
.A(n_2501),
.Y(n_3251)
);

AND2x4_ASAP7_75t_L g3252 ( 
.A(n_2579),
.B(n_1422),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2543),
.B(n_1577),
.Y(n_3253)
);

AOI22xp33_ASAP7_75t_L g3254 ( 
.A1(n_2586),
.A2(n_1583),
.B1(n_1585),
.B2(n_1579),
.Y(n_3254)
);

NOR2xp33_ASAP7_75t_L g3255 ( 
.A(n_2615),
.B(n_1586),
.Y(n_3255)
);

BUFx3_ASAP7_75t_L g3256 ( 
.A(n_2644),
.Y(n_3256)
);

BUFx3_ASAP7_75t_L g3257 ( 
.A(n_2644),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2504),
.Y(n_3258)
);

AND2x6_ASAP7_75t_L g3259 ( 
.A(n_2607),
.B(n_1150),
.Y(n_3259)
);

NOR2xp33_ASAP7_75t_L g3260 ( 
.A(n_2623),
.B(n_1589),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2664),
.Y(n_3261)
);

NAND2xp5_ASAP7_75t_SL g3262 ( 
.A(n_2607),
.B(n_2619),
.Y(n_3262)
);

INVx1_ASAP7_75t_L g3263 ( 
.A(n_2535),
.Y(n_3263)
);

NOR2xp33_ASAP7_75t_L g3264 ( 
.A(n_2629),
.B(n_2497),
.Y(n_3264)
);

CKINVDCx20_ASAP7_75t_R g3265 ( 
.A(n_2710),
.Y(n_3265)
);

NAND2xp5_ASAP7_75t_L g3266 ( 
.A(n_2551),
.B(n_1590),
.Y(n_3266)
);

INVx3_ASAP7_75t_L g3267 ( 
.A(n_2619),
.Y(n_3267)
);

BUFx6f_ASAP7_75t_L g3268 ( 
.A(n_2621),
.Y(n_3268)
);

INVx3_ASAP7_75t_L g3269 ( 
.A(n_2621),
.Y(n_3269)
);

INVx1_ASAP7_75t_L g3270 ( 
.A(n_2485),
.Y(n_3270)
);

INVx2_ASAP7_75t_L g3271 ( 
.A(n_2485),
.Y(n_3271)
);

INVx3_ASAP7_75t_L g3272 ( 
.A(n_2660),
.Y(n_3272)
);

AND2x6_ASAP7_75t_L g3273 ( 
.A(n_2713),
.B(n_1150),
.Y(n_3273)
);

INVxp33_ASAP7_75t_L g3274 ( 
.A(n_2723),
.Y(n_3274)
);

INVx4_ASAP7_75t_L g3275 ( 
.A(n_2570),
.Y(n_3275)
);

BUFx3_ASAP7_75t_L g3276 ( 
.A(n_2659),
.Y(n_3276)
);

INVx2_ASAP7_75t_L g3277 ( 
.A(n_2405),
.Y(n_3277)
);

INVx2_ASAP7_75t_L g3278 ( 
.A(n_2405),
.Y(n_3278)
);

INVx3_ASAP7_75t_L g3279 ( 
.A(n_2404),
.Y(n_3279)
);

INVx1_ASAP7_75t_L g3280 ( 
.A(n_2480),
.Y(n_3280)
);

INVx4_ASAP7_75t_L g3281 ( 
.A(n_2659),
.Y(n_3281)
);

AND3x4_ASAP7_75t_L g3282 ( 
.A(n_2580),
.B(n_1246),
.C(n_1223),
.Y(n_3282)
);

AND2x2_ASAP7_75t_SL g3283 ( 
.A(n_2413),
.B(n_1246),
.Y(n_3283)
);

INVx3_ASAP7_75t_L g3284 ( 
.A(n_2404),
.Y(n_3284)
);

OAI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_2423),
.A2(n_1596),
.B1(n_1597),
.B2(n_1594),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_2480),
.Y(n_3286)
);

NAND2xp5_ASAP7_75t_L g3287 ( 
.A(n_2642),
.B(n_1598),
.Y(n_3287)
);

OR2x2_ASAP7_75t_L g3288 ( 
.A(n_2764),
.B(n_1599),
.Y(n_3288)
);

BUFx4f_ASAP7_75t_L g3289 ( 
.A(n_2675),
.Y(n_3289)
);

BUFx3_ASAP7_75t_L g3290 ( 
.A(n_2659),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_SL g3291 ( 
.A(n_2631),
.B(n_1605),
.Y(n_3291)
);

NAND2xp5_ASAP7_75t_SL g3292 ( 
.A(n_2631),
.B(n_1607),
.Y(n_3292)
);

AND2x2_ASAP7_75t_L g3293 ( 
.A(n_2764),
.B(n_1608),
.Y(n_3293)
);

BUFx6f_ASAP7_75t_L g3294 ( 
.A(n_2404),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_L g3295 ( 
.A(n_2459),
.B(n_1611),
.Y(n_3295)
);

INVx4_ASAP7_75t_L g3296 ( 
.A(n_2659),
.Y(n_3296)
);

INVx3_ASAP7_75t_L g3297 ( 
.A(n_2404),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_2480),
.Y(n_3298)
);

NAND2xp5_ASAP7_75t_L g3299 ( 
.A(n_2642),
.B(n_1612),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_SL g3300 ( 
.A(n_2631),
.B(n_1614),
.Y(n_3300)
);

AND2x2_ASAP7_75t_L g3301 ( 
.A(n_2764),
.B(n_1615),
.Y(n_3301)
);

AOI22xp33_ASAP7_75t_L g3302 ( 
.A1(n_2420),
.A2(n_1625),
.B1(n_1626),
.B2(n_1617),
.Y(n_3302)
);

INVx3_ASAP7_75t_L g3303 ( 
.A(n_2404),
.Y(n_3303)
);

BUFx6f_ASAP7_75t_L g3304 ( 
.A(n_2404),
.Y(n_3304)
);

INVx1_ASAP7_75t_SL g3305 ( 
.A(n_2406),
.Y(n_3305)
);

INVxp67_ASAP7_75t_L g3306 ( 
.A(n_2406),
.Y(n_3306)
);

OAI22xp33_ASAP7_75t_SL g3307 ( 
.A1(n_2413),
.A2(n_1630),
.B1(n_1633),
.B2(n_1628),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_2480),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_2642),
.B(n_1636),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2642),
.B(n_1637),
.Y(n_3310)
);

NAND2xp5_ASAP7_75t_L g3311 ( 
.A(n_2642),
.B(n_1641),
.Y(n_3311)
);

INVx2_ASAP7_75t_SL g3312 ( 
.A(n_2659),
.Y(n_3312)
);

INVx1_ASAP7_75t_SL g3313 ( 
.A(n_2406),
.Y(n_3313)
);

NAND2xp5_ASAP7_75t_L g3314 ( 
.A(n_2642),
.B(n_1644),
.Y(n_3314)
);

INVx1_ASAP7_75t_SL g3315 ( 
.A(n_2406),
.Y(n_3315)
);

NAND2xp5_ASAP7_75t_L g3316 ( 
.A(n_2642),
.B(n_1651),
.Y(n_3316)
);

INVx3_ASAP7_75t_L g3317 ( 
.A(n_2404),
.Y(n_3317)
);

BUFx10_ASAP7_75t_L g3318 ( 
.A(n_2560),
.Y(n_3318)
);

NAND2xp5_ASAP7_75t_L g3319 ( 
.A(n_2642),
.B(n_1652),
.Y(n_3319)
);

NOR2xp33_ASAP7_75t_L g3320 ( 
.A(n_2459),
.B(n_1655),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2480),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_2480),
.Y(n_3322)
);

INVx3_ASAP7_75t_L g3323 ( 
.A(n_2404),
.Y(n_3323)
);

NAND2xp5_ASAP7_75t_SL g3324 ( 
.A(n_2631),
.B(n_1658),
.Y(n_3324)
);

INVx3_ASAP7_75t_L g3325 ( 
.A(n_2404),
.Y(n_3325)
);

OR2x2_ASAP7_75t_L g3326 ( 
.A(n_2764),
.B(n_1659),
.Y(n_3326)
);

INVx4_ASAP7_75t_L g3327 ( 
.A(n_2659),
.Y(n_3327)
);

INVx3_ASAP7_75t_L g3328 ( 
.A(n_2404),
.Y(n_3328)
);

INVx2_ASAP7_75t_L g3329 ( 
.A(n_2405),
.Y(n_3329)
);

BUFx3_ASAP7_75t_L g3330 ( 
.A(n_2659),
.Y(n_3330)
);

NAND2xp5_ASAP7_75t_L g3331 ( 
.A(n_2642),
.B(n_1660),
.Y(n_3331)
);

INVx1_ASAP7_75t_L g3332 ( 
.A(n_2480),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2642),
.B(n_1662),
.Y(n_3333)
);

CKINVDCx5p33_ASAP7_75t_R g3334 ( 
.A(n_2706),
.Y(n_3334)
);

AND2x4_ASAP7_75t_L g3335 ( 
.A(n_2642),
.B(n_1427),
.Y(n_3335)
);

BUFx3_ASAP7_75t_L g3336 ( 
.A(n_2659),
.Y(n_3336)
);

INVx1_ASAP7_75t_L g3337 ( 
.A(n_2480),
.Y(n_3337)
);

CKINVDCx20_ASAP7_75t_R g3338 ( 
.A(n_2706),
.Y(n_3338)
);

NOR2xp33_ASAP7_75t_L g3339 ( 
.A(n_2459),
.B(n_1664),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_2480),
.Y(n_3340)
);

NAND3xp33_ASAP7_75t_L g3341 ( 
.A(n_2678),
.B(n_1712),
.C(n_1704),
.Y(n_3341)
);

INVx4_ASAP7_75t_L g3342 ( 
.A(n_2659),
.Y(n_3342)
);

OAI221xp5_ASAP7_75t_L g3343 ( 
.A1(n_2764),
.A2(n_1668),
.B1(n_1670),
.B2(n_1666),
.C(n_1665),
.Y(n_3343)
);

AND2x2_ASAP7_75t_L g3344 ( 
.A(n_2764),
.B(n_1678),
.Y(n_3344)
);

INVx2_ASAP7_75t_L g3345 ( 
.A(n_2405),
.Y(n_3345)
);

INVx5_ASAP7_75t_L g3346 ( 
.A(n_2560),
.Y(n_3346)
);

INVx3_ASAP7_75t_L g3347 ( 
.A(n_2404),
.Y(n_3347)
);

INVx3_ASAP7_75t_L g3348 ( 
.A(n_2404),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_2480),
.Y(n_3349)
);

INVxp33_ASAP7_75t_L g3350 ( 
.A(n_2406),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2642),
.B(n_1679),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_2405),
.Y(n_3352)
);

INVx2_ASAP7_75t_SL g3353 ( 
.A(n_2659),
.Y(n_3353)
);

INVx3_ASAP7_75t_L g3354 ( 
.A(n_2404),
.Y(n_3354)
);

OR2x2_ASAP7_75t_L g3355 ( 
.A(n_2764),
.B(n_1687),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_SL g3356 ( 
.A(n_2631),
.B(n_1688),
.Y(n_3356)
);

BUFx6f_ASAP7_75t_L g3357 ( 
.A(n_2404),
.Y(n_3357)
);

NOR2x1p5_ASAP7_75t_L g3358 ( 
.A(n_2735),
.B(n_1690),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_2480),
.Y(n_3359)
);

INVx1_ASAP7_75t_L g3360 ( 
.A(n_2480),
.Y(n_3360)
);

CKINVDCx5p33_ASAP7_75t_R g3361 ( 
.A(n_2706),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_2480),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_2480),
.Y(n_3363)
);

HB1xp67_ASAP7_75t_L g3364 ( 
.A(n_2560),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_SL g3365 ( 
.A(n_2631),
.B(n_1695),
.Y(n_3365)
);

INVx2_ASAP7_75t_L g3366 ( 
.A(n_2405),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_2480),
.Y(n_3367)
);

INVx4_ASAP7_75t_SL g3368 ( 
.A(n_2580),
.Y(n_3368)
);

BUFx6f_ASAP7_75t_L g3369 ( 
.A(n_2404),
.Y(n_3369)
);

NOR2x1p5_ASAP7_75t_L g3370 ( 
.A(n_2735),
.B(n_1696),
.Y(n_3370)
);

AND2x6_ASAP7_75t_L g3371 ( 
.A(n_2588),
.B(n_1150),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_2480),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_2764),
.B(n_1697),
.Y(n_3373)
);

INVx1_ASAP7_75t_L g3374 ( 
.A(n_2480),
.Y(n_3374)
);

INVx1_ASAP7_75t_L g3375 ( 
.A(n_2480),
.Y(n_3375)
);

BUFx3_ASAP7_75t_L g3376 ( 
.A(n_2659),
.Y(n_3376)
);

INVx2_ASAP7_75t_L g3377 ( 
.A(n_2405),
.Y(n_3377)
);

INVx2_ASAP7_75t_L g3378 ( 
.A(n_2405),
.Y(n_3378)
);

CKINVDCx5p33_ASAP7_75t_R g3379 ( 
.A(n_2706),
.Y(n_3379)
);

INVx2_ASAP7_75t_L g3380 ( 
.A(n_2405),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_2480),
.Y(n_3381)
);

NAND2xp5_ASAP7_75t_L g3382 ( 
.A(n_2642),
.B(n_1717),
.Y(n_3382)
);

CKINVDCx16_ASAP7_75t_R g3383 ( 
.A(n_2560),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_2480),
.Y(n_3384)
);

INVx2_ASAP7_75t_L g3385 ( 
.A(n_2405),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_2420),
.A2(n_1722),
.B1(n_1718),
.B2(n_1441),
.Y(n_3386)
);

OAI22xp33_ASAP7_75t_SL g3387 ( 
.A1(n_2413),
.A2(n_1442),
.B1(n_1444),
.B2(n_1428),
.Y(n_3387)
);

INVx8_ASAP7_75t_L g3388 ( 
.A(n_2659),
.Y(n_3388)
);

BUFx2_ASAP7_75t_L g3389 ( 
.A(n_2560),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_2573),
.Y(n_3390)
);

AND2x6_ASAP7_75t_L g3391 ( 
.A(n_2588),
.B(n_1190),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2405),
.Y(n_3392)
);

BUFx6f_ASAP7_75t_L g3393 ( 
.A(n_2404),
.Y(n_3393)
);

AND2x4_ASAP7_75t_L g3394 ( 
.A(n_2642),
.B(n_1448),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2573),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_SL g3396 ( 
.A(n_2631),
.B(n_1277),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_2642),
.B(n_1456),
.Y(n_3397)
);

HB1xp67_ASAP7_75t_L g3398 ( 
.A(n_2560),
.Y(n_3398)
);

CKINVDCx5p33_ASAP7_75t_R g3399 ( 
.A(n_2706),
.Y(n_3399)
);

BUFx3_ASAP7_75t_L g3400 ( 
.A(n_2659),
.Y(n_3400)
);

CKINVDCx20_ASAP7_75t_R g3401 ( 
.A(n_2706),
.Y(n_3401)
);

INVx1_ASAP7_75t_SL g3402 ( 
.A(n_2406),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_2642),
.B(n_1461),
.Y(n_3403)
);

INVxp67_ASAP7_75t_SL g3404 ( 
.A(n_2404),
.Y(n_3404)
);

INVx1_ASAP7_75t_L g3405 ( 
.A(n_2573),
.Y(n_3405)
);

INVx4_ASAP7_75t_SL g3406 ( 
.A(n_2580),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2573),
.Y(n_3407)
);

BUFx3_ASAP7_75t_L g3408 ( 
.A(n_2659),
.Y(n_3408)
);

BUFx6f_ASAP7_75t_L g3409 ( 
.A(n_2404),
.Y(n_3409)
);

NOR2xp33_ASAP7_75t_L g3410 ( 
.A(n_2459),
.B(n_1466),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_2404),
.Y(n_3411)
);

BUFx3_ASAP7_75t_L g3412 ( 
.A(n_2659),
.Y(n_3412)
);

NOR2xp33_ASAP7_75t_L g3413 ( 
.A(n_2459),
.B(n_1467),
.Y(n_3413)
);

NOR2xp33_ASAP7_75t_L g3414 ( 
.A(n_2459),
.B(n_1470),
.Y(n_3414)
);

INVx1_ASAP7_75t_L g3415 ( 
.A(n_2573),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_2405),
.Y(n_3416)
);

INVx5_ASAP7_75t_L g3417 ( 
.A(n_2560),
.Y(n_3417)
);

AOI22xp33_ASAP7_75t_L g3418 ( 
.A1(n_2420),
.A2(n_1486),
.B1(n_1488),
.B2(n_1478),
.Y(n_3418)
);

BUFx4f_ASAP7_75t_L g3419 ( 
.A(n_2675),
.Y(n_3419)
);

CKINVDCx5p33_ASAP7_75t_R g3420 ( 
.A(n_2706),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2573),
.Y(n_3421)
);

INVx2_ASAP7_75t_L g3422 ( 
.A(n_2405),
.Y(n_3422)
);

NAND2xp5_ASAP7_75t_L g3423 ( 
.A(n_2642),
.B(n_1490),
.Y(n_3423)
);

INVx2_ASAP7_75t_L g3424 ( 
.A(n_2405),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_2573),
.Y(n_3425)
);

NOR2x1p5_ASAP7_75t_L g3426 ( 
.A(n_2735),
.B(n_1691),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_2573),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_2642),
.B(n_1496),
.Y(n_3428)
);

INVx1_ASAP7_75t_L g3429 ( 
.A(n_2573),
.Y(n_3429)
);

INVx1_ASAP7_75t_L g3430 ( 
.A(n_2573),
.Y(n_3430)
);

INVxp67_ASAP7_75t_SL g3431 ( 
.A(n_2404),
.Y(n_3431)
);

INVx4_ASAP7_75t_SL g3432 ( 
.A(n_2580),
.Y(n_3432)
);

NAND2xp33_ASAP7_75t_L g3433 ( 
.A(n_2565),
.B(n_1190),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_SL g3434 ( 
.A(n_2631),
.B(n_1698),
.Y(n_3434)
);

AND2x2_ASAP7_75t_L g3435 ( 
.A(n_2764),
.B(n_1497),
.Y(n_3435)
);

NAND3xp33_ASAP7_75t_L g3436 ( 
.A(n_2678),
.B(n_1226),
.C(n_1190),
.Y(n_3436)
);

AO22x2_ASAP7_75t_L g3437 ( 
.A1(n_2512),
.A2(n_1500),
.B1(n_1501),
.B2(n_1499),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_2405),
.Y(n_3438)
);

INVx4_ASAP7_75t_L g3439 ( 
.A(n_2659),
.Y(n_3439)
);

INVx2_ASAP7_75t_L g3440 ( 
.A(n_2405),
.Y(n_3440)
);

NOR2xp33_ASAP7_75t_L g3441 ( 
.A(n_2459),
.B(n_1504),
.Y(n_3441)
);

NAND2xp5_ASAP7_75t_SL g3442 ( 
.A(n_2631),
.B(n_1277),
.Y(n_3442)
);

INVx1_ASAP7_75t_SL g3443 ( 
.A(n_2406),
.Y(n_3443)
);

INVx2_ASAP7_75t_L g3444 ( 
.A(n_2405),
.Y(n_3444)
);

BUFx6f_ASAP7_75t_L g3445 ( 
.A(n_2404),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_2459),
.B(n_1505),
.Y(n_3446)
);

BUFx6f_ASAP7_75t_L g3447 ( 
.A(n_2404),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_2459),
.B(n_1514),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_2573),
.Y(n_3449)
);

BUFx3_ASAP7_75t_L g3450 ( 
.A(n_2659),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_2642),
.B(n_1516),
.Y(n_3451)
);

AO22x2_ASAP7_75t_L g3452 ( 
.A1(n_2512),
.A2(n_1521),
.B1(n_1526),
.B2(n_1517),
.Y(n_3452)
);

NAND2xp5_ASAP7_75t_L g3453 ( 
.A(n_2642),
.B(n_1527),
.Y(n_3453)
);

AOI22xp5_ASAP7_75t_L g3454 ( 
.A1(n_2471),
.A2(n_1539),
.B1(n_1540),
.B2(n_1529),
.Y(n_3454)
);

AND2x4_ASAP7_75t_L g3455 ( 
.A(n_2642),
.B(n_1541),
.Y(n_3455)
);

NOR2xp33_ASAP7_75t_L g3456 ( 
.A(n_2459),
.B(n_1542),
.Y(n_3456)
);

AND2x6_ASAP7_75t_L g3457 ( 
.A(n_2588),
.B(n_1190),
.Y(n_3457)
);

BUFx6f_ASAP7_75t_L g3458 ( 
.A(n_2404),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_2573),
.Y(n_3459)
);

INVx1_ASAP7_75t_L g3460 ( 
.A(n_3129),
.Y(n_3460)
);

NAND2xp5_ASAP7_75t_L g3461 ( 
.A(n_3001),
.B(n_1552),
.Y(n_3461)
);

NAND2xp5_ASAP7_75t_L g3462 ( 
.A(n_3001),
.B(n_1557),
.Y(n_3462)
);

INVx3_ASAP7_75t_L g3463 ( 
.A(n_3189),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_2861),
.Y(n_3464)
);

INVx8_ASAP7_75t_L g3465 ( 
.A(n_3388),
.Y(n_3465)
);

BUFx6f_ASAP7_75t_L g3466 ( 
.A(n_2834),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_2849),
.Y(n_3467)
);

NOR2xp33_ASAP7_75t_SL g3468 ( 
.A(n_3038),
.B(n_1278),
.Y(n_3468)
);

NOR3xp33_ASAP7_75t_L g3469 ( 
.A(n_3038),
.B(n_1563),
.C(n_1558),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3010),
.B(n_1566),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_SL g3471 ( 
.A(n_3383),
.B(n_1226),
.Y(n_3471)
);

OAI22xp33_ASAP7_75t_L g3472 ( 
.A1(n_3168),
.A2(n_1582),
.B1(n_1584),
.B2(n_1581),
.Y(n_3472)
);

NOR2xp67_ASAP7_75t_L g3473 ( 
.A(n_2829),
.B(n_45),
.Y(n_3473)
);

NAND2xp5_ASAP7_75t_L g3474 ( 
.A(n_3010),
.B(n_1588),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3280),
.Y(n_3475)
);

NAND2xp5_ASAP7_75t_L g3476 ( 
.A(n_2823),
.B(n_1600),
.Y(n_3476)
);

AOI22xp5_ASAP7_75t_L g3477 ( 
.A1(n_3187),
.A2(n_1609),
.B1(n_1613),
.B2(n_1604),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_3058),
.B(n_1616),
.Y(n_3478)
);

NAND2xp5_ASAP7_75t_SL g3479 ( 
.A(n_2829),
.B(n_1226),
.Y(n_3479)
);

INVx1_ASAP7_75t_L g3480 ( 
.A(n_3286),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_2853),
.B(n_1619),
.Y(n_3481)
);

NAND2xp5_ASAP7_75t_SL g3482 ( 
.A(n_2829),
.B(n_1226),
.Y(n_3482)
);

INVx2_ASAP7_75t_L g3483 ( 
.A(n_3188),
.Y(n_3483)
);

NOR2xp33_ASAP7_75t_SL g3484 ( 
.A(n_2993),
.B(n_1278),
.Y(n_3484)
);

NAND2xp5_ASAP7_75t_L g3485 ( 
.A(n_2940),
.B(n_1622),
.Y(n_3485)
);

NOR2xp33_ASAP7_75t_L g3486 ( 
.A(n_2929),
.B(n_2856),
.Y(n_3486)
);

INVx1_ASAP7_75t_L g3487 ( 
.A(n_3298),
.Y(n_3487)
);

AOI21xp5_ASAP7_75t_L g3488 ( 
.A1(n_3262),
.A2(n_1332),
.B(n_1331),
.Y(n_3488)
);

INVx2_ASAP7_75t_L g3489 ( 
.A(n_3188),
.Y(n_3489)
);

NAND2xp5_ASAP7_75t_L g3490 ( 
.A(n_3142),
.B(n_1624),
.Y(n_3490)
);

NAND2xp33_ASAP7_75t_L g3491 ( 
.A(n_2993),
.B(n_1227),
.Y(n_3491)
);

AOI22xp33_ASAP7_75t_L g3492 ( 
.A1(n_3055),
.A2(n_1309),
.B1(n_1318),
.B2(n_1227),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3192),
.Y(n_3493)
);

NAND2xp5_ASAP7_75t_SL g3494 ( 
.A(n_3346),
.B(n_1227),
.Y(n_3494)
);

OAI22xp5_ASAP7_75t_SL g3495 ( 
.A1(n_3282),
.A2(n_1634),
.B1(n_1640),
.B2(n_1629),
.Y(n_3495)
);

NOR2x1p5_ASAP7_75t_L g3496 ( 
.A(n_2826),
.B(n_1331),
.Y(n_3496)
);

INVx3_ASAP7_75t_L g3497 ( 
.A(n_3189),
.Y(n_3497)
);

NAND2xp5_ASAP7_75t_L g3498 ( 
.A(n_2869),
.B(n_1642),
.Y(n_3498)
);

NAND2xp5_ASAP7_75t_SL g3499 ( 
.A(n_3346),
.B(n_1227),
.Y(n_3499)
);

AND2x2_ASAP7_75t_L g3500 ( 
.A(n_2944),
.B(n_1649),
.Y(n_3500)
);

NAND2xp5_ASAP7_75t_L g3501 ( 
.A(n_3020),
.B(n_1653),
.Y(n_3501)
);

AOI22xp33_ASAP7_75t_L g3502 ( 
.A1(n_3217),
.A2(n_1318),
.B1(n_1363),
.B2(n_1309),
.Y(n_3502)
);

NOR2xp33_ASAP7_75t_L g3503 ( 
.A(n_3031),
.B(n_1654),
.Y(n_3503)
);

NAND2xp5_ASAP7_75t_SL g3504 ( 
.A(n_3346),
.B(n_1309),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3020),
.B(n_1656),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_SL g3506 ( 
.A(n_3417),
.B(n_1309),
.Y(n_3506)
);

AOI22xp5_ASAP7_75t_L g3507 ( 
.A1(n_2938),
.A2(n_1661),
.B1(n_1667),
.B2(n_1657),
.Y(n_3507)
);

OR2x2_ASAP7_75t_L g3508 ( 
.A(n_2804),
.B(n_1707),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3192),
.Y(n_3509)
);

OAI22xp5_ASAP7_75t_L g3510 ( 
.A1(n_3437),
.A2(n_1332),
.B1(n_1361),
.B2(n_1338),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3021),
.B(n_1669),
.Y(n_3511)
);

INVx2_ASAP7_75t_SL g3512 ( 
.A(n_3388),
.Y(n_3512)
);

NAND2xp5_ASAP7_75t_L g3513 ( 
.A(n_3021),
.B(n_1674),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_R g3514 ( 
.A(n_3338),
.B(n_3401),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3043),
.B(n_3045),
.Y(n_3515)
);

NAND2x1p5_ASAP7_75t_L g3516 ( 
.A(n_3026),
.B(n_1318),
.Y(n_3516)
);

INVx2_ASAP7_75t_L g3517 ( 
.A(n_3205),
.Y(n_3517)
);

NAND2xp5_ASAP7_75t_SL g3518 ( 
.A(n_3417),
.B(n_1318),
.Y(n_3518)
);

NAND2xp5_ASAP7_75t_L g3519 ( 
.A(n_3043),
.B(n_1676),
.Y(n_3519)
);

AND2x2_ASAP7_75t_L g3520 ( 
.A(n_2900),
.B(n_1680),
.Y(n_3520)
);

NOR2xp33_ASAP7_75t_L g3521 ( 
.A(n_2902),
.B(n_1686),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_3417),
.B(n_1363),
.Y(n_3522)
);

BUFx6f_ASAP7_75t_SL g3523 ( 
.A(n_3008),
.Y(n_3523)
);

NAND3xp33_ASAP7_75t_L g3524 ( 
.A(n_3436),
.B(n_1480),
.C(n_1363),
.Y(n_3524)
);

BUFx3_ASAP7_75t_L g3525 ( 
.A(n_3276),
.Y(n_3525)
);

INVx2_ASAP7_75t_SL g3526 ( 
.A(n_2888),
.Y(n_3526)
);

BUFx3_ASAP7_75t_L g3527 ( 
.A(n_3290),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3045),
.B(n_1689),
.Y(n_3528)
);

INVx2_ASAP7_75t_SL g3529 ( 
.A(n_2888),
.Y(n_3529)
);

NAND2xp5_ASAP7_75t_SL g3530 ( 
.A(n_3283),
.B(n_1363),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3308),
.Y(n_3531)
);

A2O1A1Ixp33_ASAP7_75t_L g3532 ( 
.A1(n_3095),
.A2(n_1361),
.B(n_1362),
.C(n_1338),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3321),
.Y(n_3533)
);

NOR2xp33_ASAP7_75t_L g3534 ( 
.A(n_3350),
.B(n_1693),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3205),
.Y(n_3535)
);

INVx1_ASAP7_75t_L g3536 ( 
.A(n_3322),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3050),
.B(n_1694),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3332),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3050),
.B(n_1702),
.Y(n_3539)
);

INVx2_ASAP7_75t_L g3540 ( 
.A(n_3060),
.Y(n_3540)
);

INVx1_ASAP7_75t_L g3541 ( 
.A(n_3337),
.Y(n_3541)
);

INVx2_ASAP7_75t_SL g3542 ( 
.A(n_3289),
.Y(n_3542)
);

NAND2xp5_ASAP7_75t_L g3543 ( 
.A(n_3060),
.B(n_1710),
.Y(n_3543)
);

NAND2xp5_ASAP7_75t_L g3544 ( 
.A(n_3064),
.B(n_1716),
.Y(n_3544)
);

INVx2_ASAP7_75t_L g3545 ( 
.A(n_3064),
.Y(n_3545)
);

INVx1_ASAP7_75t_L g3546 ( 
.A(n_3340),
.Y(n_3546)
);

NAND2xp33_ASAP7_75t_L g3547 ( 
.A(n_2993),
.B(n_1480),
.Y(n_3547)
);

BUFx6f_ASAP7_75t_L g3548 ( 
.A(n_2834),
.Y(n_3548)
);

INVx1_ASAP7_75t_L g3549 ( 
.A(n_3349),
.Y(n_3549)
);

INVx3_ASAP7_75t_L g3550 ( 
.A(n_3189),
.Y(n_3550)
);

NAND2xp5_ASAP7_75t_L g3551 ( 
.A(n_3065),
.B(n_1721),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_2885),
.B(n_2981),
.Y(n_3552)
);

NAND2xp5_ASAP7_75t_SL g3553 ( 
.A(n_2850),
.B(n_1480),
.Y(n_3553)
);

NAND2xp5_ASAP7_75t_SL g3554 ( 
.A(n_3268),
.B(n_1480),
.Y(n_3554)
);

NAND2xp5_ASAP7_75t_L g3555 ( 
.A(n_3065),
.B(n_1724),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3066),
.B(n_1725),
.Y(n_3556)
);

OR2x6_ASAP7_75t_L g3557 ( 
.A(n_3102),
.B(n_1362),
.Y(n_3557)
);

NOR2x1p5_ASAP7_75t_L g3558 ( 
.A(n_2799),
.B(n_1377),
.Y(n_3558)
);

INVx2_ASAP7_75t_L g3559 ( 
.A(n_3066),
.Y(n_3559)
);

NAND2xp5_ASAP7_75t_SL g3560 ( 
.A(n_3268),
.B(n_1519),
.Y(n_3560)
);

CKINVDCx5p33_ASAP7_75t_R g3561 ( 
.A(n_3042),
.Y(n_3561)
);

INVx1_ASAP7_75t_L g3562 ( 
.A(n_3359),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_3285),
.B(n_1726),
.Y(n_3563)
);

HB1xp67_ASAP7_75t_L g3564 ( 
.A(n_2876),
.Y(n_3564)
);

INVx2_ASAP7_75t_L g3565 ( 
.A(n_3077),
.Y(n_3565)
);

INVx2_ASAP7_75t_L g3566 ( 
.A(n_3077),
.Y(n_3566)
);

INVx2_ASAP7_75t_L g3567 ( 
.A(n_3185),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3185),
.B(n_1377),
.Y(n_3568)
);

INVx2_ASAP7_75t_L g3569 ( 
.A(n_2806),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_SL g3570 ( 
.A(n_3268),
.B(n_1519),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3335),
.B(n_1379),
.Y(n_3571)
);

BUFx3_ASAP7_75t_L g3572 ( 
.A(n_3330),
.Y(n_3572)
);

NAND2xp5_ASAP7_75t_L g3573 ( 
.A(n_3335),
.B(n_1379),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3360),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_2941),
.B(n_1384),
.Y(n_3575)
);

NOR2xp33_ASAP7_75t_L g3576 ( 
.A(n_3034),
.B(n_1384),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_SL g3577 ( 
.A(n_2892),
.B(n_1519),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_SL g3578 ( 
.A(n_3318),
.B(n_2925),
.Y(n_3578)
);

NOR2xp33_ASAP7_75t_L g3579 ( 
.A(n_2918),
.B(n_1403),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_L g3580 ( 
.A(n_3394),
.B(n_1403),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_SL g3581 ( 
.A(n_3318),
.B(n_1519),
.Y(n_3581)
);

NAND2xp5_ASAP7_75t_L g3582 ( 
.A(n_3394),
.B(n_3455),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3362),
.Y(n_3583)
);

AO22x2_ASAP7_75t_L g3584 ( 
.A1(n_3270),
.A2(n_1530),
.B1(n_1545),
.B2(n_1440),
.Y(n_3584)
);

INVx1_ASAP7_75t_L g3585 ( 
.A(n_3363),
.Y(n_3585)
);

NAND2xp5_ASAP7_75t_SL g3586 ( 
.A(n_3026),
.B(n_1543),
.Y(n_3586)
);

AOI22xp5_ASAP7_75t_L g3587 ( 
.A1(n_2938),
.A2(n_1530),
.B1(n_1545),
.B2(n_1440),
.Y(n_3587)
);

NAND2xp5_ASAP7_75t_L g3588 ( 
.A(n_3455),
.B(n_1559),
.Y(n_3588)
);

NOR2xp67_ASAP7_75t_L g3589 ( 
.A(n_2814),
.B(n_45),
.Y(n_3589)
);

INVx2_ASAP7_75t_L g3590 ( 
.A(n_2809),
.Y(n_3590)
);

AND2x4_ASAP7_75t_L g3591 ( 
.A(n_3189),
.B(n_1559),
.Y(n_3591)
);

NOR2xp67_ASAP7_75t_L g3592 ( 
.A(n_2814),
.B(n_46),
.Y(n_3592)
);

NOR2xp33_ASAP7_75t_L g3593 ( 
.A(n_3160),
.B(n_1602),
.Y(n_3593)
);

NAND2xp5_ASAP7_75t_L g3594 ( 
.A(n_2936),
.B(n_1602),
.Y(n_3594)
);

NAND2xp5_ASAP7_75t_L g3595 ( 
.A(n_3159),
.B(n_1639),
.Y(n_3595)
);

NOR2xp33_ASAP7_75t_L g3596 ( 
.A(n_3124),
.B(n_1639),
.Y(n_3596)
);

INVx1_ASAP7_75t_L g3597 ( 
.A(n_3367),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_2928),
.B(n_1643),
.Y(n_3598)
);

NAND2xp5_ASAP7_75t_SL g3599 ( 
.A(n_3026),
.B(n_1543),
.Y(n_3599)
);

INVx8_ASAP7_75t_L g3600 ( 
.A(n_3102),
.Y(n_3600)
);

INVx1_ASAP7_75t_L g3601 ( 
.A(n_3372),
.Y(n_3601)
);

AND2x2_ASAP7_75t_L g3602 ( 
.A(n_3435),
.B(n_1643),
.Y(n_3602)
);

NOR2xp33_ASAP7_75t_L g3603 ( 
.A(n_2883),
.B(n_2801),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3374),
.Y(n_3604)
);

INVx2_ASAP7_75t_L g3605 ( 
.A(n_3277),
.Y(n_3605)
);

AOI22xp33_ASAP7_75t_L g3606 ( 
.A1(n_3295),
.A2(n_1580),
.B1(n_1601),
.B2(n_1543),
.Y(n_3606)
);

AOI22xp5_ASAP7_75t_L g3607 ( 
.A1(n_2993),
.A2(n_1648),
.B1(n_1663),
.B2(n_1647),
.Y(n_3607)
);

NAND2xp5_ASAP7_75t_L g3608 ( 
.A(n_2802),
.B(n_1647),
.Y(n_3608)
);

NOR2xp33_ASAP7_75t_L g3609 ( 
.A(n_3320),
.B(n_3339),
.Y(n_3609)
);

INVx2_ASAP7_75t_L g3610 ( 
.A(n_3278),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_SL g3611 ( 
.A(n_3044),
.B(n_1543),
.Y(n_3611)
);

NAND2xp5_ASAP7_75t_SL g3612 ( 
.A(n_3044),
.B(n_3047),
.Y(n_3612)
);

INVx2_ASAP7_75t_SL g3613 ( 
.A(n_3289),
.Y(n_3613)
);

BUFx2_ASAP7_75t_L g3614 ( 
.A(n_2846),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3375),
.Y(n_3615)
);

INVx1_ASAP7_75t_L g3616 ( 
.A(n_3381),
.Y(n_3616)
);

BUFx3_ASAP7_75t_L g3617 ( 
.A(n_3336),
.Y(n_3617)
);

INVx2_ASAP7_75t_SL g3618 ( 
.A(n_3419),
.Y(n_3618)
);

INVx1_ASAP7_75t_L g3619 ( 
.A(n_3384),
.Y(n_3619)
);

INVx1_ASAP7_75t_L g3620 ( 
.A(n_2862),
.Y(n_3620)
);

AO22x2_ASAP7_75t_L g3621 ( 
.A1(n_3263),
.A2(n_1663),
.B1(n_1677),
.B2(n_1648),
.Y(n_3621)
);

NAND2xp5_ASAP7_75t_L g3622 ( 
.A(n_2802),
.B(n_1677),
.Y(n_3622)
);

INVx1_ASAP7_75t_L g3623 ( 
.A(n_2863),
.Y(n_3623)
);

NAND2xp33_ASAP7_75t_L g3624 ( 
.A(n_3004),
.B(n_1601),
.Y(n_3624)
);

AOI22xp33_ASAP7_75t_L g3625 ( 
.A1(n_3016),
.A2(n_1601),
.B1(n_1603),
.B2(n_1580),
.Y(n_3625)
);

NAND2xp5_ASAP7_75t_SL g3626 ( 
.A(n_3044),
.B(n_1580),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3047),
.B(n_1580),
.Y(n_3627)
);

NAND2xp5_ASAP7_75t_L g3628 ( 
.A(n_2807),
.B(n_1698),
.Y(n_3628)
);

NOR2xp67_ASAP7_75t_L g3629 ( 
.A(n_2815),
.B(n_46),
.Y(n_3629)
);

AOI22xp5_ASAP7_75t_L g3630 ( 
.A1(n_3004),
.A2(n_3081),
.B1(n_3413),
.B2(n_3410),
.Y(n_3630)
);

NAND2xp5_ASAP7_75t_L g3631 ( 
.A(n_2807),
.B(n_1703),
.Y(n_3631)
);

AOI21xp5_ASAP7_75t_L g3632 ( 
.A1(n_3148),
.A2(n_1703),
.B(n_1603),
.Y(n_3632)
);

NAND2xp5_ASAP7_75t_L g3633 ( 
.A(n_2810),
.B(n_46),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_2810),
.B(n_47),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_2864),
.Y(n_3635)
);

INVx2_ASAP7_75t_L g3636 ( 
.A(n_3329),
.Y(n_3636)
);

NOR2xp33_ASAP7_75t_L g3637 ( 
.A(n_2854),
.B(n_47),
.Y(n_3637)
);

NAND2xp5_ASAP7_75t_L g3638 ( 
.A(n_2817),
.B(n_3390),
.Y(n_3638)
);

NAND2xp5_ASAP7_75t_L g3639 ( 
.A(n_2817),
.B(n_48),
.Y(n_3639)
);

NAND2xp5_ASAP7_75t_SL g3640 ( 
.A(n_3047),
.B(n_1601),
.Y(n_3640)
);

HB1xp67_ASAP7_75t_L g3641 ( 
.A(n_2898),
.Y(n_3641)
);

INVx2_ASAP7_75t_L g3642 ( 
.A(n_3345),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_2872),
.Y(n_3643)
);

NOR2xp33_ASAP7_75t_L g3644 ( 
.A(n_3305),
.B(n_48),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3352),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_2879),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_L g3647 ( 
.A(n_3244),
.B(n_1645),
.C(n_1603),
.Y(n_3647)
);

NAND2xp5_ASAP7_75t_L g3648 ( 
.A(n_3390),
.B(n_49),
.Y(n_3648)
);

AOI22xp5_ASAP7_75t_L g3649 ( 
.A1(n_3004),
.A2(n_1645),
.B1(n_1708),
.B2(n_1603),
.Y(n_3649)
);

AND2x4_ASAP7_75t_L g3650 ( 
.A(n_3004),
.B(n_49),
.Y(n_3650)
);

NOR2xp33_ASAP7_75t_L g3651 ( 
.A(n_3313),
.B(n_49),
.Y(n_3651)
);

NOR2xp33_ASAP7_75t_L g3652 ( 
.A(n_3315),
.B(n_50),
.Y(n_3652)
);

NOR2xp33_ASAP7_75t_L g3653 ( 
.A(n_3402),
.B(n_50),
.Y(n_3653)
);

INVxp67_ASAP7_75t_SL g3654 ( 
.A(n_3433),
.Y(n_3654)
);

NOR2xp33_ASAP7_75t_L g3655 ( 
.A(n_3443),
.B(n_50),
.Y(n_3655)
);

NOR2xp33_ASAP7_75t_L g3656 ( 
.A(n_3306),
.B(n_51),
.Y(n_3656)
);

NAND2xp5_ASAP7_75t_L g3657 ( 
.A(n_3395),
.B(n_51),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3395),
.B(n_51),
.Y(n_3658)
);

NAND2xp5_ASAP7_75t_SL g3659 ( 
.A(n_2845),
.B(n_1645),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3081),
.A2(n_1708),
.B1(n_1711),
.B2(n_1645),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_2884),
.Y(n_3661)
);

NAND2xp5_ASAP7_75t_SL g3662 ( 
.A(n_3389),
.B(n_1708),
.Y(n_3662)
);

NAND2xp5_ASAP7_75t_L g3663 ( 
.A(n_3405),
.B(n_52),
.Y(n_3663)
);

AO22x1_ASAP7_75t_L g3664 ( 
.A1(n_3334),
.A2(n_1711),
.B1(n_1708),
.B2(n_1082),
.Y(n_3664)
);

NAND3xp33_ASAP7_75t_L g3665 ( 
.A(n_3414),
.B(n_1711),
.C(n_53),
.Y(n_3665)
);

AOI22xp33_ASAP7_75t_L g3666 ( 
.A1(n_2926),
.A2(n_1711),
.B1(n_53),
.B2(n_54),
.Y(n_3666)
);

INVx2_ASAP7_75t_L g3667 ( 
.A(n_3366),
.Y(n_3667)
);

INVx2_ASAP7_75t_L g3668 ( 
.A(n_3377),
.Y(n_3668)
);

NAND2x1_ASAP7_75t_L g3669 ( 
.A(n_3081),
.B(n_52),
.Y(n_3669)
);

NAND2xp5_ASAP7_75t_SL g3670 ( 
.A(n_3134),
.B(n_3267),
.Y(n_3670)
);

NOR2xp33_ASAP7_75t_L g3671 ( 
.A(n_2958),
.B(n_53),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3405),
.B(n_54),
.Y(n_3672)
);

NAND2xp5_ASAP7_75t_L g3673 ( 
.A(n_3459),
.B(n_55),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_2891),
.Y(n_3674)
);

NOR2xp33_ASAP7_75t_L g3675 ( 
.A(n_3213),
.B(n_55),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3459),
.B(n_55),
.Y(n_3676)
);

AND2x2_ASAP7_75t_L g3677 ( 
.A(n_3293),
.B(n_56),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_SL g3678 ( 
.A(n_3081),
.B(n_56),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_L g3679 ( 
.A(n_3407),
.B(n_56),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_2895),
.Y(n_3680)
);

INVxp67_ASAP7_75t_L g3681 ( 
.A(n_2875),
.Y(n_3681)
);

NAND2xp5_ASAP7_75t_L g3682 ( 
.A(n_3407),
.B(n_3415),
.Y(n_3682)
);

NAND2xp5_ASAP7_75t_L g3683 ( 
.A(n_3415),
.B(n_57),
.Y(n_3683)
);

INVx1_ASAP7_75t_L g3684 ( 
.A(n_2899),
.Y(n_3684)
);

INVxp67_ASAP7_75t_SL g3685 ( 
.A(n_3267),
.Y(n_3685)
);

NAND2xp5_ASAP7_75t_L g3686 ( 
.A(n_3421),
.B(n_57),
.Y(n_3686)
);

INVx2_ASAP7_75t_SL g3687 ( 
.A(n_3419),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3378),
.Y(n_3688)
);

NAND2xp5_ASAP7_75t_SL g3689 ( 
.A(n_3134),
.B(n_58),
.Y(n_3689)
);

AOI22xp33_ASAP7_75t_L g3690 ( 
.A1(n_2995),
.A2(n_59),
.B1(n_60),
.B2(n_58),
.Y(n_3690)
);

AOI22xp33_ASAP7_75t_L g3691 ( 
.A1(n_3441),
.A2(n_59),
.B1(n_60),
.B2(n_58),
.Y(n_3691)
);

A2O1A1Ixp33_ASAP7_75t_L g3692 ( 
.A1(n_3269),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3692)
);

INVx2_ASAP7_75t_SL g3693 ( 
.A(n_3089),
.Y(n_3693)
);

NAND2xp5_ASAP7_75t_L g3694 ( 
.A(n_3421),
.B(n_59),
.Y(n_3694)
);

INVx2_ASAP7_75t_L g3695 ( 
.A(n_3380),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3425),
.B(n_60),
.Y(n_3696)
);

NAND2xp5_ASAP7_75t_L g3697 ( 
.A(n_3425),
.B(n_61),
.Y(n_3697)
);

A2O1A1Ixp33_ASAP7_75t_L g3698 ( 
.A1(n_3269),
.A2(n_3),
.B(n_1),
.C(n_2),
.Y(n_3698)
);

NAND2xp5_ASAP7_75t_L g3699 ( 
.A(n_3427),
.B(n_61),
.Y(n_3699)
);

NAND2xp5_ASAP7_75t_SL g3700 ( 
.A(n_2811),
.B(n_62),
.Y(n_3700)
);

NAND2xp33_ASAP7_75t_L g3701 ( 
.A(n_2952),
.B(n_62),
.Y(n_3701)
);

NAND2xp5_ASAP7_75t_SL g3702 ( 
.A(n_2811),
.B(n_63),
.Y(n_3702)
);

NOR2xp33_ASAP7_75t_SL g3703 ( 
.A(n_2952),
.B(n_2959),
.Y(n_3703)
);

INVx2_ASAP7_75t_L g3704 ( 
.A(n_3385),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3392),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3427),
.B(n_63),
.Y(n_3706)
);

NAND2xp5_ASAP7_75t_L g3707 ( 
.A(n_3429),
.B(n_64),
.Y(n_3707)
);

INVx2_ASAP7_75t_L g3708 ( 
.A(n_3416),
.Y(n_3708)
);

NAND2xp5_ASAP7_75t_SL g3709 ( 
.A(n_2811),
.B(n_64),
.Y(n_3709)
);

NAND2xp5_ASAP7_75t_SL g3710 ( 
.A(n_2812),
.B(n_64),
.Y(n_3710)
);

OR2x2_ASAP7_75t_L g3711 ( 
.A(n_3288),
.B(n_66),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_L g3712 ( 
.A(n_3429),
.B(n_66),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_2903),
.Y(n_3713)
);

NAND2xp5_ASAP7_75t_SL g3714 ( 
.A(n_2812),
.B(n_66),
.Y(n_3714)
);

AOI22xp5_ASAP7_75t_L g3715 ( 
.A1(n_3446),
.A2(n_3448),
.B1(n_3456),
.B2(n_3452),
.Y(n_3715)
);

NOR2xp33_ASAP7_75t_L g3716 ( 
.A(n_2841),
.B(n_67),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_L g3717 ( 
.A(n_3430),
.B(n_67),
.Y(n_3717)
);

BUFx5_ASAP7_75t_L g3718 ( 
.A(n_2917),
.Y(n_3718)
);

INVxp67_ASAP7_75t_L g3719 ( 
.A(n_3301),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_2910),
.Y(n_3720)
);

INVx2_ASAP7_75t_SL g3721 ( 
.A(n_3089),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_L g3722 ( 
.A(n_3430),
.B(n_67),
.Y(n_3722)
);

NOR2xp33_ASAP7_75t_L g3723 ( 
.A(n_2948),
.B(n_68),
.Y(n_3723)
);

INVx2_ASAP7_75t_L g3724 ( 
.A(n_3422),
.Y(n_3724)
);

NAND2xp5_ASAP7_75t_L g3725 ( 
.A(n_3449),
.B(n_68),
.Y(n_3725)
);

OAI221xp5_ASAP7_75t_L g3726 ( 
.A1(n_3418),
.A2(n_70),
.B1(n_71),
.B2(n_69),
.C(n_68),
.Y(n_3726)
);

AND2x2_ASAP7_75t_L g3727 ( 
.A(n_3344),
.B(n_69),
.Y(n_3727)
);

OR2x6_ASAP7_75t_L g3728 ( 
.A(n_2815),
.B(n_69),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_2946),
.Y(n_3729)
);

NOR2xp33_ASAP7_75t_L g3730 ( 
.A(n_3274),
.B(n_70),
.Y(n_3730)
);

NAND2xp5_ASAP7_75t_L g3731 ( 
.A(n_3449),
.B(n_71),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_2950),
.Y(n_3732)
);

AOI22xp33_ASAP7_75t_L g3733 ( 
.A1(n_2932),
.A2(n_73),
.B1(n_74),
.B2(n_72),
.Y(n_3733)
);

NAND2xp5_ASAP7_75t_L g3734 ( 
.A(n_2851),
.B(n_72),
.Y(n_3734)
);

AND2x6_ASAP7_75t_L g3735 ( 
.A(n_2821),
.B(n_72),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_2857),
.B(n_74),
.Y(n_3736)
);

AND2x6_ASAP7_75t_SL g3737 ( 
.A(n_3224),
.B(n_75),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_2812),
.B(n_75),
.Y(n_3738)
);

NAND2xp5_ASAP7_75t_L g3739 ( 
.A(n_2969),
.B(n_75),
.Y(n_3739)
);

INVx2_ASAP7_75t_L g3740 ( 
.A(n_3424),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3438),
.Y(n_3741)
);

NAND2xp5_ASAP7_75t_L g3742 ( 
.A(n_2973),
.B(n_2978),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3440),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3373),
.B(n_76),
.Y(n_3744)
);

INVx2_ASAP7_75t_L g3745 ( 
.A(n_3444),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_2953),
.Y(n_3746)
);

BUFx3_ASAP7_75t_L g3747 ( 
.A(n_3376),
.Y(n_3747)
);

NAND2xp5_ASAP7_75t_L g3748 ( 
.A(n_2979),
.B(n_2896),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_2957),
.Y(n_3749)
);

BUFx8_ASAP7_75t_L g3750 ( 
.A(n_2933),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3126),
.Y(n_3751)
);

INVx2_ASAP7_75t_L g3752 ( 
.A(n_2982),
.Y(n_3752)
);

NOR2xp33_ASAP7_75t_L g3753 ( 
.A(n_3343),
.B(n_76),
.Y(n_3753)
);

NAND2xp5_ASAP7_75t_SL g3754 ( 
.A(n_3294),
.B(n_76),
.Y(n_3754)
);

NAND3xp33_ASAP7_75t_L g3755 ( 
.A(n_3224),
.B(n_78),
.C(n_77),
.Y(n_3755)
);

INVx2_ASAP7_75t_SL g3756 ( 
.A(n_3089),
.Y(n_3756)
);

NAND2xp5_ASAP7_75t_SL g3757 ( 
.A(n_3294),
.B(n_78),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_2896),
.B(n_79),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3059),
.B(n_79),
.Y(n_3759)
);

INVx1_ASAP7_75t_L g3760 ( 
.A(n_2960),
.Y(n_3760)
);

NOR2xp33_ASAP7_75t_L g3761 ( 
.A(n_3364),
.B(n_79),
.Y(n_3761)
);

NAND2xp5_ASAP7_75t_SL g3762 ( 
.A(n_3294),
.B(n_80),
.Y(n_3762)
);

NOR2x1p5_ASAP7_75t_L g3763 ( 
.A(n_3361),
.B(n_80),
.Y(n_3763)
);

INVx2_ASAP7_75t_SL g3764 ( 
.A(n_2887),
.Y(n_3764)
);

INVx2_ASAP7_75t_SL g3765 ( 
.A(n_2887),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3400),
.Y(n_3766)
);

OAI22xp5_ASAP7_75t_L g3767 ( 
.A1(n_3437),
.A2(n_81),
.B1(n_82),
.B2(n_80),
.Y(n_3767)
);

NAND3xp33_ASAP7_75t_L g3768 ( 
.A(n_3177),
.B(n_82),
.C(n_81),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3454),
.B(n_81),
.Y(n_3769)
);

INVx2_ASAP7_75t_L g3770 ( 
.A(n_3127),
.Y(n_3770)
);

INVx2_ASAP7_75t_L g3771 ( 
.A(n_3137),
.Y(n_3771)
);

NAND3xp33_ASAP7_75t_L g3772 ( 
.A(n_3183),
.B(n_83),
.C(n_82),
.Y(n_3772)
);

INVx2_ASAP7_75t_SL g3773 ( 
.A(n_3408),
.Y(n_3773)
);

NAND2xp5_ASAP7_75t_SL g3774 ( 
.A(n_3304),
.B(n_83),
.Y(n_3774)
);

INVx2_ASAP7_75t_L g3775 ( 
.A(n_3143),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_2821),
.B(n_84),
.Y(n_3776)
);

BUFx6f_ASAP7_75t_L g3777 ( 
.A(n_2834),
.Y(n_3777)
);

BUFx12f_ASAP7_75t_SL g3778 ( 
.A(n_3281),
.Y(n_3778)
);

INVx2_ASAP7_75t_L g3779 ( 
.A(n_3144),
.Y(n_3779)
);

NAND2xp5_ASAP7_75t_L g3780 ( 
.A(n_2822),
.B(n_84),
.Y(n_3780)
);

INVx2_ASAP7_75t_L g3781 ( 
.A(n_3147),
.Y(n_3781)
);

NAND2xp5_ASAP7_75t_L g3782 ( 
.A(n_2822),
.B(n_85),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_2961),
.Y(n_3783)
);

INVx2_ASAP7_75t_L g3784 ( 
.A(n_3152),
.Y(n_3784)
);

OAI22xp33_ASAP7_75t_L g3785 ( 
.A1(n_3126),
.A2(n_86),
.B1(n_87),
.B2(n_85),
.Y(n_3785)
);

NAND2xp5_ASAP7_75t_L g3786 ( 
.A(n_2825),
.B(n_86),
.Y(n_3786)
);

INVx3_ASAP7_75t_L g3787 ( 
.A(n_2947),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3398),
.B(n_86),
.Y(n_3788)
);

INVx2_ASAP7_75t_L g3789 ( 
.A(n_3154),
.Y(n_3789)
);

NAND2xp33_ASAP7_75t_L g3790 ( 
.A(n_2952),
.B(n_87),
.Y(n_3790)
);

NOR3xp33_ASAP7_75t_L g3791 ( 
.A(n_3387),
.B(n_88),
.C(n_87),
.Y(n_3791)
);

BUFx6f_ASAP7_75t_L g3792 ( 
.A(n_2866),
.Y(n_3792)
);

NAND2xp33_ASAP7_75t_SL g3793 ( 
.A(n_2848),
.B(n_88),
.Y(n_3793)
);

INVx2_ASAP7_75t_L g3794 ( 
.A(n_2825),
.Y(n_3794)
);

INVx1_ASAP7_75t_L g3795 ( 
.A(n_3138),
.Y(n_3795)
);

NAND2xp5_ASAP7_75t_SL g3796 ( 
.A(n_3304),
.B(n_89),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3452),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3186),
.Y(n_3798)
);

O2A1O1Ixp5_ASAP7_75t_L g3799 ( 
.A1(n_3275),
.A2(n_90),
.B(n_91),
.C(n_89),
.Y(n_3799)
);

NAND2xp5_ASAP7_75t_L g3800 ( 
.A(n_2827),
.B(n_89),
.Y(n_3800)
);

NAND2x1p5_ASAP7_75t_L g3801 ( 
.A(n_2994),
.B(n_2904),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_SL g3802 ( 
.A(n_3304),
.B(n_90),
.Y(n_3802)
);

INVx1_ASAP7_75t_L g3803 ( 
.A(n_3202),
.Y(n_3803)
);

INVx4_ASAP7_75t_L g3804 ( 
.A(n_3281),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_2827),
.Y(n_3805)
);

O2A1O1Ixp5_ASAP7_75t_L g3806 ( 
.A1(n_3275),
.A2(n_92),
.B(n_93),
.C(n_91),
.Y(n_3806)
);

AND2x4_ASAP7_75t_L g3807 ( 
.A(n_2904),
.B(n_91),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_2830),
.B(n_92),
.Y(n_3808)
);

NOR2xp33_ASAP7_75t_L g3809 ( 
.A(n_2912),
.B(n_92),
.Y(n_3809)
);

AOI21xp5_ASAP7_75t_L g3810 ( 
.A1(n_3070),
.A2(n_94),
.B(n_93),
.Y(n_3810)
);

AOI22xp5_ASAP7_75t_L g3811 ( 
.A1(n_2798),
.A2(n_1074),
.B1(n_1075),
.B2(n_1073),
.Y(n_3811)
);

INVx2_ASAP7_75t_L g3812 ( 
.A(n_2830),
.Y(n_3812)
);

NAND2xp5_ASAP7_75t_SL g3813 ( 
.A(n_3357),
.B(n_93),
.Y(n_3813)
);

INVx4_ASAP7_75t_L g3814 ( 
.A(n_3296),
.Y(n_3814)
);

AOI22xp33_ASAP7_75t_L g3815 ( 
.A1(n_3056),
.A2(n_95),
.B1(n_96),
.B2(n_94),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_2831),
.B(n_2832),
.Y(n_3816)
);

NAND2xp5_ASAP7_75t_L g3817 ( 
.A(n_2831),
.B(n_94),
.Y(n_3817)
);

INVxp33_ASAP7_75t_SL g3818 ( 
.A(n_3011),
.Y(n_3818)
);

HB1xp67_ASAP7_75t_L g3819 ( 
.A(n_3018),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_2832),
.B(n_96),
.Y(n_3820)
);

NAND2xp5_ASAP7_75t_L g3821 ( 
.A(n_2837),
.B(n_97),
.Y(n_3821)
);

INVxp33_ASAP7_75t_L g3822 ( 
.A(n_3178),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_2984),
.Y(n_3823)
);

NOR2xp33_ASAP7_75t_L g3824 ( 
.A(n_2954),
.B(n_97),
.Y(n_3824)
);

NOR2xp33_ASAP7_75t_L g3825 ( 
.A(n_3027),
.B(n_97),
.Y(n_3825)
);

INVx2_ASAP7_75t_L g3826 ( 
.A(n_2837),
.Y(n_3826)
);

NAND2xp5_ASAP7_75t_L g3827 ( 
.A(n_2839),
.B(n_98),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_2987),
.Y(n_3828)
);

NOR2xp67_ASAP7_75t_L g3829 ( 
.A(n_3296),
.B(n_98),
.Y(n_3829)
);

AOI21xp5_ASAP7_75t_L g3830 ( 
.A1(n_3199),
.A2(n_100),
.B(n_99),
.Y(n_3830)
);

NAND2xp33_ASAP7_75t_L g3831 ( 
.A(n_2952),
.B(n_99),
.Y(n_3831)
);

INVx2_ASAP7_75t_L g3832 ( 
.A(n_2839),
.Y(n_3832)
);

NAND2xp5_ASAP7_75t_L g3833 ( 
.A(n_2844),
.B(n_99),
.Y(n_3833)
);

O2A1O1Ixp33_ASAP7_75t_L g3834 ( 
.A1(n_3169),
.A2(n_101),
.B(n_102),
.C(n_100),
.Y(n_3834)
);

NOR2xp33_ASAP7_75t_L g3835 ( 
.A(n_3052),
.B(n_100),
.Y(n_3835)
);

NAND2xp5_ASAP7_75t_L g3836 ( 
.A(n_2844),
.B(n_101),
.Y(n_3836)
);

CKINVDCx20_ASAP7_75t_R g3837 ( 
.A(n_3379),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_2935),
.B(n_101),
.Y(n_3838)
);

AOI22xp5_ASAP7_75t_L g3839 ( 
.A1(n_3196),
.A2(n_1082),
.B1(n_103),
.B2(n_104),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3214),
.Y(n_3840)
);

NAND2xp5_ASAP7_75t_L g3841 ( 
.A(n_2935),
.B(n_102),
.Y(n_3841)
);

OAI22xp5_ASAP7_75t_L g3842 ( 
.A1(n_2939),
.A2(n_2943),
.B1(n_3196),
.B2(n_3397),
.Y(n_3842)
);

INVx2_ASAP7_75t_L g3843 ( 
.A(n_2939),
.Y(n_3843)
);

INVx4_ASAP7_75t_L g3844 ( 
.A(n_3327),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3426),
.A2(n_1082),
.B1(n_103),
.B2(n_104),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3357),
.B(n_102),
.Y(n_3846)
);

NAND2xp5_ASAP7_75t_SL g3847 ( 
.A(n_3357),
.B(n_103),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_2943),
.B(n_104),
.Y(n_3848)
);

INVx2_ASAP7_75t_L g3849 ( 
.A(n_2855),
.Y(n_3849)
);

AND2x2_ASAP7_75t_L g3850 ( 
.A(n_2897),
.B(n_105),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_SL g3851 ( 
.A(n_3369),
.B(n_105),
.Y(n_3851)
);

NAND2xp5_ASAP7_75t_L g3852 ( 
.A(n_2966),
.B(n_106),
.Y(n_3852)
);

INVx1_ASAP7_75t_L g3853 ( 
.A(n_3215),
.Y(n_3853)
);

NAND2xp5_ASAP7_75t_SL g3854 ( 
.A(n_3369),
.B(n_106),
.Y(n_3854)
);

NOR2xp33_ASAP7_75t_L g3855 ( 
.A(n_2865),
.B(n_2890),
.Y(n_3855)
);

BUFx3_ASAP7_75t_L g3856 ( 
.A(n_3412),
.Y(n_3856)
);

INVx2_ASAP7_75t_L g3857 ( 
.A(n_2858),
.Y(n_3857)
);

INVx8_ASAP7_75t_L g3858 ( 
.A(n_2994),
.Y(n_3858)
);

NOR2x1_ASAP7_75t_L g3859 ( 
.A(n_3327),
.B(n_1070),
.Y(n_3859)
);

OR2x2_ASAP7_75t_L g3860 ( 
.A(n_3326),
.B(n_106),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_2966),
.B(n_107),
.Y(n_3861)
);

NAND2xp5_ASAP7_75t_L g3862 ( 
.A(n_2914),
.B(n_2915),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3218),
.Y(n_3863)
);

O2A1O1Ixp33_ASAP7_75t_L g3864 ( 
.A1(n_3206),
.A2(n_108),
.B(n_109),
.C(n_107),
.Y(n_3864)
);

NAND2xp5_ASAP7_75t_SL g3865 ( 
.A(n_3369),
.B(n_107),
.Y(n_3865)
);

AND2x2_ASAP7_75t_L g3866 ( 
.A(n_3163),
.B(n_108),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_2859),
.Y(n_3867)
);

NAND2xp33_ASAP7_75t_L g3868 ( 
.A(n_2959),
.B(n_110),
.Y(n_3868)
);

NOR2xp33_ASAP7_75t_L g3869 ( 
.A(n_3355),
.B(n_110),
.Y(n_3869)
);

AND2x4_ASAP7_75t_L g3870 ( 
.A(n_2994),
.B(n_111),
.Y(n_3870)
);

INVx2_ASAP7_75t_L g3871 ( 
.A(n_2873),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3079),
.Y(n_3872)
);

NAND2xp5_ASAP7_75t_L g3873 ( 
.A(n_2914),
.B(n_111),
.Y(n_3873)
);

NAND2xp33_ASAP7_75t_L g3874 ( 
.A(n_2959),
.B(n_112),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_2915),
.B(n_112),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_2901),
.Y(n_3876)
);

NAND2xp5_ASAP7_75t_SL g3877 ( 
.A(n_3393),
.B(n_113),
.Y(n_3877)
);

NOR2xp33_ASAP7_75t_L g3878 ( 
.A(n_2836),
.B(n_113),
.Y(n_3878)
);

INVx1_ASAP7_75t_SL g3879 ( 
.A(n_2955),
.Y(n_3879)
);

AOI22xp5_ASAP7_75t_L g3880 ( 
.A1(n_3227),
.A2(n_1079),
.B1(n_1080),
.B2(n_1078),
.Y(n_3880)
);

INVx2_ASAP7_75t_L g3881 ( 
.A(n_2907),
.Y(n_3881)
);

INVx2_ASAP7_75t_L g3882 ( 
.A(n_2911),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3079),
.Y(n_3883)
);

INVx2_ASAP7_75t_L g3884 ( 
.A(n_2913),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_L g3885 ( 
.A(n_2930),
.B(n_114),
.Y(n_3885)
);

INVx1_ASAP7_75t_L g3886 ( 
.A(n_3080),
.Y(n_3886)
);

INVxp67_ASAP7_75t_SL g3887 ( 
.A(n_2955),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_L g3888 ( 
.A(n_2930),
.B(n_114),
.Y(n_3888)
);

NOR2xp33_ASAP7_75t_L g3889 ( 
.A(n_3173),
.B(n_114),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_L g3890 ( 
.A(n_2874),
.B(n_2927),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_L g3891 ( 
.A(n_3166),
.B(n_115),
.Y(n_3891)
);

NOR2x1p5_ASAP7_75t_L g3892 ( 
.A(n_3399),
.B(n_115),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3393),
.B(n_115),
.Y(n_3893)
);

NAND2x1_ASAP7_75t_L g3894 ( 
.A(n_3371),
.B(n_116),
.Y(n_3894)
);

NAND2xp5_ASAP7_75t_L g3895 ( 
.A(n_3193),
.B(n_116),
.Y(n_3895)
);

INVxp67_ASAP7_75t_L g3896 ( 
.A(n_3106),
.Y(n_3896)
);

AND2x4_ASAP7_75t_SL g3897 ( 
.A(n_3342),
.B(n_116),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_2920),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_2924),
.Y(n_3899)
);

NOR2xp33_ASAP7_75t_L g3900 ( 
.A(n_3173),
.B(n_117),
.Y(n_3900)
);

OR2x2_ASAP7_75t_L g3901 ( 
.A(n_3175),
.B(n_117),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3080),
.Y(n_3902)
);

BUFx3_ASAP7_75t_L g3903 ( 
.A(n_3450),
.Y(n_3903)
);

INVx2_ASAP7_75t_L g3904 ( 
.A(n_2937),
.Y(n_3904)
);

NOR2xp33_ASAP7_75t_L g3905 ( 
.A(n_3135),
.B(n_118),
.Y(n_3905)
);

INVx2_ASAP7_75t_L g3906 ( 
.A(n_2964),
.Y(n_3906)
);

NAND2xp5_ASAP7_75t_L g3907 ( 
.A(n_2805),
.B(n_118),
.Y(n_3907)
);

AOI22xp33_ASAP7_75t_L g3908 ( 
.A1(n_3208),
.A2(n_119),
.B1(n_120),
.B2(n_118),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3057),
.A2(n_120),
.B1(n_121),
.B2(n_119),
.Y(n_3909)
);

INVx2_ASAP7_75t_L g3910 ( 
.A(n_2985),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_3393),
.B(n_120),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_L g3912 ( 
.A(n_2813),
.B(n_121),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_L g3913 ( 
.A(n_2828),
.B(n_122),
.Y(n_3913)
);

NAND2xp5_ASAP7_75t_L g3914 ( 
.A(n_3287),
.B(n_122),
.Y(n_3914)
);

INVx2_ASAP7_75t_L g3915 ( 
.A(n_3002),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_L g3916 ( 
.A(n_3299),
.B(n_122),
.Y(n_3916)
);

INVx2_ASAP7_75t_SL g3917 ( 
.A(n_3049),
.Y(n_3917)
);

INVxp67_ASAP7_75t_L g3918 ( 
.A(n_2967),
.Y(n_3918)
);

INVx2_ASAP7_75t_L g3919 ( 
.A(n_3051),
.Y(n_3919)
);

INVx2_ASAP7_75t_L g3920 ( 
.A(n_3063),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_SL g3921 ( 
.A(n_3409),
.B(n_123),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_3409),
.B(n_3445),
.Y(n_3922)
);

NOR2xp33_ASAP7_75t_L g3923 ( 
.A(n_3190),
.B(n_124),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3409),
.B(n_124),
.Y(n_3924)
);

NOR2xp33_ASAP7_75t_L g3925 ( 
.A(n_3201),
.B(n_124),
.Y(n_3925)
);

INVx2_ASAP7_75t_L g3926 ( 
.A(n_3086),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_3445),
.B(n_125),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_2980),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3309),
.B(n_125),
.Y(n_3929)
);

NAND2xp5_ASAP7_75t_L g3930 ( 
.A(n_3310),
.B(n_3311),
.Y(n_3930)
);

BUFx6f_ASAP7_75t_L g3931 ( 
.A(n_2866),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_L g3932 ( 
.A(n_3314),
.B(n_125),
.Y(n_3932)
);

NOR2xp33_ASAP7_75t_L g3933 ( 
.A(n_3211),
.B(n_126),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_L g3934 ( 
.A(n_3316),
.B(n_126),
.Y(n_3934)
);

INVx2_ASAP7_75t_L g3935 ( 
.A(n_3108),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_L g3936 ( 
.A(n_3319),
.B(n_126),
.Y(n_3936)
);

AOI22x1_ASAP7_75t_SL g3937 ( 
.A1(n_3420),
.A2(n_128),
.B1(n_129),
.B2(n_127),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_SL g3938 ( 
.A(n_3445),
.B(n_127),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3447),
.B(n_127),
.Y(n_3939)
);

NAND2xp5_ASAP7_75t_SL g3940 ( 
.A(n_3447),
.B(n_128),
.Y(n_3940)
);

CKINVDCx16_ASAP7_75t_R g3941 ( 
.A(n_3101),
.Y(n_3941)
);

NOR2xp33_ASAP7_75t_L g3942 ( 
.A(n_3211),
.B(n_129),
.Y(n_3942)
);

HB1xp67_ASAP7_75t_L g3943 ( 
.A(n_3018),
.Y(n_3943)
);

OAI22xp5_ASAP7_75t_L g3944 ( 
.A1(n_3403),
.A2(n_130),
.B1(n_131),
.B2(n_129),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3014),
.Y(n_3945)
);

NOR3xp33_ASAP7_75t_L g3946 ( 
.A(n_3307),
.B(n_131),
.C(n_130),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3331),
.B(n_131),
.Y(n_3947)
);

AOI22xp5_ASAP7_75t_L g3948 ( 
.A1(n_3000),
.A2(n_1081),
.B1(n_1080),
.B2(n_133),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_L g3949 ( 
.A(n_3333),
.B(n_132),
.Y(n_3949)
);

INVx2_ASAP7_75t_L g3950 ( 
.A(n_3120),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3220),
.Y(n_3951)
);

NAND2xp5_ASAP7_75t_L g3952 ( 
.A(n_3351),
.B(n_132),
.Y(n_3952)
);

INVx1_ASAP7_75t_L g3953 ( 
.A(n_2997),
.Y(n_3953)
);

INVx2_ASAP7_75t_SL g3954 ( 
.A(n_3049),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_2999),
.Y(n_3955)
);

NOR2xp67_ASAP7_75t_SL g3956 ( 
.A(n_2992),
.B(n_132),
.Y(n_3956)
);

INVx2_ASAP7_75t_L g3957 ( 
.A(n_3122),
.Y(n_3957)
);

NOR2xp33_ASAP7_75t_L g3958 ( 
.A(n_2840),
.B(n_133),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_L g3959 ( 
.A(n_3382),
.B(n_134),
.Y(n_3959)
);

INVx1_ASAP7_75t_L g3960 ( 
.A(n_3088),
.Y(n_3960)
);

INVx2_ASAP7_75t_L g3961 ( 
.A(n_3123),
.Y(n_3961)
);

NAND2xp5_ASAP7_75t_SL g3962 ( 
.A(n_3447),
.B(n_134),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3165),
.Y(n_3963)
);

AOI221xp5_ASAP7_75t_L g3964 ( 
.A1(n_3386),
.A2(n_136),
.B1(n_137),
.B2(n_135),
.C(n_134),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_L g3965 ( 
.A(n_2894),
.B(n_135),
.Y(n_3965)
);

BUFx6f_ASAP7_75t_L g3966 ( 
.A(n_2866),
.Y(n_3966)
);

INVx1_ASAP7_75t_L g3967 ( 
.A(n_3091),
.Y(n_3967)
);

NOR2xp33_ASAP7_75t_SL g3968 ( 
.A(n_2959),
.B(n_135),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_2894),
.B(n_136),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_L g3970 ( 
.A(n_3423),
.B(n_137),
.Y(n_3970)
);

NAND2xp5_ASAP7_75t_L g3971 ( 
.A(n_3428),
.B(n_3451),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_SL g3972 ( 
.A(n_3458),
.B(n_137),
.Y(n_3972)
);

NAND2xp5_ASAP7_75t_L g3973 ( 
.A(n_3453),
.B(n_138),
.Y(n_3973)
);

INVx2_ASAP7_75t_SL g3974 ( 
.A(n_3342),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_2956),
.B(n_138),
.Y(n_3975)
);

INVx4_ASAP7_75t_L g3976 ( 
.A(n_3439),
.Y(n_3976)
);

HB1xp67_ASAP7_75t_L g3977 ( 
.A(n_2889),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_L g3978 ( 
.A(n_3083),
.B(n_139),
.Y(n_3978)
);

NOR2xp33_ASAP7_75t_L g3979 ( 
.A(n_2833),
.B(n_139),
.Y(n_3979)
);

AND2x2_ASAP7_75t_L g3980 ( 
.A(n_3085),
.B(n_140),
.Y(n_3980)
);

BUFx3_ASAP7_75t_L g3981 ( 
.A(n_2905),
.Y(n_3981)
);

OR2x2_ASAP7_75t_L g3982 ( 
.A(n_3180),
.B(n_140),
.Y(n_3982)
);

AO221x1_ASAP7_75t_L g3983 ( 
.A1(n_3067),
.A2(n_142),
.B1(n_143),
.B2(n_141),
.C(n_140),
.Y(n_3983)
);

AND2x2_ASAP7_75t_L g3984 ( 
.A(n_3180),
.B(n_141),
.Y(n_3984)
);

NAND2xp5_ASAP7_75t_L g3985 ( 
.A(n_3130),
.B(n_142),
.Y(n_3985)
);

NAND2xp5_ASAP7_75t_L g3986 ( 
.A(n_3130),
.B(n_142),
.Y(n_3986)
);

INVx1_ASAP7_75t_L g3987 ( 
.A(n_3093),
.Y(n_3987)
);

OAI22xp33_ASAP7_75t_L g3988 ( 
.A1(n_2893),
.A2(n_144),
.B1(n_145),
.B2(n_143),
.Y(n_3988)
);

CKINVDCx5p33_ASAP7_75t_R g3989 ( 
.A(n_2808),
.Y(n_3989)
);

NAND2xp5_ASAP7_75t_SL g3990 ( 
.A(n_3458),
.B(n_144),
.Y(n_3990)
);

BUFx6f_ASAP7_75t_L g3991 ( 
.A(n_2931),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3096),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_L g3993 ( 
.A(n_3131),
.B(n_3040),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_L g3994 ( 
.A(n_3131),
.B(n_145),
.Y(n_3994)
);

NAND2xp5_ASAP7_75t_L g3995 ( 
.A(n_3140),
.B(n_146),
.Y(n_3995)
);

AOI22xp33_ASAP7_75t_L g3996 ( 
.A1(n_3057),
.A2(n_147),
.B1(n_148),
.B2(n_146),
.Y(n_3996)
);

INVxp67_ASAP7_75t_L g3997 ( 
.A(n_2945),
.Y(n_3997)
);

INVx2_ASAP7_75t_L g3998 ( 
.A(n_3167),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3097),
.Y(n_3999)
);

NOR2xp33_ASAP7_75t_L g4000 ( 
.A(n_3341),
.B(n_147),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3458),
.B(n_2860),
.Y(n_4001)
);

INVx1_ASAP7_75t_L g4002 ( 
.A(n_3107),
.Y(n_4002)
);

NOR2xp33_ASAP7_75t_L g4003 ( 
.A(n_3200),
.B(n_149),
.Y(n_4003)
);

NAND2xp5_ASAP7_75t_L g4004 ( 
.A(n_3072),
.B(n_149),
.Y(n_4004)
);

AOI21xp5_ASAP7_75t_L g4005 ( 
.A1(n_2868),
.A2(n_151),
.B(n_150),
.Y(n_4005)
);

NOR2xp33_ASAP7_75t_L g4006 ( 
.A(n_3030),
.B(n_150),
.Y(n_4006)
);

NOR3xp33_ASAP7_75t_L g4007 ( 
.A(n_3396),
.B(n_152),
.C(n_150),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_L g4008 ( 
.A(n_3233),
.B(n_152),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_2867),
.B(n_2947),
.Y(n_4009)
);

INVx2_ASAP7_75t_L g4010 ( 
.A(n_3109),
.Y(n_4010)
);

AOI22xp33_ASAP7_75t_SL g4011 ( 
.A1(n_3067),
.A2(n_153),
.B1(n_154),
.B2(n_152),
.Y(n_4011)
);

AOI22xp33_ASAP7_75t_L g4012 ( 
.A1(n_3250),
.A2(n_154),
.B1(n_155),
.B2(n_153),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_L g4013 ( 
.A(n_2909),
.B(n_153),
.Y(n_4013)
);

NAND3xp33_ASAP7_75t_L g4014 ( 
.A(n_3271),
.B(n_156),
.C(n_155),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_L g4015 ( 
.A(n_3302),
.B(n_156),
.Y(n_4015)
);

INVx1_ASAP7_75t_L g4016 ( 
.A(n_3110),
.Y(n_4016)
);

NOR2xp67_ASAP7_75t_L g4017 ( 
.A(n_3439),
.B(n_156),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3111),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3116),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3117),
.Y(n_4020)
);

NAND2xp5_ASAP7_75t_L g4021 ( 
.A(n_3184),
.B(n_157),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_L g4022 ( 
.A(n_3100),
.B(n_157),
.Y(n_4022)
);

INVx1_ASAP7_75t_SL g4023 ( 
.A(n_2955),
.Y(n_4023)
);

INVx1_ASAP7_75t_L g4024 ( 
.A(n_3136),
.Y(n_4024)
);

AOI22xp5_ASAP7_75t_L g4025 ( 
.A1(n_3252),
.A2(n_1074),
.B1(n_1075),
.B2(n_1073),
.Y(n_4025)
);

AND2x2_ASAP7_75t_L g4026 ( 
.A(n_3203),
.B(n_157),
.Y(n_4026)
);

INVxp67_ASAP7_75t_L g4027 ( 
.A(n_2886),
.Y(n_4027)
);

INVx1_ASAP7_75t_L g4028 ( 
.A(n_3156),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3235),
.Y(n_4029)
);

NOR2xp33_ASAP7_75t_L g4030 ( 
.A(n_3115),
.B(n_158),
.Y(n_4030)
);

AO221x1_ASAP7_75t_L g4031 ( 
.A1(n_2947),
.A2(n_160),
.B1(n_161),
.B2(n_159),
.C(n_158),
.Y(n_4031)
);

OAI22xp33_ASAP7_75t_SL g4032 ( 
.A1(n_3434),
.A2(n_160),
.B1(n_161),
.B2(n_159),
.Y(n_4032)
);

NAND2xp5_ASAP7_75t_L g4033 ( 
.A(n_3104),
.B(n_159),
.Y(n_4033)
);

O2A1O1Ixp33_ASAP7_75t_L g4034 ( 
.A1(n_3071),
.A2(n_3074),
.B(n_3132),
.C(n_3112),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_L g4035 ( 
.A(n_3128),
.B(n_160),
.Y(n_4035)
);

INVx2_ASAP7_75t_SL g4036 ( 
.A(n_3465),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_L g4037 ( 
.A(n_3715),
.B(n_3170),
.Y(n_4037)
);

INVx1_ASAP7_75t_L g4038 ( 
.A(n_3620),
.Y(n_4038)
);

INVx2_ASAP7_75t_SL g4039 ( 
.A(n_3465),
.Y(n_4039)
);

NOR2xp33_ASAP7_75t_L g4040 ( 
.A(n_3552),
.B(n_3918),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_L g4041 ( 
.A(n_3715),
.B(n_3252),
.Y(n_4041)
);

NAND2x1p5_ASAP7_75t_L g4042 ( 
.A(n_3804),
.B(n_3098),
.Y(n_4042)
);

INVx1_ASAP7_75t_L g4043 ( 
.A(n_3623),
.Y(n_4043)
);

OAI22xp5_ASAP7_75t_L g4044 ( 
.A1(n_3630),
.A2(n_2838),
.B1(n_3358),
.B2(n_2842),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3467),
.Y(n_4045)
);

CKINVDCx5p33_ASAP7_75t_R g4046 ( 
.A(n_3514),
.Y(n_4046)
);

INVx2_ASAP7_75t_L g4047 ( 
.A(n_3483),
.Y(n_4047)
);

INVx2_ASAP7_75t_L g4048 ( 
.A(n_3489),
.Y(n_4048)
);

NOR2xp33_ASAP7_75t_L g4049 ( 
.A(n_4027),
.B(n_3149),
.Y(n_4049)
);

INVx1_ASAP7_75t_L g4050 ( 
.A(n_3475),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_3493),
.Y(n_4051)
);

NOR2xp33_ASAP7_75t_L g4052 ( 
.A(n_3997),
.B(n_2970),
.Y(n_4052)
);

AND2x2_ASAP7_75t_L g4053 ( 
.A(n_3677),
.B(n_2975),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3727),
.B(n_2975),
.Y(n_4054)
);

NAND2xp5_ASAP7_75t_SL g4055 ( 
.A(n_3484),
.B(n_2867),
.Y(n_4055)
);

NOR2xp33_ASAP7_75t_L g4056 ( 
.A(n_3719),
.B(n_2986),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3480),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3509),
.Y(n_4058)
);

INVx2_ASAP7_75t_SL g4059 ( 
.A(n_3465),
.Y(n_4059)
);

NAND2xp5_ASAP7_75t_L g4060 ( 
.A(n_3928),
.B(n_3945),
.Y(n_4060)
);

INVx1_ASAP7_75t_L g4061 ( 
.A(n_3487),
.Y(n_4061)
);

OAI22xp5_ASAP7_75t_L g4062 ( 
.A1(n_3630),
.A2(n_3370),
.B1(n_3442),
.B2(n_2852),
.Y(n_4062)
);

NAND2xp5_ASAP7_75t_SL g4063 ( 
.A(n_3484),
.B(n_3101),
.Y(n_4063)
);

AND2x2_ASAP7_75t_L g4064 ( 
.A(n_3744),
.B(n_3114),
.Y(n_4064)
);

AOI21xp5_ASAP7_75t_L g4065 ( 
.A1(n_3491),
.A2(n_2923),
.B(n_2931),
.Y(n_4065)
);

NAND2xp5_ASAP7_75t_L g4066 ( 
.A(n_3500),
.B(n_3028),
.Y(n_4066)
);

NAND2xp5_ASAP7_75t_L g4067 ( 
.A(n_3579),
.B(n_3046),
.Y(n_4067)
);

AOI22xp5_ASAP7_75t_L g4068 ( 
.A1(n_3495),
.A2(n_3264),
.B1(n_3232),
.B2(n_3255),
.Y(n_4068)
);

INVx3_ASAP7_75t_L g4069 ( 
.A(n_3858),
.Y(n_4069)
);

INVx1_ASAP7_75t_L g4070 ( 
.A(n_3531),
.Y(n_4070)
);

OAI22xp5_ASAP7_75t_L g4071 ( 
.A1(n_3507),
.A2(n_3113),
.B1(n_3035),
.B2(n_2949),
.Y(n_4071)
);

INVx1_ASAP7_75t_SL g4072 ( 
.A(n_3981),
.Y(n_4072)
);

BUFx6f_ASAP7_75t_L g4073 ( 
.A(n_3858),
.Y(n_4073)
);

INVx3_ASAP7_75t_L g4074 ( 
.A(n_3858),
.Y(n_4074)
);

INVx5_ASAP7_75t_L g4075 ( 
.A(n_3600),
.Y(n_4075)
);

INVx3_ASAP7_75t_L g4076 ( 
.A(n_3801),
.Y(n_4076)
);

INVx2_ASAP7_75t_SL g4077 ( 
.A(n_3600),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3678),
.B(n_3113),
.Y(n_4078)
);

BUFx3_ASAP7_75t_L g4079 ( 
.A(n_3600),
.Y(n_4079)
);

INVx3_ASAP7_75t_L g4080 ( 
.A(n_3801),
.Y(n_4080)
);

OR2x2_ASAP7_75t_L g4081 ( 
.A(n_3582),
.B(n_3614),
.Y(n_4081)
);

BUFx2_ASAP7_75t_L g4082 ( 
.A(n_3557),
.Y(n_4082)
);

NOR3xp33_ASAP7_75t_SL g4083 ( 
.A(n_3561),
.B(n_2882),
.C(n_2877),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_L g4084 ( 
.A(n_3520),
.B(n_3090),
.Y(n_4084)
);

NAND2xp5_ASAP7_75t_L g4085 ( 
.A(n_3602),
.B(n_3103),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3890),
.B(n_3221),
.Y(n_4086)
);

INVx1_ASAP7_75t_L g4087 ( 
.A(n_3533),
.Y(n_4087)
);

AND3x1_ASAP7_75t_L g4088 ( 
.A(n_3716),
.B(n_3037),
.C(n_3015),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3536),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_L g4090 ( 
.A(n_3486),
.B(n_3507),
.Y(n_4090)
);

NAND2xp5_ASAP7_75t_L g4091 ( 
.A(n_3598),
.B(n_3508),
.Y(n_4091)
);

BUFx6f_ASAP7_75t_L g4092 ( 
.A(n_3466),
.Y(n_4092)
);

HB1xp67_ASAP7_75t_L g4093 ( 
.A(n_3557),
.Y(n_4093)
);

INVx3_ASAP7_75t_L g4094 ( 
.A(n_3804),
.Y(n_4094)
);

INVx1_ASAP7_75t_SL g4095 ( 
.A(n_3525),
.Y(n_4095)
);

AND2x6_ASAP7_75t_L g4096 ( 
.A(n_3463),
.B(n_2931),
.Y(n_4096)
);

NOR2xp33_ASAP7_75t_L g4097 ( 
.A(n_3495),
.B(n_3032),
.Y(n_4097)
);

INVx2_ASAP7_75t_L g4098 ( 
.A(n_3517),
.Y(n_4098)
);

INVx1_ASAP7_75t_L g4099 ( 
.A(n_3538),
.Y(n_4099)
);

HB1xp67_ASAP7_75t_L g4100 ( 
.A(n_3557),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3541),
.Y(n_4101)
);

INVx2_ASAP7_75t_L g4102 ( 
.A(n_3535),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3546),
.Y(n_4103)
);

INVx2_ASAP7_75t_SL g4104 ( 
.A(n_3814),
.Y(n_4104)
);

AOI22xp33_ASAP7_75t_L g4105 ( 
.A1(n_3603),
.A2(n_3221),
.B1(n_3226),
.B2(n_3273),
.Y(n_4105)
);

BUFx2_ASAP7_75t_L g4106 ( 
.A(n_3778),
.Y(n_4106)
);

INVx1_ASAP7_75t_L g4107 ( 
.A(n_3549),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_L g4108 ( 
.A(n_3464),
.B(n_3226),
.Y(n_4108)
);

AOI21xp5_ASAP7_75t_L g4109 ( 
.A1(n_3547),
.A2(n_2934),
.B(n_2824),
.Y(n_4109)
);

AND2x4_ASAP7_75t_SL g4110 ( 
.A(n_3814),
.B(n_3098),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3678),
.B(n_2848),
.Y(n_4111)
);

AO21x1_ASAP7_75t_L g4112 ( 
.A1(n_3510),
.A2(n_2983),
.B(n_3243),
.Y(n_4112)
);

OR2x2_ASAP7_75t_L g4113 ( 
.A(n_3711),
.B(n_3860),
.Y(n_4113)
);

INVxp67_ASAP7_75t_L g4114 ( 
.A(n_3564),
.Y(n_4114)
);

NOR2x1_ASAP7_75t_R g4115 ( 
.A(n_3844),
.B(n_2971),
.Y(n_4115)
);

AOI22xp5_ASAP7_75t_L g4116 ( 
.A1(n_3609),
.A2(n_3468),
.B1(n_3587),
.B2(n_3472),
.Y(n_4116)
);

AOI22xp33_ASAP7_75t_L g4117 ( 
.A1(n_3946),
.A2(n_3273),
.B1(n_3128),
.B2(n_3259),
.Y(n_4117)
);

CKINVDCx6p67_ASAP7_75t_R g4118 ( 
.A(n_3523),
.Y(n_4118)
);

HB1xp67_ASAP7_75t_L g4119 ( 
.A(n_3896),
.Y(n_4119)
);

BUFx12f_ASAP7_75t_L g4120 ( 
.A(n_3750),
.Y(n_4120)
);

NOR2xp67_ASAP7_75t_L g4121 ( 
.A(n_3844),
.B(n_3976),
.Y(n_4121)
);

INVx3_ASAP7_75t_L g4122 ( 
.A(n_3976),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3930),
.B(n_3078),
.Y(n_4123)
);

AOI22xp5_ASAP7_75t_L g4124 ( 
.A1(n_3468),
.A2(n_3587),
.B1(n_3469),
.B2(n_3791),
.Y(n_4124)
);

AOI22xp5_ASAP7_75t_L g4125 ( 
.A1(n_3728),
.A2(n_3239),
.B1(n_3260),
.B2(n_3024),
.Y(n_4125)
);

AND2x2_ASAP7_75t_L g4126 ( 
.A(n_3866),
.B(n_3161),
.Y(n_4126)
);

NOR2xp33_ASAP7_75t_L g4127 ( 
.A(n_3822),
.B(n_3818),
.Y(n_4127)
);

BUFx3_ASAP7_75t_L g4128 ( 
.A(n_3527),
.Y(n_4128)
);

OAI21x1_ASAP7_75t_L g4129 ( 
.A1(n_3516),
.A2(n_2847),
.B(n_2820),
.Y(n_4129)
);

BUFx3_ASAP7_75t_L g4130 ( 
.A(n_3572),
.Y(n_4130)
);

OR2x6_ASAP7_75t_L g4131 ( 
.A(n_3728),
.B(n_3006),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_3463),
.B(n_2816),
.Y(n_4132)
);

AND2x2_ASAP7_75t_SL g4133 ( 
.A(n_3624),
.B(n_3006),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_3562),
.Y(n_4134)
);

AOI22xp33_ASAP7_75t_L g4135 ( 
.A1(n_3671),
.A2(n_3273),
.B1(n_3128),
.B2(n_3259),
.Y(n_4135)
);

NOR2xp33_ASAP7_75t_L g4136 ( 
.A(n_3819),
.B(n_3265),
.Y(n_4136)
);

INVx2_ASAP7_75t_L g4137 ( 
.A(n_3540),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_L g4138 ( 
.A(n_4030),
.B(n_2880),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_3850),
.B(n_3194),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3923),
.B(n_2919),
.Y(n_4140)
);

HB1xp67_ASAP7_75t_L g4141 ( 
.A(n_3641),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_SL g4142 ( 
.A(n_3968),
.B(n_3062),
.Y(n_4142)
);

AND2x4_ASAP7_75t_L g4143 ( 
.A(n_3497),
.B(n_2816),
.Y(n_4143)
);

AND2x2_ASAP7_75t_L g4144 ( 
.A(n_3980),
.B(n_3182),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_3574),
.Y(n_4145)
);

NOR2x1p5_ASAP7_75t_L g4146 ( 
.A(n_3669),
.B(n_2908),
.Y(n_4146)
);

AOI22xp5_ASAP7_75t_L g4147 ( 
.A1(n_3728),
.A2(n_3041),
.B1(n_3291),
.B2(n_2803),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_3583),
.Y(n_4148)
);

NAND2xp5_ASAP7_75t_SL g4149 ( 
.A(n_3968),
.B(n_3062),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_3585),
.Y(n_4150)
);

BUFx2_ASAP7_75t_L g4151 ( 
.A(n_3977),
.Y(n_4151)
);

NOR2xp33_ASAP7_75t_L g4152 ( 
.A(n_3943),
.B(n_3862),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_3597),
.Y(n_4153)
);

INVx4_ASAP7_75t_SL g4154 ( 
.A(n_3523),
.Y(n_4154)
);

NOR2xp33_ASAP7_75t_R g4155 ( 
.A(n_3941),
.B(n_2942),
.Y(n_4155)
);

INVx2_ASAP7_75t_SL g4156 ( 
.A(n_3617),
.Y(n_4156)
);

BUFx2_ASAP7_75t_L g4157 ( 
.A(n_3747),
.Y(n_4157)
);

NOR2xp33_ASAP7_75t_L g4158 ( 
.A(n_3751),
.B(n_3084),
.Y(n_4158)
);

INVx4_ASAP7_75t_L g4159 ( 
.A(n_3766),
.Y(n_4159)
);

AO21x1_ASAP7_75t_L g4160 ( 
.A1(n_3510),
.A2(n_3246),
.B(n_3243),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_3601),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3503),
.B(n_2922),
.Y(n_4162)
);

INVx1_ASAP7_75t_L g4163 ( 
.A(n_3604),
.Y(n_4163)
);

INVx2_ASAP7_75t_L g4164 ( 
.A(n_3545),
.Y(n_4164)
);

OR2x2_ASAP7_75t_L g4165 ( 
.A(n_3982),
.B(n_3237),
.Y(n_4165)
);

BUFx6f_ASAP7_75t_L g4166 ( 
.A(n_3466),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_3615),
.Y(n_4167)
);

NOR2xp33_ASAP7_75t_L g4168 ( 
.A(n_3681),
.B(n_3013),
.Y(n_4168)
);

INVx2_ASAP7_75t_L g4169 ( 
.A(n_3559),
.Y(n_4169)
);

NOR2xp33_ASAP7_75t_R g4170 ( 
.A(n_3837),
.B(n_2933),
.Y(n_4170)
);

BUFx6f_ASAP7_75t_L g4171 ( 
.A(n_3466),
.Y(n_4171)
);

NOR2xp33_ASAP7_75t_L g4172 ( 
.A(n_3855),
.B(n_3048),
.Y(n_4172)
);

AND2x2_ASAP7_75t_L g4173 ( 
.A(n_3984),
.B(n_2819),
.Y(n_4173)
);

AOI22xp33_ASAP7_75t_L g4174 ( 
.A1(n_3755),
.A2(n_3273),
.B1(n_3128),
.B2(n_3259),
.Y(n_4174)
);

INVx2_ASAP7_75t_L g4175 ( 
.A(n_3565),
.Y(n_4175)
);

A2O1A1Ixp33_ASAP7_75t_L g4176 ( 
.A1(n_3793),
.A2(n_3164),
.B(n_3191),
.C(n_3272),
.Y(n_4176)
);

NAND2xp5_ASAP7_75t_SL g4177 ( 
.A(n_3703),
.B(n_3062),
.Y(n_4177)
);

INVx1_ASAP7_75t_L g4178 ( 
.A(n_3616),
.Y(n_4178)
);

NAND2xp5_ASAP7_75t_L g4179 ( 
.A(n_3476),
.B(n_2951),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_3619),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_3460),
.Y(n_4181)
);

INVx2_ASAP7_75t_L g4182 ( 
.A(n_3566),
.Y(n_4182)
);

HB1xp67_ASAP7_75t_L g4183 ( 
.A(n_3798),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_3635),
.Y(n_4184)
);

NAND2xp5_ASAP7_75t_SL g4185 ( 
.A(n_3703),
.B(n_3125),
.Y(n_4185)
);

NAND2xp5_ASAP7_75t_L g4186 ( 
.A(n_3478),
.B(n_3840),
.Y(n_4186)
);

CKINVDCx5p33_ASAP7_75t_R g4187 ( 
.A(n_3750),
.Y(n_4187)
);

INVx1_ASAP7_75t_L g4188 ( 
.A(n_3643),
.Y(n_4188)
);

NAND2xp5_ASAP7_75t_SL g4189 ( 
.A(n_3650),
.B(n_3125),
.Y(n_4189)
);

HB1xp67_ASAP7_75t_L g4190 ( 
.A(n_3578),
.Y(n_4190)
);

CKINVDCx5p33_ASAP7_75t_R g4191 ( 
.A(n_3989),
.Y(n_4191)
);

INVx2_ASAP7_75t_SL g4192 ( 
.A(n_3856),
.Y(n_4192)
);

HB1xp67_ASAP7_75t_L g4193 ( 
.A(n_4010),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_3646),
.Y(n_4194)
);

NAND2xp5_ASAP7_75t_L g4195 ( 
.A(n_3853),
.B(n_3863),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_3661),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_3567),
.Y(n_4197)
);

HB1xp67_ASAP7_75t_L g4198 ( 
.A(n_4019),
.Y(n_4198)
);

NAND3xp33_ASAP7_75t_SL g4199 ( 
.A(n_3845),
.B(n_3300),
.C(n_3292),
.Y(n_4199)
);

NAND2xp5_ASAP7_75t_L g4200 ( 
.A(n_3481),
.B(n_3017),
.Y(n_4200)
);

NAND2x1p5_ASAP7_75t_L g4201 ( 
.A(n_3512),
.B(n_2835),
.Y(n_4201)
);

INVx3_ASAP7_75t_L g4202 ( 
.A(n_3497),
.Y(n_4202)
);

INVx2_ASAP7_75t_SL g4203 ( 
.A(n_3903),
.Y(n_4203)
);

NAND3xp33_ASAP7_75t_SL g4204 ( 
.A(n_3845),
.B(n_3365),
.C(n_3356),
.Y(n_4204)
);

NAND2xp5_ASAP7_75t_SL g4205 ( 
.A(n_3650),
.B(n_3125),
.Y(n_4205)
);

AOI22xp5_ASAP7_75t_L g4206 ( 
.A1(n_4006),
.A2(n_3324),
.B1(n_3053),
.B2(n_3158),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_3674),
.Y(n_4207)
);

INVx2_ASAP7_75t_L g4208 ( 
.A(n_3569),
.Y(n_4208)
);

BUFx6f_ASAP7_75t_L g4209 ( 
.A(n_3548),
.Y(n_4209)
);

AOI21xp33_ASAP7_75t_L g4210 ( 
.A1(n_3842),
.A2(n_3431),
.B(n_3404),
.Y(n_4210)
);

AND2x2_ASAP7_75t_SL g4211 ( 
.A(n_3897),
.B(n_3150),
.Y(n_4211)
);

NAND3xp33_ASAP7_75t_SL g4212 ( 
.A(n_3880),
.B(n_3254),
.C(n_3230),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_3498),
.B(n_3485),
.Y(n_4213)
);

AOI22xp5_ASAP7_75t_L g4214 ( 
.A1(n_3842),
.A2(n_3247),
.B1(n_3146),
.B2(n_3139),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_SL g4215 ( 
.A(n_3607),
.B(n_3157),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_3993),
.B(n_2972),
.Y(n_4216)
);

AOI21xp33_ASAP7_75t_L g4217 ( 
.A1(n_3596),
.A2(n_3118),
.B(n_2800),
.Y(n_4217)
);

INVx1_ASAP7_75t_L g4218 ( 
.A(n_3680),
.Y(n_4218)
);

OAI21xp5_ASAP7_75t_L g4219 ( 
.A1(n_3665),
.A2(n_3971),
.B(n_4034),
.Y(n_4219)
);

OAI22xp5_ASAP7_75t_SL g4220 ( 
.A1(n_3889),
.A2(n_2988),
.B1(n_3099),
.B2(n_2878),
.Y(n_4220)
);

BUFx3_ASAP7_75t_L g4221 ( 
.A(n_3974),
.Y(n_4221)
);

INVx3_ASAP7_75t_L g4222 ( 
.A(n_3550),
.Y(n_4222)
);

NAND2x1_ASAP7_75t_SL g4223 ( 
.A(n_3880),
.B(n_3153),
.Y(n_4223)
);

AOI22xp5_ASAP7_75t_L g4224 ( 
.A1(n_3824),
.A2(n_2968),
.B1(n_3019),
.B2(n_2916),
.Y(n_4224)
);

AND2x6_ASAP7_75t_SL g4225 ( 
.A(n_4003),
.B(n_2818),
.Y(n_4225)
);

NAND2xp5_ASAP7_75t_L g4226 ( 
.A(n_3563),
.B(n_3007),
.Y(n_4226)
);

INVx1_ASAP7_75t_L g4227 ( 
.A(n_3684),
.Y(n_4227)
);

AND2x2_ASAP7_75t_SL g4228 ( 
.A(n_3701),
.B(n_3150),
.Y(n_4228)
);

AOI21xp5_ASAP7_75t_L g4229 ( 
.A1(n_3654),
.A2(n_2934),
.B(n_2974),
.Y(n_4229)
);

CKINVDCx5p33_ASAP7_75t_R g4230 ( 
.A(n_3763),
.Y(n_4230)
);

AND2x4_ASAP7_75t_L g4231 ( 
.A(n_3550),
.B(n_2843),
.Y(n_4231)
);

AOI22xp5_ASAP7_75t_L g4232 ( 
.A1(n_3869),
.A2(n_3753),
.B1(n_3825),
.B2(n_3900),
.Y(n_4232)
);

AND2x6_ASAP7_75t_L g4233 ( 
.A(n_3607),
.B(n_2934),
.Y(n_4233)
);

HB1xp67_ASAP7_75t_L g4234 ( 
.A(n_4020),
.Y(n_4234)
);

OAI22xp5_ASAP7_75t_L g4235 ( 
.A1(n_3477),
.A2(n_2976),
.B1(n_3248),
.B2(n_3246),
.Y(n_4235)
);

AOI22xp33_ASAP7_75t_L g4236 ( 
.A1(n_3755),
.A2(n_3259),
.B1(n_3236),
.B2(n_3272),
.Y(n_4236)
);

NAND2xp5_ASAP7_75t_L g4237 ( 
.A(n_3477),
.B(n_3022),
.Y(n_4237)
);

INVx1_ASAP7_75t_L g4238 ( 
.A(n_3713),
.Y(n_4238)
);

INVx5_ASAP7_75t_L g4239 ( 
.A(n_3735),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_3516),
.Y(n_4240)
);

NAND2xp5_ASAP7_75t_L g4241 ( 
.A(n_3769),
.B(n_3575),
.Y(n_4241)
);

BUFx12f_ASAP7_75t_SL g4242 ( 
.A(n_3807),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_3742),
.B(n_3033),
.Y(n_4243)
);

AND2x4_ASAP7_75t_L g4244 ( 
.A(n_3794),
.B(n_2843),
.Y(n_4244)
);

AND2x6_ASAP7_75t_SL g4245 ( 
.A(n_3807),
.B(n_3933),
.Y(n_4245)
);

INVx3_ASAP7_75t_L g4246 ( 
.A(n_3591),
.Y(n_4246)
);

INVx2_ASAP7_75t_SL g4247 ( 
.A(n_3773),
.Y(n_4247)
);

INVx2_ASAP7_75t_L g4248 ( 
.A(n_3590),
.Y(n_4248)
);

BUFx2_ASAP7_75t_L g4249 ( 
.A(n_3693),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_3605),
.Y(n_4250)
);

INVx3_ASAP7_75t_L g4251 ( 
.A(n_3591),
.Y(n_4251)
);

INVx1_ASAP7_75t_SL g4252 ( 
.A(n_3764),
.Y(n_4252)
);

INVx1_ASAP7_75t_L g4253 ( 
.A(n_3720),
.Y(n_4253)
);

INVxp67_ASAP7_75t_L g4254 ( 
.A(n_3905),
.Y(n_4254)
);

AND2x2_ASAP7_75t_L g4255 ( 
.A(n_4026),
.B(n_3197),
.Y(n_4255)
);

INVx1_ASAP7_75t_L g4256 ( 
.A(n_3729),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_3732),
.Y(n_4257)
);

INVx2_ASAP7_75t_L g4258 ( 
.A(n_3610),
.Y(n_4258)
);

INVx1_ASAP7_75t_L g4259 ( 
.A(n_3746),
.Y(n_4259)
);

INVx1_ASAP7_75t_L g4260 ( 
.A(n_3749),
.Y(n_4260)
);

OR2x2_ASAP7_75t_L g4261 ( 
.A(n_3901),
.B(n_3241),
.Y(n_4261)
);

HB1xp67_ASAP7_75t_L g4262 ( 
.A(n_3803),
.Y(n_4262)
);

NOR2x1_ASAP7_75t_L g4263 ( 
.A(n_3496),
.B(n_2988),
.Y(n_4263)
);

NAND2xp5_ASAP7_75t_L g4264 ( 
.A(n_3748),
.B(n_3039),
.Y(n_4264)
);

AND2x6_ASAP7_75t_L g4265 ( 
.A(n_3649),
.B(n_3328),
.Y(n_4265)
);

INVx2_ASAP7_75t_L g4266 ( 
.A(n_3636),
.Y(n_4266)
);

CKINVDCx5p33_ASAP7_75t_R g4267 ( 
.A(n_3892),
.Y(n_4267)
);

NAND2xp5_ASAP7_75t_SL g4268 ( 
.A(n_3649),
.B(n_3157),
.Y(n_4268)
);

NAND2xp5_ASAP7_75t_L g4269 ( 
.A(n_3490),
.B(n_3082),
.Y(n_4269)
);

INVx8_ASAP7_75t_L g4270 ( 
.A(n_3870),
.Y(n_4270)
);

NAND2xp5_ASAP7_75t_L g4271 ( 
.A(n_3805),
.B(n_3092),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_3812),
.B(n_3826),
.Y(n_4272)
);

OR2x6_ASAP7_75t_L g4273 ( 
.A(n_3526),
.B(n_3529),
.Y(n_4273)
);

INVx2_ASAP7_75t_L g4274 ( 
.A(n_3642),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_3832),
.B(n_3238),
.Y(n_4275)
);

O2A1O1Ixp33_ASAP7_75t_L g4276 ( 
.A1(n_4021),
.A2(n_3225),
.B(n_3023),
.C(n_3209),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_SL g4277 ( 
.A(n_3660),
.B(n_3157),
.Y(n_4277)
);

AND2x6_ASAP7_75t_SL g4278 ( 
.A(n_3942),
.B(n_3835),
.Y(n_4278)
);

NAND3xp33_ASAP7_75t_SL g4279 ( 
.A(n_3839),
.B(n_3153),
.C(n_3253),
.Y(n_4279)
);

AND2x2_ASAP7_75t_L g4280 ( 
.A(n_3811),
.B(n_3249),
.Y(n_4280)
);

AND2x4_ASAP7_75t_L g4281 ( 
.A(n_3843),
.B(n_2800),
.Y(n_4281)
);

INVx2_ASAP7_75t_L g4282 ( 
.A(n_3645),
.Y(n_4282)
);

AOI22xp33_ASAP7_75t_L g4283 ( 
.A1(n_4007),
.A2(n_3236),
.B1(n_3248),
.B2(n_2870),
.Y(n_4283)
);

OAI22xp33_ASAP7_75t_L g4284 ( 
.A1(n_3839),
.A2(n_3257),
.B1(n_3256),
.B2(n_3069),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_3760),
.Y(n_4285)
);

CKINVDCx20_ASAP7_75t_R g4286 ( 
.A(n_3542),
.Y(n_4286)
);

INVx2_ASAP7_75t_L g4287 ( 
.A(n_3667),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_3737),
.B(n_3005),
.Y(n_4288)
);

INVx1_ASAP7_75t_L g4289 ( 
.A(n_3783),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_3872),
.B(n_3258),
.Y(n_4290)
);

BUFx3_ASAP7_75t_L g4291 ( 
.A(n_3765),
.Y(n_4291)
);

INVx2_ASAP7_75t_L g4292 ( 
.A(n_3668),
.Y(n_4292)
);

NOR2xp67_ASAP7_75t_L g4293 ( 
.A(n_3721),
.B(n_3312),
.Y(n_4293)
);

INVx1_ASAP7_75t_L g4294 ( 
.A(n_3795),
.Y(n_4294)
);

AOI22xp5_ASAP7_75t_L g4295 ( 
.A1(n_3735),
.A2(n_3223),
.B1(n_3266),
.B2(n_3171),
.Y(n_4295)
);

INVx2_ASAP7_75t_L g4296 ( 
.A(n_3688),
.Y(n_4296)
);

NAND2xp5_ASAP7_75t_L g4297 ( 
.A(n_3883),
.B(n_3261),
.Y(n_4297)
);

AND2x2_ASAP7_75t_SL g4298 ( 
.A(n_3790),
.B(n_2996),
.Y(n_4298)
);

INVx2_ASAP7_75t_L g4299 ( 
.A(n_3695),
.Y(n_4299)
);

AOI22xp33_ASAP7_75t_L g4300 ( 
.A1(n_3797),
.A2(n_3236),
.B1(n_2870),
.B2(n_2881),
.Y(n_4300)
);

BUFx3_ASAP7_75t_L g4301 ( 
.A(n_3756),
.Y(n_4301)
);

AND2x4_ASAP7_75t_L g4302 ( 
.A(n_3670),
.B(n_3752),
.Y(n_4302)
);

INVx3_ASAP7_75t_L g4303 ( 
.A(n_3870),
.Y(n_4303)
);

BUFx3_ASAP7_75t_L g4304 ( 
.A(n_3613),
.Y(n_4304)
);

INVx2_ASAP7_75t_SL g4305 ( 
.A(n_3618),
.Y(n_4305)
);

AND3x2_ASAP7_75t_SL g4306 ( 
.A(n_3737),
.B(n_3068),
.C(n_2818),
.Y(n_4306)
);

AOI22xp5_ASAP7_75t_L g4307 ( 
.A1(n_3735),
.A2(n_3236),
.B1(n_3231),
.B2(n_3234),
.Y(n_4307)
);

A2O1A1Ixp33_ASAP7_75t_L g4308 ( 
.A1(n_3948),
.A2(n_3284),
.B(n_3297),
.C(n_3279),
.Y(n_4308)
);

BUFx3_ASAP7_75t_L g4309 ( 
.A(n_3687),
.Y(n_4309)
);

OAI21xp33_ASAP7_75t_L g4310 ( 
.A1(n_4025),
.A2(n_3073),
.B(n_3212),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_3811),
.B(n_3029),
.Y(n_4311)
);

AO22x1_ASAP7_75t_L g4312 ( 
.A1(n_3735),
.A2(n_2917),
.B1(n_2871),
.B2(n_2881),
.Y(n_4312)
);

NOR2xp33_ASAP7_75t_SL g4313 ( 
.A(n_3956),
.B(n_3008),
.Y(n_4313)
);

INVx3_ASAP7_75t_L g4314 ( 
.A(n_3718),
.Y(n_4314)
);

INVx2_ASAP7_75t_L g4315 ( 
.A(n_3704),
.Y(n_4315)
);

HB1xp67_ASAP7_75t_L g4316 ( 
.A(n_3849),
.Y(n_4316)
);

AOI22xp5_ASAP7_75t_L g4317 ( 
.A1(n_3730),
.A2(n_2871),
.B1(n_2881),
.B2(n_2870),
.Y(n_4317)
);

BUFx3_ASAP7_75t_L g4318 ( 
.A(n_3917),
.Y(n_4318)
);

INVx1_ASAP7_75t_SL g4319 ( 
.A(n_3954),
.Y(n_4319)
);

INVx2_ASAP7_75t_L g4320 ( 
.A(n_3705),
.Y(n_4320)
);

AOI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_3809),
.A2(n_2871),
.B1(n_2881),
.B2(n_2870),
.Y(n_4321)
);

BUFx2_ASAP7_75t_L g4322 ( 
.A(n_3787),
.Y(n_4322)
);

INVx1_ASAP7_75t_L g4323 ( 
.A(n_3823),
.Y(n_4323)
);

INVx2_ASAP7_75t_L g4324 ( 
.A(n_3708),
.Y(n_4324)
);

OAI22xp33_ASAP7_75t_L g4325 ( 
.A1(n_4025),
.A2(n_3075),
.B1(n_3069),
.B2(n_2906),
.Y(n_4325)
);

NAND2x1p5_ASAP7_75t_L g4326 ( 
.A(n_3894),
.B(n_2963),
.Y(n_4326)
);

BUFx3_ASAP7_75t_L g4327 ( 
.A(n_3787),
.Y(n_4327)
);

INVx2_ASAP7_75t_L g4328 ( 
.A(n_3724),
.Y(n_4328)
);

INVx1_ASAP7_75t_L g4329 ( 
.A(n_3828),
.Y(n_4329)
);

BUFx6f_ASAP7_75t_L g4330 ( 
.A(n_3548),
.Y(n_4330)
);

NAND2xp5_ASAP7_75t_L g4331 ( 
.A(n_3886),
.B(n_3222),
.Y(n_4331)
);

NAND2xp33_ASAP7_75t_L g4332 ( 
.A(n_3718),
.B(n_2871),
.Y(n_4332)
);

HB1xp67_ASAP7_75t_L g4333 ( 
.A(n_3857),
.Y(n_4333)
);

INVx1_ASAP7_75t_L g4334 ( 
.A(n_3951),
.Y(n_4334)
);

AND2x6_ASAP7_75t_SL g4335 ( 
.A(n_3637),
.B(n_3368),
.Y(n_4335)
);

INVx2_ASAP7_75t_SL g4336 ( 
.A(n_3558),
.Y(n_4336)
);

OR2x2_ASAP7_75t_L g4337 ( 
.A(n_3758),
.B(n_3133),
.Y(n_4337)
);

NAND2xp5_ASAP7_75t_L g4338 ( 
.A(n_3902),
.B(n_3228),
.Y(n_4338)
);

INVx1_ASAP7_75t_L g4339 ( 
.A(n_3953),
.Y(n_4339)
);

AOI21xp5_ASAP7_75t_L g4340 ( 
.A1(n_3647),
.A2(n_3284),
.B(n_3279),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_3955),
.Y(n_4341)
);

INVx3_ASAP7_75t_L g4342 ( 
.A(n_3718),
.Y(n_4342)
);

INVx2_ASAP7_75t_SL g4343 ( 
.A(n_4009),
.Y(n_4343)
);

INVx2_ASAP7_75t_SL g4344 ( 
.A(n_3577),
.Y(n_4344)
);

NAND2xp5_ASAP7_75t_SL g4345 ( 
.A(n_3660),
.B(n_3094),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_3960),
.Y(n_4346)
);

AOI22xp5_ASAP7_75t_L g4347 ( 
.A1(n_3958),
.A2(n_2906),
.B1(n_3155),
.B2(n_3176),
.Y(n_4347)
);

AO22x1_ASAP7_75t_L g4348 ( 
.A1(n_3767),
.A2(n_2917),
.B1(n_3391),
.B2(n_3371),
.Y(n_4348)
);

BUFx3_ASAP7_75t_L g4349 ( 
.A(n_3867),
.Y(n_4349)
);

NAND2xp5_ASAP7_75t_SL g4350 ( 
.A(n_3718),
.B(n_3948),
.Y(n_4350)
);

INVx1_ASAP7_75t_L g4351 ( 
.A(n_3967),
.Y(n_4351)
);

INVx1_ASAP7_75t_L g4352 ( 
.A(n_3987),
.Y(n_4352)
);

NAND2xp5_ASAP7_75t_L g4353 ( 
.A(n_3595),
.B(n_3229),
.Y(n_4353)
);

INVx2_ASAP7_75t_L g4354 ( 
.A(n_3740),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_3992),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_3999),
.Y(n_4356)
);

NAND2xp5_ASAP7_75t_SL g4357 ( 
.A(n_3718),
.B(n_3094),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_L g4358 ( 
.A(n_3461),
.B(n_3245),
.Y(n_4358)
);

NAND2xp5_ASAP7_75t_L g4359 ( 
.A(n_3462),
.B(n_3251),
.Y(n_4359)
);

INVx1_ASAP7_75t_L g4360 ( 
.A(n_4002),
.Y(n_4360)
);

NAND2xp5_ASAP7_75t_L g4361 ( 
.A(n_3470),
.B(n_3141),
.Y(n_4361)
);

INVx1_ASAP7_75t_L g4362 ( 
.A(n_4016),
.Y(n_4362)
);

HB1xp67_ASAP7_75t_L g4363 ( 
.A(n_3871),
.Y(n_4363)
);

INVx2_ASAP7_75t_L g4364 ( 
.A(n_3741),
.Y(n_4364)
);

INVx1_ASAP7_75t_L g4365 ( 
.A(n_4018),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4028),
.Y(n_4366)
);

INVx1_ASAP7_75t_SL g4367 ( 
.A(n_3471),
.Y(n_4367)
);

OR2x6_ASAP7_75t_L g4368 ( 
.A(n_3589),
.B(n_2963),
.Y(n_4368)
);

NAND2xp5_ASAP7_75t_L g4369 ( 
.A(n_3474),
.B(n_3141),
.Y(n_4369)
);

INVx2_ASAP7_75t_L g4370 ( 
.A(n_3743),
.Y(n_4370)
);

INVx1_ASAP7_75t_L g4371 ( 
.A(n_4029),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4024),
.Y(n_4372)
);

INVx2_ASAP7_75t_L g4373 ( 
.A(n_3745),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_3876),
.Y(n_4374)
);

AND2x2_ASAP7_75t_L g4375 ( 
.A(n_3723),
.B(n_3198),
.Y(n_4375)
);

AOI22xp33_ASAP7_75t_L g4376 ( 
.A1(n_3983),
.A2(n_3155),
.B1(n_3179),
.B2(n_3219),
.Y(n_4376)
);

INVxp67_ASAP7_75t_L g4377 ( 
.A(n_3656),
.Y(n_4377)
);

INVx1_ASAP7_75t_L g4378 ( 
.A(n_3881),
.Y(n_4378)
);

HB1xp67_ASAP7_75t_L g4379 ( 
.A(n_3882),
.Y(n_4379)
);

NAND2xp5_ASAP7_75t_L g4380 ( 
.A(n_3515),
.B(n_3174),
.Y(n_4380)
);

INVx2_ASAP7_75t_L g4381 ( 
.A(n_3770),
.Y(n_4381)
);

NAND2xp5_ASAP7_75t_SL g4382 ( 
.A(n_3665),
.B(n_3297),
.Y(n_4382)
);

INVx1_ASAP7_75t_L g4383 ( 
.A(n_3884),
.Y(n_4383)
);

AND2x4_ASAP7_75t_L g4384 ( 
.A(n_3638),
.B(n_3303),
.Y(n_4384)
);

AOI22xp5_ASAP7_75t_L g4385 ( 
.A1(n_3675),
.A2(n_3353),
.B1(n_3012),
.B2(n_3121),
.Y(n_4385)
);

NOR2xp33_ASAP7_75t_SL g4386 ( 
.A(n_3767),
.B(n_2963),
.Y(n_4386)
);

AOI22xp33_ASAP7_75t_L g4387 ( 
.A1(n_3979),
.A2(n_3242),
.B1(n_3219),
.B2(n_3195),
.Y(n_4387)
);

CKINVDCx5p33_ASAP7_75t_R g4388 ( 
.A(n_3937),
.Y(n_4388)
);

NAND3xp33_ASAP7_75t_L g4389 ( 
.A(n_3799),
.B(n_3172),
.C(n_3162),
.Y(n_4389)
);

NAND2xp5_ASAP7_75t_L g4390 ( 
.A(n_3534),
.B(n_3181),
.Y(n_4390)
);

INVx2_ASAP7_75t_SL g4391 ( 
.A(n_3859),
.Y(n_4391)
);

INVx2_ASAP7_75t_L g4392 ( 
.A(n_3771),
.Y(n_4392)
);

INVx2_ASAP7_75t_L g4393 ( 
.A(n_3775),
.Y(n_4393)
);

CKINVDCx5p33_ASAP7_75t_R g4394 ( 
.A(n_3664),
.Y(n_4394)
);

INVx2_ASAP7_75t_L g4395 ( 
.A(n_3779),
.Y(n_4395)
);

AND2x6_ASAP7_75t_L g4396 ( 
.A(n_3548),
.B(n_3411),
.Y(n_4396)
);

BUFx3_ASAP7_75t_L g4397 ( 
.A(n_3898),
.Y(n_4397)
);

CKINVDCx5p33_ASAP7_75t_R g4398 ( 
.A(n_3644),
.Y(n_4398)
);

NAND2xp5_ASAP7_75t_L g4399 ( 
.A(n_3576),
.B(n_3204),
.Y(n_4399)
);

CKINVDCx5p33_ASAP7_75t_R g4400 ( 
.A(n_3651),
.Y(n_4400)
);

NAND2xp5_ASAP7_75t_L g4401 ( 
.A(n_3521),
.B(n_3105),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_3899),
.Y(n_4402)
);

AOI22xp33_ASAP7_75t_L g4403 ( 
.A1(n_4000),
.A2(n_3242),
.B1(n_3076),
.B2(n_3172),
.Y(n_4403)
);

CKINVDCx5p33_ASAP7_75t_R g4404 ( 
.A(n_3652),
.Y(n_4404)
);

AOI21xp5_ASAP7_75t_L g4405 ( 
.A1(n_3647),
.A2(n_3317),
.B(n_3303),
.Y(n_4405)
);

NOR2xp33_ASAP7_75t_L g4406 ( 
.A(n_3530),
.B(n_2921),
.Y(n_4406)
);

BUFx2_ASAP7_75t_L g4407 ( 
.A(n_3781),
.Y(n_4407)
);

INVx3_ASAP7_75t_L g4408 ( 
.A(n_3777),
.Y(n_4408)
);

OR2x6_ASAP7_75t_L g4409 ( 
.A(n_3592),
.B(n_2965),
.Y(n_4409)
);

A2O1A1Ixp33_ASAP7_75t_L g4410 ( 
.A1(n_3831),
.A2(n_3323),
.B(n_3325),
.C(n_3317),
.Y(n_4410)
);

NAND2xp5_ASAP7_75t_L g4411 ( 
.A(n_3759),
.B(n_3210),
.Y(n_4411)
);

NAND2xp5_ASAP7_75t_L g4412 ( 
.A(n_3970),
.B(n_3210),
.Y(n_4412)
);

INVx2_ASAP7_75t_L g4413 ( 
.A(n_3784),
.Y(n_4413)
);

AO22x1_ASAP7_75t_L g4414 ( 
.A1(n_3944),
.A2(n_2917),
.B1(n_3391),
.B2(n_3371),
.Y(n_4414)
);

AOI22xp5_ASAP7_75t_L g4415 ( 
.A1(n_3925),
.A2(n_3121),
.B1(n_3076),
.B2(n_3198),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_L g4416 ( 
.A(n_3891),
.B(n_2990),
.Y(n_4416)
);

NAND2x1p5_ASAP7_75t_L g4417 ( 
.A(n_3473),
.B(n_2965),
.Y(n_4417)
);

NAND2xp5_ASAP7_75t_SL g4418 ( 
.A(n_3553),
.B(n_3323),
.Y(n_4418)
);

INVx3_ASAP7_75t_L g4419 ( 
.A(n_3777),
.Y(n_4419)
);

INVx3_ASAP7_75t_L g4420 ( 
.A(n_3777),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_3904),
.Y(n_4421)
);

AND2x4_ASAP7_75t_L g4422 ( 
.A(n_3682),
.B(n_3325),
.Y(n_4422)
);

CKINVDCx20_ASAP7_75t_R g4423 ( 
.A(n_3653),
.Y(n_4423)
);

NAND2xp5_ASAP7_75t_SL g4424 ( 
.A(n_3629),
.B(n_3328),
.Y(n_4424)
);

INVx2_ASAP7_75t_L g4425 ( 
.A(n_3789),
.Y(n_4425)
);

AOI22xp33_ASAP7_75t_L g4426 ( 
.A1(n_3988),
.A2(n_3172),
.B1(n_3162),
.B2(n_3207),
.Y(n_4426)
);

INVx3_ASAP7_75t_L g4427 ( 
.A(n_3792),
.Y(n_4427)
);

NAND2xp5_ASAP7_75t_SL g4428 ( 
.A(n_3829),
.B(n_3347),
.Y(n_4428)
);

BUFx2_ASAP7_75t_L g4429 ( 
.A(n_3906),
.Y(n_4429)
);

INVx8_ASAP7_75t_L g4430 ( 
.A(n_3792),
.Y(n_4430)
);

BUFx12f_ASAP7_75t_L g4431 ( 
.A(n_3792),
.Y(n_4431)
);

OAI22xp5_ASAP7_75t_SL g4432 ( 
.A1(n_4011),
.A2(n_3068),
.B1(n_3003),
.B2(n_3009),
.Y(n_4432)
);

NOR3xp33_ASAP7_75t_L g4433 ( 
.A(n_3878),
.B(n_3216),
.C(n_3145),
.Y(n_4433)
);

AOI22xp33_ASAP7_75t_L g4434 ( 
.A1(n_3689),
.A2(n_3162),
.B1(n_3207),
.B2(n_3210),
.Y(n_4434)
);

NAND2xp5_ASAP7_75t_SL g4435 ( 
.A(n_4017),
.B(n_3347),
.Y(n_4435)
);

NAND2xp5_ASAP7_75t_L g4436 ( 
.A(n_3973),
.B(n_3216),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_3910),
.Y(n_4437)
);

NAND2xp5_ASAP7_75t_L g4438 ( 
.A(n_3895),
.B(n_3069),
.Y(n_4438)
);

BUFx12f_ASAP7_75t_L g4439 ( 
.A(n_3931),
.Y(n_4439)
);

INVx4_ASAP7_75t_L g4440 ( 
.A(n_3931),
.Y(n_4440)
);

NAND2xp5_ASAP7_75t_SL g4441 ( 
.A(n_4014),
.B(n_3348),
.Y(n_4441)
);

INVxp33_ASAP7_75t_L g4442 ( 
.A(n_3655),
.Y(n_4442)
);

INVx1_ASAP7_75t_L g4443 ( 
.A(n_3915),
.Y(n_4443)
);

AND2x2_ASAP7_75t_L g4444 ( 
.A(n_3909),
.B(n_3075),
.Y(n_4444)
);

AND2x2_ASAP7_75t_L g4445 ( 
.A(n_3996),
.B(n_3075),
.Y(n_4445)
);

INVx2_ASAP7_75t_L g4446 ( 
.A(n_3919),
.Y(n_4446)
);

INVx1_ASAP7_75t_L g4447 ( 
.A(n_3920),
.Y(n_4447)
);

AND2x4_ASAP7_75t_L g4448 ( 
.A(n_3816),
.B(n_3348),
.Y(n_4448)
);

BUFx4f_ASAP7_75t_L g4449 ( 
.A(n_3926),
.Y(n_4449)
);

INVx2_ASAP7_75t_SL g4450 ( 
.A(n_3935),
.Y(n_4450)
);

INVx2_ASAP7_75t_L g4451 ( 
.A(n_3950),
.Y(n_4451)
);

INVx1_ASAP7_75t_L g4452 ( 
.A(n_3957),
.Y(n_4452)
);

AOI22xp33_ASAP7_75t_L g4453 ( 
.A1(n_3492),
.A2(n_3207),
.B1(n_3061),
.B2(n_3145),
.Y(n_4453)
);

INVx2_ASAP7_75t_SL g4454 ( 
.A(n_3961),
.Y(n_4454)
);

AOI22xp33_ASAP7_75t_L g4455 ( 
.A1(n_3964),
.A2(n_3061),
.B1(n_3151),
.B2(n_3133),
.Y(n_4455)
);

AND2x6_ASAP7_75t_L g4456 ( 
.A(n_3931),
.B(n_3354),
.Y(n_4456)
);

AND2x4_ASAP7_75t_L g4457 ( 
.A(n_3685),
.B(n_3354),
.Y(n_4457)
);

BUFx5_ASAP7_75t_L g4458 ( 
.A(n_3966),
.Y(n_4458)
);

INVx2_ASAP7_75t_L g4459 ( 
.A(n_3963),
.Y(n_4459)
);

NAND2x1p5_ASAP7_75t_L g4460 ( 
.A(n_3581),
.B(n_2965),
.Y(n_4460)
);

INVx5_ASAP7_75t_L g4461 ( 
.A(n_3966),
.Y(n_4461)
);

A2O1A1Ixp33_ASAP7_75t_L g4462 ( 
.A1(n_3868),
.A2(n_3411),
.B(n_3151),
.C(n_2998),
.Y(n_4462)
);

INVx2_ASAP7_75t_L g4463 ( 
.A(n_3998),
.Y(n_4463)
);

INVx4_ASAP7_75t_L g4464 ( 
.A(n_3966),
.Y(n_4464)
);

CKINVDCx5p33_ASAP7_75t_R g4465 ( 
.A(n_3761),
.Y(n_4465)
);

NOR2xp33_ASAP7_75t_L g4466 ( 
.A(n_3978),
.B(n_3995),
.Y(n_4466)
);

NAND2xp33_ASAP7_75t_L g4467 ( 
.A(n_3502),
.B(n_3371),
.Y(n_4467)
);

AOI22xp33_ASAP7_75t_L g4468 ( 
.A1(n_3726),
.A2(n_3666),
.B1(n_4015),
.B2(n_4013),
.Y(n_4468)
);

AOI22xp33_ASAP7_75t_L g4469 ( 
.A1(n_4031),
.A2(n_3061),
.B1(n_2998),
.B2(n_3025),
.Y(n_4469)
);

HB1xp67_ASAP7_75t_L g4470 ( 
.A(n_3873),
.Y(n_4470)
);

AND2x2_ASAP7_75t_L g4471 ( 
.A(n_3571),
.B(n_3240),
.Y(n_4471)
);

NOR2xp33_ASAP7_75t_L g4472 ( 
.A(n_4008),
.B(n_3087),
.Y(n_4472)
);

AND2x2_ASAP7_75t_L g4473 ( 
.A(n_3573),
.B(n_3240),
.Y(n_4473)
);

BUFx6f_ASAP7_75t_L g4474 ( 
.A(n_3991),
.Y(n_4474)
);

BUFx6f_ASAP7_75t_L g4475 ( 
.A(n_3991),
.Y(n_4475)
);

NOR2xp33_ASAP7_75t_L g4476 ( 
.A(n_3965),
.B(n_3087),
.Y(n_4476)
);

NAND2xp5_ASAP7_75t_SL g4477 ( 
.A(n_4014),
.B(n_3119),
.Y(n_4477)
);

BUFx8_ASAP7_75t_L g4478 ( 
.A(n_3991),
.Y(n_4478)
);

NOR2xp33_ASAP7_75t_L g4479 ( 
.A(n_3969),
.B(n_3119),
.Y(n_4479)
);

AOI21xp5_ASAP7_75t_L g4480 ( 
.A1(n_3874),
.A2(n_3025),
.B(n_2962),
.Y(n_4480)
);

AOI22xp5_ASAP7_75t_L g4481 ( 
.A1(n_3788),
.A2(n_3036),
.B1(n_3054),
.B2(n_2962),
.Y(n_4481)
);

INVx1_ASAP7_75t_L g4482 ( 
.A(n_3734),
.Y(n_4482)
);

INVx3_ASAP7_75t_L g4483 ( 
.A(n_3879),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_3736),
.Y(n_4484)
);

NAND2xp5_ASAP7_75t_L g4485 ( 
.A(n_3907),
.B(n_3036),
.Y(n_4485)
);

INVx3_ASAP7_75t_L g4486 ( 
.A(n_3879),
.Y(n_4486)
);

INVx2_ASAP7_75t_L g4487 ( 
.A(n_3633),
.Y(n_4487)
);

OAI21xp33_ASAP7_75t_SL g4488 ( 
.A1(n_3700),
.A2(n_3054),
.B(n_3391),
.Y(n_4488)
);

AOI21xp33_ASAP7_75t_L g4489 ( 
.A1(n_4022),
.A2(n_3003),
.B(n_2996),
.Y(n_4489)
);

INVx2_ASAP7_75t_L g4490 ( 
.A(n_3634),
.Y(n_4490)
);

INVx2_ASAP7_75t_SL g4491 ( 
.A(n_4001),
.Y(n_4491)
);

AND2x6_ASAP7_75t_SL g4492 ( 
.A(n_3593),
.B(n_3368),
.Y(n_4492)
);

AND2x4_ASAP7_75t_L g4493 ( 
.A(n_3612),
.B(n_3391),
.Y(n_4493)
);

NAND2xp5_ASAP7_75t_L g4494 ( 
.A(n_3912),
.B(n_2977),
.Y(n_4494)
);

NAND2xp5_ASAP7_75t_L g4495 ( 
.A(n_3913),
.B(n_2977),
.Y(n_4495)
);

OR2x4_ASAP7_75t_L g4496 ( 
.A(n_3875),
.B(n_2996),
.Y(n_4496)
);

NAND2xp5_ASAP7_75t_L g4497 ( 
.A(n_3914),
.B(n_2977),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_3916),
.B(n_3929),
.Y(n_4498)
);

INVx1_ASAP7_75t_L g4499 ( 
.A(n_3739),
.Y(n_4499)
);

O2A1O1Ixp33_ASAP7_75t_L g4500 ( 
.A1(n_4033),
.A2(n_3432),
.B(n_3406),
.C(n_162),
.Y(n_4500)
);

BUFx2_ASAP7_75t_L g4501 ( 
.A(n_3584),
.Y(n_4501)
);

INVx1_ASAP7_75t_L g4502 ( 
.A(n_3852),
.Y(n_4502)
);

OR2x6_ASAP7_75t_L g4503 ( 
.A(n_3944),
.B(n_2989),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_3861),
.Y(n_4504)
);

NAND2x1p5_ASAP7_75t_L g4505 ( 
.A(n_3479),
.B(n_2989),
.Y(n_4505)
);

INVx2_ASAP7_75t_L g4506 ( 
.A(n_3639),
.Y(n_4506)
);

AOI22xp33_ASAP7_75t_L g4507 ( 
.A1(n_4012),
.A2(n_3457),
.B1(n_3009),
.B2(n_3003),
.Y(n_4507)
);

INVx2_ASAP7_75t_L g4508 ( 
.A(n_3648),
.Y(n_4508)
);

INVx1_ASAP7_75t_L g4509 ( 
.A(n_3657),
.Y(n_4509)
);

INVx2_ASAP7_75t_L g4510 ( 
.A(n_3658),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_3932),
.B(n_2989),
.Y(n_4511)
);

NAND2xp5_ASAP7_75t_SL g4512 ( 
.A(n_4032),
.B(n_3009),
.Y(n_4512)
);

NOR2xp33_ASAP7_75t_L g4513 ( 
.A(n_3885),
.B(n_2991),
.Y(n_4513)
);

BUFx3_ASAP7_75t_L g4514 ( 
.A(n_4023),
.Y(n_4514)
);

NAND2xp5_ASAP7_75t_L g4515 ( 
.A(n_3934),
.B(n_2991),
.Y(n_4515)
);

INVxp67_ASAP7_75t_L g4516 ( 
.A(n_3584),
.Y(n_4516)
);

NAND2xp5_ASAP7_75t_L g4517 ( 
.A(n_3936),
.B(n_2991),
.Y(n_4517)
);

NAND2xp5_ASAP7_75t_L g4518 ( 
.A(n_3947),
.B(n_3949),
.Y(n_4518)
);

AND2x4_ASAP7_75t_L g4519 ( 
.A(n_4023),
.B(n_3457),
.Y(n_4519)
);

OR2x2_ASAP7_75t_L g4520 ( 
.A(n_3580),
.B(n_161),
.Y(n_4520)
);

AOI22xp5_ASAP7_75t_L g4521 ( 
.A1(n_4035),
.A2(n_3457),
.B1(n_3432),
.B2(n_3406),
.Y(n_4521)
);

NAND2xp5_ASAP7_75t_L g4522 ( 
.A(n_3952),
.B(n_162),
.Y(n_4522)
);

BUFx2_ASAP7_75t_L g4523 ( 
.A(n_3621),
.Y(n_4523)
);

NOR2xp33_ASAP7_75t_L g4524 ( 
.A(n_3888),
.B(n_163),
.Y(n_4524)
);

NAND2xp5_ASAP7_75t_SL g4525 ( 
.A(n_4032),
.B(n_3457),
.Y(n_4525)
);

NAND2xp5_ASAP7_75t_L g4526 ( 
.A(n_3959),
.B(n_163),
.Y(n_4526)
);

AOI22xp5_ASAP7_75t_L g4527 ( 
.A1(n_3785),
.A2(n_164),
.B1(n_165),
.B2(n_163),
.Y(n_4527)
);

BUFx2_ASAP7_75t_L g4528 ( 
.A(n_3621),
.Y(n_4528)
);

NOR3xp33_ASAP7_75t_SL g4529 ( 
.A(n_3532),
.B(n_1081),
.C(n_165),
.Y(n_4529)
);

INVx1_ASAP7_75t_L g4530 ( 
.A(n_3663),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_SL g4531 ( 
.A(n_3768),
.B(n_164),
.Y(n_4531)
);

BUFx2_ASAP7_75t_L g4532 ( 
.A(n_3887),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_3975),
.B(n_165),
.Y(n_4533)
);

INVx2_ASAP7_75t_L g4534 ( 
.A(n_3672),
.Y(n_4534)
);

AOI22xp33_ASAP7_75t_L g4535 ( 
.A1(n_3815),
.A2(n_167),
.B1(n_168),
.B2(n_166),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_SL g4536 ( 
.A(n_3768),
.B(n_166),
.Y(n_4536)
);

INVx2_ASAP7_75t_L g4537 ( 
.A(n_3673),
.Y(n_4537)
);

NAND2xp5_ASAP7_75t_L g4538 ( 
.A(n_3588),
.B(n_167),
.Y(n_4538)
);

INVx2_ASAP7_75t_SL g4539 ( 
.A(n_3985),
.Y(n_4539)
);

NOR2xp33_ASAP7_75t_L g4540 ( 
.A(n_3986),
.B(n_3994),
.Y(n_4540)
);

INVx3_ASAP7_75t_L g4541 ( 
.A(n_3676),
.Y(n_4541)
);

INVx1_ASAP7_75t_L g4542 ( 
.A(n_3679),
.Y(n_4542)
);

INVx1_ASAP7_75t_L g4543 ( 
.A(n_3683),
.Y(n_4543)
);

NAND2xp5_ASAP7_75t_L g4544 ( 
.A(n_3594),
.B(n_167),
.Y(n_4544)
);

NAND2xp5_ASAP7_75t_L g4545 ( 
.A(n_3501),
.B(n_168),
.Y(n_4545)
);

INVx3_ASAP7_75t_L g4546 ( 
.A(n_3686),
.Y(n_4546)
);

NOR2xp33_ASAP7_75t_L g4547 ( 
.A(n_3505),
.B(n_168),
.Y(n_4547)
);

BUFx6f_ASAP7_75t_L g4548 ( 
.A(n_3922),
.Y(n_4548)
);

NOR2xp33_ASAP7_75t_L g4549 ( 
.A(n_3511),
.B(n_169),
.Y(n_4549)
);

AND2x4_ASAP7_75t_L g4550 ( 
.A(n_3694),
.B(n_169),
.Y(n_4550)
);

INVx2_ASAP7_75t_L g4551 ( 
.A(n_3696),
.Y(n_4551)
);

NAND2xp5_ASAP7_75t_SL g4552 ( 
.A(n_3772),
.B(n_169),
.Y(n_4552)
);

OAI22xp5_ASAP7_75t_L g4553 ( 
.A1(n_3908),
.A2(n_171),
.B1(n_172),
.B2(n_170),
.Y(n_4553)
);

NAND2xp5_ASAP7_75t_L g4554 ( 
.A(n_3513),
.B(n_170),
.Y(n_4554)
);

BUFx2_ASAP7_75t_L g4555 ( 
.A(n_3697),
.Y(n_4555)
);

INVx2_ASAP7_75t_L g4556 ( 
.A(n_3699),
.Y(n_4556)
);

AND2x4_ASAP7_75t_L g4557 ( 
.A(n_3706),
.B(n_170),
.Y(n_4557)
);

OR2x6_ASAP7_75t_L g4558 ( 
.A(n_3810),
.B(n_171),
.Y(n_4558)
);

NAND2xp5_ASAP7_75t_L g4559 ( 
.A(n_3519),
.B(n_172),
.Y(n_4559)
);

NAND2xp5_ASAP7_75t_L g4560 ( 
.A(n_3528),
.B(n_172),
.Y(n_4560)
);

BUFx6f_ASAP7_75t_L g4561 ( 
.A(n_3482),
.Y(n_4561)
);

NOR2x1p5_ASAP7_75t_L g4562 ( 
.A(n_3772),
.B(n_173),
.Y(n_4562)
);

INVx2_ASAP7_75t_L g4563 ( 
.A(n_3707),
.Y(n_4563)
);

AND2x4_ASAP7_75t_L g4564 ( 
.A(n_3712),
.B(n_173),
.Y(n_4564)
);

INVx1_ASAP7_75t_L g4565 ( 
.A(n_3717),
.Y(n_4565)
);

NAND2xp5_ASAP7_75t_L g4566 ( 
.A(n_3537),
.B(n_173),
.Y(n_4566)
);

AOI22xp33_ASAP7_75t_L g4567 ( 
.A1(n_3690),
.A2(n_3691),
.B1(n_3733),
.B2(n_3709),
.Y(n_4567)
);

AOI22xp33_ASAP7_75t_SL g4568 ( 
.A1(n_3722),
.A2(n_175),
.B1(n_176),
.B2(n_174),
.Y(n_4568)
);

INVx1_ASAP7_75t_L g4569 ( 
.A(n_3725),
.Y(n_4569)
);

AOI22xp5_ASAP7_75t_L g4570 ( 
.A1(n_4004),
.A2(n_175),
.B1(n_176),
.B2(n_174),
.Y(n_4570)
);

CKINVDCx5p33_ASAP7_75t_R g4571 ( 
.A(n_3731),
.Y(n_4571)
);

NOR2xp33_ASAP7_75t_L g4572 ( 
.A(n_3539),
.B(n_3543),
.Y(n_4572)
);

NAND2xp33_ASAP7_75t_L g4573 ( 
.A(n_3692),
.B(n_175),
.Y(n_4573)
);

AND2x4_ASAP7_75t_L g4574 ( 
.A(n_3776),
.B(n_176),
.Y(n_4574)
);

NAND2xp5_ASAP7_75t_L g4575 ( 
.A(n_3544),
.B(n_177),
.Y(n_4575)
);

BUFx3_ASAP7_75t_L g4576 ( 
.A(n_3780),
.Y(n_4576)
);

INVx2_ASAP7_75t_L g4577 ( 
.A(n_3782),
.Y(n_4577)
);

AOI22xp33_ASAP7_75t_L g4578 ( 
.A1(n_3702),
.A2(n_179),
.B1(n_180),
.B2(n_178),
.Y(n_4578)
);

NAND2xp33_ASAP7_75t_L g4579 ( 
.A(n_3698),
.B(n_178),
.Y(n_4579)
);

HB1xp67_ASAP7_75t_L g4580 ( 
.A(n_3786),
.Y(n_4580)
);

INVxp67_ASAP7_75t_L g4581 ( 
.A(n_3800),
.Y(n_4581)
);

NAND2xp5_ASAP7_75t_L g4582 ( 
.A(n_3551),
.B(n_3555),
.Y(n_4582)
);

NAND2x1p5_ASAP7_75t_L g4583 ( 
.A(n_3494),
.B(n_183),
.Y(n_4583)
);

NAND2xp5_ASAP7_75t_SL g4584 ( 
.A(n_3864),
.B(n_179),
.Y(n_4584)
);

INVx1_ASAP7_75t_L g4585 ( 
.A(n_3808),
.Y(n_4585)
);

INVx4_ASAP7_75t_L g4586 ( 
.A(n_3499),
.Y(n_4586)
);

INVx2_ASAP7_75t_L g4587 ( 
.A(n_3817),
.Y(n_4587)
);

AND2x4_ASAP7_75t_L g4588 ( 
.A(n_3820),
.B(n_180),
.Y(n_4588)
);

BUFx3_ASAP7_75t_L g4589 ( 
.A(n_3821),
.Y(n_4589)
);

NAND2xp5_ASAP7_75t_SL g4590 ( 
.A(n_3504),
.B(n_180),
.Y(n_4590)
);

INVx4_ASAP7_75t_L g4591 ( 
.A(n_3506),
.Y(n_4591)
);

NAND2xp5_ASAP7_75t_L g4592 ( 
.A(n_3556),
.B(n_181),
.Y(n_4592)
);

CKINVDCx6p67_ASAP7_75t_R g4593 ( 
.A(n_3659),
.Y(n_4593)
);

INVx1_ASAP7_75t_L g4594 ( 
.A(n_3827),
.Y(n_4594)
);

NOR2x1p5_ASAP7_75t_L g4595 ( 
.A(n_3833),
.B(n_181),
.Y(n_4595)
);

NAND2xp5_ASAP7_75t_L g4596 ( 
.A(n_3836),
.B(n_181),
.Y(n_4596)
);

INVx1_ASAP7_75t_L g4597 ( 
.A(n_3838),
.Y(n_4597)
);

NAND2xp5_ASAP7_75t_L g4598 ( 
.A(n_3841),
.B(n_182),
.Y(n_4598)
);

NAND2xp5_ASAP7_75t_L g4599 ( 
.A(n_3848),
.B(n_182),
.Y(n_4599)
);

AND2x4_ASAP7_75t_SL g4600 ( 
.A(n_3606),
.B(n_183),
.Y(n_4600)
);

AND2x4_ASAP7_75t_L g4601 ( 
.A(n_3710),
.B(n_184),
.Y(n_4601)
);

INVx5_ASAP7_75t_L g4602 ( 
.A(n_3518),
.Y(n_4602)
);

NAND2xp5_ASAP7_75t_L g4603 ( 
.A(n_3568),
.B(n_184),
.Y(n_4603)
);

INVx2_ASAP7_75t_SL g4604 ( 
.A(n_4075),
.Y(n_4604)
);

AND2x2_ASAP7_75t_L g4605 ( 
.A(n_4064),
.B(n_4053),
.Y(n_4605)
);

NAND2xp5_ASAP7_75t_SL g4606 ( 
.A(n_4133),
.B(n_3806),
.Y(n_4606)
);

AOI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_4312),
.A2(n_3560),
.B(n_3554),
.Y(n_4607)
);

AND2x2_ASAP7_75t_L g4608 ( 
.A(n_4054),
.B(n_4139),
.Y(n_4608)
);

NAND2xp5_ASAP7_75t_SL g4609 ( 
.A(n_4239),
.B(n_3834),
.Y(n_4609)
);

AOI21x1_ASAP7_75t_L g4610 ( 
.A1(n_4312),
.A2(n_3522),
.B(n_3586),
.Y(n_4610)
);

INVx2_ASAP7_75t_L g4611 ( 
.A(n_4381),
.Y(n_4611)
);

INVx1_ASAP7_75t_L g4612 ( 
.A(n_4181),
.Y(n_4612)
);

NAND2xp5_ASAP7_75t_L g4613 ( 
.A(n_4060),
.B(n_3608),
.Y(n_4613)
);

AOI21xp5_ASAP7_75t_L g4614 ( 
.A1(n_4414),
.A2(n_3570),
.B(n_3599),
.Y(n_4614)
);

NAND2xp5_ASAP7_75t_SL g4615 ( 
.A(n_4239),
.B(n_3662),
.Y(n_4615)
);

OR2x6_ASAP7_75t_SL g4616 ( 
.A(n_4230),
.B(n_3622),
.Y(n_4616)
);

NAND2xp5_ASAP7_75t_L g4617 ( 
.A(n_4502),
.B(n_3628),
.Y(n_4617)
);

AOI21xp5_ASAP7_75t_L g4618 ( 
.A1(n_4348),
.A2(n_3626),
.B(n_3611),
.Y(n_4618)
);

O2A1O1Ixp5_ASAP7_75t_L g4619 ( 
.A1(n_4348),
.A2(n_3865),
.B(n_3877),
.C(n_3854),
.Y(n_4619)
);

INVx1_ASAP7_75t_L g4620 ( 
.A(n_4038),
.Y(n_4620)
);

NAND2xp5_ASAP7_75t_L g4621 ( 
.A(n_4504),
.B(n_3631),
.Y(n_4621)
);

NAND2xp5_ASAP7_75t_L g4622 ( 
.A(n_4091),
.B(n_3830),
.Y(n_4622)
);

OAI21xp5_ASAP7_75t_L g4623 ( 
.A1(n_4214),
.A2(n_4005),
.B(n_3625),
.Y(n_4623)
);

AOI21xp5_ASAP7_75t_L g4624 ( 
.A1(n_4332),
.A2(n_3640),
.B(n_3627),
.Y(n_4624)
);

AND2x2_ASAP7_75t_L g4625 ( 
.A(n_4193),
.B(n_4198),
.Y(n_4625)
);

NAND2xp5_ASAP7_75t_L g4626 ( 
.A(n_4090),
.B(n_3488),
.Y(n_4626)
);

OAI21xp5_ASAP7_75t_L g4627 ( 
.A1(n_4116),
.A2(n_3632),
.B(n_3714),
.Y(n_4627)
);

NAND2x1_ASAP7_75t_L g4628 ( 
.A(n_4265),
.B(n_3524),
.Y(n_4628)
);

BUFx6f_ASAP7_75t_L g4629 ( 
.A(n_4073),
.Y(n_4629)
);

NAND2xp5_ASAP7_75t_SL g4630 ( 
.A(n_4239),
.B(n_3962),
.Y(n_4630)
);

NAND2xp5_ASAP7_75t_SL g4631 ( 
.A(n_4228),
.B(n_3972),
.Y(n_4631)
);

OR2x6_ASAP7_75t_L g4632 ( 
.A(n_4131),
.B(n_3990),
.Y(n_4632)
);

HB1xp67_ASAP7_75t_L g4633 ( 
.A(n_4407),
.Y(n_4633)
);

BUFx6f_ASAP7_75t_L g4634 ( 
.A(n_4073),
.Y(n_4634)
);

AOI21xp5_ASAP7_75t_L g4635 ( 
.A1(n_4467),
.A2(n_3524),
.B(n_3738),
.Y(n_4635)
);

NAND2xp5_ASAP7_75t_L g4636 ( 
.A(n_4186),
.B(n_3796),
.Y(n_4636)
);

NOR2xp67_ASAP7_75t_L g4637 ( 
.A(n_4075),
.B(n_189),
.Y(n_4637)
);

AOI21xp5_ASAP7_75t_L g4638 ( 
.A1(n_4142),
.A2(n_3757),
.B(n_3754),
.Y(n_4638)
);

NAND2xp5_ASAP7_75t_L g4639 ( 
.A(n_4043),
.B(n_3846),
.Y(n_4639)
);

NAND2xp5_ASAP7_75t_L g4640 ( 
.A(n_4045),
.B(n_3847),
.Y(n_4640)
);

BUFx2_ASAP7_75t_L g4641 ( 
.A(n_4242),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4050),
.Y(n_4642)
);

A2O1A1Ixp33_ASAP7_75t_L g4643 ( 
.A1(n_4500),
.A2(n_3774),
.B(n_3802),
.C(n_3762),
.Y(n_4643)
);

NAND2xp5_ASAP7_75t_L g4644 ( 
.A(n_4057),
.B(n_3921),
.Y(n_4644)
);

O2A1O1Ixp5_ASAP7_75t_L g4645 ( 
.A1(n_4525),
.A2(n_3927),
.B(n_3938),
.C(n_3924),
.Y(n_4645)
);

AOI22xp33_ASAP7_75t_L g4646 ( 
.A1(n_4212),
.A2(n_3851),
.B1(n_3893),
.B2(n_3813),
.Y(n_4646)
);

O2A1O1Ixp5_ASAP7_75t_L g4647 ( 
.A1(n_4345),
.A2(n_3939),
.B(n_3940),
.C(n_3911),
.Y(n_4647)
);

NAND2xp5_ASAP7_75t_L g4648 ( 
.A(n_4061),
.B(n_185),
.Y(n_4648)
);

NOR2xp33_ASAP7_75t_SL g4649 ( 
.A(n_4075),
.B(n_1070),
.Y(n_4649)
);

NAND2xp5_ASAP7_75t_L g4650 ( 
.A(n_4070),
.B(n_185),
.Y(n_4650)
);

NAND2xp5_ASAP7_75t_L g4651 ( 
.A(n_4087),
.B(n_186),
.Y(n_4651)
);

AOI22xp5_ASAP7_75t_L g4652 ( 
.A1(n_4124),
.A2(n_4044),
.B1(n_4232),
.B2(n_4071),
.Y(n_4652)
);

AOI21x1_ASAP7_75t_L g4653 ( 
.A1(n_4112),
.A2(n_187),
.B(n_186),
.Y(n_4653)
);

NOR2xp33_ASAP7_75t_L g4654 ( 
.A(n_4097),
.B(n_187),
.Y(n_4654)
);

AOI21xp5_ASAP7_75t_L g4655 ( 
.A1(n_4149),
.A2(n_188),
.B(n_187),
.Y(n_4655)
);

NOR2x1_ASAP7_75t_L g4656 ( 
.A(n_4146),
.B(n_188),
.Y(n_4656)
);

OR2x2_ASAP7_75t_L g4657 ( 
.A(n_4234),
.B(n_188),
.Y(n_4657)
);

O2A1O1Ixp33_ASAP7_75t_L g4658 ( 
.A1(n_4226),
.A2(n_190),
.B(n_191),
.C(n_189),
.Y(n_4658)
);

A2O1A1Ixp33_ASAP7_75t_L g4659 ( 
.A1(n_4121),
.A2(n_190),
.B(n_191),
.C(n_189),
.Y(n_4659)
);

NOR2xp33_ASAP7_75t_L g4660 ( 
.A(n_4442),
.B(n_190),
.Y(n_4660)
);

NAND2xp5_ASAP7_75t_L g4661 ( 
.A(n_4089),
.B(n_192),
.Y(n_4661)
);

OAI21xp5_ASAP7_75t_L g4662 ( 
.A1(n_4219),
.A2(n_193),
.B(n_192),
.Y(n_4662)
);

AOI21x1_ASAP7_75t_L g4663 ( 
.A1(n_4078),
.A2(n_194),
.B(n_192),
.Y(n_4663)
);

OAI21xp5_ASAP7_75t_L g4664 ( 
.A1(n_4531),
.A2(n_195),
.B(n_194),
.Y(n_4664)
);

INVx2_ASAP7_75t_L g4665 ( 
.A(n_4392),
.Y(n_4665)
);

NAND2xp5_ASAP7_75t_L g4666 ( 
.A(n_4099),
.B(n_194),
.Y(n_4666)
);

OAI21xp5_ASAP7_75t_L g4667 ( 
.A1(n_4536),
.A2(n_196),
.B(n_195),
.Y(n_4667)
);

AOI21xp5_ASAP7_75t_L g4668 ( 
.A1(n_4268),
.A2(n_197),
.B(n_196),
.Y(n_4668)
);

O2A1O1Ixp33_ASAP7_75t_L g4669 ( 
.A1(n_4062),
.A2(n_197),
.B(n_198),
.C(n_196),
.Y(n_4669)
);

AOI21x1_ASAP7_75t_L g4670 ( 
.A1(n_4477),
.A2(n_199),
.B(n_198),
.Y(n_4670)
);

NAND2xp5_ASAP7_75t_L g4671 ( 
.A(n_4101),
.B(n_198),
.Y(n_4671)
);

AOI21xp5_ASAP7_75t_L g4672 ( 
.A1(n_4277),
.A2(n_200),
.B(n_199),
.Y(n_4672)
);

BUFx6f_ASAP7_75t_L g4673 ( 
.A(n_4073),
.Y(n_4673)
);

NOR2xp33_ASAP7_75t_L g4674 ( 
.A(n_4571),
.B(n_199),
.Y(n_4674)
);

NAND3xp33_ASAP7_75t_L g4675 ( 
.A(n_4516),
.B(n_201),
.C(n_200),
.Y(n_4675)
);

NAND2xp5_ASAP7_75t_L g4676 ( 
.A(n_4103),
.B(n_200),
.Y(n_4676)
);

BUFx2_ASAP7_75t_L g4677 ( 
.A(n_4478),
.Y(n_4677)
);

AOI21xp5_ASAP7_75t_L g4678 ( 
.A1(n_4109),
.A2(n_4065),
.B(n_4111),
.Y(n_4678)
);

AOI21xp5_ASAP7_75t_L g4679 ( 
.A1(n_4350),
.A2(n_202),
.B(n_201),
.Y(n_4679)
);

NAND2xp5_ASAP7_75t_L g4680 ( 
.A(n_4107),
.B(n_201),
.Y(n_4680)
);

HB1xp67_ASAP7_75t_L g4681 ( 
.A(n_4262),
.Y(n_4681)
);

INVxp67_ASAP7_75t_L g4682 ( 
.A(n_4151),
.Y(n_4682)
);

NAND2xp5_ASAP7_75t_SL g4683 ( 
.A(n_4298),
.B(n_202),
.Y(n_4683)
);

OAI22xp5_ASAP7_75t_L g4684 ( 
.A1(n_4131),
.A2(n_4595),
.B1(n_4105),
.B2(n_4503),
.Y(n_4684)
);

OAI321xp33_ASAP7_75t_L g4685 ( 
.A1(n_4279),
.A2(n_3),
.A3(n_5),
.B1(n_1),
.B2(n_2),
.C(n_4),
.Y(n_4685)
);

AOI21xp5_ASAP7_75t_L g4686 ( 
.A1(n_4340),
.A2(n_203),
.B(n_202),
.Y(n_4686)
);

NAND2xp5_ASAP7_75t_L g4687 ( 
.A(n_4134),
.B(n_4145),
.Y(n_4687)
);

NAND2xp5_ASAP7_75t_SL g4688 ( 
.A(n_4094),
.B(n_204),
.Y(n_4688)
);

AOI21x1_ASAP7_75t_L g4689 ( 
.A1(n_4357),
.A2(n_205),
.B(n_204),
.Y(n_4689)
);

AOI21xp5_ASAP7_75t_L g4690 ( 
.A1(n_4405),
.A2(n_205),
.B(n_204),
.Y(n_4690)
);

OAI21xp33_ASAP7_75t_L g4691 ( 
.A1(n_4386),
.A2(n_206),
.B(n_205),
.Y(n_4691)
);

OAI21xp5_ASAP7_75t_L g4692 ( 
.A1(n_4552),
.A2(n_207),
.B(n_206),
.Y(n_4692)
);

AND2x2_ASAP7_75t_L g4693 ( 
.A(n_4429),
.B(n_206),
.Y(n_4693)
);

A2O1A1Ixp33_ASAP7_75t_L g4694 ( 
.A1(n_4223),
.A2(n_208),
.B(n_209),
.C(n_207),
.Y(n_4694)
);

INVx3_ASAP7_75t_L g4695 ( 
.A(n_4076),
.Y(n_4695)
);

INVx1_ASAP7_75t_L g4696 ( 
.A(n_4148),
.Y(n_4696)
);

INVx1_ASAP7_75t_L g4697 ( 
.A(n_4150),
.Y(n_4697)
);

OAI321xp33_ASAP7_75t_L g4698 ( 
.A1(n_4432),
.A2(n_3),
.A3(n_5),
.B1(n_1),
.B2(n_2),
.C(n_4),
.Y(n_4698)
);

O2A1O1Ixp5_ASAP7_75t_L g4699 ( 
.A1(n_4160),
.A2(n_208),
.B(n_209),
.C(n_207),
.Y(n_4699)
);

AND2x2_ASAP7_75t_L g4700 ( 
.A(n_4173),
.B(n_208),
.Y(n_4700)
);

AOI21xp5_ASAP7_75t_L g4701 ( 
.A1(n_4441),
.A2(n_210),
.B(n_209),
.Y(n_4701)
);

AND2x2_ASAP7_75t_L g4702 ( 
.A(n_4349),
.B(n_210),
.Y(n_4702)
);

INVx1_ASAP7_75t_L g4703 ( 
.A(n_4153),
.Y(n_4703)
);

O2A1O1Ixp33_ASAP7_75t_L g4704 ( 
.A1(n_4138),
.A2(n_212),
.B(n_213),
.C(n_211),
.Y(n_4704)
);

OAI22xp5_ASAP7_75t_L g4705 ( 
.A1(n_4503),
.A2(n_212),
.B1(n_213),
.B2(n_211),
.Y(n_4705)
);

AOI21xp5_ASAP7_75t_L g4706 ( 
.A1(n_4382),
.A2(n_212),
.B(n_211),
.Y(n_4706)
);

NAND2xp5_ASAP7_75t_L g4707 ( 
.A(n_4161),
.B(n_213),
.Y(n_4707)
);

A2O1A1Ixp33_ASAP7_75t_L g4708 ( 
.A1(n_4529),
.A2(n_215),
.B(n_216),
.C(n_214),
.Y(n_4708)
);

AOI21xp5_ASAP7_75t_L g4709 ( 
.A1(n_4177),
.A2(n_215),
.B(n_214),
.Y(n_4709)
);

BUFx3_ASAP7_75t_L g4710 ( 
.A(n_4079),
.Y(n_4710)
);

CKINVDCx10_ASAP7_75t_R g4711 ( 
.A(n_4273),
.Y(n_4711)
);

O2A1O1Ixp33_ASAP7_75t_L g4712 ( 
.A1(n_4140),
.A2(n_216),
.B(n_217),
.C(n_214),
.Y(n_4712)
);

NOR2xp33_ASAP7_75t_R g4713 ( 
.A(n_4187),
.B(n_1072),
.Y(n_4713)
);

NAND2xp5_ASAP7_75t_L g4714 ( 
.A(n_4163),
.B(n_217),
.Y(n_4714)
);

OAI22xp5_ASAP7_75t_L g4715 ( 
.A1(n_4174),
.A2(n_219),
.B1(n_220),
.B2(n_218),
.Y(n_4715)
);

NAND2x1p5_ASAP7_75t_L g4716 ( 
.A(n_4106),
.B(n_4211),
.Y(n_4716)
);

BUFx6f_ASAP7_75t_L g4717 ( 
.A(n_4431),
.Y(n_4717)
);

NAND2xp5_ASAP7_75t_L g4718 ( 
.A(n_4167),
.B(n_4178),
.Y(n_4718)
);

NAND2xp5_ASAP7_75t_L g4719 ( 
.A(n_4180),
.B(n_218),
.Y(n_4719)
);

INVx3_ASAP7_75t_L g4720 ( 
.A(n_4076),
.Y(n_4720)
);

CKINVDCx6p67_ASAP7_75t_R g4721 ( 
.A(n_4120),
.Y(n_4721)
);

AOI21xp5_ASAP7_75t_L g4722 ( 
.A1(n_4185),
.A2(n_220),
.B(n_219),
.Y(n_4722)
);

AOI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4501),
.A2(n_221),
.B(n_219),
.Y(n_4723)
);

OAI22xp5_ASAP7_75t_L g4724 ( 
.A1(n_4041),
.A2(n_222),
.B1(n_223),
.B2(n_221),
.Y(n_4724)
);

OAI21xp5_ASAP7_75t_L g4725 ( 
.A1(n_4584),
.A2(n_223),
.B(n_222),
.Y(n_4725)
);

NOR2xp33_ASAP7_75t_L g4726 ( 
.A(n_4288),
.B(n_4398),
.Y(n_4726)
);

AOI22xp5_ASAP7_75t_L g4727 ( 
.A1(n_4068),
.A2(n_1079),
.B1(n_1080),
.B2(n_1078),
.Y(n_4727)
);

NAND2xp5_ASAP7_75t_L g4728 ( 
.A(n_4184),
.B(n_222),
.Y(n_4728)
);

NOR2xp67_ASAP7_75t_SL g4729 ( 
.A(n_4069),
.B(n_223),
.Y(n_4729)
);

NOR2xp67_ASAP7_75t_SL g4730 ( 
.A(n_4069),
.B(n_224),
.Y(n_4730)
);

AOI21xp5_ASAP7_75t_L g4731 ( 
.A1(n_4215),
.A2(n_225),
.B(n_224),
.Y(n_4731)
);

BUFx3_ASAP7_75t_L g4732 ( 
.A(n_4128),
.Y(n_4732)
);

AOI22xp5_ASAP7_75t_L g4733 ( 
.A1(n_4572),
.A2(n_226),
.B1(n_227),
.B2(n_225),
.Y(n_4733)
);

AOI21xp5_ASAP7_75t_L g4734 ( 
.A1(n_4308),
.A2(n_226),
.B(n_225),
.Y(n_4734)
);

OAI22xp5_ASAP7_75t_L g4735 ( 
.A1(n_4117),
.A2(n_227),
.B1(n_228),
.B2(n_226),
.Y(n_4735)
);

NAND2xp33_ASAP7_75t_SL g4736 ( 
.A(n_4562),
.B(n_228),
.Y(n_4736)
);

AOI21xp5_ASAP7_75t_L g4737 ( 
.A1(n_4325),
.A2(n_230),
.B(n_229),
.Y(n_4737)
);

AOI22xp5_ASAP7_75t_L g4738 ( 
.A1(n_4311),
.A2(n_1070),
.B1(n_1071),
.B2(n_1069),
.Y(n_4738)
);

NAND3xp33_ASAP7_75t_SL g4739 ( 
.A(n_4313),
.B(n_4),
.C(n_5),
.Y(n_4739)
);

AOI21xp5_ASAP7_75t_L g4740 ( 
.A1(n_4189),
.A2(n_231),
.B(n_230),
.Y(n_4740)
);

INVxp67_ASAP7_75t_SL g4741 ( 
.A(n_4316),
.Y(n_4741)
);

NAND2xp5_ASAP7_75t_L g4742 ( 
.A(n_4188),
.B(n_4194),
.Y(n_4742)
);

NAND2xp5_ASAP7_75t_SL g4743 ( 
.A(n_4094),
.B(n_231),
.Y(n_4743)
);

AOI21xp5_ASAP7_75t_L g4744 ( 
.A1(n_4205),
.A2(n_232),
.B(n_231),
.Y(n_4744)
);

NOR2x1_ASAP7_75t_L g4745 ( 
.A(n_4122),
.B(n_232),
.Y(n_4745)
);

OAI21xp5_ASAP7_75t_L g4746 ( 
.A1(n_4067),
.A2(n_234),
.B(n_233),
.Y(n_4746)
);

NAND3xp33_ASAP7_75t_L g4747 ( 
.A(n_4466),
.B(n_234),
.C(n_233),
.Y(n_4747)
);

NAND2xp5_ASAP7_75t_L g4748 ( 
.A(n_4196),
.B(n_233),
.Y(n_4748)
);

NAND2xp5_ASAP7_75t_SL g4749 ( 
.A(n_4122),
.B(n_235),
.Y(n_4749)
);

AOI21xp5_ASAP7_75t_L g4750 ( 
.A1(n_4488),
.A2(n_236),
.B(n_235),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4393),
.Y(n_4751)
);

NAND2xp5_ASAP7_75t_L g4752 ( 
.A(n_4207),
.B(n_236),
.Y(n_4752)
);

INVx1_ASAP7_75t_L g4753 ( 
.A(n_4218),
.Y(n_4753)
);

NAND2xp5_ASAP7_75t_L g4754 ( 
.A(n_4227),
.B(n_236),
.Y(n_4754)
);

NAND2xp5_ASAP7_75t_L g4755 ( 
.A(n_4238),
.B(n_4253),
.Y(n_4755)
);

OAI21x1_ASAP7_75t_L g4756 ( 
.A1(n_4314),
.A2(n_238),
.B(n_237),
.Y(n_4756)
);

OR2x6_ASAP7_75t_SL g4757 ( 
.A(n_4267),
.B(n_1078),
.Y(n_4757)
);

NOR2xp33_ASAP7_75t_SL g4758 ( 
.A(n_4115),
.B(n_1081),
.Y(n_4758)
);

O2A1O1Ixp33_ASAP7_75t_L g4759 ( 
.A1(n_4241),
.A2(n_238),
.B(n_239),
.C(n_237),
.Y(n_4759)
);

NAND2xp5_ASAP7_75t_L g4760 ( 
.A(n_4256),
.B(n_237),
.Y(n_4760)
);

AOI22xp33_ASAP7_75t_L g4761 ( 
.A1(n_4523),
.A2(n_4528),
.B1(n_4589),
.B2(n_4576),
.Y(n_4761)
);

INVx1_ASAP7_75t_L g4762 ( 
.A(n_4257),
.Y(n_4762)
);

AOI21xp5_ASAP7_75t_L g4763 ( 
.A1(n_4480),
.A2(n_240),
.B(n_239),
.Y(n_4763)
);

AOI21xp5_ASAP7_75t_L g4764 ( 
.A1(n_4229),
.A2(n_240),
.B(n_239),
.Y(n_4764)
);

NOR2xp33_ASAP7_75t_L g4765 ( 
.A(n_4400),
.B(n_240),
.Y(n_4765)
);

OAI21xp5_ASAP7_75t_L g4766 ( 
.A1(n_4310),
.A2(n_242),
.B(n_241),
.Y(n_4766)
);

AOI21xp33_ASAP7_75t_L g4767 ( 
.A1(n_4498),
.A2(n_243),
.B(n_242),
.Y(n_4767)
);

BUFx2_ASAP7_75t_L g4768 ( 
.A(n_4478),
.Y(n_4768)
);

NAND2x1p5_ASAP7_75t_L g4769 ( 
.A(n_4159),
.B(n_4074),
.Y(n_4769)
);

AOI21xp5_ASAP7_75t_L g4770 ( 
.A1(n_4135),
.A2(n_243),
.B(n_242),
.Y(n_4770)
);

INVx1_ASAP7_75t_L g4771 ( 
.A(n_4259),
.Y(n_4771)
);

NAND3xp33_ASAP7_75t_SL g4772 ( 
.A(n_4394),
.B(n_4),
.C(n_5),
.Y(n_4772)
);

AOI221xp5_ASAP7_75t_L g4773 ( 
.A1(n_4547),
.A2(n_246),
.B1(n_247),
.B2(n_245),
.C(n_244),
.Y(n_4773)
);

OAI21xp33_ASAP7_75t_L g4774 ( 
.A1(n_4377),
.A2(n_245),
.B(n_244),
.Y(n_4774)
);

CKINVDCx5p33_ASAP7_75t_R g4775 ( 
.A(n_4155),
.Y(n_4775)
);

INVx1_ASAP7_75t_L g4776 ( 
.A(n_4260),
.Y(n_4776)
);

O2A1O1Ixp33_ASAP7_75t_SL g4777 ( 
.A1(n_4063),
.A2(n_245),
.B(n_246),
.C(n_244),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_SL g4778 ( 
.A(n_4469),
.B(n_247),
.Y(n_4778)
);

AOI21xp5_ASAP7_75t_L g4779 ( 
.A1(n_4389),
.A2(n_249),
.B(n_248),
.Y(n_4779)
);

AOI21xp5_ASAP7_75t_L g4780 ( 
.A1(n_4240),
.A2(n_4418),
.B(n_4462),
.Y(n_4780)
);

NAND2xp5_ASAP7_75t_L g4781 ( 
.A(n_4285),
.B(n_248),
.Y(n_4781)
);

INVx2_ASAP7_75t_L g4782 ( 
.A(n_4395),
.Y(n_4782)
);

NOR2xp33_ASAP7_75t_L g4783 ( 
.A(n_4404),
.B(n_249),
.Y(n_4783)
);

AOI21xp5_ASAP7_75t_L g4784 ( 
.A1(n_4240),
.A2(n_251),
.B(n_250),
.Y(n_4784)
);

NAND2xp5_ASAP7_75t_L g4785 ( 
.A(n_4289),
.B(n_251),
.Y(n_4785)
);

NAND2xp5_ASAP7_75t_L g4786 ( 
.A(n_4294),
.B(n_252),
.Y(n_4786)
);

AOI21xp5_ASAP7_75t_L g4787 ( 
.A1(n_4272),
.A2(n_254),
.B(n_253),
.Y(n_4787)
);

AND2x4_ASAP7_75t_L g4788 ( 
.A(n_4246),
.B(n_254),
.Y(n_4788)
);

AND2x4_ASAP7_75t_L g4789 ( 
.A(n_4246),
.B(n_4251),
.Y(n_4789)
);

AND2x2_ASAP7_75t_L g4790 ( 
.A(n_4397),
.B(n_255),
.Y(n_4790)
);

INVx3_ASAP7_75t_L g4791 ( 
.A(n_4080),
.Y(n_4791)
);

NOR2xp33_ASAP7_75t_L g4792 ( 
.A(n_4245),
.B(n_255),
.Y(n_4792)
);

AND2x4_ASAP7_75t_L g4793 ( 
.A(n_4251),
.B(n_4303),
.Y(n_4793)
);

AOI21xp5_ASAP7_75t_L g4794 ( 
.A1(n_4410),
.A2(n_256),
.B(n_255),
.Y(n_4794)
);

AOI22xp5_ASAP7_75t_L g4795 ( 
.A1(n_4254),
.A2(n_4423),
.B1(n_4540),
.B2(n_4237),
.Y(n_4795)
);

NOR2xp33_ASAP7_75t_SL g4796 ( 
.A(n_4118),
.B(n_1066),
.Y(n_4796)
);

INVx1_ASAP7_75t_L g4797 ( 
.A(n_4323),
.Y(n_4797)
);

AND2x2_ASAP7_75t_SL g4798 ( 
.A(n_4449),
.B(n_256),
.Y(n_4798)
);

NAND2xp5_ASAP7_75t_L g4799 ( 
.A(n_4329),
.B(n_256),
.Y(n_4799)
);

AOI21xp5_ASAP7_75t_L g4800 ( 
.A1(n_4086),
.A2(n_258),
.B(n_257),
.Y(n_4800)
);

NAND2xp5_ASAP7_75t_L g4801 ( 
.A(n_4334),
.B(n_257),
.Y(n_4801)
);

O2A1O1Ixp33_ASAP7_75t_SL g4802 ( 
.A1(n_4055),
.A2(n_258),
.B(n_259),
.C(n_257),
.Y(n_4802)
);

NAND2xp5_ASAP7_75t_SL g4803 ( 
.A(n_4104),
.B(n_258),
.Y(n_4803)
);

AOI21x1_ASAP7_75t_L g4804 ( 
.A1(n_4512),
.A2(n_260),
.B(n_259),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_SL g4805 ( 
.A(n_4080),
.B(n_260),
.Y(n_4805)
);

CKINVDCx16_ASAP7_75t_R g4806 ( 
.A(n_4170),
.Y(n_4806)
);

AOI22xp5_ASAP7_75t_L g4807 ( 
.A1(n_4125),
.A2(n_1072),
.B1(n_1074),
.B2(n_1071),
.Y(n_4807)
);

NAND2xp5_ASAP7_75t_L g4808 ( 
.A(n_4339),
.B(n_261),
.Y(n_4808)
);

AOI21xp5_ASAP7_75t_L g4809 ( 
.A1(n_4235),
.A2(n_262),
.B(n_261),
.Y(n_4809)
);

AND2x2_ASAP7_75t_SL g4810 ( 
.A(n_4082),
.B(n_262),
.Y(n_4810)
);

BUFx12f_ASAP7_75t_L g4811 ( 
.A(n_4046),
.Y(n_4811)
);

BUFx2_ASAP7_75t_L g4812 ( 
.A(n_4439),
.Y(n_4812)
);

O2A1O1Ixp33_ASAP7_75t_L g4813 ( 
.A1(n_4162),
.A2(n_263),
.B(n_264),
.C(n_262),
.Y(n_4813)
);

AOI21xp5_ASAP7_75t_L g4814 ( 
.A1(n_4236),
.A2(n_264),
.B(n_263),
.Y(n_4814)
);

O2A1O1Ixp33_ASAP7_75t_SL g4815 ( 
.A1(n_4521),
.A2(n_265),
.B(n_266),
.C(n_263),
.Y(n_4815)
);

OA22x2_ASAP7_75t_L g4816 ( 
.A1(n_4388),
.A2(n_266),
.B1(n_267),
.B2(n_265),
.Y(n_4816)
);

AND2x2_ASAP7_75t_L g4817 ( 
.A(n_4144),
.B(n_265),
.Y(n_4817)
);

OAI21xp5_ASAP7_75t_L g4818 ( 
.A1(n_4176),
.A2(n_268),
.B(n_267),
.Y(n_4818)
);

AOI21xp5_ASAP7_75t_L g4819 ( 
.A1(n_4284),
.A2(n_269),
.B(n_268),
.Y(n_4819)
);

OAI21xp5_ASAP7_75t_L g4820 ( 
.A1(n_4276),
.A2(n_269),
.B(n_268),
.Y(n_4820)
);

NAND2xp5_ASAP7_75t_L g4821 ( 
.A(n_4341),
.B(n_271),
.Y(n_4821)
);

AOI22xp5_ASAP7_75t_L g4822 ( 
.A1(n_4037),
.A2(n_1063),
.B1(n_1065),
.B2(n_1062),
.Y(n_4822)
);

NAND2xp5_ASAP7_75t_L g4823 ( 
.A(n_4346),
.B(n_271),
.Y(n_4823)
);

BUFx6f_ASAP7_75t_L g4824 ( 
.A(n_4074),
.Y(n_4824)
);

O2A1O1Ixp5_ASAP7_75t_L g4825 ( 
.A1(n_4586),
.A2(n_272),
.B(n_273),
.C(n_271),
.Y(n_4825)
);

A2O1A1Ixp33_ASAP7_75t_L g4826 ( 
.A1(n_4307),
.A2(n_273),
.B(n_274),
.C(n_272),
.Y(n_4826)
);

NAND2xp5_ASAP7_75t_L g4827 ( 
.A(n_4351),
.B(n_272),
.Y(n_4827)
);

BUFx8_ASAP7_75t_SL g4828 ( 
.A(n_4191),
.Y(n_4828)
);

AND2x2_ASAP7_75t_L g4829 ( 
.A(n_4333),
.B(n_273),
.Y(n_4829)
);

AND2x2_ASAP7_75t_L g4830 ( 
.A(n_4363),
.B(n_274),
.Y(n_4830)
);

AOI21xp5_ASAP7_75t_L g4831 ( 
.A1(n_4424),
.A2(n_275),
.B(n_274),
.Y(n_4831)
);

INVx4_ASAP7_75t_L g4832 ( 
.A(n_4110),
.Y(n_4832)
);

A2O1A1Ixp33_ASAP7_75t_L g4833 ( 
.A1(n_4573),
.A2(n_276),
.B(n_277),
.C(n_275),
.Y(n_4833)
);

NAND2xp5_ASAP7_75t_L g4834 ( 
.A(n_4352),
.B(n_277),
.Y(n_4834)
);

INVx1_ASAP7_75t_L g4835 ( 
.A(n_4355),
.Y(n_4835)
);

AOI21x1_ASAP7_75t_L g4836 ( 
.A1(n_4493),
.A2(n_279),
.B(n_278),
.Y(n_4836)
);

NAND2xp5_ASAP7_75t_L g4837 ( 
.A(n_4356),
.B(n_278),
.Y(n_4837)
);

NAND2xp5_ASAP7_75t_SL g4838 ( 
.A(n_4493),
.B(n_278),
.Y(n_4838)
);

CKINVDCx14_ASAP7_75t_R g4839 ( 
.A(n_4286),
.Y(n_4839)
);

NOR2xp33_ASAP7_75t_L g4840 ( 
.A(n_4465),
.B(n_279),
.Y(n_4840)
);

AND2x2_ASAP7_75t_L g4841 ( 
.A(n_4379),
.B(n_280),
.Y(n_4841)
);

NAND2xp5_ASAP7_75t_L g4842 ( 
.A(n_4360),
.B(n_4362),
.Y(n_4842)
);

NAND2x1p5_ASAP7_75t_L g4843 ( 
.A(n_4159),
.B(n_280),
.Y(n_4843)
);

AOI21xp5_ASAP7_75t_L g4844 ( 
.A1(n_4428),
.A2(n_281),
.B(n_280),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4365),
.Y(n_4845)
);

NOR2x1p5_ASAP7_75t_SL g4846 ( 
.A(n_4458),
.B(n_281),
.Y(n_4846)
);

NAND2xp5_ASAP7_75t_L g4847 ( 
.A(n_4366),
.B(n_4371),
.Y(n_4847)
);

O2A1O1Ixp33_ASAP7_75t_SL g4848 ( 
.A1(n_4093),
.A2(n_282),
.B(n_283),
.C(n_281),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_SL g4849 ( 
.A(n_4602),
.B(n_282),
.Y(n_4849)
);

NAND2xp5_ASAP7_75t_L g4850 ( 
.A(n_4372),
.B(n_282),
.Y(n_4850)
);

INVx1_ASAP7_75t_L g4851 ( 
.A(n_4195),
.Y(n_4851)
);

O2A1O1Ixp33_ASAP7_75t_L g4852 ( 
.A1(n_4518),
.A2(n_284),
.B(n_285),
.C(n_283),
.Y(n_4852)
);

OAI22xp5_ASAP7_75t_L g4853 ( 
.A1(n_4270),
.A2(n_285),
.B1(n_286),
.B2(n_284),
.Y(n_4853)
);

NAND2xp5_ASAP7_75t_SL g4854 ( 
.A(n_4602),
.B(n_284),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4183),
.Y(n_4855)
);

AND2x4_ASAP7_75t_L g4856 ( 
.A(n_4303),
.B(n_285),
.Y(n_4856)
);

BUFx12f_ASAP7_75t_SL g4857 ( 
.A(n_4273),
.Y(n_4857)
);

OAI21x1_ASAP7_75t_L g4858 ( 
.A1(n_4314),
.A2(n_287),
.B(n_286),
.Y(n_4858)
);

AOI21xp5_ASAP7_75t_L g4859 ( 
.A1(n_4435),
.A2(n_288),
.B(n_286),
.Y(n_4859)
);

NAND2xp5_ASAP7_75t_L g4860 ( 
.A(n_4482),
.B(n_288),
.Y(n_4860)
);

NAND2xp5_ASAP7_75t_L g4861 ( 
.A(n_4484),
.B(n_288),
.Y(n_4861)
);

AOI22xp5_ASAP7_75t_L g4862 ( 
.A1(n_4280),
.A2(n_1066),
.B1(n_1067),
.B2(n_1065),
.Y(n_4862)
);

OAI21x1_ASAP7_75t_L g4863 ( 
.A1(n_4342),
.A2(n_290),
.B(n_289),
.Y(n_4863)
);

NOR2xp33_ASAP7_75t_L g4864 ( 
.A(n_4401),
.B(n_289),
.Y(n_4864)
);

NAND2xp5_ASAP7_75t_L g4865 ( 
.A(n_4499),
.B(n_290),
.Y(n_4865)
);

BUFx2_ASAP7_75t_L g4866 ( 
.A(n_4496),
.Y(n_4866)
);

OAI22xp5_ASAP7_75t_L g4867 ( 
.A1(n_4270),
.A2(n_291),
.B1(n_292),
.B2(n_290),
.Y(n_4867)
);

NOR2xp33_ASAP7_75t_L g4868 ( 
.A(n_4095),
.B(n_291),
.Y(n_4868)
);

NAND2xp33_ASAP7_75t_L g4869 ( 
.A(n_4265),
.B(n_291),
.Y(n_4869)
);

OAI21x1_ASAP7_75t_L g4870 ( 
.A1(n_4342),
.A2(n_293),
.B(n_292),
.Y(n_4870)
);

AOI21xp5_ASAP7_75t_L g4871 ( 
.A1(n_4519),
.A2(n_293),
.B(n_292),
.Y(n_4871)
);

OAI321xp33_ASAP7_75t_L g4872 ( 
.A1(n_4527),
.A2(n_8),
.A3(n_10),
.B1(n_6),
.B2(n_7),
.C(n_9),
.Y(n_4872)
);

BUFx2_ASAP7_75t_L g4873 ( 
.A(n_4221),
.Y(n_4873)
);

NOR2x1p5_ASAP7_75t_SL g4874 ( 
.A(n_4458),
.B(n_294),
.Y(n_4874)
);

BUFx2_ASAP7_75t_L g4875 ( 
.A(n_4042),
.Y(n_4875)
);

NOR2xp33_ASAP7_75t_L g4876 ( 
.A(n_4049),
.B(n_294),
.Y(n_4876)
);

AOI21xp5_ASAP7_75t_L g4877 ( 
.A1(n_4519),
.A2(n_295),
.B(n_294),
.Y(n_4877)
);

INVx1_ASAP7_75t_L g4878 ( 
.A(n_4374),
.Y(n_4878)
);

AOI21xp5_ASAP7_75t_L g4879 ( 
.A1(n_4129),
.A2(n_296),
.B(n_295),
.Y(n_4879)
);

NAND2xp5_ASAP7_75t_SL g4880 ( 
.A(n_4602),
.B(n_295),
.Y(n_4880)
);

AOI22xp5_ASAP7_75t_L g4881 ( 
.A1(n_4199),
.A2(n_1077),
.B1(n_1079),
.B2(n_1076),
.Y(n_4881)
);

BUFx8_ASAP7_75t_L g4882 ( 
.A(n_4036),
.Y(n_4882)
);

NAND2xp5_ASAP7_75t_SL g4883 ( 
.A(n_4461),
.B(n_296),
.Y(n_4883)
);

NOR2xp33_ASAP7_75t_L g4884 ( 
.A(n_4072),
.B(n_296),
.Y(n_4884)
);

OAI22xp5_ASAP7_75t_L g4885 ( 
.A1(n_4283),
.A2(n_298),
.B1(n_299),
.B2(n_297),
.Y(n_4885)
);

AOI21xp5_ASAP7_75t_L g4886 ( 
.A1(n_4300),
.A2(n_299),
.B(n_298),
.Y(n_4886)
);

AOI21xp5_ASAP7_75t_L g4887 ( 
.A1(n_4579),
.A2(n_300),
.B(n_299),
.Y(n_4887)
);

INVx2_ASAP7_75t_L g4888 ( 
.A(n_4413),
.Y(n_4888)
);

NOR2xp33_ASAP7_75t_L g4889 ( 
.A(n_4168),
.B(n_300),
.Y(n_4889)
);

NAND2xp5_ASAP7_75t_L g4890 ( 
.A(n_4470),
.B(n_300),
.Y(n_4890)
);

INVx2_ASAP7_75t_L g4891 ( 
.A(n_4425),
.Y(n_4891)
);

AOI21xp5_ASAP7_75t_L g4892 ( 
.A1(n_4210),
.A2(n_4048),
.B(n_4047),
.Y(n_4892)
);

NOR2xp33_ASAP7_75t_L g4893 ( 
.A(n_4278),
.B(n_301),
.Y(n_4893)
);

CKINVDCx5p33_ASAP7_75t_R g4894 ( 
.A(n_4083),
.Y(n_4894)
);

NAND2xp5_ASAP7_75t_L g4895 ( 
.A(n_4509),
.B(n_301),
.Y(n_4895)
);

OAI21x1_ASAP7_75t_L g4896 ( 
.A1(n_4408),
.A2(n_302),
.B(n_301),
.Y(n_4896)
);

AOI22xp33_ASAP7_75t_L g4897 ( 
.A1(n_4204),
.A2(n_304),
.B1(n_305),
.B2(n_303),
.Y(n_4897)
);

AOI22xp33_ASAP7_75t_L g4898 ( 
.A1(n_4555),
.A2(n_306),
.B1(n_307),
.B2(n_305),
.Y(n_4898)
);

NAND2xp5_ASAP7_75t_L g4899 ( 
.A(n_4530),
.B(n_306),
.Y(n_4899)
);

OAI22xp5_ASAP7_75t_L g4900 ( 
.A1(n_4567),
.A2(n_308),
.B1(n_309),
.B2(n_306),
.Y(n_4900)
);

NAND2xp5_ASAP7_75t_L g4901 ( 
.A(n_4542),
.B(n_308),
.Y(n_4901)
);

AO22x1_ASAP7_75t_L g4902 ( 
.A1(n_4265),
.A2(n_310),
.B1(n_311),
.B2(n_309),
.Y(n_4902)
);

BUFx12f_ASAP7_75t_L g4903 ( 
.A(n_4039),
.Y(n_4903)
);

INVx2_ASAP7_75t_L g4904 ( 
.A(n_4208),
.Y(n_4904)
);

NOR2xp33_ASAP7_75t_L g4905 ( 
.A(n_4336),
.B(n_4052),
.Y(n_4905)
);

INVx2_ASAP7_75t_L g4906 ( 
.A(n_4248),
.Y(n_4906)
);

NOR2xp33_ASAP7_75t_L g4907 ( 
.A(n_4136),
.B(n_310),
.Y(n_4907)
);

NAND2xp5_ASAP7_75t_L g4908 ( 
.A(n_4543),
.B(n_310),
.Y(n_4908)
);

NOR2xp33_ASAP7_75t_L g4909 ( 
.A(n_4172),
.B(n_312),
.Y(n_4909)
);

NAND2xp5_ASAP7_75t_L g4910 ( 
.A(n_4565),
.B(n_313),
.Y(n_4910)
);

AOI21xp5_ASAP7_75t_L g4911 ( 
.A1(n_4051),
.A2(n_314),
.B(n_313),
.Y(n_4911)
);

BUFx2_ASAP7_75t_SL g4912 ( 
.A(n_4077),
.Y(n_4912)
);

NAND3xp33_ASAP7_75t_L g4913 ( 
.A(n_4568),
.B(n_315),
.C(n_314),
.Y(n_4913)
);

AOI21xp5_ASAP7_75t_L g4914 ( 
.A1(n_4058),
.A2(n_315),
.B(n_314),
.Y(n_4914)
);

OAI21xp33_ASAP7_75t_L g4915 ( 
.A1(n_4066),
.A2(n_316),
.B(n_315),
.Y(n_4915)
);

NAND2xp5_ASAP7_75t_SL g4916 ( 
.A(n_4461),
.B(n_317),
.Y(n_4916)
);

INVx2_ASAP7_75t_L g4917 ( 
.A(n_4250),
.Y(n_4917)
);

INVx1_ASAP7_75t_L g4918 ( 
.A(n_4378),
.Y(n_4918)
);

NOR2xp33_ASAP7_75t_L g4919 ( 
.A(n_4059),
.B(n_317),
.Y(n_4919)
);

OAI21xp5_ASAP7_75t_L g4920 ( 
.A1(n_4581),
.A2(n_318),
.B(n_317),
.Y(n_4920)
);

AOI21xp5_ASAP7_75t_L g4921 ( 
.A1(n_4098),
.A2(n_4137),
.B(n_4102),
.Y(n_4921)
);

NAND2xp5_ASAP7_75t_L g4922 ( 
.A(n_4569),
.B(n_318),
.Y(n_4922)
);

OAI21xp5_ASAP7_75t_L g4923 ( 
.A1(n_4269),
.A2(n_319),
.B(n_318),
.Y(n_4923)
);

NAND2xp5_ASAP7_75t_L g4924 ( 
.A(n_4585),
.B(n_319),
.Y(n_4924)
);

AND2x2_ASAP7_75t_L g4925 ( 
.A(n_4123),
.B(n_319),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4383),
.Y(n_4926)
);

OAI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4455),
.A2(n_321),
.B1(n_322),
.B2(n_320),
.Y(n_4927)
);

OAI21xp5_ASAP7_75t_L g4928 ( 
.A1(n_4549),
.A2(n_322),
.B(n_321),
.Y(n_4928)
);

NAND2xp5_ASAP7_75t_L g4929 ( 
.A(n_4594),
.B(n_321),
.Y(n_4929)
);

AOI21xp5_ASAP7_75t_L g4930 ( 
.A1(n_4164),
.A2(n_323),
.B(n_322),
.Y(n_4930)
);

INVx1_ASAP7_75t_L g4931 ( 
.A(n_4402),
.Y(n_4931)
);

CKINVDCx6p67_ASAP7_75t_R g4932 ( 
.A(n_4130),
.Y(n_4932)
);

INVx3_ASAP7_75t_L g4933 ( 
.A(n_4096),
.Y(n_4933)
);

OAI21x1_ASAP7_75t_L g4934 ( 
.A1(n_4408),
.A2(n_4420),
.B(n_4419),
.Y(n_4934)
);

INVx2_ASAP7_75t_L g4935 ( 
.A(n_4258),
.Y(n_4935)
);

INVx2_ASAP7_75t_L g4936 ( 
.A(n_4266),
.Y(n_4936)
);

NAND2xp5_ASAP7_75t_L g4937 ( 
.A(n_4597),
.B(n_323),
.Y(n_4937)
);

CKINVDCx10_ASAP7_75t_R g4938 ( 
.A(n_4306),
.Y(n_4938)
);

O2A1O1Ixp5_ASAP7_75t_L g4939 ( 
.A1(n_4586),
.A2(n_324),
.B(n_325),
.C(n_323),
.Y(n_4939)
);

O2A1O1Ixp33_ASAP7_75t_L g4940 ( 
.A1(n_4179),
.A2(n_4580),
.B(n_4213),
.C(n_4582),
.Y(n_4940)
);

AOI22xp5_ASAP7_75t_L g4941 ( 
.A1(n_4255),
.A2(n_1072),
.B1(n_1075),
.B2(n_1069),
.Y(n_4941)
);

AOI21xp5_ASAP7_75t_L g4942 ( 
.A1(n_4169),
.A2(n_326),
.B(n_324),
.Y(n_4942)
);

AOI22xp5_ASAP7_75t_L g4943 ( 
.A1(n_4040),
.A2(n_1076),
.B1(n_1077),
.B2(n_1069),
.Y(n_4943)
);

NOR2x1_ASAP7_75t_L g4944 ( 
.A(n_4301),
.B(n_324),
.Y(n_4944)
);

NAND2xp5_ASAP7_75t_SL g4945 ( 
.A(n_4461),
.B(n_326),
.Y(n_4945)
);

AOI21xp5_ASAP7_75t_L g4946 ( 
.A1(n_4175),
.A2(n_328),
.B(n_327),
.Y(n_4946)
);

OAI21xp5_ASAP7_75t_L g4947 ( 
.A1(n_4553),
.A2(n_4468),
.B(n_4570),
.Y(n_4947)
);

NAND2xp33_ASAP7_75t_L g4948 ( 
.A(n_4265),
.B(n_327),
.Y(n_4948)
);

AOI21xp5_ASAP7_75t_L g4949 ( 
.A1(n_4182),
.A2(n_328),
.B(n_327),
.Y(n_4949)
);

OAI22xp5_ASAP7_75t_L g4950 ( 
.A1(n_4100),
.A2(n_330),
.B1(n_331),
.B2(n_329),
.Y(n_4950)
);

O2A1O1Ixp33_ASAP7_75t_SL g4951 ( 
.A1(n_4367),
.A2(n_330),
.B(n_331),
.C(n_329),
.Y(n_4951)
);

AOI21xp5_ASAP7_75t_L g4952 ( 
.A1(n_4197),
.A2(n_330),
.B(n_329),
.Y(n_4952)
);

NAND2xp5_ASAP7_75t_L g4953 ( 
.A(n_4113),
.B(n_331),
.Y(n_4953)
);

AOI22xp5_ASAP7_75t_L g4954 ( 
.A1(n_4084),
.A2(n_1060),
.B1(n_1061),
.B2(n_1059),
.Y(n_4954)
);

A2O1A1Ixp33_ASAP7_75t_L g4955 ( 
.A1(n_4600),
.A2(n_333),
.B(n_334),
.C(n_332),
.Y(n_4955)
);

AOI21xp5_ASAP7_75t_L g4956 ( 
.A1(n_4275),
.A2(n_333),
.B(n_332),
.Y(n_4956)
);

OAI21x1_ASAP7_75t_L g4957 ( 
.A1(n_4419),
.A2(n_335),
.B(n_334),
.Y(n_4957)
);

OAI22xp5_ASAP7_75t_SL g4958 ( 
.A1(n_4220),
.A2(n_335),
.B1(n_336),
.B2(n_334),
.Y(n_4958)
);

INVx1_ASAP7_75t_L g4959 ( 
.A(n_4421),
.Y(n_4959)
);

BUFx4f_ASAP7_75t_L g4960 ( 
.A(n_4201),
.Y(n_4960)
);

NAND2xp5_ASAP7_75t_L g4961 ( 
.A(n_4152),
.B(n_4141),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4437),
.B(n_335),
.Y(n_4962)
);

NAND2xp5_ASAP7_75t_L g4963 ( 
.A(n_4443),
.B(n_336),
.Y(n_4963)
);

OAI21x1_ASAP7_75t_L g4964 ( 
.A1(n_4420),
.A2(n_338),
.B(n_337),
.Y(n_4964)
);

AOI21xp5_ASAP7_75t_L g4965 ( 
.A1(n_4450),
.A2(n_338),
.B(n_337),
.Y(n_4965)
);

INVx4_ASAP7_75t_L g4966 ( 
.A(n_4154),
.Y(n_4966)
);

NOR2x1_ASAP7_75t_L g4967 ( 
.A(n_4249),
.B(n_337),
.Y(n_4967)
);

NAND2xp5_ASAP7_75t_L g4968 ( 
.A(n_4447),
.B(n_338),
.Y(n_4968)
);

NAND2xp5_ASAP7_75t_L g4969 ( 
.A(n_4452),
.B(n_339),
.Y(n_4969)
);

INVx1_ASAP7_75t_L g4970 ( 
.A(n_4274),
.Y(n_4970)
);

INVx1_ASAP7_75t_L g4971 ( 
.A(n_4282),
.Y(n_4971)
);

AOI21xp5_ASAP7_75t_L g4972 ( 
.A1(n_4454),
.A2(n_340),
.B(n_339),
.Y(n_4972)
);

NOR2xp33_ASAP7_75t_L g4973 ( 
.A(n_4416),
.B(n_340),
.Y(n_4973)
);

NAND2xp5_ASAP7_75t_L g4974 ( 
.A(n_4539),
.B(n_341),
.Y(n_4974)
);

INVx2_ASAP7_75t_L g4975 ( 
.A(n_4287),
.Y(n_4975)
);

A2O1A1Ixp33_ASAP7_75t_L g4976 ( 
.A1(n_4147),
.A2(n_342),
.B(n_343),
.C(n_341),
.Y(n_4976)
);

NAND2xp5_ASAP7_75t_L g4977 ( 
.A(n_4487),
.B(n_4490),
.Y(n_4977)
);

AOI21xp5_ASAP7_75t_L g4978 ( 
.A1(n_4427),
.A2(n_342),
.B(n_341),
.Y(n_4978)
);

NAND2xp5_ASAP7_75t_L g4979 ( 
.A(n_4506),
.B(n_342),
.Y(n_4979)
);

AOI21xp5_ASAP7_75t_L g4980 ( 
.A1(n_4427),
.A2(n_344),
.B(n_343),
.Y(n_4980)
);

NOR2xp33_ASAP7_75t_SL g4981 ( 
.A(n_4263),
.B(n_1055),
.Y(n_4981)
);

NAND2xp5_ASAP7_75t_L g4982 ( 
.A(n_4508),
.B(n_343),
.Y(n_4982)
);

BUFx4f_ASAP7_75t_L g4983 ( 
.A(n_4368),
.Y(n_4983)
);

A2O1A1Ixp33_ASAP7_75t_L g4984 ( 
.A1(n_4317),
.A2(n_345),
.B(n_346),
.C(n_344),
.Y(n_4984)
);

AOI22xp5_ASAP7_75t_L g4985 ( 
.A1(n_4126),
.A2(n_1058),
.B1(n_1059),
.B2(n_1057),
.Y(n_4985)
);

INVx2_ASAP7_75t_L g4986 ( 
.A(n_4292),
.Y(n_4986)
);

NAND2xp5_ASAP7_75t_L g4987 ( 
.A(n_4510),
.B(n_346),
.Y(n_4987)
);

OAI21xp5_ASAP7_75t_L g4988 ( 
.A1(n_4224),
.A2(n_347),
.B(n_346),
.Y(n_4988)
);

NAND2xp5_ASAP7_75t_SL g4989 ( 
.A(n_4088),
.B(n_347),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4534),
.B(n_347),
.Y(n_4990)
);

INVx3_ASAP7_75t_L g4991 ( 
.A(n_4096),
.Y(n_4991)
);

AND2x2_ASAP7_75t_L g4992 ( 
.A(n_4261),
.B(n_348),
.Y(n_4992)
);

AOI22xp5_ASAP7_75t_L g4993 ( 
.A1(n_4524),
.A2(n_1060),
.B1(n_1062),
.B2(n_1059),
.Y(n_4993)
);

AOI21xp5_ASAP7_75t_L g4994 ( 
.A1(n_4457),
.A2(n_349),
.B(n_348),
.Y(n_4994)
);

OAI22xp5_ASAP7_75t_L g4995 ( 
.A1(n_4426),
.A2(n_350),
.B1(n_351),
.B2(n_348),
.Y(n_4995)
);

A2O1A1Ixp33_ASAP7_75t_L g4996 ( 
.A1(n_4391),
.A2(n_351),
.B(n_352),
.C(n_350),
.Y(n_4996)
);

AOI21xp5_ASAP7_75t_L g4997 ( 
.A1(n_4457),
.A2(n_351),
.B(n_350),
.Y(n_4997)
);

NOR2xp33_ASAP7_75t_L g4998 ( 
.A(n_4158),
.B(n_352),
.Y(n_4998)
);

NOR2xp33_ASAP7_75t_L g4999 ( 
.A(n_4157),
.B(n_352),
.Y(n_4999)
);

AND2x2_ASAP7_75t_L g5000 ( 
.A(n_4081),
.B(n_353),
.Y(n_5000)
);

INVx1_ASAP7_75t_L g5001 ( 
.A(n_4296),
.Y(n_5001)
);

INVx1_ASAP7_75t_L g5002 ( 
.A(n_4299),
.Y(n_5002)
);

INVx2_ASAP7_75t_L g5003 ( 
.A(n_4315),
.Y(n_5003)
);

AOI21xp5_ASAP7_75t_L g5004 ( 
.A1(n_4331),
.A2(n_354),
.B(n_353),
.Y(n_5004)
);

NAND2xp5_ASAP7_75t_L g5005 ( 
.A(n_4537),
.B(n_354),
.Y(n_5005)
);

AOI21xp5_ASAP7_75t_L g5006 ( 
.A1(n_4338),
.A2(n_4297),
.B(n_4290),
.Y(n_5006)
);

NAND2xp5_ASAP7_75t_SL g5007 ( 
.A(n_4591),
.B(n_354),
.Y(n_5007)
);

NAND2xp5_ASAP7_75t_L g5008 ( 
.A(n_4551),
.B(n_355),
.Y(n_5008)
);

NAND2xp5_ASAP7_75t_L g5009 ( 
.A(n_4556),
.B(n_355),
.Y(n_5009)
);

AOI21xp5_ASAP7_75t_L g5010 ( 
.A1(n_4563),
.A2(n_357),
.B(n_356),
.Y(n_5010)
);

AOI21xp5_ASAP7_75t_L g5011 ( 
.A1(n_4577),
.A2(n_358),
.B(n_356),
.Y(n_5011)
);

AOI21xp5_ASAP7_75t_L g5012 ( 
.A1(n_4587),
.A2(n_359),
.B(n_356),
.Y(n_5012)
);

AOI22xp5_ASAP7_75t_L g5013 ( 
.A1(n_4085),
.A2(n_1055),
.B1(n_1056),
.B2(n_1054),
.Y(n_5013)
);

AOI21xp5_ASAP7_75t_L g5014 ( 
.A1(n_4384),
.A2(n_360),
.B(n_359),
.Y(n_5014)
);

NAND2xp33_ASAP7_75t_L g5015 ( 
.A(n_4233),
.B(n_360),
.Y(n_5015)
);

NAND2xp5_ASAP7_75t_SL g5016 ( 
.A(n_4591),
.B(n_361),
.Y(n_5016)
);

AOI21x1_ASAP7_75t_L g5017 ( 
.A1(n_4532),
.A2(n_362),
.B(n_361),
.Y(n_5017)
);

AND2x2_ASAP7_75t_L g5018 ( 
.A(n_4471),
.B(n_362),
.Y(n_5018)
);

AOI22xp33_ASAP7_75t_L g5019 ( 
.A1(n_4541),
.A2(n_364),
.B1(n_365),
.B2(n_363),
.Y(n_5019)
);

OAI22xp5_ASAP7_75t_L g5020 ( 
.A1(n_4507),
.A2(n_4558),
.B1(n_4321),
.B2(n_4593),
.Y(n_5020)
);

NAND2xp5_ASAP7_75t_L g5021 ( 
.A(n_4119),
.B(n_363),
.Y(n_5021)
);

AOI22xp33_ASAP7_75t_L g5022 ( 
.A1(n_4541),
.A2(n_364),
.B1(n_365),
.B2(n_363),
.Y(n_5022)
);

NAND2xp5_ASAP7_75t_SL g5023 ( 
.A(n_4293),
.B(n_364),
.Y(n_5023)
);

NOR2xp67_ASAP7_75t_L g5024 ( 
.A(n_4156),
.B(n_4192),
.Y(n_5024)
);

AOI22xp33_ASAP7_75t_L g5025 ( 
.A1(n_4546),
.A2(n_366),
.B1(n_367),
.B2(n_365),
.Y(n_5025)
);

NAND2xp5_ASAP7_75t_SL g5026 ( 
.A(n_4440),
.B(n_366),
.Y(n_5026)
);

AOI21xp5_ASAP7_75t_L g5027 ( 
.A1(n_4384),
.A2(n_368),
.B(n_367),
.Y(n_5027)
);

OAI22xp5_ASAP7_75t_L g5028 ( 
.A1(n_4558),
.A2(n_4546),
.B1(n_4347),
.B2(n_4601),
.Y(n_5028)
);

NAND3xp33_ASAP7_75t_SL g5029 ( 
.A(n_4206),
.B(n_6),
.C(n_7),
.Y(n_5029)
);

OAI21xp5_ASAP7_75t_L g5030 ( 
.A1(n_4535),
.A2(n_368),
.B(n_367),
.Y(n_5030)
);

AOI21xp5_ASAP7_75t_L g5031 ( 
.A1(n_4422),
.A2(n_369),
.B(n_368),
.Y(n_5031)
);

NOR2xp67_ASAP7_75t_L g5032 ( 
.A(n_4203),
.B(n_370),
.Y(n_5032)
);

INVx3_ASAP7_75t_L g5033 ( 
.A(n_4096),
.Y(n_5033)
);

NOR2xp33_ASAP7_75t_SL g5034 ( 
.A(n_4127),
.B(n_369),
.Y(n_5034)
);

OAI21xp33_ASAP7_75t_L g5035 ( 
.A1(n_4522),
.A2(n_370),
.B(n_369),
.Y(n_5035)
);

BUFx8_ASAP7_75t_SL g5036 ( 
.A(n_4304),
.Y(n_5036)
);

INVx2_ASAP7_75t_L g5037 ( 
.A(n_4320),
.Y(n_5037)
);

OAI21x1_ASAP7_75t_L g5038 ( 
.A1(n_4202),
.A2(n_371),
.B(n_370),
.Y(n_5038)
);

NAND2xp5_ASAP7_75t_SL g5039 ( 
.A(n_4440),
.B(n_371),
.Y(n_5039)
);

INVx2_ASAP7_75t_L g5040 ( 
.A(n_4324),
.Y(n_5040)
);

AOI21xp5_ASAP7_75t_L g5041 ( 
.A1(n_4422),
.A2(n_372),
.B(n_371),
.Y(n_5041)
);

NOR2xp67_ASAP7_75t_L g5042 ( 
.A(n_4247),
.B(n_373),
.Y(n_5042)
);

NOR2xp33_ASAP7_75t_L g5043 ( 
.A(n_4056),
.B(n_372),
.Y(n_5043)
);

INVx1_ASAP7_75t_L g5044 ( 
.A(n_4328),
.Y(n_5044)
);

AOI21xp5_ASAP7_75t_L g5045 ( 
.A1(n_4448),
.A2(n_375),
.B(n_374),
.Y(n_5045)
);

AOI21xp33_ASAP7_75t_L g5046 ( 
.A1(n_4344),
.A2(n_375),
.B(n_374),
.Y(n_5046)
);

NAND2xp5_ASAP7_75t_L g5047 ( 
.A(n_4216),
.B(n_374),
.Y(n_5047)
);

BUFx6f_ASAP7_75t_L g5048 ( 
.A(n_4430),
.Y(n_5048)
);

CKINVDCx10_ASAP7_75t_R g5049 ( 
.A(n_4154),
.Y(n_5049)
);

NAND2xp5_ASAP7_75t_L g5050 ( 
.A(n_4243),
.B(n_376),
.Y(n_5050)
);

O2A1O1Ixp33_ASAP7_75t_SL g5051 ( 
.A1(n_4190),
.A2(n_4590),
.B(n_4217),
.C(n_4489),
.Y(n_5051)
);

INVx1_ASAP7_75t_L g5052 ( 
.A(n_4354),
.Y(n_5052)
);

INVx2_ASAP7_75t_SL g5053 ( 
.A(n_4309),
.Y(n_5053)
);

INVx2_ASAP7_75t_L g5054 ( 
.A(n_4364),
.Y(n_5054)
);

CKINVDCx5p33_ASAP7_75t_R g5055 ( 
.A(n_4225),
.Y(n_5055)
);

AOI21xp5_ASAP7_75t_L g5056 ( 
.A1(n_4448),
.A2(n_4485),
.B(n_4373),
.Y(n_5056)
);

NAND2xp5_ASAP7_75t_SL g5057 ( 
.A(n_4464),
.B(n_376),
.Y(n_5057)
);

INVx5_ASAP7_75t_L g5058 ( 
.A(n_4430),
.Y(n_5058)
);

INVx2_ASAP7_75t_L g5059 ( 
.A(n_4370),
.Y(n_5059)
);

AOI21xp5_ASAP7_75t_L g5060 ( 
.A1(n_4446),
.A2(n_377),
.B(n_376),
.Y(n_5060)
);

AOI21xp5_ASAP7_75t_L g5061 ( 
.A1(n_4451),
.A2(n_379),
.B(n_378),
.Y(n_5061)
);

NOR3xp33_ASAP7_75t_L g5062 ( 
.A(n_4472),
.B(n_387),
.C(n_379),
.Y(n_5062)
);

A2O1A1Ixp33_ASAP7_75t_L g5063 ( 
.A1(n_4601),
.A2(n_379),
.B(n_380),
.C(n_378),
.Y(n_5063)
);

NAND2xp5_ASAP7_75t_L g5064 ( 
.A(n_4108),
.B(n_378),
.Y(n_5064)
);

AOI21xp5_ASAP7_75t_L g5065 ( 
.A1(n_4459),
.A2(n_381),
.B(n_380),
.Y(n_5065)
);

INVx2_ASAP7_75t_SL g5066 ( 
.A(n_4291),
.Y(n_5066)
);

BUFx8_ASAP7_75t_L g5067 ( 
.A(n_4305),
.Y(n_5067)
);

OAI22xp5_ASAP7_75t_L g5068 ( 
.A1(n_4295),
.A2(n_381),
.B1(n_382),
.B2(n_380),
.Y(n_5068)
);

AOI21xp5_ASAP7_75t_L g5069 ( 
.A1(n_4463),
.A2(n_383),
.B(n_382),
.Y(n_5069)
);

INVx4_ASAP7_75t_L g5070 ( 
.A(n_4368),
.Y(n_5070)
);

INVx1_ASAP7_75t_L g5071 ( 
.A(n_4380),
.Y(n_5071)
);

OAI21xp5_ASAP7_75t_L g5072 ( 
.A1(n_4526),
.A2(n_383),
.B(n_382),
.Y(n_5072)
);

OAI22xp5_ASAP7_75t_L g5073 ( 
.A1(n_4578),
.A2(n_4387),
.B1(n_4361),
.B2(n_4369),
.Y(n_5073)
);

NAND2xp5_ASAP7_75t_L g5074 ( 
.A(n_4114),
.B(n_4550),
.Y(n_5074)
);

AOI21x1_ASAP7_75t_L g5075 ( 
.A1(n_4322),
.A2(n_385),
.B(n_384),
.Y(n_5075)
);

A2O1A1Ixp33_ASAP7_75t_L g5076 ( 
.A1(n_4406),
.A2(n_4415),
.B(n_4479),
.C(n_4476),
.Y(n_5076)
);

OAI22xp5_ASAP7_75t_L g5077 ( 
.A1(n_4412),
.A2(n_4434),
.B1(n_4165),
.B2(n_4390),
.Y(n_5077)
);

NAND2xp5_ASAP7_75t_SL g5078 ( 
.A(n_4464),
.B(n_384),
.Y(n_5078)
);

O2A1O1Ixp33_ASAP7_75t_L g5079 ( 
.A1(n_4533),
.A2(n_4264),
.B(n_4554),
.C(n_4545),
.Y(n_5079)
);

OAI21xp5_ASAP7_75t_L g5080 ( 
.A1(n_4544),
.A2(n_387),
.B(n_386),
.Y(n_5080)
);

OAI21x1_ASAP7_75t_L g5081 ( 
.A1(n_4678),
.A2(n_4486),
.B(n_4483),
.Y(n_5081)
);

AO21x2_ASAP7_75t_L g5082 ( 
.A1(n_4653),
.A2(n_4411),
.B(n_4438),
.Y(n_5082)
);

CKINVDCx6p67_ASAP7_75t_R g5083 ( 
.A(n_5049),
.Y(n_5083)
);

AOI21xp33_ASAP7_75t_L g5084 ( 
.A1(n_4684),
.A2(n_4598),
.B(n_4596),
.Y(n_5084)
);

INVx8_ASAP7_75t_L g5085 ( 
.A(n_4903),
.Y(n_5085)
);

OAI21x1_ASAP7_75t_L g5086 ( 
.A1(n_4628),
.A2(n_4486),
.B(n_4483),
.Y(n_5086)
);

INVx1_ASAP7_75t_L g5087 ( 
.A(n_4681),
.Y(n_5087)
);

OR2x2_ASAP7_75t_L g5088 ( 
.A(n_4741),
.B(n_4200),
.Y(n_5088)
);

OAI21x1_ASAP7_75t_L g5089 ( 
.A1(n_4618),
.A2(n_4222),
.B(n_4202),
.Y(n_5089)
);

OAI22x1_ASAP7_75t_L g5090 ( 
.A1(n_4832),
.A2(n_4252),
.B1(n_4343),
.B2(n_4417),
.Y(n_5090)
);

INVx2_ASAP7_75t_L g5091 ( 
.A(n_4611),
.Y(n_5091)
);

INVx1_ASAP7_75t_L g5092 ( 
.A(n_4620),
.Y(n_5092)
);

OAI21x1_ASAP7_75t_L g5093 ( 
.A1(n_4610),
.A2(n_4222),
.B(n_4326),
.Y(n_5093)
);

OAI21x1_ASAP7_75t_L g5094 ( 
.A1(n_4614),
.A2(n_4607),
.B(n_4934),
.Y(n_5094)
);

NAND2xp5_ASAP7_75t_SL g5095 ( 
.A(n_4832),
.B(n_4561),
.Y(n_5095)
);

AOI21xp5_ASAP7_75t_L g5096 ( 
.A1(n_4869),
.A2(n_4491),
.B(n_4453),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_L g5097 ( 
.A(n_4625),
.B(n_4550),
.Y(n_5097)
);

NAND2xp5_ASAP7_75t_L g5098 ( 
.A(n_4851),
.B(n_4557),
.Y(n_5098)
);

OAI21xp5_ASAP7_75t_L g5099 ( 
.A1(n_4747),
.A2(n_4599),
.B(n_4564),
.Y(n_5099)
);

NAND2xp5_ASAP7_75t_L g5100 ( 
.A(n_5071),
.B(n_4557),
.Y(n_5100)
);

AO31x2_ASAP7_75t_L g5101 ( 
.A1(n_5020),
.A2(n_4513),
.A3(n_4436),
.B(n_4603),
.Y(n_5101)
);

AO21x1_ASAP7_75t_L g5102 ( 
.A1(n_4736),
.A2(n_4302),
.B(n_4564),
.Y(n_5102)
);

AOI21xp5_ASAP7_75t_L g5103 ( 
.A1(n_4948),
.A2(n_4561),
.B(n_4359),
.Y(n_5103)
);

NAND2xp5_ASAP7_75t_L g5104 ( 
.A(n_4633),
.B(n_4574),
.Y(n_5104)
);

A2O1A1Ixp33_ASAP7_75t_L g5105 ( 
.A1(n_5032),
.A2(n_4433),
.B(n_4375),
.C(n_4318),
.Y(n_5105)
);

AOI21x1_ASAP7_75t_L g5106 ( 
.A1(n_4902),
.A2(n_4409),
.B(n_4302),
.Y(n_5106)
);

OA22x2_ASAP7_75t_L g5107 ( 
.A1(n_4652),
.A2(n_4409),
.B1(n_4385),
.B2(n_4319),
.Y(n_5107)
);

AOI21xp5_ASAP7_75t_L g5108 ( 
.A1(n_5015),
.A2(n_4561),
.B(n_4358),
.Y(n_5108)
);

OAI21xp5_ASAP7_75t_L g5109 ( 
.A1(n_4955),
.A2(n_4588),
.B(n_4574),
.Y(n_5109)
);

AOI21xp5_ASAP7_75t_L g5110 ( 
.A1(n_4606),
.A2(n_4166),
.B(n_4092),
.Y(n_5110)
);

NAND2xp5_ASAP7_75t_L g5111 ( 
.A(n_4940),
.B(n_4588),
.Y(n_5111)
);

AO21x1_ASAP7_75t_L g5112 ( 
.A1(n_5028),
.A2(n_4583),
.B(n_4244),
.Y(n_5112)
);

AND2x4_ASAP7_75t_L g5113 ( 
.A(n_4866),
.B(n_4514),
.Y(n_5113)
);

AOI21xp5_ASAP7_75t_L g5114 ( 
.A1(n_4635),
.A2(n_4166),
.B(n_4092),
.Y(n_5114)
);

OAI22x1_ASAP7_75t_L g5115 ( 
.A1(n_4873),
.A2(n_4641),
.B1(n_4716),
.B2(n_4966),
.Y(n_5115)
);

AND2x2_ASAP7_75t_L g5116 ( 
.A(n_4608),
.B(n_4281),
.Y(n_5116)
);

BUFx6f_ASAP7_75t_L g5117 ( 
.A(n_4960),
.Y(n_5117)
);

INVx1_ASAP7_75t_L g5118 ( 
.A(n_4642),
.Y(n_5118)
);

INVx1_ASAP7_75t_L g5119 ( 
.A(n_4696),
.Y(n_5119)
);

INVx1_ASAP7_75t_L g5120 ( 
.A(n_4697),
.Y(n_5120)
);

AND2x2_ASAP7_75t_L g5121 ( 
.A(n_4605),
.B(n_4700),
.Y(n_5121)
);

AO21x2_ASAP7_75t_L g5122 ( 
.A1(n_4723),
.A2(n_4495),
.B(n_4494),
.Y(n_5122)
);

OAI21x1_ASAP7_75t_L g5123 ( 
.A1(n_4780),
.A2(n_4460),
.B(n_4403),
.Y(n_5123)
);

INVx4_ASAP7_75t_L g5124 ( 
.A(n_4960),
.Y(n_5124)
);

OAI21xp5_ASAP7_75t_L g5125 ( 
.A1(n_5042),
.A2(n_4560),
.B(n_4559),
.Y(n_5125)
);

OAI21xp5_ASAP7_75t_L g5126 ( 
.A1(n_4685),
.A2(n_4575),
.B(n_4566),
.Y(n_5126)
);

AO21x1_ASAP7_75t_L g5127 ( 
.A1(n_4758),
.A2(n_4244),
.B(n_4281),
.Y(n_5127)
);

AOI21x1_ASAP7_75t_L g5128 ( 
.A1(n_5017),
.A2(n_4143),
.B(n_4132),
.Y(n_5128)
);

OAI21x1_ASAP7_75t_L g5129 ( 
.A1(n_4892),
.A2(n_4505),
.B(n_4376),
.Y(n_5129)
);

OAI21x1_ASAP7_75t_L g5130 ( 
.A1(n_4624),
.A2(n_4445),
.B(n_4444),
.Y(n_5130)
);

O2A1O1Ixp5_ASAP7_75t_L g5131 ( 
.A1(n_4989),
.A2(n_4538),
.B(n_4592),
.C(n_4497),
.Y(n_5131)
);

OAI21x1_ASAP7_75t_L g5132 ( 
.A1(n_4619),
.A2(n_4515),
.B(n_4511),
.Y(n_5132)
);

NOR2xp33_ASAP7_75t_L g5133 ( 
.A(n_4710),
.B(n_4335),
.Y(n_5133)
);

AND2x2_ASAP7_75t_L g5134 ( 
.A(n_4855),
.B(n_4473),
.Y(n_5134)
);

OAI21x1_ASAP7_75t_L g5135 ( 
.A1(n_4779),
.A2(n_4517),
.B(n_4337),
.Y(n_5135)
);

AOI21xp5_ASAP7_75t_L g5136 ( 
.A1(n_5051),
.A2(n_4166),
.B(n_4092),
.Y(n_5136)
);

NAND2x1_ASAP7_75t_L g5137 ( 
.A(n_4966),
.B(n_4233),
.Y(n_5137)
);

INVx2_ASAP7_75t_L g5138 ( 
.A(n_4665),
.Y(n_5138)
);

OAI21x1_ASAP7_75t_L g5139 ( 
.A1(n_4804),
.A2(n_4481),
.B(n_4271),
.Y(n_5139)
);

AOI21x1_ASAP7_75t_L g5140 ( 
.A1(n_5075),
.A2(n_4143),
.B(n_4132),
.Y(n_5140)
);

AND2x4_ASAP7_75t_L g5141 ( 
.A(n_4933),
.B(n_4233),
.Y(n_5141)
);

OAI22x1_ASAP7_75t_L g5142 ( 
.A1(n_4682),
.A2(n_4656),
.B1(n_4792),
.B2(n_5055),
.Y(n_5142)
);

AOI21xp5_ASAP7_75t_L g5143 ( 
.A1(n_4609),
.A2(n_4209),
.B(n_4171),
.Y(n_5143)
);

A2O1A1Ixp33_ASAP7_75t_L g5144 ( 
.A1(n_4669),
.A2(n_4399),
.B(n_4520),
.C(n_4327),
.Y(n_5144)
);

OAI21x1_ASAP7_75t_L g5145 ( 
.A1(n_4699),
.A2(n_4353),
.B(n_4233),
.Y(n_5145)
);

NAND2xp5_ASAP7_75t_L g5146 ( 
.A(n_4612),
.B(n_4231),
.Y(n_5146)
);

INVx4_ASAP7_75t_L g5147 ( 
.A(n_4717),
.Y(n_5147)
);

NAND2xp5_ASAP7_75t_L g5148 ( 
.A(n_4977),
.B(n_4231),
.Y(n_5148)
);

OAI21x1_ASAP7_75t_L g5149 ( 
.A1(n_4638),
.A2(n_4096),
.B(n_4458),
.Y(n_5149)
);

OAI21x1_ASAP7_75t_L g5150 ( 
.A1(n_4663),
.A2(n_4458),
.B(n_4209),
.Y(n_5150)
);

OAI21x1_ASAP7_75t_L g5151 ( 
.A1(n_4933),
.A2(n_5033),
.B(n_4991),
.Y(n_5151)
);

AOI21xp5_ASAP7_75t_L g5152 ( 
.A1(n_4630),
.A2(n_4209),
.B(n_4171),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_L g5153 ( 
.A(n_4878),
.B(n_4492),
.Y(n_5153)
);

A2O1A1Ixp33_ASAP7_75t_L g5154 ( 
.A1(n_4691),
.A2(n_4548),
.B(n_4330),
.C(n_4474),
.Y(n_5154)
);

OAI21x1_ASAP7_75t_L g5155 ( 
.A1(n_4991),
.A2(n_4330),
.B(n_4171),
.Y(n_5155)
);

NAND2xp5_ASAP7_75t_SL g5156 ( 
.A(n_4983),
.B(n_4548),
.Y(n_5156)
);

NAND2xp5_ASAP7_75t_L g5157 ( 
.A(n_4918),
.B(n_4548),
.Y(n_5157)
);

OR2x6_ASAP7_75t_L g5158 ( 
.A(n_4677),
.B(n_4474),
.Y(n_5158)
);

NAND2xp5_ASAP7_75t_L g5159 ( 
.A(n_4926),
.B(n_4396),
.Y(n_5159)
);

OAI21x1_ASAP7_75t_L g5160 ( 
.A1(n_5033),
.A2(n_4474),
.B(n_4330),
.Y(n_5160)
);

NAND2xp5_ASAP7_75t_L g5161 ( 
.A(n_4931),
.B(n_4396),
.Y(n_5161)
);

OAI21xp5_ASAP7_75t_L g5162 ( 
.A1(n_4739),
.A2(n_4456),
.B(n_4396),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_4959),
.B(n_4396),
.Y(n_5163)
);

AND2x2_ASAP7_75t_L g5164 ( 
.A(n_4961),
.B(n_4475),
.Y(n_5164)
);

OAI21x1_ASAP7_75t_L g5165 ( 
.A1(n_4645),
.A2(n_4475),
.B(n_4456),
.Y(n_5165)
);

NAND2xp5_ASAP7_75t_L g5166 ( 
.A(n_4703),
.B(n_4753),
.Y(n_5166)
);

AO221x2_ASAP7_75t_L g5167 ( 
.A1(n_4958),
.A2(n_390),
.B1(n_391),
.B2(n_388),
.C(n_386),
.Y(n_5167)
);

AND2x2_ASAP7_75t_L g5168 ( 
.A(n_5018),
.B(n_4475),
.Y(n_5168)
);

NAND3xp33_ASAP7_75t_SL g5169 ( 
.A(n_4713),
.B(n_388),
.C(n_386),
.Y(n_5169)
);

INVx1_ASAP7_75t_L g5170 ( 
.A(n_4762),
.Y(n_5170)
);

NAND2xp5_ASAP7_75t_L g5171 ( 
.A(n_4771),
.B(n_4456),
.Y(n_5171)
);

INVx1_ASAP7_75t_L g5172 ( 
.A(n_4776),
.Y(n_5172)
);

INVxp67_ASAP7_75t_SL g5173 ( 
.A(n_5056),
.Y(n_5173)
);

OAI21x1_ASAP7_75t_L g5174 ( 
.A1(n_4647),
.A2(n_4456),
.B(n_390),
.Y(n_5174)
);

AO31x2_ASAP7_75t_L g5175 ( 
.A1(n_5077),
.A2(n_391),
.A3(n_392),
.B(n_388),
.Y(n_5175)
);

NAND2xp5_ASAP7_75t_L g5176 ( 
.A(n_4797),
.B(n_391),
.Y(n_5176)
);

AOI21xp5_ASAP7_75t_L g5177 ( 
.A1(n_4631),
.A2(n_393),
.B(n_392),
.Y(n_5177)
);

AO21x1_ASAP7_75t_L g5178 ( 
.A1(n_4649),
.A2(n_393),
.B(n_392),
.Y(n_5178)
);

OAI22xp5_ASAP7_75t_L g5179 ( 
.A1(n_4810),
.A2(n_394),
.B1(n_395),
.B2(n_393),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_L g5180 ( 
.A(n_4835),
.B(n_394),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_4845),
.B(n_394),
.Y(n_5181)
);

NAND2xp5_ASAP7_75t_L g5182 ( 
.A(n_4970),
.B(n_4971),
.Y(n_5182)
);

NOR2xp33_ASAP7_75t_L g5183 ( 
.A(n_4732),
.B(n_6),
.Y(n_5183)
);

AND2x2_ASAP7_75t_L g5184 ( 
.A(n_4817),
.B(n_7),
.Y(n_5184)
);

AOI21xp5_ASAP7_75t_SL g5185 ( 
.A1(n_4694),
.A2(n_396),
.B(n_395),
.Y(n_5185)
);

AND2x4_ASAP7_75t_L g5186 ( 
.A(n_4789),
.B(n_395),
.Y(n_5186)
);

AOI21xp5_ASAP7_75t_L g5187 ( 
.A1(n_4615),
.A2(n_5006),
.B(n_4643),
.Y(n_5187)
);

OAI21x1_ASAP7_75t_L g5188 ( 
.A1(n_4921),
.A2(n_397),
.B(n_396),
.Y(n_5188)
);

O2A1O1Ixp5_ASAP7_75t_L g5189 ( 
.A1(n_4683),
.A2(n_397),
.B(n_398),
.C(n_396),
.Y(n_5189)
);

INVx1_ASAP7_75t_L g5190 ( 
.A(n_4687),
.Y(n_5190)
);

NAND2xp5_ASAP7_75t_L g5191 ( 
.A(n_5001),
.B(n_397),
.Y(n_5191)
);

INVx5_ASAP7_75t_L g5192 ( 
.A(n_5036),
.Y(n_5192)
);

NAND2xp5_ASAP7_75t_L g5193 ( 
.A(n_5002),
.B(n_398),
.Y(n_5193)
);

OAI21x1_ASAP7_75t_L g5194 ( 
.A1(n_4689),
.A2(n_400),
.B(n_399),
.Y(n_5194)
);

OAI22xp5_ASAP7_75t_L g5195 ( 
.A1(n_4738),
.A2(n_400),
.B1(n_401),
.B2(n_399),
.Y(n_5195)
);

O2A1O1Ixp5_ASAP7_75t_L g5196 ( 
.A1(n_4729),
.A2(n_4730),
.B(n_4983),
.C(n_4867),
.Y(n_5196)
);

OAI21x1_ASAP7_75t_L g5197 ( 
.A1(n_4756),
.A2(n_401),
.B(n_400),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_4718),
.Y(n_5198)
);

BUFx2_ASAP7_75t_L g5199 ( 
.A(n_4857),
.Y(n_5199)
);

A2O1A1Ixp33_ASAP7_75t_L g5200 ( 
.A1(n_4798),
.A2(n_402),
.B(n_403),
.C(n_401),
.Y(n_5200)
);

OAI21x1_ASAP7_75t_L g5201 ( 
.A1(n_4858),
.A2(n_403),
.B(n_402),
.Y(n_5201)
);

OAI21x1_ASAP7_75t_L g5202 ( 
.A1(n_4863),
.A2(n_404),
.B(n_403),
.Y(n_5202)
);

INVx2_ASAP7_75t_L g5203 ( 
.A(n_4751),
.Y(n_5203)
);

INVx8_ASAP7_75t_L g5204 ( 
.A(n_4717),
.Y(n_5204)
);

INVx3_ASAP7_75t_L g5205 ( 
.A(n_4882),
.Y(n_5205)
);

OAI21x1_ASAP7_75t_L g5206 ( 
.A1(n_4870),
.A2(n_405),
.B(n_404),
.Y(n_5206)
);

A2O1A1Ixp33_ASAP7_75t_L g5207 ( 
.A1(n_4658),
.A2(n_406),
.B(n_407),
.C(n_405),
.Y(n_5207)
);

BUFx2_ASAP7_75t_R g5208 ( 
.A(n_4775),
.Y(n_5208)
);

CKINVDCx5p33_ASAP7_75t_R g5209 ( 
.A(n_4721),
.Y(n_5209)
);

OAI21xp5_ASAP7_75t_L g5210 ( 
.A1(n_4659),
.A2(n_406),
.B(n_405),
.Y(n_5210)
);

AO31x2_ASAP7_75t_L g5211 ( 
.A1(n_4705),
.A2(n_407),
.A3(n_408),
.B(n_406),
.Y(n_5211)
);

AOI21xp5_ASAP7_75t_L g5212 ( 
.A1(n_4627),
.A2(n_408),
.B(n_407),
.Y(n_5212)
);

INVx2_ASAP7_75t_SL g5213 ( 
.A(n_4882),
.Y(n_5213)
);

BUFx6f_ASAP7_75t_L g5214 ( 
.A(n_5048),
.Y(n_5214)
);

OAI21x1_ASAP7_75t_SL g5215 ( 
.A1(n_5070),
.A2(n_409),
.B(n_408),
.Y(n_5215)
);

OAI21x1_ASAP7_75t_L g5216 ( 
.A1(n_4769),
.A2(n_410),
.B(n_409),
.Y(n_5216)
);

INVx3_ASAP7_75t_L g5217 ( 
.A(n_5067),
.Y(n_5217)
);

AOI21xp5_ASAP7_75t_L g5218 ( 
.A1(n_4623),
.A2(n_410),
.B(n_409),
.Y(n_5218)
);

NOR2x1_ASAP7_75t_SL g5219 ( 
.A(n_4632),
.B(n_410),
.Y(n_5219)
);

AOI21xp5_ASAP7_75t_L g5220 ( 
.A1(n_4734),
.A2(n_412),
.B(n_411),
.Y(n_5220)
);

AOI21x1_ASAP7_75t_SL g5221 ( 
.A1(n_5050),
.A2(n_413),
.B(n_412),
.Y(n_5221)
);

INVx1_ASAP7_75t_L g5222 ( 
.A(n_4742),
.Y(n_5222)
);

OAI21x1_ASAP7_75t_L g5223 ( 
.A1(n_4670),
.A2(n_414),
.B(n_413),
.Y(n_5223)
);

NAND2xp5_ASAP7_75t_SL g5224 ( 
.A(n_5024),
.B(n_414),
.Y(n_5224)
);

HAxp5_ASAP7_75t_L g5225 ( 
.A(n_4757),
.B(n_7),
.CON(n_5225),
.SN(n_5225)
);

NAND2xp5_ASAP7_75t_SL g5226 ( 
.A(n_5070),
.B(n_414),
.Y(n_5226)
);

AOI21xp33_ASAP7_75t_L g5227 ( 
.A1(n_5079),
.A2(n_416),
.B(n_415),
.Y(n_5227)
);

HB1xp67_ASAP7_75t_L g5228 ( 
.A(n_4782),
.Y(n_5228)
);

NAND2xp5_ASAP7_75t_L g5229 ( 
.A(n_5044),
.B(n_415),
.Y(n_5229)
);

INVx2_ASAP7_75t_SL g5230 ( 
.A(n_5067),
.Y(n_5230)
);

OAI21x1_ASAP7_75t_L g5231 ( 
.A1(n_4836),
.A2(n_417),
.B(n_416),
.Y(n_5231)
);

BUFx2_ASAP7_75t_L g5232 ( 
.A(n_4789),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_4755),
.Y(n_5233)
);

NOR3xp33_ASAP7_75t_L g5234 ( 
.A(n_4772),
.B(n_4698),
.C(n_5029),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_4842),
.Y(n_5235)
);

OAI21x1_ASAP7_75t_L g5236 ( 
.A1(n_4896),
.A2(n_418),
.B(n_417),
.Y(n_5236)
);

A2O1A1Ixp33_ASAP7_75t_L g5237 ( 
.A1(n_4637),
.A2(n_420),
.B(n_421),
.C(n_419),
.Y(n_5237)
);

NAND2xp5_ASAP7_75t_L g5238 ( 
.A(n_5052),
.B(n_419),
.Y(n_5238)
);

BUFx4f_ASAP7_75t_SL g5239 ( 
.A(n_4932),
.Y(n_5239)
);

OAI21xp5_ASAP7_75t_L g5240 ( 
.A1(n_5063),
.A2(n_421),
.B(n_420),
.Y(n_5240)
);

BUFx4f_ASAP7_75t_L g5241 ( 
.A(n_4768),
.Y(n_5241)
);

AOI21x1_ASAP7_75t_L g5242 ( 
.A1(n_4875),
.A2(n_5016),
.B(n_5007),
.Y(n_5242)
);

BUFx6f_ASAP7_75t_L g5243 ( 
.A(n_5048),
.Y(n_5243)
);

NAND3xp33_ASAP7_75t_L g5244 ( 
.A(n_5034),
.B(n_5062),
.C(n_4909),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_4847),
.B(n_420),
.Y(n_5245)
);

AOI21xp5_ASAP7_75t_L g5246 ( 
.A1(n_4626),
.A2(n_423),
.B(n_422),
.Y(n_5246)
);

AOI211x1_ASAP7_75t_L g5247 ( 
.A1(n_4928),
.A2(n_423),
.B(n_424),
.C(n_422),
.Y(n_5247)
);

NAND2xp5_ASAP7_75t_L g5248 ( 
.A(n_4888),
.B(n_422),
.Y(n_5248)
);

OAI21x1_ASAP7_75t_L g5249 ( 
.A1(n_4957),
.A2(n_424),
.B(n_423),
.Y(n_5249)
);

NAND2xp5_ASAP7_75t_L g5250 ( 
.A(n_4891),
.B(n_425),
.Y(n_5250)
);

AOI21xp5_ASAP7_75t_L g5251 ( 
.A1(n_4766),
.A2(n_427),
.B(n_425),
.Y(n_5251)
);

OAI21x1_ASAP7_75t_L g5252 ( 
.A1(n_4964),
.A2(n_427),
.B(n_425),
.Y(n_5252)
);

AOI21xp5_ASAP7_75t_L g5253 ( 
.A1(n_4750),
.A2(n_428),
.B(n_427),
.Y(n_5253)
);

INVx2_ASAP7_75t_L g5254 ( 
.A(n_4904),
.Y(n_5254)
);

OAI22xp5_ASAP7_75t_L g5255 ( 
.A1(n_4616),
.A2(n_429),
.B1(n_430),
.B2(n_428),
.Y(n_5255)
);

CKINVDCx8_ASAP7_75t_R g5256 ( 
.A(n_4938),
.Y(n_5256)
);

OAI21x1_ASAP7_75t_L g5257 ( 
.A1(n_5038),
.A2(n_429),
.B(n_428),
.Y(n_5257)
);

OAI21x1_ASAP7_75t_L g5258 ( 
.A1(n_4679),
.A2(n_430),
.B(n_429),
.Y(n_5258)
);

NAND2xp5_ASAP7_75t_SL g5259 ( 
.A(n_4824),
.B(n_431),
.Y(n_5259)
);

BUFx12f_ASAP7_75t_L g5260 ( 
.A(n_4717),
.Y(n_5260)
);

OAI22xp5_ASAP7_75t_L g5261 ( 
.A1(n_4862),
.A2(n_432),
.B1(n_433),
.B2(n_431),
.Y(n_5261)
);

NOR2xp33_ASAP7_75t_L g5262 ( 
.A(n_5066),
.B(n_8),
.Y(n_5262)
);

O2A1O1Ixp5_ASAP7_75t_L g5263 ( 
.A1(n_4853),
.A2(n_432),
.B(n_433),
.C(n_431),
.Y(n_5263)
);

NAND2xp5_ASAP7_75t_L g5264 ( 
.A(n_4906),
.B(n_432),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_4917),
.Y(n_5265)
);

OAI21x1_ASAP7_75t_L g5266 ( 
.A1(n_4745),
.A2(n_434),
.B(n_433),
.Y(n_5266)
);

AO31x2_ASAP7_75t_L g5267 ( 
.A1(n_5073),
.A2(n_435),
.A3(n_436),
.B(n_434),
.Y(n_5267)
);

OAI21x1_ASAP7_75t_L g5268 ( 
.A1(n_4668),
.A2(n_436),
.B(n_435),
.Y(n_5268)
);

AOI21xp5_ASAP7_75t_L g5269 ( 
.A1(n_4809),
.A2(n_437),
.B(n_436),
.Y(n_5269)
);

NAND2xp5_ASAP7_75t_SL g5270 ( 
.A(n_4824),
.B(n_437),
.Y(n_5270)
);

AOI221x1_ASAP7_75t_L g5271 ( 
.A1(n_4774),
.A2(n_439),
.B1(n_440),
.B2(n_438),
.C(n_437),
.Y(n_5271)
);

AOI21xp5_ASAP7_75t_L g5272 ( 
.A1(n_4819),
.A2(n_439),
.B(n_438),
.Y(n_5272)
);

OAI21xp33_ASAP7_75t_L g5273 ( 
.A1(n_4796),
.A2(n_441),
.B(n_440),
.Y(n_5273)
);

OAI21xp5_ASAP7_75t_L g5274 ( 
.A1(n_4825),
.A2(n_441),
.B(n_440),
.Y(n_5274)
);

AOI221xp5_ASAP7_75t_L g5275 ( 
.A1(n_4660),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.C(n_11),
.Y(n_5275)
);

AOI21xp5_ASAP7_75t_SL g5276 ( 
.A1(n_4818),
.A2(n_442),
.B(n_441),
.Y(n_5276)
);

AOI21x1_ASAP7_75t_L g5277 ( 
.A1(n_4849),
.A2(n_443),
.B(n_442),
.Y(n_5277)
);

OAI21x1_ASAP7_75t_L g5278 ( 
.A1(n_4672),
.A2(n_444),
.B(n_442),
.Y(n_5278)
);

AOI22xp33_ASAP7_75t_L g5279 ( 
.A1(n_4947),
.A2(n_445),
.B1(n_446),
.B2(n_444),
.Y(n_5279)
);

A2O1A1Ixp33_ASAP7_75t_L g5280 ( 
.A1(n_4846),
.A2(n_445),
.B(n_446),
.C(n_444),
.Y(n_5280)
);

AOI22xp5_ASAP7_75t_SL g5281 ( 
.A1(n_4806),
.A2(n_448),
.B1(n_449),
.B2(n_447),
.Y(n_5281)
);

OAI21x1_ASAP7_75t_L g5282 ( 
.A1(n_4695),
.A2(n_449),
.B(n_448),
.Y(n_5282)
);

A2O1A1Ixp33_ASAP7_75t_L g5283 ( 
.A1(n_4874),
.A2(n_450),
.B(n_451),
.C(n_449),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_4935),
.Y(n_5284)
);

OAI21x1_ASAP7_75t_SL g5285 ( 
.A1(n_4761),
.A2(n_451),
.B(n_450),
.Y(n_5285)
);

AOI22xp33_ASAP7_75t_L g5286 ( 
.A1(n_4654),
.A2(n_452),
.B1(n_453),
.B2(n_450),
.Y(n_5286)
);

AND2x2_ASAP7_75t_L g5287 ( 
.A(n_4992),
.B(n_8),
.Y(n_5287)
);

OAI21x1_ASAP7_75t_L g5288 ( 
.A1(n_4695),
.A2(n_453),
.B(n_452),
.Y(n_5288)
);

NAND2xp5_ASAP7_75t_L g5289 ( 
.A(n_4936),
.B(n_452),
.Y(n_5289)
);

NOR2x1_ASAP7_75t_R g5290 ( 
.A(n_4912),
.B(n_453),
.Y(n_5290)
);

OAI21xp33_ASAP7_75t_L g5291 ( 
.A1(n_4893),
.A2(n_455),
.B(n_454),
.Y(n_5291)
);

OAI21x1_ASAP7_75t_L g5292 ( 
.A1(n_4720),
.A2(n_456),
.B(n_455),
.Y(n_5292)
);

OAI21xp5_ASAP7_75t_L g5293 ( 
.A1(n_4939),
.A2(n_458),
.B(n_457),
.Y(n_5293)
);

INVx2_ASAP7_75t_L g5294 ( 
.A(n_4975),
.Y(n_5294)
);

OAI21xp5_ASAP7_75t_L g5295 ( 
.A1(n_4675),
.A2(n_4976),
.B(n_4852),
.Y(n_5295)
);

NAND2xp5_ASAP7_75t_L g5296 ( 
.A(n_4986),
.B(n_457),
.Y(n_5296)
);

NAND2xp5_ASAP7_75t_L g5297 ( 
.A(n_5003),
.B(n_457),
.Y(n_5297)
);

NOR2xp67_ASAP7_75t_L g5298 ( 
.A(n_4604),
.B(n_462),
.Y(n_5298)
);

OAI21xp5_ASAP7_75t_L g5299 ( 
.A1(n_4704),
.A2(n_459),
.B(n_458),
.Y(n_5299)
);

INVx1_ASAP7_75t_L g5300 ( 
.A(n_5037),
.Y(n_5300)
);

NAND2xp5_ASAP7_75t_L g5301 ( 
.A(n_5040),
.B(n_5054),
.Y(n_5301)
);

AO31x2_ASAP7_75t_L g5302 ( 
.A1(n_4984),
.A2(n_460),
.A3(n_461),
.B(n_458),
.Y(n_5302)
);

OAI21x1_ASAP7_75t_L g5303 ( 
.A1(n_4720),
.A2(n_461),
.B(n_460),
.Y(n_5303)
);

NAND2xp5_ASAP7_75t_L g5304 ( 
.A(n_5059),
.B(n_460),
.Y(n_5304)
);

AND2x2_ASAP7_75t_L g5305 ( 
.A(n_4702),
.B(n_9),
.Y(n_5305)
);

AOI21xp5_ASAP7_75t_L g5306 ( 
.A1(n_4838),
.A2(n_462),
.B(n_461),
.Y(n_5306)
);

OAI21x1_ASAP7_75t_L g5307 ( 
.A1(n_4791),
.A2(n_463),
.B(n_462),
.Y(n_5307)
);

OAI21x1_ASAP7_75t_L g5308 ( 
.A1(n_4791),
.A2(n_465),
.B(n_464),
.Y(n_5308)
);

INVx2_ASAP7_75t_SL g5309 ( 
.A(n_4711),
.Y(n_5309)
);

OAI21x1_ASAP7_75t_SL g5310 ( 
.A1(n_4920),
.A2(n_465),
.B(n_464),
.Y(n_5310)
);

OAI21x1_ASAP7_75t_L g5311 ( 
.A1(n_4794),
.A2(n_465),
.B(n_464),
.Y(n_5311)
);

OAI21x1_ASAP7_75t_L g5312 ( 
.A1(n_4639),
.A2(n_467),
.B(n_466),
.Y(n_5312)
);

NAND2xp5_ASAP7_75t_L g5313 ( 
.A(n_5000),
.B(n_466),
.Y(n_5313)
);

INVx2_ASAP7_75t_L g5314 ( 
.A(n_4629),
.Y(n_5314)
);

AOI21xp5_ASAP7_75t_L g5315 ( 
.A1(n_4778),
.A2(n_467),
.B(n_466),
.Y(n_5315)
);

AND2x2_ASAP7_75t_L g5316 ( 
.A(n_4790),
.B(n_9),
.Y(n_5316)
);

INVx2_ASAP7_75t_L g5317 ( 
.A(n_4629),
.Y(n_5317)
);

OAI21x1_ASAP7_75t_L g5318 ( 
.A1(n_4640),
.A2(n_4644),
.B(n_4820),
.Y(n_5318)
);

OAI21x1_ASAP7_75t_L g5319 ( 
.A1(n_4763),
.A2(n_468),
.B(n_467),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_5074),
.B(n_10),
.Y(n_5320)
);

BUFx6f_ASAP7_75t_L g5321 ( 
.A(n_5048),
.Y(n_5321)
);

AOI21xp5_ASAP7_75t_L g5322 ( 
.A1(n_4622),
.A2(n_469),
.B(n_468),
.Y(n_5322)
);

OAI21xp5_ASAP7_75t_L g5323 ( 
.A1(n_4712),
.A2(n_469),
.B(n_468),
.Y(n_5323)
);

NAND2xp5_ASAP7_75t_L g5324 ( 
.A(n_4829),
.B(n_469),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_4830),
.B(n_470),
.Y(n_5325)
);

BUFx6f_ASAP7_75t_L g5326 ( 
.A(n_4629),
.Y(n_5326)
);

OAI21x1_ASAP7_75t_L g5327 ( 
.A1(n_4737),
.A2(n_471),
.B(n_470),
.Y(n_5327)
);

NAND3xp33_ASAP7_75t_SL g5328 ( 
.A(n_4843),
.B(n_471),
.C(n_470),
.Y(n_5328)
);

NAND2xp5_ASAP7_75t_SL g5329 ( 
.A(n_4824),
.B(n_471),
.Y(n_5329)
);

OAI21x1_ASAP7_75t_L g5330 ( 
.A1(n_4731),
.A2(n_473),
.B(n_472),
.Y(n_5330)
);

AND2x2_ASAP7_75t_L g5331 ( 
.A(n_4693),
.B(n_10),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_4841),
.B(n_472),
.Y(n_5332)
);

INVx3_ASAP7_75t_L g5333 ( 
.A(n_4634),
.Y(n_5333)
);

NAND2xp5_ASAP7_75t_L g5334 ( 
.A(n_4925),
.B(n_472),
.Y(n_5334)
);

AOI21x1_ASAP7_75t_SL g5335 ( 
.A1(n_4788),
.A2(n_474),
.B(n_473),
.Y(n_5335)
);

NAND2xp5_ASAP7_75t_L g5336 ( 
.A(n_4795),
.B(n_474),
.Y(n_5336)
);

OAI21x1_ASAP7_75t_L g5337 ( 
.A1(n_4764),
.A2(n_475),
.B(n_474),
.Y(n_5337)
);

A2O1A1Ixp33_ASAP7_75t_L g5338 ( 
.A1(n_4759),
.A2(n_476),
.B(n_477),
.C(n_475),
.Y(n_5338)
);

AOI21xp5_ASAP7_75t_L g5339 ( 
.A1(n_4613),
.A2(n_476),
.B(n_475),
.Y(n_5339)
);

OAI21xp5_ASAP7_75t_L g5340 ( 
.A1(n_4913),
.A2(n_478),
.B(n_477),
.Y(n_5340)
);

AOI22xp5_ASAP7_75t_L g5341 ( 
.A1(n_4973),
.A2(n_4981),
.B1(n_4900),
.B2(n_4889),
.Y(n_5341)
);

NAND2xp5_ASAP7_75t_L g5342 ( 
.A(n_4617),
.B(n_477),
.Y(n_5342)
);

BUFx6f_ASAP7_75t_L g5343 ( 
.A(n_4634),
.Y(n_5343)
);

AND2x2_ASAP7_75t_L g5344 ( 
.A(n_4788),
.B(n_11),
.Y(n_5344)
);

AOI21xp5_ASAP7_75t_L g5345 ( 
.A1(n_4632),
.A2(n_479),
.B(n_478),
.Y(n_5345)
);

NAND3xp33_ASAP7_75t_L g5346 ( 
.A(n_4967),
.B(n_479),
.C(n_478),
.Y(n_5346)
);

OAI21xp5_ASAP7_75t_L g5347 ( 
.A1(n_4813),
.A2(n_480),
.B(n_479),
.Y(n_5347)
);

OAI21x1_ASAP7_75t_L g5348 ( 
.A1(n_4646),
.A2(n_481),
.B(n_480),
.Y(n_5348)
);

INVx1_ASAP7_75t_L g5349 ( 
.A(n_4657),
.Y(n_5349)
);

OAI21x1_ASAP7_75t_L g5350 ( 
.A1(n_4879),
.A2(n_482),
.B(n_481),
.Y(n_5350)
);

OAI21x1_ASAP7_75t_L g5351 ( 
.A1(n_4686),
.A2(n_482),
.B(n_481),
.Y(n_5351)
);

OAI21x1_ASAP7_75t_L g5352 ( 
.A1(n_4690),
.A2(n_483),
.B(n_482),
.Y(n_5352)
);

AOI21xp5_ASAP7_75t_L g5353 ( 
.A1(n_4815),
.A2(n_484),
.B(n_483),
.Y(n_5353)
);

AOI21x1_ASAP7_75t_L g5354 ( 
.A1(n_4854),
.A2(n_485),
.B(n_484),
.Y(n_5354)
);

INVx2_ASAP7_75t_SL g5355 ( 
.A(n_4812),
.Y(n_5355)
);

NAND3xp33_ASAP7_75t_L g5356 ( 
.A(n_4944),
.B(n_485),
.C(n_484),
.Y(n_5356)
);

AOI21x1_ASAP7_75t_L g5357 ( 
.A1(n_4880),
.A2(n_487),
.B(n_486),
.Y(n_5357)
);

AOI21xp5_ASAP7_75t_L g5358 ( 
.A1(n_4802),
.A2(n_487),
.B(n_486),
.Y(n_5358)
);

NOR2x1_ASAP7_75t_R g5359 ( 
.A(n_4811),
.B(n_486),
.Y(n_5359)
);

NAND2xp5_ASAP7_75t_L g5360 ( 
.A(n_4621),
.B(n_487),
.Y(n_5360)
);

AOI21xp5_ASAP7_75t_L g5361 ( 
.A1(n_4688),
.A2(n_489),
.B(n_488),
.Y(n_5361)
);

A2O1A1Ixp33_ASAP7_75t_L g5362 ( 
.A1(n_4708),
.A2(n_489),
.B(n_490),
.C(n_488),
.Y(n_5362)
);

AOI21xp5_ASAP7_75t_L g5363 ( 
.A1(n_4743),
.A2(n_490),
.B(n_488),
.Y(n_5363)
);

INVx1_ASAP7_75t_L g5364 ( 
.A(n_4890),
.Y(n_5364)
);

INVx1_ASAP7_75t_L g5365 ( 
.A(n_4648),
.Y(n_5365)
);

AOI21xp33_ASAP7_75t_L g5366 ( 
.A1(n_4915),
.A2(n_491),
.B(n_490),
.Y(n_5366)
);

INVxp67_ASAP7_75t_SL g5367 ( 
.A(n_4749),
.Y(n_5367)
);

AOI21xp5_ASAP7_75t_L g5368 ( 
.A1(n_4777),
.A2(n_492),
.B(n_491),
.Y(n_5368)
);

BUFx3_ASAP7_75t_L g5369 ( 
.A(n_5053),
.Y(n_5369)
);

INVx2_ASAP7_75t_SL g5370 ( 
.A(n_5058),
.Y(n_5370)
);

OAI21x1_ASAP7_75t_L g5371 ( 
.A1(n_4770),
.A2(n_493),
.B(n_491),
.Y(n_5371)
);

INVx1_ASAP7_75t_SL g5372 ( 
.A(n_4634),
.Y(n_5372)
);

AOI22xp5_ASAP7_75t_L g5373 ( 
.A1(n_4674),
.A2(n_494),
.B1(n_495),
.B2(n_493),
.Y(n_5373)
);

AND2x2_ASAP7_75t_L g5374 ( 
.A(n_4856),
.B(n_11),
.Y(n_5374)
);

AND3x4_ASAP7_75t_L g5375 ( 
.A(n_4839),
.B(n_494),
.C(n_493),
.Y(n_5375)
);

AOI211x1_ASAP7_75t_L g5376 ( 
.A1(n_5021),
.A2(n_4988),
.B(n_4746),
.C(n_4953),
.Y(n_5376)
);

CKINVDCx5p33_ASAP7_75t_R g5377 ( 
.A(n_4828),
.Y(n_5377)
);

NAND2xp5_ASAP7_75t_SL g5378 ( 
.A(n_4673),
.B(n_494),
.Y(n_5378)
);

OAI21x1_ASAP7_75t_L g5379 ( 
.A1(n_4725),
.A2(n_497),
.B(n_496),
.Y(n_5379)
);

AOI21xp5_ASAP7_75t_L g5380 ( 
.A1(n_4887),
.A2(n_497),
.B(n_496),
.Y(n_5380)
);

OAI21x1_ASAP7_75t_L g5381 ( 
.A1(n_4886),
.A2(n_497),
.B(n_496),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_L g5382 ( 
.A(n_5047),
.B(n_498),
.Y(n_5382)
);

OAI21xp5_ASAP7_75t_L g5383 ( 
.A1(n_4833),
.A2(n_4996),
.B(n_4826),
.Y(n_5383)
);

AOI21xp5_ASAP7_75t_L g5384 ( 
.A1(n_4636),
.A2(n_499),
.B(n_498),
.Y(n_5384)
);

INVx3_ASAP7_75t_L g5385 ( 
.A(n_4673),
.Y(n_5385)
);

OAI21xp5_ASAP7_75t_L g5386 ( 
.A1(n_4662),
.A2(n_499),
.B(n_498),
.Y(n_5386)
);

AOI21xp5_ASAP7_75t_L g5387 ( 
.A1(n_5026),
.A2(n_501),
.B(n_500),
.Y(n_5387)
);

INVx3_ASAP7_75t_L g5388 ( 
.A(n_4673),
.Y(n_5388)
);

NAND2x1p5_ASAP7_75t_L g5389 ( 
.A(n_5058),
.B(n_500),
.Y(n_5389)
);

AOI21xp5_ASAP7_75t_L g5390 ( 
.A1(n_5039),
.A2(n_501),
.B(n_500),
.Y(n_5390)
);

AOI21x1_ASAP7_75t_SL g5391 ( 
.A1(n_4856),
.A2(n_502),
.B(n_501),
.Y(n_5391)
);

BUFx3_ASAP7_75t_L g5392 ( 
.A(n_5058),
.Y(n_5392)
);

OAI21x1_ASAP7_75t_L g5393 ( 
.A1(n_4814),
.A2(n_503),
.B(n_502),
.Y(n_5393)
);

AO21x1_ASAP7_75t_L g5394 ( 
.A1(n_4999),
.A2(n_504),
.B(n_502),
.Y(n_5394)
);

INVx1_ASAP7_75t_L g5395 ( 
.A(n_4650),
.Y(n_5395)
);

AND2x6_ASAP7_75t_L g5396 ( 
.A(n_4793),
.B(n_504),
.Y(n_5396)
);

OAI21xp5_ASAP7_75t_SL g5397 ( 
.A1(n_4881),
.A2(n_505),
.B(n_504),
.Y(n_5397)
);

OAI21x1_ASAP7_75t_L g5398 ( 
.A1(n_4655),
.A2(n_5078),
.B(n_5057),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_4651),
.Y(n_5399)
);

AOI21xp5_ASAP7_75t_L g5400 ( 
.A1(n_5076),
.A2(n_506),
.B(n_505),
.Y(n_5400)
);

INVx2_ASAP7_75t_SL g5401 ( 
.A(n_5204),
.Y(n_5401)
);

BUFx3_ASAP7_75t_L g5402 ( 
.A(n_5260),
.Y(n_5402)
);

INVx2_ASAP7_75t_L g5403 ( 
.A(n_5228),
.Y(n_5403)
);

NAND2xp5_ASAP7_75t_L g5404 ( 
.A(n_5190),
.B(n_5198),
.Y(n_5404)
);

INVx3_ASAP7_75t_SL g5405 ( 
.A(n_5085),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5092),
.Y(n_5406)
);

BUFx3_ASAP7_75t_L g5407 ( 
.A(n_5085),
.Y(n_5407)
);

CKINVDCx20_ASAP7_75t_R g5408 ( 
.A(n_5239),
.Y(n_5408)
);

BUFx3_ASAP7_75t_L g5409 ( 
.A(n_5241),
.Y(n_5409)
);

BUFx3_ASAP7_75t_L g5410 ( 
.A(n_5204),
.Y(n_5410)
);

INVx3_ASAP7_75t_SL g5411 ( 
.A(n_5209),
.Y(n_5411)
);

OR2x2_ASAP7_75t_L g5412 ( 
.A(n_5088),
.B(n_4979),
.Y(n_5412)
);

INVx3_ASAP7_75t_SL g5413 ( 
.A(n_5205),
.Y(n_5413)
);

AND2x4_ASAP7_75t_L g5414 ( 
.A(n_5113),
.B(n_4793),
.Y(n_5414)
);

INVx1_ASAP7_75t_L g5415 ( 
.A(n_5118),
.Y(n_5415)
);

BUFx12f_ASAP7_75t_L g5416 ( 
.A(n_5213),
.Y(n_5416)
);

BUFx3_ASAP7_75t_L g5417 ( 
.A(n_5217),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5119),
.Y(n_5418)
);

NAND2x1p5_ASAP7_75t_L g5419 ( 
.A(n_5124),
.B(n_5023),
.Y(n_5419)
);

NAND2xp5_ASAP7_75t_L g5420 ( 
.A(n_5222),
.B(n_5233),
.Y(n_5420)
);

INVx1_ASAP7_75t_SL g5421 ( 
.A(n_5369),
.Y(n_5421)
);

BUFx3_ASAP7_75t_L g5422 ( 
.A(n_5117),
.Y(n_5422)
);

INVx3_ASAP7_75t_L g5423 ( 
.A(n_5147),
.Y(n_5423)
);

INVx2_ASAP7_75t_L g5424 ( 
.A(n_5091),
.Y(n_5424)
);

BUFx6f_ASAP7_75t_L g5425 ( 
.A(n_5214),
.Y(n_5425)
);

INVx1_ASAP7_75t_SL g5426 ( 
.A(n_5230),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5138),
.Y(n_5427)
);

NOR2xp33_ASAP7_75t_L g5428 ( 
.A(n_5309),
.B(n_4726),
.Y(n_5428)
);

BUFx6f_ASAP7_75t_L g5429 ( 
.A(n_5214),
.Y(n_5429)
);

INVx1_ASAP7_75t_SL g5430 ( 
.A(n_5355),
.Y(n_5430)
);

NAND2xp5_ASAP7_75t_L g5431 ( 
.A(n_5235),
.B(n_4864),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_5120),
.Y(n_5432)
);

INVx1_ASAP7_75t_SL g5433 ( 
.A(n_5199),
.Y(n_5433)
);

INVx2_ASAP7_75t_SL g5434 ( 
.A(n_5192),
.Y(n_5434)
);

BUFx3_ASAP7_75t_L g5435 ( 
.A(n_5117),
.Y(n_5435)
);

INVx2_ASAP7_75t_L g5436 ( 
.A(n_5203),
.Y(n_5436)
);

INVx1_ASAP7_75t_L g5437 ( 
.A(n_5170),
.Y(n_5437)
);

INVx1_ASAP7_75t_L g5438 ( 
.A(n_5172),
.Y(n_5438)
);

BUFx3_ASAP7_75t_L g5439 ( 
.A(n_5192),
.Y(n_5439)
);

INVx3_ASAP7_75t_L g5440 ( 
.A(n_5243),
.Y(n_5440)
);

INVx1_ASAP7_75t_L g5441 ( 
.A(n_5166),
.Y(n_5441)
);

INVx4_ASAP7_75t_L g5442 ( 
.A(n_5192),
.Y(n_5442)
);

HB1xp67_ASAP7_75t_L g5443 ( 
.A(n_5116),
.Y(n_5443)
);

NAND2xp5_ASAP7_75t_L g5444 ( 
.A(n_5349),
.B(n_4998),
.Y(n_5444)
);

INVx8_ASAP7_75t_L g5445 ( 
.A(n_5158),
.Y(n_5445)
);

NAND2x1p5_ASAP7_75t_L g5446 ( 
.A(n_5392),
.B(n_4883),
.Y(n_5446)
);

INVx1_ASAP7_75t_SL g5447 ( 
.A(n_5243),
.Y(n_5447)
);

INVx4_ASAP7_75t_L g5448 ( 
.A(n_5321),
.Y(n_5448)
);

BUFx2_ASAP7_75t_SL g5449 ( 
.A(n_5298),
.Y(n_5449)
);

INVx8_ASAP7_75t_L g5450 ( 
.A(n_5321),
.Y(n_5450)
);

AND2x2_ASAP7_75t_L g5451 ( 
.A(n_5164),
.B(n_4905),
.Y(n_5451)
);

BUFx4_ASAP7_75t_SL g5452 ( 
.A(n_5377),
.Y(n_5452)
);

BUFx10_ASAP7_75t_L g5453 ( 
.A(n_5133),
.Y(n_5453)
);

INVx1_ASAP7_75t_SL g5454 ( 
.A(n_5121),
.Y(n_5454)
);

INVx1_ASAP7_75t_L g5455 ( 
.A(n_5087),
.Y(n_5455)
);

CKINVDCx6p67_ASAP7_75t_R g5456 ( 
.A(n_5083),
.Y(n_5456)
);

BUFx6f_ASAP7_75t_L g5457 ( 
.A(n_5326),
.Y(n_5457)
);

NOR2xp67_ASAP7_75t_SL g5458 ( 
.A(n_5276),
.B(n_4994),
.Y(n_5458)
);

BUFx12f_ASAP7_75t_L g5459 ( 
.A(n_5389),
.Y(n_5459)
);

CKINVDCx5p33_ASAP7_75t_R g5460 ( 
.A(n_5256),
.Y(n_5460)
);

BUFx6f_ASAP7_75t_L g5461 ( 
.A(n_5326),
.Y(n_5461)
);

AND2x4_ASAP7_75t_L g5462 ( 
.A(n_5113),
.B(n_4894),
.Y(n_5462)
);

BUFx2_ASAP7_75t_L g5463 ( 
.A(n_5158),
.Y(n_5463)
);

INVx3_ASAP7_75t_L g5464 ( 
.A(n_5370),
.Y(n_5464)
);

INVx5_ASAP7_75t_L g5465 ( 
.A(n_5396),
.Y(n_5465)
);

BUFx3_ASAP7_75t_L g5466 ( 
.A(n_5168),
.Y(n_5466)
);

BUFx3_ASAP7_75t_L g5467 ( 
.A(n_5115),
.Y(n_5467)
);

INVx2_ASAP7_75t_L g5468 ( 
.A(n_5254),
.Y(n_5468)
);

INVx2_ASAP7_75t_L g5469 ( 
.A(n_5265),
.Y(n_5469)
);

INVx8_ASAP7_75t_L g5470 ( 
.A(n_5396),
.Y(n_5470)
);

BUFx6f_ASAP7_75t_L g5471 ( 
.A(n_5343),
.Y(n_5471)
);

BUFx2_ASAP7_75t_L g5472 ( 
.A(n_5232),
.Y(n_5472)
);

INVx4_ASAP7_75t_L g5473 ( 
.A(n_5375),
.Y(n_5473)
);

INVx5_ASAP7_75t_SL g5474 ( 
.A(n_5186),
.Y(n_5474)
);

INVx1_ASAP7_75t_SL g5475 ( 
.A(n_5208),
.Y(n_5475)
);

INVxp67_ASAP7_75t_SL g5476 ( 
.A(n_5173),
.Y(n_5476)
);

AOI22xp33_ASAP7_75t_L g5477 ( 
.A1(n_5167),
.A2(n_4816),
.B1(n_5068),
.B2(n_5035),
.Y(n_5477)
);

INVx3_ASAP7_75t_L g5478 ( 
.A(n_5137),
.Y(n_5478)
);

BUFx2_ASAP7_75t_L g5479 ( 
.A(n_5232),
.Y(n_5479)
);

INVx1_ASAP7_75t_SL g5480 ( 
.A(n_5372),
.Y(n_5480)
);

INVxp67_ASAP7_75t_SL g5481 ( 
.A(n_5111),
.Y(n_5481)
);

CKINVDCx5p33_ASAP7_75t_R g5482 ( 
.A(n_5142),
.Y(n_5482)
);

BUFx6f_ASAP7_75t_L g5483 ( 
.A(n_5343),
.Y(n_5483)
);

INVxp33_ASAP7_75t_L g5484 ( 
.A(n_5290),
.Y(n_5484)
);

BUFx6f_ASAP7_75t_L g5485 ( 
.A(n_5333),
.Y(n_5485)
);

NOR2xp33_ASAP7_75t_L g5486 ( 
.A(n_5359),
.B(n_4876),
.Y(n_5486)
);

CKINVDCx8_ASAP7_75t_R g5487 ( 
.A(n_5396),
.Y(n_5487)
);

INVx8_ASAP7_75t_L g5488 ( 
.A(n_5186),
.Y(n_5488)
);

BUFx3_ASAP7_75t_L g5489 ( 
.A(n_5385),
.Y(n_5489)
);

CKINVDCx5p33_ASAP7_75t_R g5490 ( 
.A(n_5183),
.Y(n_5490)
);

INVx3_ASAP7_75t_SL g5491 ( 
.A(n_5095),
.Y(n_5491)
);

BUFx5_ASAP7_75t_L g5492 ( 
.A(n_5141),
.Y(n_5492)
);

INVx4_ASAP7_75t_L g5493 ( 
.A(n_5388),
.Y(n_5493)
);

BUFx6f_ASAP7_75t_L g5494 ( 
.A(n_5314),
.Y(n_5494)
);

INVx2_ASAP7_75t_SL g5495 ( 
.A(n_5090),
.Y(n_5495)
);

CKINVDCx14_ASAP7_75t_R g5496 ( 
.A(n_5184),
.Y(n_5496)
);

BUFx3_ASAP7_75t_L g5497 ( 
.A(n_5134),
.Y(n_5497)
);

CKINVDCx11_ASAP7_75t_R g5498 ( 
.A(n_5317),
.Y(n_5498)
);

BUFx3_ASAP7_75t_L g5499 ( 
.A(n_5344),
.Y(n_5499)
);

INVx3_ASAP7_75t_L g5500 ( 
.A(n_5141),
.Y(n_5500)
);

BUFx2_ASAP7_75t_SL g5501 ( 
.A(n_5127),
.Y(n_5501)
);

INVx2_ASAP7_75t_L g5502 ( 
.A(n_5294),
.Y(n_5502)
);

BUFx5_ASAP7_75t_L g5503 ( 
.A(n_5284),
.Y(n_5503)
);

BUFx24_ASAP7_75t_L g5504 ( 
.A(n_5225),
.Y(n_5504)
);

AOI22xp33_ASAP7_75t_L g5505 ( 
.A1(n_5167),
.A2(n_4735),
.B1(n_4715),
.B2(n_4907),
.Y(n_5505)
);

BUFx2_ASAP7_75t_L g5506 ( 
.A(n_5104),
.Y(n_5506)
);

HB1xp67_ASAP7_75t_L g5507 ( 
.A(n_5182),
.Y(n_5507)
);

INVx1_ASAP7_75t_L g5508 ( 
.A(n_5300),
.Y(n_5508)
);

INVx1_ASAP7_75t_SL g5509 ( 
.A(n_5374),
.Y(n_5509)
);

INVx1_ASAP7_75t_SL g5510 ( 
.A(n_5153),
.Y(n_5510)
);

NAND2x1p5_ASAP7_75t_L g5511 ( 
.A(n_5281),
.B(n_4916),
.Y(n_5511)
);

NAND2xp5_ASAP7_75t_L g5512 ( 
.A(n_5365),
.B(n_4822),
.Y(n_5512)
);

INVx4_ASAP7_75t_L g5513 ( 
.A(n_5305),
.Y(n_5513)
);

BUFx6f_ASAP7_75t_L g5514 ( 
.A(n_5156),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5301),
.Y(n_5515)
);

INVx1_ASAP7_75t_SL g5516 ( 
.A(n_5316),
.Y(n_5516)
);

NAND2xp5_ASAP7_75t_L g5517 ( 
.A(n_5395),
.B(n_4860),
.Y(n_5517)
);

INVx4_ASAP7_75t_L g5518 ( 
.A(n_5107),
.Y(n_5518)
);

AND2x2_ASAP7_75t_L g5519 ( 
.A(n_5097),
.B(n_4868),
.Y(n_5519)
);

BUFx2_ASAP7_75t_L g5520 ( 
.A(n_5151),
.Y(n_5520)
);

CKINVDCx8_ASAP7_75t_R g5521 ( 
.A(n_5262),
.Y(n_5521)
);

BUFx12f_ASAP7_75t_L g5522 ( 
.A(n_5287),
.Y(n_5522)
);

INVx1_ASAP7_75t_L g5523 ( 
.A(n_5098),
.Y(n_5523)
);

INVx6_ASAP7_75t_SL g5524 ( 
.A(n_5219),
.Y(n_5524)
);

HB1xp67_ASAP7_75t_L g5525 ( 
.A(n_5148),
.Y(n_5525)
);

INVx1_ASAP7_75t_L g5526 ( 
.A(n_5146),
.Y(n_5526)
);

BUFx2_ASAP7_75t_L g5527 ( 
.A(n_5155),
.Y(n_5527)
);

NAND2xp5_ASAP7_75t_L g5528 ( 
.A(n_5399),
.B(n_4861),
.Y(n_5528)
);

NOR2xp33_ASAP7_75t_L g5529 ( 
.A(n_5364),
.B(n_4765),
.Y(n_5529)
);

INVx1_ASAP7_75t_L g5530 ( 
.A(n_5157),
.Y(n_5530)
);

INVx3_ASAP7_75t_L g5531 ( 
.A(n_5106),
.Y(n_5531)
);

BUFx6f_ASAP7_75t_L g5532 ( 
.A(n_5160),
.Y(n_5532)
);

INVx4_ASAP7_75t_L g5533 ( 
.A(n_5331),
.Y(n_5533)
);

INVx4_ASAP7_75t_L g5534 ( 
.A(n_5320),
.Y(n_5534)
);

BUFx2_ASAP7_75t_L g5535 ( 
.A(n_5162),
.Y(n_5535)
);

INVx2_ASAP7_75t_SL g5536 ( 
.A(n_5100),
.Y(n_5536)
);

BUFx5_ASAP7_75t_L g5537 ( 
.A(n_5335),
.Y(n_5537)
);

BUFx4_ASAP7_75t_SL g5538 ( 
.A(n_5244),
.Y(n_5538)
);

INVx1_ASAP7_75t_SL g5539 ( 
.A(n_5313),
.Y(n_5539)
);

INVx2_ASAP7_75t_L g5540 ( 
.A(n_5171),
.Y(n_5540)
);

BUFx12f_ASAP7_75t_L g5541 ( 
.A(n_5169),
.Y(n_5541)
);

INVx1_ASAP7_75t_L g5542 ( 
.A(n_5159),
.Y(n_5542)
);

INVx1_ASAP7_75t_SL g5543 ( 
.A(n_5224),
.Y(n_5543)
);

INVx1_ASAP7_75t_L g5544 ( 
.A(n_5161),
.Y(n_5544)
);

INVx6_ASAP7_75t_SL g5545 ( 
.A(n_5196),
.Y(n_5545)
);

INVx2_ASAP7_75t_SL g5546 ( 
.A(n_5163),
.Y(n_5546)
);

BUFx2_ASAP7_75t_L g5547 ( 
.A(n_5149),
.Y(n_5547)
);

INVxp67_ASAP7_75t_SL g5548 ( 
.A(n_5102),
.Y(n_5548)
);

NOR2xp33_ASAP7_75t_L g5549 ( 
.A(n_5334),
.B(n_4783),
.Y(n_5549)
);

INVx4_ASAP7_75t_L g5550 ( 
.A(n_5122),
.Y(n_5550)
);

BUFx3_ASAP7_75t_L g5551 ( 
.A(n_5216),
.Y(n_5551)
);

INVx1_ASAP7_75t_L g5552 ( 
.A(n_5176),
.Y(n_5552)
);

BUFx2_ASAP7_75t_SL g5553 ( 
.A(n_5112),
.Y(n_5553)
);

BUFx8_ASAP7_75t_L g5554 ( 
.A(n_5273),
.Y(n_5554)
);

NAND2x1p5_ASAP7_75t_L g5555 ( 
.A(n_5226),
.B(n_4945),
.Y(n_5555)
);

OR2x6_ASAP7_75t_L g5556 ( 
.A(n_5109),
.B(n_4884),
.Y(n_5556)
);

BUFx6f_ASAP7_75t_L g5557 ( 
.A(n_5242),
.Y(n_5557)
);

AOI22xp33_ASAP7_75t_SL g5558 ( 
.A1(n_5255),
.A2(n_4923),
.B1(n_4840),
.B2(n_5072),
.Y(n_5558)
);

INVx1_ASAP7_75t_L g5559 ( 
.A(n_5180),
.Y(n_5559)
);

BUFx2_ASAP7_75t_L g5560 ( 
.A(n_5367),
.Y(n_5560)
);

CKINVDCx5p33_ASAP7_75t_R g5561 ( 
.A(n_5179),
.Y(n_5561)
);

INVx5_ASAP7_75t_L g5562 ( 
.A(n_5328),
.Y(n_5562)
);

HB1xp67_ASAP7_75t_L g5563 ( 
.A(n_5132),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_5081),
.Y(n_5564)
);

BUFx6f_ASAP7_75t_L g5565 ( 
.A(n_5165),
.Y(n_5565)
);

INVx2_ASAP7_75t_SL g5566 ( 
.A(n_5324),
.Y(n_5566)
);

INVx3_ASAP7_75t_L g5567 ( 
.A(n_5140),
.Y(n_5567)
);

BUFx3_ASAP7_75t_L g5568 ( 
.A(n_5325),
.Y(n_5568)
);

INVx4_ASAP7_75t_L g5569 ( 
.A(n_5082),
.Y(n_5569)
);

INVx2_ASAP7_75t_L g5570 ( 
.A(n_5130),
.Y(n_5570)
);

INVx6_ASAP7_75t_L g5571 ( 
.A(n_5105),
.Y(n_5571)
);

BUFx12f_ASAP7_75t_L g5572 ( 
.A(n_5200),
.Y(n_5572)
);

INVx3_ASAP7_75t_L g5573 ( 
.A(n_5128),
.Y(n_5573)
);

INVx2_ASAP7_75t_L g5574 ( 
.A(n_5089),
.Y(n_5574)
);

BUFx12f_ASAP7_75t_L g5575 ( 
.A(n_5178),
.Y(n_5575)
);

INVx5_ASAP7_75t_L g5576 ( 
.A(n_5391),
.Y(n_5576)
);

BUFx2_ASAP7_75t_SL g5577 ( 
.A(n_5394),
.Y(n_5577)
);

INVx1_ASAP7_75t_L g5578 ( 
.A(n_5181),
.Y(n_5578)
);

INVx2_ASAP7_75t_L g5579 ( 
.A(n_5101),
.Y(n_5579)
);

BUFx3_ASAP7_75t_L g5580 ( 
.A(n_5332),
.Y(n_5580)
);

INVx3_ASAP7_75t_L g5581 ( 
.A(n_5277),
.Y(n_5581)
);

BUFx3_ASAP7_75t_L g5582 ( 
.A(n_5215),
.Y(n_5582)
);

INVx1_ASAP7_75t_L g5583 ( 
.A(n_5191),
.Y(n_5583)
);

NAND2xp5_ASAP7_75t_L g5584 ( 
.A(n_5101),
.B(n_4865),
.Y(n_5584)
);

BUFx4f_ASAP7_75t_SL g5585 ( 
.A(n_5259),
.Y(n_5585)
);

BUFx5_ASAP7_75t_L g5586 ( 
.A(n_5221),
.Y(n_5586)
);

BUFx6f_ASAP7_75t_L g5587 ( 
.A(n_5093),
.Y(n_5587)
);

INVx3_ASAP7_75t_L g5588 ( 
.A(n_5354),
.Y(n_5588)
);

CKINVDCx20_ASAP7_75t_R g5589 ( 
.A(n_5336),
.Y(n_5589)
);

AOI22xp33_ASAP7_75t_L g5590 ( 
.A1(n_5234),
.A2(n_4885),
.B1(n_5043),
.B2(n_4995),
.Y(n_5590)
);

INVx1_ASAP7_75t_SL g5591 ( 
.A(n_5342),
.Y(n_5591)
);

BUFx3_ASAP7_75t_L g5592 ( 
.A(n_5193),
.Y(n_5592)
);

INVx5_ASAP7_75t_SL g5593 ( 
.A(n_5291),
.Y(n_5593)
);

HB1xp67_ASAP7_75t_L g5594 ( 
.A(n_5403),
.Y(n_5594)
);

CKINVDCx20_ASAP7_75t_R g5595 ( 
.A(n_5408),
.Y(n_5595)
);

AND2x2_ASAP7_75t_L g5596 ( 
.A(n_5542),
.B(n_5086),
.Y(n_5596)
);

AND2x2_ASAP7_75t_L g5597 ( 
.A(n_5544),
.B(n_5094),
.Y(n_5597)
);

AO21x2_ASAP7_75t_L g5598 ( 
.A1(n_5548),
.A2(n_5187),
.B(n_5125),
.Y(n_5598)
);

HB1xp67_ASAP7_75t_L g5599 ( 
.A(n_5454),
.Y(n_5599)
);

INVx1_ASAP7_75t_SL g5600 ( 
.A(n_5413),
.Y(n_5600)
);

HB1xp67_ASAP7_75t_L g5601 ( 
.A(n_5497),
.Y(n_5601)
);

OAI221xp5_ASAP7_75t_L g5602 ( 
.A1(n_5511),
.A2(n_5397),
.B1(n_5341),
.B2(n_5295),
.C(n_5084),
.Y(n_5602)
);

AND2x4_ASAP7_75t_L g5603 ( 
.A(n_5466),
.B(n_5136),
.Y(n_5603)
);

INVx2_ASAP7_75t_L g5604 ( 
.A(n_5503),
.Y(n_5604)
);

OAI21x1_ASAP7_75t_L g5605 ( 
.A1(n_5567),
.A2(n_5129),
.B(n_5150),
.Y(n_5605)
);

NOR2xp67_ASAP7_75t_L g5606 ( 
.A(n_5442),
.B(n_5346),
.Y(n_5606)
);

INVx1_ASAP7_75t_SL g5607 ( 
.A(n_5405),
.Y(n_5607)
);

OAI21x1_ASAP7_75t_L g5608 ( 
.A1(n_5573),
.A2(n_5143),
.B(n_5123),
.Y(n_5608)
);

AO21x2_ASAP7_75t_L g5609 ( 
.A1(n_5563),
.A2(n_5227),
.B(n_5110),
.Y(n_5609)
);

INVx2_ASAP7_75t_SL g5610 ( 
.A(n_5402),
.Y(n_5610)
);

NAND2xp5_ASAP7_75t_L g5611 ( 
.A(n_5507),
.B(n_5318),
.Y(n_5611)
);

INVx2_ASAP7_75t_L g5612 ( 
.A(n_5503),
.Y(n_5612)
);

OAI21x1_ASAP7_75t_L g5613 ( 
.A1(n_5531),
.A2(n_5579),
.B(n_5570),
.Y(n_5613)
);

NAND2x1p5_ASAP7_75t_L g5614 ( 
.A(n_5407),
.B(n_5270),
.Y(n_5614)
);

OAI21xp5_ASAP7_75t_L g5615 ( 
.A1(n_5484),
.A2(n_5263),
.B(n_5356),
.Y(n_5615)
);

NOR2xp33_ASAP7_75t_L g5616 ( 
.A(n_5456),
.B(n_5382),
.Y(n_5616)
);

AND2x4_ASAP7_75t_L g5617 ( 
.A(n_5414),
.B(n_5152),
.Y(n_5617)
);

OAI21x1_ASAP7_75t_L g5618 ( 
.A1(n_5478),
.A2(n_5103),
.B(n_5108),
.Y(n_5618)
);

OAI21x1_ASAP7_75t_L g5619 ( 
.A1(n_5574),
.A2(n_5114),
.B(n_5139),
.Y(n_5619)
);

INVx1_ASAP7_75t_L g5620 ( 
.A(n_5406),
.Y(n_5620)
);

OAI21x1_ASAP7_75t_L g5621 ( 
.A1(n_5476),
.A2(n_5096),
.B(n_5174),
.Y(n_5621)
);

OAI21x1_ASAP7_75t_SL g5622 ( 
.A1(n_5495),
.A2(n_5310),
.B(n_5285),
.Y(n_5622)
);

NAND2xp5_ASAP7_75t_L g5623 ( 
.A(n_5481),
.B(n_5175),
.Y(n_5623)
);

INVx1_ASAP7_75t_L g5624 ( 
.A(n_5415),
.Y(n_5624)
);

NAND2xp5_ASAP7_75t_L g5625 ( 
.A(n_5523),
.B(n_5175),
.Y(n_5625)
);

OAI21xp5_ASAP7_75t_L g5626 ( 
.A1(n_5473),
.A2(n_5189),
.B(n_5237),
.Y(n_5626)
);

INVx3_ASAP7_75t_SL g5627 ( 
.A(n_5411),
.Y(n_5627)
);

AO31x2_ASAP7_75t_L g5628 ( 
.A1(n_5550),
.A2(n_5154),
.A3(n_5271),
.B(n_5280),
.Y(n_5628)
);

NAND2xp5_ASAP7_75t_L g5629 ( 
.A(n_5441),
.B(n_5267),
.Y(n_5629)
);

OAI22xp5_ASAP7_75t_L g5630 ( 
.A1(n_5487),
.A2(n_5283),
.B1(n_5376),
.B2(n_5247),
.Y(n_5630)
);

OAI21x1_ASAP7_75t_L g5631 ( 
.A1(n_5564),
.A2(n_5145),
.B(n_5135),
.Y(n_5631)
);

BUFx6f_ASAP7_75t_L g5632 ( 
.A(n_5410),
.Y(n_5632)
);

HB1xp67_ASAP7_75t_L g5633 ( 
.A(n_5472),
.Y(n_5633)
);

AO31x2_ASAP7_75t_L g5634 ( 
.A1(n_5569),
.A2(n_5245),
.A3(n_5144),
.B(n_5238),
.Y(n_5634)
);

NAND3xp33_ASAP7_75t_L g5635 ( 
.A(n_5584),
.B(n_5131),
.C(n_5218),
.Y(n_5635)
);

AOI22xp33_ASAP7_75t_L g5636 ( 
.A1(n_5572),
.A2(n_5299),
.B1(n_5347),
.B2(n_5323),
.Y(n_5636)
);

AND2x6_ASAP7_75t_L g5637 ( 
.A(n_5474),
.B(n_4919),
.Y(n_5637)
);

OA21x2_ASAP7_75t_L g5638 ( 
.A1(n_5535),
.A2(n_5398),
.B(n_5099),
.Y(n_5638)
);

AOI22xp33_ASAP7_75t_L g5639 ( 
.A1(n_5541),
.A2(n_5212),
.B1(n_5240),
.B2(n_5195),
.Y(n_5639)
);

AND2x2_ASAP7_75t_L g5640 ( 
.A(n_5540),
.B(n_5267),
.Y(n_5640)
);

OA21x2_ASAP7_75t_L g5641 ( 
.A1(n_5482),
.A2(n_5520),
.B(n_5547),
.Y(n_5641)
);

AO21x2_ASAP7_75t_L g5642 ( 
.A1(n_5455),
.A2(n_5420),
.B(n_5404),
.Y(n_5642)
);

INVx1_ASAP7_75t_L g5643 ( 
.A(n_5418),
.Y(n_5643)
);

BUFx3_ASAP7_75t_L g5644 ( 
.A(n_5409),
.Y(n_5644)
);

AOI21xp33_ASAP7_75t_L g5645 ( 
.A1(n_5554),
.A2(n_5575),
.B(n_5577),
.Y(n_5645)
);

OAI21x1_ASAP7_75t_L g5646 ( 
.A1(n_5581),
.A2(n_5357),
.B(n_5231),
.Y(n_5646)
);

BUFx2_ASAP7_75t_L g5647 ( 
.A(n_5423),
.Y(n_5647)
);

OAI21x1_ASAP7_75t_L g5648 ( 
.A1(n_5588),
.A2(n_5188),
.B(n_5223),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5515),
.B(n_5360),
.Y(n_5649)
);

NAND2x1p5_ASAP7_75t_L g5650 ( 
.A(n_5422),
.B(n_5329),
.Y(n_5650)
);

INVx1_ASAP7_75t_L g5651 ( 
.A(n_5432),
.Y(n_5651)
);

AND2x4_ASAP7_75t_L g5652 ( 
.A(n_5465),
.B(n_5378),
.Y(n_5652)
);

NAND2xp5_ASAP7_75t_L g5653 ( 
.A(n_5526),
.B(n_5229),
.Y(n_5653)
);

AO31x2_ASAP7_75t_L g5654 ( 
.A1(n_5527),
.A2(n_5250),
.A3(n_5264),
.B(n_5248),
.Y(n_5654)
);

AO21x2_ASAP7_75t_L g5655 ( 
.A1(n_5552),
.A2(n_5345),
.B(n_5293),
.Y(n_5655)
);

BUFx3_ASAP7_75t_L g5656 ( 
.A(n_5416),
.Y(n_5656)
);

INVx6_ASAP7_75t_L g5657 ( 
.A(n_5459),
.Y(n_5657)
);

INVx1_ASAP7_75t_L g5658 ( 
.A(n_5437),
.Y(n_5658)
);

AOI21xp5_ASAP7_75t_L g5659 ( 
.A1(n_5470),
.A2(n_5185),
.B(n_5251),
.Y(n_5659)
);

OAI22xp5_ASAP7_75t_L g5660 ( 
.A1(n_5465),
.A2(n_5373),
.B1(n_5286),
.B2(n_5338),
.Y(n_5660)
);

OAI22xp5_ASAP7_75t_L g5661 ( 
.A1(n_5593),
.A2(n_5207),
.B1(n_4985),
.B2(n_5279),
.Y(n_5661)
);

INVx2_ASAP7_75t_L g5662 ( 
.A(n_5503),
.Y(n_5662)
);

INVx2_ASAP7_75t_L g5663 ( 
.A(n_5479),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5438),
.Y(n_5664)
);

NOR2xp33_ASAP7_75t_L g5665 ( 
.A(n_5426),
.B(n_4974),
.Y(n_5665)
);

INVx4_ASAP7_75t_L g5666 ( 
.A(n_5417),
.Y(n_5666)
);

NAND2x1p5_ASAP7_75t_L g5667 ( 
.A(n_5435),
.B(n_5282),
.Y(n_5667)
);

AO31x2_ASAP7_75t_L g5668 ( 
.A1(n_5518),
.A2(n_5296),
.A3(n_5297),
.B(n_5289),
.Y(n_5668)
);

AND2x4_ASAP7_75t_L g5669 ( 
.A(n_5500),
.B(n_5304),
.Y(n_5669)
);

BUFx12f_ASAP7_75t_SL g5670 ( 
.A(n_5513),
.Y(n_5670)
);

AO31x2_ASAP7_75t_L g5671 ( 
.A1(n_5463),
.A2(n_5322),
.A3(n_4666),
.B(n_4671),
.Y(n_5671)
);

AOI22x1_ASAP7_75t_L g5672 ( 
.A1(n_5553),
.A2(n_5400),
.B1(n_5177),
.B2(n_5353),
.Y(n_5672)
);

BUFx2_ASAP7_75t_L g5673 ( 
.A(n_5560),
.Y(n_5673)
);

AO21x2_ASAP7_75t_L g5674 ( 
.A1(n_5559),
.A2(n_5578),
.B(n_5528),
.Y(n_5674)
);

AOI222xp33_ASAP7_75t_L g5675 ( 
.A1(n_5562),
.A2(n_5275),
.B1(n_5261),
.B2(n_5340),
.C1(n_5126),
.C2(n_5386),
.Y(n_5675)
);

AO21x2_ASAP7_75t_L g5676 ( 
.A1(n_5517),
.A2(n_5274),
.B(n_5366),
.Y(n_5676)
);

CKINVDCx20_ASAP7_75t_R g5677 ( 
.A(n_5460),
.Y(n_5677)
);

INVx1_ASAP7_75t_L g5678 ( 
.A(n_5508),
.Y(n_5678)
);

NOR2xp33_ASAP7_75t_L g5679 ( 
.A(n_5496),
.B(n_4895),
.Y(n_5679)
);

INVx1_ASAP7_75t_L g5680 ( 
.A(n_5525),
.Y(n_5680)
);

NAND2xp5_ASAP7_75t_SL g5681 ( 
.A(n_5467),
.B(n_5210),
.Y(n_5681)
);

AND2x4_ASAP7_75t_L g5682 ( 
.A(n_5439),
.B(n_5312),
.Y(n_5682)
);

OAI21x1_ASAP7_75t_L g5683 ( 
.A1(n_5464),
.A2(n_5194),
.B(n_5266),
.Y(n_5683)
);

AO31x2_ASAP7_75t_L g5684 ( 
.A1(n_5506),
.A2(n_4676),
.A3(n_4680),
.B(n_4661),
.Y(n_5684)
);

OAI21x1_ASAP7_75t_L g5685 ( 
.A1(n_5446),
.A2(n_5292),
.B(n_5288),
.Y(n_5685)
);

INVx1_ASAP7_75t_L g5686 ( 
.A(n_5530),
.Y(n_5686)
);

OAI21xp5_ASAP7_75t_L g5687 ( 
.A1(n_5562),
.A2(n_5339),
.B(n_5358),
.Y(n_5687)
);

CKINVDCx5p33_ASAP7_75t_R g5688 ( 
.A(n_5452),
.Y(n_5688)
);

INVx3_ASAP7_75t_L g5689 ( 
.A(n_5524),
.Y(n_5689)
);

HB1xp67_ASAP7_75t_L g5690 ( 
.A(n_5443),
.Y(n_5690)
);

OAI21x1_ASAP7_75t_L g5691 ( 
.A1(n_5555),
.A2(n_5307),
.B(n_5303),
.Y(n_5691)
);

AOI22xp33_ASAP7_75t_L g5692 ( 
.A1(n_5458),
.A2(n_5383),
.B1(n_5246),
.B2(n_5272),
.Y(n_5692)
);

NOR2xp33_ASAP7_75t_L g5693 ( 
.A(n_5434),
.B(n_5475),
.Y(n_5693)
);

OAI21x1_ASAP7_75t_SL g5694 ( 
.A1(n_5533),
.A2(n_5368),
.B(n_4667),
.Y(n_5694)
);

NAND2xp5_ASAP7_75t_L g5695 ( 
.A(n_5583),
.B(n_5211),
.Y(n_5695)
);

AO31x2_ASAP7_75t_L g5696 ( 
.A1(n_5493),
.A2(n_4714),
.A3(n_4719),
.B(n_4707),
.Y(n_5696)
);

BUFx8_ASAP7_75t_L g5697 ( 
.A(n_5401),
.Y(n_5697)
);

AND2x4_ASAP7_75t_L g5698 ( 
.A(n_5421),
.B(n_5308),
.Y(n_5698)
);

OAI21x1_ASAP7_75t_L g5699 ( 
.A1(n_5419),
.A2(n_5201),
.B(n_5197),
.Y(n_5699)
);

OAI22xp5_ASAP7_75t_L g5700 ( 
.A1(n_5556),
.A2(n_4941),
.B1(n_5362),
.B2(n_4897),
.Y(n_5700)
);

HB1xp67_ASAP7_75t_L g5701 ( 
.A(n_5430),
.Y(n_5701)
);

OA21x2_ASAP7_75t_L g5702 ( 
.A1(n_5433),
.A2(n_5206),
.B(n_5202),
.Y(n_5702)
);

AND2x4_ASAP7_75t_L g5703 ( 
.A(n_5489),
.B(n_5546),
.Y(n_5703)
);

INVxp67_ASAP7_75t_SL g5704 ( 
.A(n_5424),
.Y(n_5704)
);

NAND2xp5_ASAP7_75t_L g5705 ( 
.A(n_5536),
.B(n_5211),
.Y(n_5705)
);

AOI21xp5_ASAP7_75t_L g5706 ( 
.A1(n_5488),
.A2(n_4848),
.B(n_4951),
.Y(n_5706)
);

OA21x2_ASAP7_75t_L g5707 ( 
.A1(n_5510),
.A2(n_5348),
.B(n_5249),
.Y(n_5707)
);

OR2x2_ASAP7_75t_L g5708 ( 
.A(n_5427),
.B(n_4982),
.Y(n_5708)
);

OAI21x1_ASAP7_75t_L g5709 ( 
.A1(n_5440),
.A2(n_5257),
.B(n_5252),
.Y(n_5709)
);

AOI22xp33_ASAP7_75t_L g5710 ( 
.A1(n_5571),
.A2(n_4724),
.B1(n_5380),
.B2(n_5384),
.Y(n_5710)
);

INVx2_ASAP7_75t_L g5711 ( 
.A(n_5436),
.Y(n_5711)
);

INVx2_ASAP7_75t_L g5712 ( 
.A(n_5468),
.Y(n_5712)
);

NAND2xp5_ASAP7_75t_L g5713 ( 
.A(n_5412),
.B(n_4899),
.Y(n_5713)
);

BUFx4f_ASAP7_75t_L g5714 ( 
.A(n_5488),
.Y(n_5714)
);

OAI22xp5_ASAP7_75t_L g5715 ( 
.A1(n_5585),
.A2(n_4727),
.B1(n_4993),
.B2(n_4733),
.Y(n_5715)
);

NAND2x1p5_ASAP7_75t_L g5716 ( 
.A(n_5448),
.B(n_4803),
.Y(n_5716)
);

NAND2xp5_ASAP7_75t_SL g5717 ( 
.A(n_5557),
.B(n_5387),
.Y(n_5717)
);

INVx2_ASAP7_75t_L g5718 ( 
.A(n_5469),
.Y(n_5718)
);

OAI21x1_ASAP7_75t_L g5719 ( 
.A1(n_5502),
.A2(n_5236),
.B(n_5350),
.Y(n_5719)
);

OAI21x1_ASAP7_75t_L g5720 ( 
.A1(n_5512),
.A2(n_5545),
.B(n_5444),
.Y(n_5720)
);

INVx2_ASAP7_75t_SL g5721 ( 
.A(n_5450),
.Y(n_5721)
);

NAND2xp5_ASAP7_75t_L g5722 ( 
.A(n_5480),
.B(n_4901),
.Y(n_5722)
);

OA21x2_ASAP7_75t_L g5723 ( 
.A1(n_5431),
.A2(n_4748),
.B(n_4728),
.Y(n_5723)
);

INVx1_ASAP7_75t_L g5724 ( 
.A(n_5451),
.Y(n_5724)
);

INVx2_ASAP7_75t_L g5725 ( 
.A(n_5494),
.Y(n_5725)
);

NAND2xp5_ASAP7_75t_SL g5726 ( 
.A(n_5557),
.B(n_5491),
.Y(n_5726)
);

AOI22xp33_ASAP7_75t_L g5727 ( 
.A1(n_5561),
.A2(n_5589),
.B1(n_5537),
.B2(n_5558),
.Y(n_5727)
);

INVx2_ASAP7_75t_L g5728 ( 
.A(n_5494),
.Y(n_5728)
);

INVx1_ASAP7_75t_L g5729 ( 
.A(n_5594),
.Y(n_5729)
);

OAI22xp5_ASAP7_75t_L g5730 ( 
.A1(n_5601),
.A2(n_5501),
.B1(n_5449),
.B2(n_5516),
.Y(n_5730)
);

INVx2_ASAP7_75t_L g5731 ( 
.A(n_5673),
.Y(n_5731)
);

BUFx2_ASAP7_75t_L g5732 ( 
.A(n_5670),
.Y(n_5732)
);

INVx2_ASAP7_75t_L g5733 ( 
.A(n_5673),
.Y(n_5733)
);

INVx1_ASAP7_75t_L g5734 ( 
.A(n_5686),
.Y(n_5734)
);

INVx1_ASAP7_75t_L g5735 ( 
.A(n_5620),
.Y(n_5735)
);

BUFx4f_ASAP7_75t_L g5736 ( 
.A(n_5657),
.Y(n_5736)
);

INVx2_ASAP7_75t_L g5737 ( 
.A(n_5599),
.Y(n_5737)
);

CKINVDCx20_ASAP7_75t_R g5738 ( 
.A(n_5595),
.Y(n_5738)
);

INVx1_ASAP7_75t_L g5739 ( 
.A(n_5624),
.Y(n_5739)
);

INVx6_ASAP7_75t_L g5740 ( 
.A(n_5697),
.Y(n_5740)
);

INVx2_ASAP7_75t_L g5741 ( 
.A(n_5690),
.Y(n_5741)
);

BUFx3_ASAP7_75t_L g5742 ( 
.A(n_5632),
.Y(n_5742)
);

AND2x2_ASAP7_75t_L g5743 ( 
.A(n_5633),
.B(n_5509),
.Y(n_5743)
);

INVx2_ASAP7_75t_L g5744 ( 
.A(n_5642),
.Y(n_5744)
);

OAI22xp5_ASAP7_75t_L g5745 ( 
.A1(n_5727),
.A2(n_5499),
.B1(n_5582),
.B2(n_5534),
.Y(n_5745)
);

INVx2_ASAP7_75t_L g5746 ( 
.A(n_5711),
.Y(n_5746)
);

BUFx3_ASAP7_75t_L g5747 ( 
.A(n_5632),
.Y(n_5747)
);

CKINVDCx11_ASAP7_75t_R g5748 ( 
.A(n_5677),
.Y(n_5748)
);

AOI22xp33_ASAP7_75t_SL g5749 ( 
.A1(n_5666),
.A2(n_5445),
.B1(n_5522),
.B2(n_5543),
.Y(n_5749)
);

BUFx6f_ASAP7_75t_L g5750 ( 
.A(n_5656),
.Y(n_5750)
);

NAND2x1p5_ASAP7_75t_L g5751 ( 
.A(n_5714),
.B(n_5425),
.Y(n_5751)
);

HB1xp67_ASAP7_75t_L g5752 ( 
.A(n_5704),
.Y(n_5752)
);

AOI22xp5_ASAP7_75t_SL g5753 ( 
.A1(n_5600),
.A2(n_5462),
.B1(n_5490),
.B2(n_5486),
.Y(n_5753)
);

HB1xp67_ASAP7_75t_L g5754 ( 
.A(n_5701),
.Y(n_5754)
);

INVx1_ASAP7_75t_L g5755 ( 
.A(n_5643),
.Y(n_5755)
);

INVx1_ASAP7_75t_L g5756 ( 
.A(n_5651),
.Y(n_5756)
);

AOI22xp33_ASAP7_75t_L g5757 ( 
.A1(n_5602),
.A2(n_5551),
.B1(n_5537),
.B2(n_5576),
.Y(n_5757)
);

INVx2_ASAP7_75t_L g5758 ( 
.A(n_5712),
.Y(n_5758)
);

INVx1_ASAP7_75t_L g5759 ( 
.A(n_5658),
.Y(n_5759)
);

AND2x4_ASAP7_75t_L g5760 ( 
.A(n_5597),
.B(n_5587),
.Y(n_5760)
);

INVx1_ASAP7_75t_L g5761 ( 
.A(n_5664),
.Y(n_5761)
);

OA21x2_ASAP7_75t_L g5762 ( 
.A1(n_5645),
.A2(n_5519),
.B(n_5591),
.Y(n_5762)
);

AO21x2_ASAP7_75t_L g5763 ( 
.A1(n_5613),
.A2(n_5529),
.B(n_5428),
.Y(n_5763)
);

OR2x2_ASAP7_75t_L g5764 ( 
.A(n_5680),
.B(n_5539),
.Y(n_5764)
);

INVx1_ASAP7_75t_L g5765 ( 
.A(n_5678),
.Y(n_5765)
);

INVx1_ASAP7_75t_L g5766 ( 
.A(n_5674),
.Y(n_5766)
);

BUFx2_ASAP7_75t_L g5767 ( 
.A(n_5647),
.Y(n_5767)
);

OAI21x1_ASAP7_75t_L g5768 ( 
.A1(n_5608),
.A2(n_5477),
.B(n_5379),
.Y(n_5768)
);

INVx1_ASAP7_75t_L g5769 ( 
.A(n_5611),
.Y(n_5769)
);

NAND2xp5_ASAP7_75t_L g5770 ( 
.A(n_5640),
.B(n_5566),
.Y(n_5770)
);

INVx2_ASAP7_75t_SL g5771 ( 
.A(n_5657),
.Y(n_5771)
);

AO21x1_ASAP7_75t_L g5772 ( 
.A1(n_5681),
.A2(n_5504),
.B(n_5549),
.Y(n_5772)
);

INVx2_ASAP7_75t_L g5773 ( 
.A(n_5718),
.Y(n_5773)
);

INVx1_ASAP7_75t_L g5774 ( 
.A(n_5724),
.Y(n_5774)
);

INVx1_ASAP7_75t_L g5775 ( 
.A(n_5695),
.Y(n_5775)
);

INVx1_ASAP7_75t_L g5776 ( 
.A(n_5708),
.Y(n_5776)
);

INVx2_ASAP7_75t_SL g5777 ( 
.A(n_5627),
.Y(n_5777)
);

INVx1_ASAP7_75t_L g5778 ( 
.A(n_5708),
.Y(n_5778)
);

NAND2x1p5_ASAP7_75t_L g5779 ( 
.A(n_5607),
.B(n_5425),
.Y(n_5779)
);

AOI22xp33_ASAP7_75t_L g5780 ( 
.A1(n_5672),
.A2(n_5537),
.B1(n_5576),
.B2(n_5568),
.Y(n_5780)
);

INVx1_ASAP7_75t_L g5781 ( 
.A(n_5629),
.Y(n_5781)
);

INVx1_ASAP7_75t_L g5782 ( 
.A(n_5649),
.Y(n_5782)
);

NAND2x1p5_ASAP7_75t_L g5783 ( 
.A(n_5689),
.B(n_5429),
.Y(n_5783)
);

OA21x2_ASAP7_75t_L g5784 ( 
.A1(n_5720),
.A2(n_5447),
.B(n_5538),
.Y(n_5784)
);

HB1xp67_ASAP7_75t_L g5785 ( 
.A(n_5663),
.Y(n_5785)
);

AND2x2_ASAP7_75t_L g5786 ( 
.A(n_5703),
.B(n_5492),
.Y(n_5786)
);

NAND2x1p5_ASAP7_75t_L g5787 ( 
.A(n_5644),
.B(n_5429),
.Y(n_5787)
);

INVx4_ASAP7_75t_SL g5788 ( 
.A(n_5637),
.Y(n_5788)
);

NAND2x1p5_ASAP7_75t_L g5789 ( 
.A(n_5610),
.B(n_5457),
.Y(n_5789)
);

INVx1_ASAP7_75t_L g5790 ( 
.A(n_5705),
.Y(n_5790)
);

INVx1_ASAP7_75t_L g5791 ( 
.A(n_5653),
.Y(n_5791)
);

INVx1_ASAP7_75t_L g5792 ( 
.A(n_5640),
.Y(n_5792)
);

HB1xp67_ASAP7_75t_L g5793 ( 
.A(n_5603),
.Y(n_5793)
);

BUFx3_ASAP7_75t_L g5794 ( 
.A(n_5688),
.Y(n_5794)
);

AND2x2_ASAP7_75t_L g5795 ( 
.A(n_5725),
.B(n_5492),
.Y(n_5795)
);

INVx1_ASAP7_75t_L g5796 ( 
.A(n_5625),
.Y(n_5796)
);

CKINVDCx11_ASAP7_75t_R g5797 ( 
.A(n_5652),
.Y(n_5797)
);

CKINVDCx11_ASAP7_75t_R g5798 ( 
.A(n_5728),
.Y(n_5798)
);

INVx1_ASAP7_75t_L g5799 ( 
.A(n_5623),
.Y(n_5799)
);

INVx1_ASAP7_75t_L g5800 ( 
.A(n_5722),
.Y(n_5800)
);

CKINVDCx5p33_ASAP7_75t_R g5801 ( 
.A(n_5693),
.Y(n_5801)
);

CKINVDCx14_ASAP7_75t_R g5802 ( 
.A(n_5637),
.Y(n_5802)
);

AND2x2_ASAP7_75t_L g5803 ( 
.A(n_5617),
.B(n_5492),
.Y(n_5803)
);

CKINVDCx20_ASAP7_75t_R g5804 ( 
.A(n_5721),
.Y(n_5804)
);

INVx2_ASAP7_75t_L g5805 ( 
.A(n_5698),
.Y(n_5805)
);

OA21x2_ASAP7_75t_L g5806 ( 
.A1(n_5618),
.A2(n_4754),
.B(n_4752),
.Y(n_5806)
);

NAND2xp5_ASAP7_75t_L g5807 ( 
.A(n_5654),
.B(n_5592),
.Y(n_5807)
);

CKINVDCx10_ASAP7_75t_R g5808 ( 
.A(n_5616),
.Y(n_5808)
);

CKINVDCx20_ASAP7_75t_R g5809 ( 
.A(n_5679),
.Y(n_5809)
);

INVx2_ASAP7_75t_L g5810 ( 
.A(n_5597),
.Y(n_5810)
);

OAI22xp5_ASAP7_75t_L g5811 ( 
.A1(n_5606),
.A2(n_5521),
.B1(n_5580),
.B2(n_5505),
.Y(n_5811)
);

AOI22xp33_ASAP7_75t_L g5812 ( 
.A1(n_5598),
.A2(n_5590),
.B1(n_5586),
.B2(n_5498),
.Y(n_5812)
);

INVx3_ASAP7_75t_L g5813 ( 
.A(n_5637),
.Y(n_5813)
);

BUFx6f_ASAP7_75t_L g5814 ( 
.A(n_5716),
.Y(n_5814)
);

AOI22xp33_ASAP7_75t_L g5815 ( 
.A1(n_5661),
.A2(n_5586),
.B1(n_5453),
.B2(n_5514),
.Y(n_5815)
);

INVx1_ASAP7_75t_L g5816 ( 
.A(n_5713),
.Y(n_5816)
);

CKINVDCx20_ASAP7_75t_R g5817 ( 
.A(n_5665),
.Y(n_5817)
);

OAI22xp5_ASAP7_75t_L g5818 ( 
.A1(n_5636),
.A2(n_5514),
.B1(n_5485),
.B2(n_5450),
.Y(n_5818)
);

OAI22xp5_ASAP7_75t_L g5819 ( 
.A1(n_5614),
.A2(n_5485),
.B1(n_5457),
.B2(n_5471),
.Y(n_5819)
);

AOI22xp33_ASAP7_75t_L g5820 ( 
.A1(n_5635),
.A2(n_5586),
.B1(n_4950),
.B2(n_5390),
.Y(n_5820)
);

BUFx10_ASAP7_75t_L g5821 ( 
.A(n_5682),
.Y(n_5821)
);

AOI22xp33_ASAP7_75t_L g5822 ( 
.A1(n_5694),
.A2(n_5080),
.B1(n_5306),
.B2(n_4767),
.Y(n_5822)
);

INVx1_ASAP7_75t_L g5823 ( 
.A(n_5596),
.Y(n_5823)
);

INVx1_ASAP7_75t_L g5824 ( 
.A(n_5596),
.Y(n_5824)
);

AOI21x1_ASAP7_75t_L g5825 ( 
.A1(n_5726),
.A2(n_4781),
.B(n_4760),
.Y(n_5825)
);

NAND2x1p5_ASAP7_75t_L g5826 ( 
.A(n_5699),
.B(n_5461),
.Y(n_5826)
);

AND2x2_ASAP7_75t_L g5827 ( 
.A(n_5641),
.B(n_5532),
.Y(n_5827)
);

AOI22xp33_ASAP7_75t_SL g5828 ( 
.A1(n_5638),
.A2(n_5565),
.B1(n_5587),
.B2(n_5532),
.Y(n_5828)
);

AND2x2_ASAP7_75t_L g5829 ( 
.A(n_5669),
.B(n_5565),
.Y(n_5829)
);

INVx1_ASAP7_75t_L g5830 ( 
.A(n_5654),
.Y(n_5830)
);

INVx1_ASAP7_75t_SL g5831 ( 
.A(n_5723),
.Y(n_5831)
);

BUFx2_ASAP7_75t_L g5832 ( 
.A(n_5702),
.Y(n_5832)
);

INVx1_ASAP7_75t_L g5833 ( 
.A(n_5684),
.Y(n_5833)
);

AO21x1_ASAP7_75t_L g5834 ( 
.A1(n_5659),
.A2(n_4877),
.B(n_4871),
.Y(n_5834)
);

INVx2_ASAP7_75t_L g5835 ( 
.A(n_5604),
.Y(n_5835)
);

NAND2xp5_ASAP7_75t_L g5836 ( 
.A(n_5684),
.B(n_5461),
.Y(n_5836)
);

AO21x2_ASAP7_75t_L g5837 ( 
.A1(n_5609),
.A2(n_5605),
.B(n_5717),
.Y(n_5837)
);

INVx1_ASAP7_75t_SL g5838 ( 
.A(n_5650),
.Y(n_5838)
);

HB1xp67_ASAP7_75t_L g5839 ( 
.A(n_5668),
.Y(n_5839)
);

HB1xp67_ASAP7_75t_L g5840 ( 
.A(n_5668),
.Y(n_5840)
);

INVx1_ASAP7_75t_L g5841 ( 
.A(n_5696),
.Y(n_5841)
);

OAI21x1_ASAP7_75t_L g5842 ( 
.A1(n_5631),
.A2(n_5363),
.B(n_5361),
.Y(n_5842)
);

INVx1_ASAP7_75t_L g5843 ( 
.A(n_5696),
.Y(n_5843)
);

BUFx12f_ASAP7_75t_L g5844 ( 
.A(n_5667),
.Y(n_5844)
);

INVx2_ASAP7_75t_L g5845 ( 
.A(n_5612),
.Y(n_5845)
);

OAI21x1_ASAP7_75t_L g5846 ( 
.A1(n_5619),
.A2(n_5327),
.B(n_4997),
.Y(n_5846)
);

INVx2_ASAP7_75t_L g5847 ( 
.A(n_5662),
.Y(n_5847)
);

OA21x2_ASAP7_75t_L g5848 ( 
.A1(n_5621),
.A2(n_4786),
.B(n_4785),
.Y(n_5848)
);

INVx2_ASAP7_75t_SL g5849 ( 
.A(n_5709),
.Y(n_5849)
);

HB1xp67_ASAP7_75t_L g5850 ( 
.A(n_5719),
.Y(n_5850)
);

BUFx3_ASAP7_75t_L g5851 ( 
.A(n_5622),
.Y(n_5851)
);

INVx1_ASAP7_75t_L g5852 ( 
.A(n_5648),
.Y(n_5852)
);

INVx1_ASAP7_75t_L g5853 ( 
.A(n_5646),
.Y(n_5853)
);

INVx2_ASAP7_75t_L g5854 ( 
.A(n_5671),
.Y(n_5854)
);

INVx2_ASAP7_75t_SL g5855 ( 
.A(n_5671),
.Y(n_5855)
);

AND2x2_ASAP7_75t_L g5856 ( 
.A(n_5634),
.B(n_5471),
.Y(n_5856)
);

INVx1_ASAP7_75t_L g5857 ( 
.A(n_5707),
.Y(n_5857)
);

HB1xp67_ASAP7_75t_L g5858 ( 
.A(n_5628),
.Y(n_5858)
);

INVxp67_ASAP7_75t_L g5859 ( 
.A(n_5615),
.Y(n_5859)
);

OA21x2_ASAP7_75t_L g5860 ( 
.A1(n_5772),
.A2(n_5691),
.B(n_5685),
.Y(n_5860)
);

CKINVDCx11_ASAP7_75t_R g5861 ( 
.A(n_5748),
.Y(n_5861)
);

CKINVDCx5p33_ASAP7_75t_R g5862 ( 
.A(n_5738),
.Y(n_5862)
);

HB1xp67_ASAP7_75t_L g5863 ( 
.A(n_5752),
.Y(n_5863)
);

AND2x2_ASAP7_75t_L g5864 ( 
.A(n_5793),
.B(n_5634),
.Y(n_5864)
);

BUFx3_ASAP7_75t_L g5865 ( 
.A(n_5740),
.Y(n_5865)
);

INVx2_ASAP7_75t_L g5866 ( 
.A(n_5767),
.Y(n_5866)
);

OA21x2_ASAP7_75t_L g5867 ( 
.A1(n_5859),
.A2(n_5687),
.B(n_5626),
.Y(n_5867)
);

AND2x2_ASAP7_75t_L g5868 ( 
.A(n_5829),
.B(n_5483),
.Y(n_5868)
);

AO31x2_ASAP7_75t_L g5869 ( 
.A1(n_5833),
.A2(n_5630),
.A3(n_5660),
.B(n_5700),
.Y(n_5869)
);

HB1xp67_ASAP7_75t_L g5870 ( 
.A(n_5767),
.Y(n_5870)
);

INVx2_ASAP7_75t_L g5871 ( 
.A(n_5754),
.Y(n_5871)
);

OAI21x1_ASAP7_75t_L g5872 ( 
.A1(n_5762),
.A2(n_5706),
.B(n_5683),
.Y(n_5872)
);

BUFx2_ASAP7_75t_L g5873 ( 
.A(n_5732),
.Y(n_5873)
);

INVx2_ASAP7_75t_SL g5874 ( 
.A(n_5740),
.Y(n_5874)
);

AOI21xp5_ASAP7_75t_L g5875 ( 
.A1(n_5732),
.A2(n_5655),
.B(n_5676),
.Y(n_5875)
);

HB1xp67_ASAP7_75t_L g5876 ( 
.A(n_5731),
.Y(n_5876)
);

BUFx12f_ASAP7_75t_L g5877 ( 
.A(n_5750),
.Y(n_5877)
);

AO21x1_ASAP7_75t_SL g5878 ( 
.A1(n_5780),
.A2(n_5639),
.B(n_5692),
.Y(n_5878)
);

INVx1_ASAP7_75t_L g5879 ( 
.A(n_5735),
.Y(n_5879)
);

INVx1_ASAP7_75t_L g5880 ( 
.A(n_5739),
.Y(n_5880)
);

INVx2_ASAP7_75t_L g5881 ( 
.A(n_5746),
.Y(n_5881)
);

INVx1_ASAP7_75t_L g5882 ( 
.A(n_5755),
.Y(n_5882)
);

INVx1_ASAP7_75t_L g5883 ( 
.A(n_5756),
.Y(n_5883)
);

INVx1_ASAP7_75t_L g5884 ( 
.A(n_5759),
.Y(n_5884)
);

HB1xp67_ASAP7_75t_L g5885 ( 
.A(n_5733),
.Y(n_5885)
);

AND2x2_ASAP7_75t_L g5886 ( 
.A(n_5821),
.B(n_5483),
.Y(n_5886)
);

OR2x2_ASAP7_75t_SL g5887 ( 
.A(n_5762),
.B(n_5628),
.Y(n_5887)
);

NAND2xp5_ASAP7_75t_L g5888 ( 
.A(n_5799),
.B(n_5675),
.Y(n_5888)
);

NAND2xp5_ASAP7_75t_L g5889 ( 
.A(n_5790),
.B(n_5710),
.Y(n_5889)
);

INVx2_ASAP7_75t_L g5890 ( 
.A(n_5758),
.Y(n_5890)
);

HB1xp67_ASAP7_75t_L g5891 ( 
.A(n_5741),
.Y(n_5891)
);

HB1xp67_ASAP7_75t_L g5892 ( 
.A(n_5737),
.Y(n_5892)
);

INVx2_ASAP7_75t_L g5893 ( 
.A(n_5773),
.Y(n_5893)
);

INVx2_ASAP7_75t_SL g5894 ( 
.A(n_5736),
.Y(n_5894)
);

OAI21x1_ASAP7_75t_L g5895 ( 
.A1(n_5730),
.A2(n_5715),
.B(n_5315),
.Y(n_5895)
);

INVx2_ASAP7_75t_L g5896 ( 
.A(n_5810),
.Y(n_5896)
);

INVx1_ASAP7_75t_L g5897 ( 
.A(n_5761),
.Y(n_5897)
);

INVx1_ASAP7_75t_L g5898 ( 
.A(n_5765),
.Y(n_5898)
);

AOI21x1_ASAP7_75t_L g5899 ( 
.A1(n_5811),
.A2(n_4805),
.B(n_4801),
.Y(n_5899)
);

INVx2_ASAP7_75t_L g5900 ( 
.A(n_5835),
.Y(n_5900)
);

INVx2_ASAP7_75t_L g5901 ( 
.A(n_5845),
.Y(n_5901)
);

INVx2_ASAP7_75t_L g5902 ( 
.A(n_5847),
.Y(n_5902)
);

BUFx2_ASAP7_75t_SL g5903 ( 
.A(n_5771),
.Y(n_5903)
);

HB1xp67_ASAP7_75t_L g5904 ( 
.A(n_5785),
.Y(n_5904)
);

INVx8_ASAP7_75t_L g5905 ( 
.A(n_5750),
.Y(n_5905)
);

HB1xp67_ASAP7_75t_L g5906 ( 
.A(n_5729),
.Y(n_5906)
);

INVx2_ASAP7_75t_L g5907 ( 
.A(n_5792),
.Y(n_5907)
);

INVx5_ASAP7_75t_SL g5908 ( 
.A(n_5814),
.Y(n_5908)
);

INVx2_ASAP7_75t_SL g5909 ( 
.A(n_5742),
.Y(n_5909)
);

INVx1_ASAP7_75t_L g5910 ( 
.A(n_5734),
.Y(n_5910)
);

OAI21x1_ASAP7_75t_L g5911 ( 
.A1(n_5857),
.A2(n_4692),
.B(n_4664),
.Y(n_5911)
);

INVx1_ASAP7_75t_L g5912 ( 
.A(n_5776),
.Y(n_5912)
);

BUFx6f_ASAP7_75t_L g5913 ( 
.A(n_5794),
.Y(n_5913)
);

AO21x1_ASAP7_75t_L g5914 ( 
.A1(n_5807),
.A2(n_5027),
.B(n_5014),
.Y(n_5914)
);

INVx1_ASAP7_75t_L g5915 ( 
.A(n_5778),
.Y(n_5915)
);

BUFx3_ASAP7_75t_L g5916 ( 
.A(n_5804),
.Y(n_5916)
);

BUFx6f_ASAP7_75t_L g5917 ( 
.A(n_5747),
.Y(n_5917)
);

INVx1_ASAP7_75t_L g5918 ( 
.A(n_5775),
.Y(n_5918)
);

OAI21x1_ASAP7_75t_L g5919 ( 
.A1(n_5827),
.A2(n_5319),
.B(n_5258),
.Y(n_5919)
);

AOI21xp5_ASAP7_75t_L g5920 ( 
.A1(n_5802),
.A2(n_4808),
.B(n_4799),
.Y(n_5920)
);

INVx2_ASAP7_75t_L g5921 ( 
.A(n_5805),
.Y(n_5921)
);

INVx1_ASAP7_75t_L g5922 ( 
.A(n_5781),
.Y(n_5922)
);

INVx3_ASAP7_75t_L g5923 ( 
.A(n_5844),
.Y(n_5923)
);

BUFx6f_ASAP7_75t_L g5924 ( 
.A(n_5777),
.Y(n_5924)
);

INVx4_ASAP7_75t_L g5925 ( 
.A(n_5788),
.Y(n_5925)
);

INVx2_ASAP7_75t_L g5926 ( 
.A(n_5852),
.Y(n_5926)
);

AO31x2_ASAP7_75t_L g5927 ( 
.A1(n_5832),
.A2(n_4821),
.A3(n_4827),
.B(n_4823),
.Y(n_5927)
);

INVx1_ASAP7_75t_L g5928 ( 
.A(n_5796),
.Y(n_5928)
);

INVx2_ASAP7_75t_L g5929 ( 
.A(n_5764),
.Y(n_5929)
);

INVx2_ASAP7_75t_L g5930 ( 
.A(n_5823),
.Y(n_5930)
);

INVx3_ASAP7_75t_L g5931 ( 
.A(n_5779),
.Y(n_5931)
);

INVx1_ASAP7_75t_L g5932 ( 
.A(n_5774),
.Y(n_5932)
);

INVx1_ASAP7_75t_L g5933 ( 
.A(n_5836),
.Y(n_5933)
);

INVx1_ASAP7_75t_L g5934 ( 
.A(n_5841),
.Y(n_5934)
);

INVx1_ASAP7_75t_L g5935 ( 
.A(n_5843),
.Y(n_5935)
);

INVx1_ASAP7_75t_L g5936 ( 
.A(n_5800),
.Y(n_5936)
);

AND2x2_ASAP7_75t_L g5937 ( 
.A(n_5803),
.B(n_5838),
.Y(n_5937)
);

INVx2_ASAP7_75t_L g5938 ( 
.A(n_5824),
.Y(n_5938)
);

OAI21x1_ASAP7_75t_L g5939 ( 
.A1(n_5744),
.A2(n_5830),
.B(n_5813),
.Y(n_5939)
);

INVx2_ASAP7_75t_L g5940 ( 
.A(n_5743),
.Y(n_5940)
);

INVx2_ASAP7_75t_L g5941 ( 
.A(n_5854),
.Y(n_5941)
);

OAI321xp33_ASAP7_75t_L g5942 ( 
.A1(n_5818),
.A2(n_4943),
.A3(n_4807),
.B1(n_4954),
.B2(n_5013),
.C(n_4908),
.Y(n_5942)
);

INVx1_ASAP7_75t_SL g5943 ( 
.A(n_5798),
.Y(n_5943)
);

AND2x4_ASAP7_75t_L g5944 ( 
.A(n_5788),
.B(n_5268),
.Y(n_5944)
);

INVx2_ASAP7_75t_SL g5945 ( 
.A(n_5787),
.Y(n_5945)
);

INVx1_ASAP7_75t_L g5946 ( 
.A(n_5770),
.Y(n_5946)
);

AND2x4_ASAP7_75t_L g5947 ( 
.A(n_5856),
.B(n_5278),
.Y(n_5947)
);

INVx1_ASAP7_75t_L g5948 ( 
.A(n_5853),
.Y(n_5948)
);

INVx2_ASAP7_75t_L g5949 ( 
.A(n_5849),
.Y(n_5949)
);

INVx1_ASAP7_75t_L g5950 ( 
.A(n_5782),
.Y(n_5950)
);

AND2x2_ASAP7_75t_L g5951 ( 
.A(n_5786),
.B(n_5302),
.Y(n_5951)
);

INVx2_ASAP7_75t_L g5952 ( 
.A(n_5855),
.Y(n_5952)
);

AND2x2_ASAP7_75t_L g5953 ( 
.A(n_5831),
.B(n_5302),
.Y(n_5953)
);

OAI221xp5_ASAP7_75t_SL g5954 ( 
.A1(n_5815),
.A2(n_4898),
.B1(n_4773),
.B2(n_5022),
.C(n_5019),
.Y(n_5954)
);

AO31x2_ASAP7_75t_L g5955 ( 
.A1(n_5832),
.A2(n_4834),
.A3(n_4850),
.B(n_4837),
.Y(n_5955)
);

INVx1_ASAP7_75t_L g5956 ( 
.A(n_5791),
.Y(n_5956)
);

INVx1_ASAP7_75t_L g5957 ( 
.A(n_5858),
.Y(n_5957)
);

INVx2_ASAP7_75t_L g5958 ( 
.A(n_5760),
.Y(n_5958)
);

OR2x2_ASAP7_75t_L g5959 ( 
.A(n_5769),
.B(n_4987),
.Y(n_5959)
);

INVx1_ASAP7_75t_L g5960 ( 
.A(n_5766),
.Y(n_5960)
);

OAI21x1_ASAP7_75t_L g5961 ( 
.A1(n_5784),
.A2(n_5789),
.B(n_5839),
.Y(n_5961)
);

INVx2_ASAP7_75t_L g5962 ( 
.A(n_5760),
.Y(n_5962)
);

BUFx2_ASAP7_75t_SL g5963 ( 
.A(n_5814),
.Y(n_5963)
);

INVx1_ASAP7_75t_L g5964 ( 
.A(n_5840),
.Y(n_5964)
);

INVx1_ASAP7_75t_L g5965 ( 
.A(n_5816),
.Y(n_5965)
);

NAND2xp5_ASAP7_75t_L g5966 ( 
.A(n_5806),
.B(n_5848),
.Y(n_5966)
);

INVx1_ASAP7_75t_L g5967 ( 
.A(n_5850),
.Y(n_5967)
);

INVx2_ASAP7_75t_L g5968 ( 
.A(n_5826),
.Y(n_5968)
);

INVx1_ASAP7_75t_L g5969 ( 
.A(n_5806),
.Y(n_5969)
);

INVx2_ASAP7_75t_L g5970 ( 
.A(n_5837),
.Y(n_5970)
);

INVx1_ASAP7_75t_L g5971 ( 
.A(n_5768),
.Y(n_5971)
);

NAND2xp5_ASAP7_75t_L g5972 ( 
.A(n_5848),
.B(n_4910),
.Y(n_5972)
);

INVx2_ASAP7_75t_L g5973 ( 
.A(n_5795),
.Y(n_5973)
);

INVx1_ASAP7_75t_L g5974 ( 
.A(n_5763),
.Y(n_5974)
);

INVx1_ASAP7_75t_L g5975 ( 
.A(n_5851),
.Y(n_5975)
);

BUFx2_ASAP7_75t_L g5976 ( 
.A(n_5784),
.Y(n_5976)
);

OAI21x1_ASAP7_75t_L g5977 ( 
.A1(n_5745),
.A2(n_5783),
.B(n_5819),
.Y(n_5977)
);

INVx2_ASAP7_75t_L g5978 ( 
.A(n_5904),
.Y(n_5978)
);

INVx1_ASAP7_75t_L g5979 ( 
.A(n_5863),
.Y(n_5979)
);

INVx2_ASAP7_75t_L g5980 ( 
.A(n_5873),
.Y(n_5980)
);

AO21x2_ASAP7_75t_L g5981 ( 
.A1(n_5875),
.A2(n_5842),
.B(n_5825),
.Y(n_5981)
);

AO21x2_ASAP7_75t_L g5982 ( 
.A1(n_5957),
.A2(n_5964),
.B(n_5970),
.Y(n_5982)
);

INVx1_ASAP7_75t_L g5983 ( 
.A(n_5873),
.Y(n_5983)
);

BUFx6f_ASAP7_75t_L g5984 ( 
.A(n_5877),
.Y(n_5984)
);

INVx2_ASAP7_75t_L g5985 ( 
.A(n_5871),
.Y(n_5985)
);

OAI21xp33_ASAP7_75t_L g5986 ( 
.A1(n_5888),
.A2(n_5971),
.B(n_5895),
.Y(n_5986)
);

INVx2_ASAP7_75t_SL g5987 ( 
.A(n_5905),
.Y(n_5987)
);

NAND2xp5_ASAP7_75t_L g5988 ( 
.A(n_5889),
.B(n_5812),
.Y(n_5988)
);

INVx2_ASAP7_75t_L g5989 ( 
.A(n_5866),
.Y(n_5989)
);

BUFx6f_ASAP7_75t_L g5990 ( 
.A(n_5861),
.Y(n_5990)
);

INVx2_ASAP7_75t_L g5991 ( 
.A(n_5900),
.Y(n_5991)
);

INVx1_ASAP7_75t_L g5992 ( 
.A(n_5918),
.Y(n_5992)
);

INVx2_ASAP7_75t_L g5993 ( 
.A(n_5901),
.Y(n_5993)
);

BUFx6f_ASAP7_75t_L g5994 ( 
.A(n_5865),
.Y(n_5994)
);

NOR2xp33_ASAP7_75t_L g5995 ( 
.A(n_5874),
.B(n_5753),
.Y(n_5995)
);

OR2x2_ASAP7_75t_L g5996 ( 
.A(n_5972),
.B(n_5757),
.Y(n_5996)
);

INVx2_ASAP7_75t_L g5997 ( 
.A(n_5902),
.Y(n_5997)
);

INVx1_ASAP7_75t_L g5998 ( 
.A(n_5906),
.Y(n_5998)
);

INVx4_ASAP7_75t_L g5999 ( 
.A(n_5905),
.Y(n_5999)
);

HB1xp67_ASAP7_75t_L g6000 ( 
.A(n_5870),
.Y(n_6000)
);

INVx2_ASAP7_75t_L g6001 ( 
.A(n_5881),
.Y(n_6001)
);

AOI22xp33_ASAP7_75t_SL g6002 ( 
.A1(n_5903),
.A2(n_5817),
.B1(n_5809),
.B2(n_5801),
.Y(n_6002)
);

INVxp67_ASAP7_75t_SL g6003 ( 
.A(n_5872),
.Y(n_6003)
);

OR2x2_ASAP7_75t_L g6004 ( 
.A(n_5922),
.B(n_5928),
.Y(n_6004)
);

INVx2_ASAP7_75t_L g6005 ( 
.A(n_5890),
.Y(n_6005)
);

NOR2xp67_ASAP7_75t_SL g6006 ( 
.A(n_5903),
.B(n_4872),
.Y(n_6006)
);

INVx1_ASAP7_75t_L g6007 ( 
.A(n_5950),
.Y(n_6007)
);

NAND2x1p5_ASAP7_75t_L g6008 ( 
.A(n_5923),
.B(n_5825),
.Y(n_6008)
);

AND2x2_ASAP7_75t_L g6009 ( 
.A(n_5937),
.B(n_5749),
.Y(n_6009)
);

INVx1_ASAP7_75t_L g6010 ( 
.A(n_5956),
.Y(n_6010)
);

HB1xp67_ASAP7_75t_L g6011 ( 
.A(n_5891),
.Y(n_6011)
);

INVx2_ASAP7_75t_SL g6012 ( 
.A(n_5916),
.Y(n_6012)
);

BUFx2_ASAP7_75t_SL g6013 ( 
.A(n_5925),
.Y(n_6013)
);

HB1xp67_ASAP7_75t_L g6014 ( 
.A(n_5892),
.Y(n_6014)
);

INVx1_ASAP7_75t_L g6015 ( 
.A(n_5965),
.Y(n_6015)
);

INVx2_ASAP7_75t_L g6016 ( 
.A(n_5893),
.Y(n_6016)
);

NAND2xp5_ASAP7_75t_L g6017 ( 
.A(n_5869),
.B(n_5834),
.Y(n_6017)
);

OA21x2_ASAP7_75t_L g6018 ( 
.A1(n_5976),
.A2(n_5846),
.B(n_5820),
.Y(n_6018)
);

AND2x2_ASAP7_75t_L g6019 ( 
.A(n_5977),
.B(n_5797),
.Y(n_6019)
);

INVx2_ASAP7_75t_L g6020 ( 
.A(n_5929),
.Y(n_6020)
);

NAND2xp5_ASAP7_75t_L g6021 ( 
.A(n_5869),
.B(n_5822),
.Y(n_6021)
);

BUFx3_ASAP7_75t_L g6022 ( 
.A(n_5917),
.Y(n_6022)
);

INVx3_ASAP7_75t_L g6023 ( 
.A(n_5924),
.Y(n_6023)
);

AND2x2_ASAP7_75t_L g6024 ( 
.A(n_5975),
.B(n_5828),
.Y(n_6024)
);

INVx2_ASAP7_75t_L g6025 ( 
.A(n_5941),
.Y(n_6025)
);

OAI211xp5_ASAP7_75t_SL g6026 ( 
.A1(n_5920),
.A2(n_5025),
.B(n_5269),
.C(n_5046),
.Y(n_6026)
);

NAND2x1p5_ASAP7_75t_L g6027 ( 
.A(n_5917),
.B(n_5751),
.Y(n_6027)
);

AND2x4_ASAP7_75t_L g6028 ( 
.A(n_5909),
.B(n_5330),
.Y(n_6028)
);

OR2x6_ASAP7_75t_L g6029 ( 
.A(n_5963),
.B(n_5031),
.Y(n_6029)
);

OR2x6_ASAP7_75t_L g6030 ( 
.A(n_5963),
.B(n_5041),
.Y(n_6030)
);

INVx1_ASAP7_75t_L g6031 ( 
.A(n_5932),
.Y(n_6031)
);

INVx1_ASAP7_75t_L g6032 ( 
.A(n_5879),
.Y(n_6032)
);

INVx2_ASAP7_75t_L g6033 ( 
.A(n_5921),
.Y(n_6033)
);

BUFx3_ASAP7_75t_L g6034 ( 
.A(n_5913),
.Y(n_6034)
);

INVx1_ASAP7_75t_L g6035 ( 
.A(n_5880),
.Y(n_6035)
);

INVx1_ASAP7_75t_L g6036 ( 
.A(n_5882),
.Y(n_6036)
);

INVx2_ASAP7_75t_L g6037 ( 
.A(n_5896),
.Y(n_6037)
);

INVx2_ASAP7_75t_L g6038 ( 
.A(n_5907),
.Y(n_6038)
);

AND2x2_ASAP7_75t_L g6039 ( 
.A(n_5945),
.B(n_5808),
.Y(n_6039)
);

INVx1_ASAP7_75t_L g6040 ( 
.A(n_5883),
.Y(n_6040)
);

INVx1_ASAP7_75t_L g6041 ( 
.A(n_5884),
.Y(n_6041)
);

AO21x2_ASAP7_75t_L g6042 ( 
.A1(n_5974),
.A2(n_4924),
.B(n_4922),
.Y(n_6042)
);

AO21x2_ASAP7_75t_L g6043 ( 
.A1(n_5967),
.A2(n_4937),
.B(n_4929),
.Y(n_6043)
);

INVx2_ASAP7_75t_SL g6044 ( 
.A(n_5924),
.Y(n_6044)
);

OAI21x1_ASAP7_75t_L g6045 ( 
.A1(n_5939),
.A2(n_5352),
.B(n_5351),
.Y(n_6045)
);

INVxp67_ASAP7_75t_L g6046 ( 
.A(n_5878),
.Y(n_6046)
);

INVx1_ASAP7_75t_L g6047 ( 
.A(n_5897),
.Y(n_6047)
);

OAI21x1_ASAP7_75t_L g6048 ( 
.A1(n_5961),
.A2(n_5337),
.B(n_5393),
.Y(n_6048)
);

INVx2_ASAP7_75t_L g6049 ( 
.A(n_5930),
.Y(n_6049)
);

INVx3_ASAP7_75t_L g6050 ( 
.A(n_5913),
.Y(n_6050)
);

INVx2_ASAP7_75t_L g6051 ( 
.A(n_5938),
.Y(n_6051)
);

NAND2xp5_ASAP7_75t_L g6052 ( 
.A(n_5869),
.B(n_4990),
.Y(n_6052)
);

INVx2_ASAP7_75t_L g6053 ( 
.A(n_5952),
.Y(n_6053)
);

INVx2_ASAP7_75t_L g6054 ( 
.A(n_5876),
.Y(n_6054)
);

INVx1_ASAP7_75t_L g6055 ( 
.A(n_5898),
.Y(n_6055)
);

INVx1_ASAP7_75t_L g6056 ( 
.A(n_5910),
.Y(n_6056)
);

INVx2_ASAP7_75t_L g6057 ( 
.A(n_5885),
.Y(n_6057)
);

AO21x2_ASAP7_75t_L g6058 ( 
.A1(n_5960),
.A2(n_5008),
.B(n_5005),
.Y(n_6058)
);

INVx1_ASAP7_75t_L g6059 ( 
.A(n_5936),
.Y(n_6059)
);

INVx2_ASAP7_75t_L g6060 ( 
.A(n_5926),
.Y(n_6060)
);

INVx2_ASAP7_75t_SL g6061 ( 
.A(n_5943),
.Y(n_6061)
);

OR2x6_ASAP7_75t_L g6062 ( 
.A(n_5894),
.B(n_5045),
.Y(n_6062)
);

INVx2_ASAP7_75t_L g6063 ( 
.A(n_5940),
.Y(n_6063)
);

OR2x6_ASAP7_75t_L g6064 ( 
.A(n_5944),
.B(n_4965),
.Y(n_6064)
);

INVx1_ASAP7_75t_L g6065 ( 
.A(n_5912),
.Y(n_6065)
);

INVx2_ASAP7_75t_L g6066 ( 
.A(n_5949),
.Y(n_6066)
);

OR2x6_ASAP7_75t_L g6067 ( 
.A(n_5944),
.B(n_5976),
.Y(n_6067)
);

INVx2_ASAP7_75t_L g6068 ( 
.A(n_5946),
.Y(n_6068)
);

NOR2xp33_ASAP7_75t_L g6069 ( 
.A(n_5862),
.B(n_5009),
.Y(n_6069)
);

INVx1_ASAP7_75t_L g6070 ( 
.A(n_5915),
.Y(n_6070)
);

INVx3_ASAP7_75t_L g6071 ( 
.A(n_5908),
.Y(n_6071)
);

NAND2xp5_ASAP7_75t_L g6072 ( 
.A(n_5927),
.B(n_4962),
.Y(n_6072)
);

INVx1_ASAP7_75t_L g6073 ( 
.A(n_5948),
.Y(n_6073)
);

HB1xp67_ASAP7_75t_L g6074 ( 
.A(n_5969),
.Y(n_6074)
);

INVx4_ASAP7_75t_L g6075 ( 
.A(n_5931),
.Y(n_6075)
);

INVx3_ASAP7_75t_L g6076 ( 
.A(n_5908),
.Y(n_6076)
);

HB1xp67_ASAP7_75t_L g6077 ( 
.A(n_5934),
.Y(n_6077)
);

HB1xp67_ASAP7_75t_L g6078 ( 
.A(n_5935),
.Y(n_6078)
);

BUFx2_ASAP7_75t_L g6079 ( 
.A(n_5860),
.Y(n_6079)
);

INVx1_ASAP7_75t_L g6080 ( 
.A(n_5959),
.Y(n_6080)
);

BUFx4f_ASAP7_75t_L g6081 ( 
.A(n_5867),
.Y(n_6081)
);

INVx1_ASAP7_75t_L g6082 ( 
.A(n_5953),
.Y(n_6082)
);

AND2x2_ASAP7_75t_L g6083 ( 
.A(n_5951),
.B(n_5064),
.Y(n_6083)
);

INVx2_ASAP7_75t_L g6084 ( 
.A(n_5933),
.Y(n_6084)
);

AO21x2_ASAP7_75t_L g6085 ( 
.A1(n_5966),
.A2(n_4968),
.B(n_4963),
.Y(n_6085)
);

BUFx2_ASAP7_75t_L g6086 ( 
.A(n_5860),
.Y(n_6086)
);

BUFx2_ASAP7_75t_L g6087 ( 
.A(n_5887),
.Y(n_6087)
);

HB1xp67_ASAP7_75t_L g6088 ( 
.A(n_5867),
.Y(n_6088)
);

INVx1_ASAP7_75t_L g6089 ( 
.A(n_5947),
.Y(n_6089)
);

HB1xp67_ASAP7_75t_L g6090 ( 
.A(n_5864),
.Y(n_6090)
);

INVx1_ASAP7_75t_L g6091 ( 
.A(n_5947),
.Y(n_6091)
);

NAND2xp5_ASAP7_75t_L g6092 ( 
.A(n_5927),
.B(n_5955),
.Y(n_6092)
);

HB1xp67_ASAP7_75t_L g6093 ( 
.A(n_5927),
.Y(n_6093)
);

INVx4_ASAP7_75t_SL g6094 ( 
.A(n_5886),
.Y(n_6094)
);

INVx1_ASAP7_75t_L g6095 ( 
.A(n_5955),
.Y(n_6095)
);

BUFx3_ASAP7_75t_L g6096 ( 
.A(n_5868),
.Y(n_6096)
);

INVx2_ASAP7_75t_L g6097 ( 
.A(n_5973),
.Y(n_6097)
);

INVx3_ASAP7_75t_L g6098 ( 
.A(n_5958),
.Y(n_6098)
);

AO21x2_ASAP7_75t_L g6099 ( 
.A1(n_5899),
.A2(n_4969),
.B(n_4844),
.Y(n_6099)
);

AND2x2_ASAP7_75t_L g6100 ( 
.A(n_5962),
.B(n_5311),
.Y(n_6100)
);

INVx2_ASAP7_75t_SL g6101 ( 
.A(n_5968),
.Y(n_6101)
);

OR2x2_ASAP7_75t_L g6102 ( 
.A(n_5955),
.B(n_11),
.Y(n_6102)
);

INVx2_ASAP7_75t_L g6103 ( 
.A(n_5919),
.Y(n_6103)
);

INVx2_ASAP7_75t_SL g6104 ( 
.A(n_5911),
.Y(n_6104)
);

OAI21xp5_ASAP7_75t_L g6105 ( 
.A1(n_5899),
.A2(n_5220),
.B(n_5253),
.Y(n_6105)
);

OR2x2_ASAP7_75t_L g6106 ( 
.A(n_5914),
.B(n_12),
.Y(n_6106)
);

HB1xp67_ASAP7_75t_L g6107 ( 
.A(n_5954),
.Y(n_6107)
);

INVx1_ASAP7_75t_L g6108 ( 
.A(n_5942),
.Y(n_6108)
);

INVx1_ASAP7_75t_L g6109 ( 
.A(n_5878),
.Y(n_6109)
);

AND2x2_ASAP7_75t_L g6110 ( 
.A(n_5873),
.B(n_5371),
.Y(n_6110)
);

INVx2_ASAP7_75t_L g6111 ( 
.A(n_5904),
.Y(n_6111)
);

NOR2xp33_ASAP7_75t_L g6112 ( 
.A(n_5865),
.B(n_506),
.Y(n_6112)
);

NAND2xp5_ASAP7_75t_L g6113 ( 
.A(n_5888),
.B(n_4706),
.Y(n_6113)
);

INVx2_ASAP7_75t_L g6114 ( 
.A(n_5904),
.Y(n_6114)
);

AND2x2_ASAP7_75t_L g6115 ( 
.A(n_5873),
.B(n_5381),
.Y(n_6115)
);

HB1xp67_ASAP7_75t_L g6116 ( 
.A(n_5863),
.Y(n_6116)
);

INVx2_ASAP7_75t_L g6117 ( 
.A(n_5904),
.Y(n_6117)
);

AND2x4_ASAP7_75t_L g6118 ( 
.A(n_5873),
.B(n_4701),
.Y(n_6118)
);

INVx1_ASAP7_75t_L g6119 ( 
.A(n_5863),
.Y(n_6119)
);

BUFx3_ASAP7_75t_L g6120 ( 
.A(n_5877),
.Y(n_6120)
);

HB1xp67_ASAP7_75t_L g6121 ( 
.A(n_5863),
.Y(n_6121)
);

INVx1_ASAP7_75t_L g6122 ( 
.A(n_5863),
.Y(n_6122)
);

INVx1_ASAP7_75t_L g6123 ( 
.A(n_5863),
.Y(n_6123)
);

HB1xp67_ASAP7_75t_L g6124 ( 
.A(n_5863),
.Y(n_6124)
);

OA21x2_ASAP7_75t_L g6125 ( 
.A1(n_5875),
.A2(n_4859),
.B(n_4831),
.Y(n_6125)
);

INVx1_ASAP7_75t_L g6126 ( 
.A(n_5863),
.Y(n_6126)
);

OA21x2_ASAP7_75t_L g6127 ( 
.A1(n_5875),
.A2(n_4722),
.B(n_4709),
.Y(n_6127)
);

INVx4_ASAP7_75t_L g6128 ( 
.A(n_5877),
.Y(n_6128)
);

INVx1_ASAP7_75t_L g6129 ( 
.A(n_5863),
.Y(n_6129)
);

AND2x2_ASAP7_75t_L g6130 ( 
.A(n_5873),
.B(n_4800),
.Y(n_6130)
);

OA21x2_ASAP7_75t_L g6131 ( 
.A1(n_5875),
.A2(n_4787),
.B(n_4978),
.Y(n_6131)
);

INVx1_ASAP7_75t_L g6132 ( 
.A(n_5863),
.Y(n_6132)
);

AO21x2_ASAP7_75t_L g6133 ( 
.A1(n_5875),
.A2(n_5030),
.B(n_4972),
.Y(n_6133)
);

BUFx2_ASAP7_75t_SL g6134 ( 
.A(n_5865),
.Y(n_6134)
);

INVx4_ASAP7_75t_L g6135 ( 
.A(n_5984),
.Y(n_6135)
);

NAND2xp33_ASAP7_75t_R g6136 ( 
.A(n_6109),
.B(n_6019),
.Y(n_6136)
);

INVx4_ASAP7_75t_L g6137 ( 
.A(n_5984),
.Y(n_6137)
);

INVx1_ASAP7_75t_L g6138 ( 
.A(n_6116),
.Y(n_6138)
);

AOI31xp33_ASAP7_75t_L g6139 ( 
.A1(n_6046),
.A2(n_4927),
.A3(n_5004),
.B(n_4956),
.Y(n_6139)
);

INVx2_ASAP7_75t_L g6140 ( 
.A(n_5980),
.Y(n_6140)
);

AND2x2_ASAP7_75t_L g6141 ( 
.A(n_6009),
.B(n_12),
.Y(n_6141)
);

INVx2_ASAP7_75t_L g6142 ( 
.A(n_6012),
.Y(n_6142)
);

AND2x2_ASAP7_75t_L g6143 ( 
.A(n_6134),
.B(n_12),
.Y(n_6143)
);

HB1xp67_ASAP7_75t_L g6144 ( 
.A(n_6121),
.Y(n_6144)
);

OR2x2_ASAP7_75t_L g6145 ( 
.A(n_5979),
.B(n_13),
.Y(n_6145)
);

HB1xp67_ASAP7_75t_L g6146 ( 
.A(n_6124),
.Y(n_6146)
);

INVx1_ASAP7_75t_L g6147 ( 
.A(n_6074),
.Y(n_6147)
);

CKINVDCx20_ASAP7_75t_R g6148 ( 
.A(n_5990),
.Y(n_6148)
);

AND2x4_ASAP7_75t_L g6149 ( 
.A(n_6039),
.B(n_4740),
.Y(n_6149)
);

HB1xp67_ASAP7_75t_L g6150 ( 
.A(n_6011),
.Y(n_6150)
);

AND2x2_ASAP7_75t_L g6151 ( 
.A(n_6134),
.B(n_13),
.Y(n_6151)
);

INVx2_ASAP7_75t_L g6152 ( 
.A(n_6014),
.Y(n_6152)
);

INVx3_ASAP7_75t_L g6153 ( 
.A(n_5994),
.Y(n_6153)
);

AND2x2_ASAP7_75t_L g6154 ( 
.A(n_5995),
.B(n_13),
.Y(n_6154)
);

AO31x2_ASAP7_75t_L g6155 ( 
.A1(n_6087),
.A2(n_4784),
.A3(n_5011),
.B(n_5010),
.Y(n_6155)
);

AND2x2_ASAP7_75t_L g6156 ( 
.A(n_6075),
.B(n_13),
.Y(n_6156)
);

AND2x4_ASAP7_75t_L g6157 ( 
.A(n_6094),
.B(n_4744),
.Y(n_6157)
);

INVx2_ASAP7_75t_L g6158 ( 
.A(n_6054),
.Y(n_6158)
);

HB1xp67_ASAP7_75t_L g6159 ( 
.A(n_6000),
.Y(n_6159)
);

INVx1_ASAP7_75t_L g6160 ( 
.A(n_5983),
.Y(n_6160)
);

AND2x2_ASAP7_75t_L g6161 ( 
.A(n_6023),
.B(n_14),
.Y(n_6161)
);

INVxp67_ASAP7_75t_L g6162 ( 
.A(n_6061),
.Y(n_6162)
);

AND2x2_ASAP7_75t_L g6163 ( 
.A(n_6094),
.B(n_14),
.Y(n_6163)
);

AND2x2_ASAP7_75t_L g6164 ( 
.A(n_6013),
.B(n_14),
.Y(n_6164)
);

AND2x4_ASAP7_75t_L g6165 ( 
.A(n_6022),
.B(n_5012),
.Y(n_6165)
);

INVx1_ASAP7_75t_L g6166 ( 
.A(n_6119),
.Y(n_6166)
);

AND2x2_ASAP7_75t_L g6167 ( 
.A(n_6013),
.B(n_14),
.Y(n_6167)
);

INVx2_ASAP7_75t_SL g6168 ( 
.A(n_5994),
.Y(n_6168)
);

AND2x2_ASAP7_75t_L g6169 ( 
.A(n_6027),
.B(n_15),
.Y(n_6169)
);

OR2x2_ASAP7_75t_L g6170 ( 
.A(n_6122),
.B(n_15),
.Y(n_6170)
);

BUFx2_ASAP7_75t_L g6171 ( 
.A(n_6071),
.Y(n_6171)
);

AND2x2_ASAP7_75t_L g6172 ( 
.A(n_6044),
.B(n_15),
.Y(n_6172)
);

OR2x2_ASAP7_75t_L g6173 ( 
.A(n_6123),
.B(n_15),
.Y(n_6173)
);

INVx2_ASAP7_75t_L g6174 ( 
.A(n_6057),
.Y(n_6174)
);

AND2x4_ASAP7_75t_SL g6175 ( 
.A(n_6128),
.B(n_16),
.Y(n_6175)
);

AND2x2_ASAP7_75t_L g6176 ( 
.A(n_6024),
.B(n_16),
.Y(n_6176)
);

AND2x2_ASAP7_75t_L g6177 ( 
.A(n_6050),
.B(n_16),
.Y(n_6177)
);

AND2x2_ASAP7_75t_L g6178 ( 
.A(n_6096),
.B(n_16),
.Y(n_6178)
);

INVx1_ASAP7_75t_L g6179 ( 
.A(n_6126),
.Y(n_6179)
);

INVx2_ASAP7_75t_L g6180 ( 
.A(n_5978),
.Y(n_6180)
);

AND2x2_ASAP7_75t_L g6181 ( 
.A(n_6130),
.B(n_17),
.Y(n_6181)
);

AND2x2_ASAP7_75t_L g6182 ( 
.A(n_6067),
.B(n_17),
.Y(n_6182)
);

INVx1_ASAP7_75t_L g6183 ( 
.A(n_6129),
.Y(n_6183)
);

HB1xp67_ASAP7_75t_L g6184 ( 
.A(n_6132),
.Y(n_6184)
);

HB1xp67_ASAP7_75t_L g6185 ( 
.A(n_6111),
.Y(n_6185)
);

AND2x2_ASAP7_75t_L g6186 ( 
.A(n_6067),
.B(n_18),
.Y(n_6186)
);

NAND2xp5_ASAP7_75t_L g6187 ( 
.A(n_6108),
.B(n_4911),
.Y(n_6187)
);

AND2x2_ASAP7_75t_L g6188 ( 
.A(n_6101),
.B(n_6076),
.Y(n_6188)
);

BUFx2_ASAP7_75t_L g6189 ( 
.A(n_5999),
.Y(n_6189)
);

NAND2xp5_ASAP7_75t_L g6190 ( 
.A(n_6021),
.B(n_6085),
.Y(n_6190)
);

HB1xp67_ASAP7_75t_L g6191 ( 
.A(n_6114),
.Y(n_6191)
);

BUFx2_ASAP7_75t_L g6192 ( 
.A(n_6008),
.Y(n_6192)
);

OAI211xp5_ASAP7_75t_SL g6193 ( 
.A1(n_6109),
.A2(n_4980),
.B(n_4930),
.C(n_4942),
.Y(n_6193)
);

AND2x2_ASAP7_75t_L g6194 ( 
.A(n_6089),
.B(n_18),
.Y(n_6194)
);

BUFx3_ASAP7_75t_L g6195 ( 
.A(n_5990),
.Y(n_6195)
);

HB1xp67_ASAP7_75t_L g6196 ( 
.A(n_6117),
.Y(n_6196)
);

AND2x2_ASAP7_75t_L g6197 ( 
.A(n_6091),
.B(n_18),
.Y(n_6197)
);

INVx4_ASAP7_75t_L g6198 ( 
.A(n_6120),
.Y(n_6198)
);

NOR2x1_ASAP7_75t_L g6199 ( 
.A(n_6106),
.B(n_4952),
.Y(n_6199)
);

INVx1_ASAP7_75t_L g6200 ( 
.A(n_5998),
.Y(n_6200)
);

INVx1_ASAP7_75t_L g6201 ( 
.A(n_6004),
.Y(n_6201)
);

INVx1_ASAP7_75t_L g6202 ( 
.A(n_6080),
.Y(n_6202)
);

AND2x2_ASAP7_75t_L g6203 ( 
.A(n_6064),
.B(n_18),
.Y(n_6203)
);

AOI22xp33_ASAP7_75t_L g6204 ( 
.A1(n_6107),
.A2(n_4946),
.B1(n_4949),
.B2(n_4914),
.Y(n_6204)
);

AO21x2_ASAP7_75t_L g6205 ( 
.A1(n_6017),
.A2(n_5061),
.B(n_5060),
.Y(n_6205)
);

INVx1_ASAP7_75t_L g6206 ( 
.A(n_6056),
.Y(n_6206)
);

OR2x2_ASAP7_75t_L g6207 ( 
.A(n_5985),
.B(n_19),
.Y(n_6207)
);

INVx1_ASAP7_75t_L g6208 ( 
.A(n_6056),
.Y(n_6208)
);

INVx2_ASAP7_75t_L g6209 ( 
.A(n_6028),
.Y(n_6209)
);

INVx1_ASAP7_75t_L g6210 ( 
.A(n_5992),
.Y(n_6210)
);

AND2x4_ASAP7_75t_L g6211 ( 
.A(n_5987),
.B(n_5065),
.Y(n_6211)
);

INVx1_ASAP7_75t_L g6212 ( 
.A(n_5992),
.Y(n_6212)
);

INVx2_ASAP7_75t_L g6213 ( 
.A(n_6028),
.Y(n_6213)
);

AND2x2_ASAP7_75t_L g6214 ( 
.A(n_6064),
.B(n_19),
.Y(n_6214)
);

NOR2xp67_ASAP7_75t_L g6215 ( 
.A(n_6088),
.B(n_19),
.Y(n_6215)
);

INVx1_ASAP7_75t_L g6216 ( 
.A(n_6077),
.Y(n_6216)
);

AND2x2_ASAP7_75t_L g6217 ( 
.A(n_6002),
.B(n_19),
.Y(n_6217)
);

INVx1_ASAP7_75t_L g6218 ( 
.A(n_6078),
.Y(n_6218)
);

AND2x2_ASAP7_75t_L g6219 ( 
.A(n_6082),
.B(n_20),
.Y(n_6219)
);

NAND2xp5_ASAP7_75t_L g6220 ( 
.A(n_6110),
.B(n_5069),
.Y(n_6220)
);

INVx2_ASAP7_75t_L g6221 ( 
.A(n_6053),
.Y(n_6221)
);

NAND2xp5_ASAP7_75t_L g6222 ( 
.A(n_6115),
.B(n_20),
.Y(n_6222)
);

INVx1_ASAP7_75t_L g6223 ( 
.A(n_6068),
.Y(n_6223)
);

BUFx3_ASAP7_75t_L g6224 ( 
.A(n_6034),
.Y(n_6224)
);

AND2x2_ASAP7_75t_L g6225 ( 
.A(n_6090),
.B(n_20),
.Y(n_6225)
);

AND2x2_ASAP7_75t_L g6226 ( 
.A(n_6020),
.B(n_6098),
.Y(n_6226)
);

AOI22xp33_ASAP7_75t_L g6227 ( 
.A1(n_5988),
.A2(n_6081),
.B1(n_5986),
.B2(n_5996),
.Y(n_6227)
);

AND2x2_ASAP7_75t_L g6228 ( 
.A(n_6083),
.B(n_21),
.Y(n_6228)
);

BUFx3_ASAP7_75t_L g6229 ( 
.A(n_6112),
.Y(n_6229)
);

AND2x2_ASAP7_75t_L g6230 ( 
.A(n_6063),
.B(n_21),
.Y(n_6230)
);

AO21x2_ASAP7_75t_L g6231 ( 
.A1(n_6003),
.A2(n_21),
.B(n_22),
.Y(n_6231)
);

NOR2xp33_ASAP7_75t_L g6232 ( 
.A(n_6113),
.B(n_22),
.Y(n_6232)
);

INVx2_ASAP7_75t_L g6233 ( 
.A(n_6100),
.Y(n_6233)
);

INVx1_ASAP7_75t_L g6234 ( 
.A(n_6007),
.Y(n_6234)
);

HB1xp67_ASAP7_75t_L g6235 ( 
.A(n_5989),
.Y(n_6235)
);

INVx2_ASAP7_75t_L g6236 ( 
.A(n_6084),
.Y(n_6236)
);

AND2x4_ASAP7_75t_L g6237 ( 
.A(n_6118),
.B(n_507),
.Y(n_6237)
);

NAND2xp5_ASAP7_75t_L g6238 ( 
.A(n_6043),
.B(n_22),
.Y(n_6238)
);

INVx2_ASAP7_75t_L g6239 ( 
.A(n_6066),
.Y(n_6239)
);

NAND2xp5_ASAP7_75t_L g6240 ( 
.A(n_6042),
.B(n_22),
.Y(n_6240)
);

INVx2_ASAP7_75t_L g6241 ( 
.A(n_6033),
.Y(n_6241)
);

AND2x2_ASAP7_75t_L g6242 ( 
.A(n_6118),
.B(n_23),
.Y(n_6242)
);

BUFx6f_ASAP7_75t_L g6243 ( 
.A(n_6048),
.Y(n_6243)
);

AND2x2_ASAP7_75t_L g6244 ( 
.A(n_6062),
.B(n_23),
.Y(n_6244)
);

BUFx3_ASAP7_75t_L g6245 ( 
.A(n_6069),
.Y(n_6245)
);

INVxp67_ASAP7_75t_SL g6246 ( 
.A(n_6006),
.Y(n_6246)
);

AOI22xp33_ASAP7_75t_L g6247 ( 
.A1(n_6087),
.A2(n_508),
.B1(n_509),
.B2(n_507),
.Y(n_6247)
);

INVx2_ASAP7_75t_L g6248 ( 
.A(n_5991),
.Y(n_6248)
);

HB1xp67_ASAP7_75t_L g6249 ( 
.A(n_6010),
.Y(n_6249)
);

AND2x2_ASAP7_75t_L g6250 ( 
.A(n_6062),
.B(n_23),
.Y(n_6250)
);

AND2x2_ASAP7_75t_L g6251 ( 
.A(n_6097),
.B(n_24),
.Y(n_6251)
);

AND2x2_ASAP7_75t_L g6252 ( 
.A(n_6104),
.B(n_24),
.Y(n_6252)
);

AOI22xp33_ASAP7_75t_L g6253 ( 
.A1(n_6006),
.A2(n_508),
.B1(n_509),
.B2(n_507),
.Y(n_6253)
);

AND2x2_ASAP7_75t_L g6254 ( 
.A(n_6029),
.B(n_24),
.Y(n_6254)
);

INVx1_ASAP7_75t_L g6255 ( 
.A(n_6015),
.Y(n_6255)
);

INVx1_ASAP7_75t_L g6256 ( 
.A(n_6059),
.Y(n_6256)
);

AND2x2_ASAP7_75t_L g6257 ( 
.A(n_6029),
.B(n_25),
.Y(n_6257)
);

AND2x2_ASAP7_75t_L g6258 ( 
.A(n_6030),
.B(n_25),
.Y(n_6258)
);

INVx1_ASAP7_75t_L g6259 ( 
.A(n_6031),
.Y(n_6259)
);

NAND2xp5_ASAP7_75t_L g6260 ( 
.A(n_6052),
.B(n_25),
.Y(n_6260)
);

AND2x2_ASAP7_75t_L g6261 ( 
.A(n_6030),
.B(n_25),
.Y(n_6261)
);

INVx1_ASAP7_75t_L g6262 ( 
.A(n_6032),
.Y(n_6262)
);

INVx1_ASAP7_75t_L g6263 ( 
.A(n_6035),
.Y(n_6263)
);

INVx2_ASAP7_75t_L g6264 ( 
.A(n_5993),
.Y(n_6264)
);

INVx1_ASAP7_75t_L g6265 ( 
.A(n_6036),
.Y(n_6265)
);

AND2x2_ASAP7_75t_L g6266 ( 
.A(n_5981),
.B(n_26),
.Y(n_6266)
);

AND2x2_ASAP7_75t_L g6267 ( 
.A(n_6103),
.B(n_26),
.Y(n_6267)
);

NAND2xp5_ASAP7_75t_L g6268 ( 
.A(n_6058),
.B(n_6072),
.Y(n_6268)
);

INVx2_ASAP7_75t_L g6269 ( 
.A(n_5997),
.Y(n_6269)
);

OR2x2_ASAP7_75t_L g6270 ( 
.A(n_6102),
.B(n_6065),
.Y(n_6270)
);

BUFx3_ASAP7_75t_L g6271 ( 
.A(n_6001),
.Y(n_6271)
);

AND2x2_ASAP7_75t_L g6272 ( 
.A(n_6018),
.B(n_26),
.Y(n_6272)
);

AND2x2_ASAP7_75t_L g6273 ( 
.A(n_6018),
.B(n_26),
.Y(n_6273)
);

INVx1_ASAP7_75t_L g6274 ( 
.A(n_6040),
.Y(n_6274)
);

INVx1_ASAP7_75t_L g6275 ( 
.A(n_6041),
.Y(n_6275)
);

AND2x2_ASAP7_75t_L g6276 ( 
.A(n_6005),
.B(n_27),
.Y(n_6276)
);

HB1xp67_ASAP7_75t_L g6277 ( 
.A(n_6047),
.Y(n_6277)
);

NAND2xp5_ASAP7_75t_L g6278 ( 
.A(n_6133),
.B(n_27),
.Y(n_6278)
);

BUFx2_ASAP7_75t_L g6279 ( 
.A(n_6079),
.Y(n_6279)
);

AND2x2_ASAP7_75t_L g6280 ( 
.A(n_6016),
.B(n_27),
.Y(n_6280)
);

BUFx6f_ASAP7_75t_L g6281 ( 
.A(n_6045),
.Y(n_6281)
);

INVx2_ASAP7_75t_L g6282 ( 
.A(n_6025),
.Y(n_6282)
);

NOR2xp33_ASAP7_75t_L g6283 ( 
.A(n_6079),
.B(n_6086),
.Y(n_6283)
);

HB1xp67_ASAP7_75t_L g6284 ( 
.A(n_6055),
.Y(n_6284)
);

INVx2_ASAP7_75t_L g6285 ( 
.A(n_6037),
.Y(n_6285)
);

INVx4_ASAP7_75t_L g6286 ( 
.A(n_6099),
.Y(n_6286)
);

AND2x2_ASAP7_75t_L g6287 ( 
.A(n_6038),
.B(n_28),
.Y(n_6287)
);

HB1xp67_ASAP7_75t_L g6288 ( 
.A(n_6060),
.Y(n_6288)
);

NAND2xp5_ASAP7_75t_L g6289 ( 
.A(n_6070),
.B(n_28),
.Y(n_6289)
);

INVx2_ASAP7_75t_L g6290 ( 
.A(n_6049),
.Y(n_6290)
);

AO21x2_ASAP7_75t_L g6291 ( 
.A1(n_6092),
.A2(n_28),
.B(n_29),
.Y(n_6291)
);

INVx2_ASAP7_75t_L g6292 ( 
.A(n_6051),
.Y(n_6292)
);

AND2x2_ASAP7_75t_L g6293 ( 
.A(n_6086),
.B(n_28),
.Y(n_6293)
);

AND2x2_ASAP7_75t_L g6294 ( 
.A(n_6095),
.B(n_29),
.Y(n_6294)
);

INVx2_ASAP7_75t_L g6295 ( 
.A(n_5982),
.Y(n_6295)
);

INVx1_ASAP7_75t_L g6296 ( 
.A(n_6073),
.Y(n_6296)
);

INVx1_ASAP7_75t_L g6297 ( 
.A(n_6093),
.Y(n_6297)
);

NAND2xp5_ASAP7_75t_L g6298 ( 
.A(n_6131),
.B(n_29),
.Y(n_6298)
);

AND2x2_ASAP7_75t_L g6299 ( 
.A(n_6125),
.B(n_29),
.Y(n_6299)
);

BUFx3_ASAP7_75t_L g6300 ( 
.A(n_6125),
.Y(n_6300)
);

AND2x2_ASAP7_75t_L g6301 ( 
.A(n_6127),
.B(n_30),
.Y(n_6301)
);

AO21x2_ASAP7_75t_L g6302 ( 
.A1(n_6105),
.A2(n_30),
.B(n_31),
.Y(n_6302)
);

AND2x2_ASAP7_75t_L g6303 ( 
.A(n_6127),
.B(n_31),
.Y(n_6303)
);

AND2x2_ASAP7_75t_L g6304 ( 
.A(n_6131),
.B(n_31),
.Y(n_6304)
);

INVx1_ASAP7_75t_L g6305 ( 
.A(n_6026),
.Y(n_6305)
);

INVx1_ASAP7_75t_L g6306 ( 
.A(n_6116),
.Y(n_6306)
);

NOR2x1_ASAP7_75t_SL g6307 ( 
.A(n_6013),
.B(n_509),
.Y(n_6307)
);

INVx1_ASAP7_75t_L g6308 ( 
.A(n_6074),
.Y(n_6308)
);

INVx2_ASAP7_75t_L g6309 ( 
.A(n_5980),
.Y(n_6309)
);

AND2x2_ASAP7_75t_L g6310 ( 
.A(n_6009),
.B(n_32),
.Y(n_6310)
);

NAND2xp5_ASAP7_75t_L g6311 ( 
.A(n_6130),
.B(n_32),
.Y(n_6311)
);

INVx1_ASAP7_75t_L g6312 ( 
.A(n_6074),
.Y(n_6312)
);

INVx2_ASAP7_75t_L g6313 ( 
.A(n_6142),
.Y(n_6313)
);

BUFx2_ASAP7_75t_L g6314 ( 
.A(n_6189),
.Y(n_6314)
);

OR2x6_ASAP7_75t_L g6315 ( 
.A(n_6198),
.B(n_510),
.Y(n_6315)
);

AND2x2_ASAP7_75t_L g6316 ( 
.A(n_6153),
.B(n_32),
.Y(n_6316)
);

BUFx3_ASAP7_75t_L g6317 ( 
.A(n_6148),
.Y(n_6317)
);

OR2x2_ASAP7_75t_L g6318 ( 
.A(n_6222),
.B(n_32),
.Y(n_6318)
);

AND2x2_ASAP7_75t_L g6319 ( 
.A(n_6153),
.B(n_33),
.Y(n_6319)
);

INVx1_ASAP7_75t_L g6320 ( 
.A(n_6150),
.Y(n_6320)
);

AND2x2_ASAP7_75t_L g6321 ( 
.A(n_6224),
.B(n_6168),
.Y(n_6321)
);

INVx2_ASAP7_75t_SL g6322 ( 
.A(n_6198),
.Y(n_6322)
);

HB1xp67_ASAP7_75t_L g6323 ( 
.A(n_6144),
.Y(n_6323)
);

AND2x2_ASAP7_75t_L g6324 ( 
.A(n_6171),
.B(n_33),
.Y(n_6324)
);

INVx1_ASAP7_75t_L g6325 ( 
.A(n_6146),
.Y(n_6325)
);

AND2x2_ASAP7_75t_L g6326 ( 
.A(n_6188),
.B(n_34),
.Y(n_6326)
);

BUFx2_ASAP7_75t_L g6327 ( 
.A(n_6162),
.Y(n_6327)
);

AND2x4_ASAP7_75t_L g6328 ( 
.A(n_6195),
.B(n_510),
.Y(n_6328)
);

AND2x2_ASAP7_75t_L g6329 ( 
.A(n_6154),
.B(n_34),
.Y(n_6329)
);

OR2x2_ASAP7_75t_L g6330 ( 
.A(n_6293),
.B(n_34),
.Y(n_6330)
);

AOI221xp5_ASAP7_75t_L g6331 ( 
.A1(n_6246),
.A2(n_36),
.B1(n_34),
.B2(n_35),
.C(n_37),
.Y(n_6331)
);

INVxp67_ASAP7_75t_L g6332 ( 
.A(n_6307),
.Y(n_6332)
);

INVx3_ASAP7_75t_L g6333 ( 
.A(n_6135),
.Y(n_6333)
);

INVx1_ASAP7_75t_L g6334 ( 
.A(n_6159),
.Y(n_6334)
);

INVx1_ASAP7_75t_L g6335 ( 
.A(n_6143),
.Y(n_6335)
);

INVx1_ASAP7_75t_L g6336 ( 
.A(n_6151),
.Y(n_6336)
);

INVx2_ASAP7_75t_L g6337 ( 
.A(n_6164),
.Y(n_6337)
);

NAND2xp5_ASAP7_75t_L g6338 ( 
.A(n_6141),
.B(n_35),
.Y(n_6338)
);

AND2x2_ASAP7_75t_L g6339 ( 
.A(n_6245),
.B(n_35),
.Y(n_6339)
);

AND2x2_ASAP7_75t_L g6340 ( 
.A(n_6267),
.B(n_35),
.Y(n_6340)
);

INVx1_ASAP7_75t_L g6341 ( 
.A(n_6167),
.Y(n_6341)
);

INVx2_ASAP7_75t_L g6342 ( 
.A(n_6271),
.Y(n_6342)
);

AND2x2_ASAP7_75t_L g6343 ( 
.A(n_6310),
.B(n_36),
.Y(n_6343)
);

INVx2_ASAP7_75t_L g6344 ( 
.A(n_6156),
.Y(n_6344)
);

AND2x4_ASAP7_75t_L g6345 ( 
.A(n_6135),
.B(n_511),
.Y(n_6345)
);

HB1xp67_ASAP7_75t_L g6346 ( 
.A(n_6147),
.Y(n_6346)
);

AND2x2_ASAP7_75t_SL g6347 ( 
.A(n_6192),
.B(n_511),
.Y(n_6347)
);

INVx1_ASAP7_75t_L g6348 ( 
.A(n_6252),
.Y(n_6348)
);

INVx3_ASAP7_75t_L g6349 ( 
.A(n_6137),
.Y(n_6349)
);

OR2x2_ASAP7_75t_L g6350 ( 
.A(n_6138),
.B(n_36),
.Y(n_6350)
);

NAND2xp5_ASAP7_75t_L g6351 ( 
.A(n_6266),
.B(n_36),
.Y(n_6351)
);

AND2x2_ASAP7_75t_L g6352 ( 
.A(n_6229),
.B(n_37),
.Y(n_6352)
);

CKINVDCx5p33_ASAP7_75t_R g6353 ( 
.A(n_6137),
.Y(n_6353)
);

NAND2x1_ASAP7_75t_L g6354 ( 
.A(n_6286),
.B(n_512),
.Y(n_6354)
);

INVx2_ASAP7_75t_L g6355 ( 
.A(n_6169),
.Y(n_6355)
);

AND2x4_ASAP7_75t_L g6356 ( 
.A(n_6149),
.B(n_512),
.Y(n_6356)
);

INVxp67_ASAP7_75t_SL g6357 ( 
.A(n_6307),
.Y(n_6357)
);

NAND2xp5_ASAP7_75t_L g6358 ( 
.A(n_6272),
.B(n_38),
.Y(n_6358)
);

NAND2xp5_ASAP7_75t_L g6359 ( 
.A(n_6273),
.B(n_6215),
.Y(n_6359)
);

CKINVDCx5p33_ASAP7_75t_R g6360 ( 
.A(n_6175),
.Y(n_6360)
);

INVx1_ASAP7_75t_L g6361 ( 
.A(n_6147),
.Y(n_6361)
);

AND2x2_ASAP7_75t_L g6362 ( 
.A(n_6182),
.B(n_38),
.Y(n_6362)
);

NAND2xp5_ASAP7_75t_L g6363 ( 
.A(n_6176),
.B(n_6305),
.Y(n_6363)
);

OR2x2_ASAP7_75t_L g6364 ( 
.A(n_6306),
.B(n_38),
.Y(n_6364)
);

NAND2xp5_ASAP7_75t_L g6365 ( 
.A(n_6181),
.B(n_38),
.Y(n_6365)
);

HB1xp67_ASAP7_75t_L g6366 ( 
.A(n_6308),
.Y(n_6366)
);

AND2x4_ASAP7_75t_L g6367 ( 
.A(n_6149),
.B(n_513),
.Y(n_6367)
);

AND2x2_ASAP7_75t_L g6368 ( 
.A(n_6186),
.B(n_39),
.Y(n_6368)
);

NAND2xp5_ASAP7_75t_L g6369 ( 
.A(n_6304),
.B(n_39),
.Y(n_6369)
);

HB1xp67_ASAP7_75t_L g6370 ( 
.A(n_6308),
.Y(n_6370)
);

NAND2xp5_ASAP7_75t_L g6371 ( 
.A(n_6299),
.B(n_39),
.Y(n_6371)
);

OR2x2_ASAP7_75t_L g6372 ( 
.A(n_6270),
.B(n_40),
.Y(n_6372)
);

INVx1_ASAP7_75t_L g6373 ( 
.A(n_6312),
.Y(n_6373)
);

INVx3_ASAP7_75t_L g6374 ( 
.A(n_6163),
.Y(n_6374)
);

NAND2xp5_ASAP7_75t_SL g6375 ( 
.A(n_6227),
.B(n_40),
.Y(n_6375)
);

INVx1_ASAP7_75t_L g6376 ( 
.A(n_6312),
.Y(n_6376)
);

AND2x2_ASAP7_75t_L g6377 ( 
.A(n_6226),
.B(n_40),
.Y(n_6377)
);

INVx2_ASAP7_75t_L g6378 ( 
.A(n_6152),
.Y(n_6378)
);

AND3x1_ASAP7_75t_L g6379 ( 
.A(n_6217),
.B(n_40),
.C(n_41),
.Y(n_6379)
);

AND2x4_ASAP7_75t_L g6380 ( 
.A(n_6157),
.B(n_513),
.Y(n_6380)
);

AND2x2_ASAP7_75t_L g6381 ( 
.A(n_6242),
.B(n_41),
.Y(n_6381)
);

INVx1_ASAP7_75t_L g6382 ( 
.A(n_6185),
.Y(n_6382)
);

INVx1_ASAP7_75t_L g6383 ( 
.A(n_6191),
.Y(n_6383)
);

INVx2_ASAP7_75t_L g6384 ( 
.A(n_6158),
.Y(n_6384)
);

INVxp67_ASAP7_75t_SL g6385 ( 
.A(n_6225),
.Y(n_6385)
);

AND2x2_ASAP7_75t_L g6386 ( 
.A(n_6294),
.B(n_41),
.Y(n_6386)
);

INVx1_ASAP7_75t_L g6387 ( 
.A(n_6196),
.Y(n_6387)
);

BUFx3_ASAP7_75t_L g6388 ( 
.A(n_6172),
.Y(n_6388)
);

INVx1_ASAP7_75t_L g6389 ( 
.A(n_6184),
.Y(n_6389)
);

INVx1_ASAP7_75t_L g6390 ( 
.A(n_6279),
.Y(n_6390)
);

INVx2_ASAP7_75t_L g6391 ( 
.A(n_6174),
.Y(n_6391)
);

AND2x2_ASAP7_75t_L g6392 ( 
.A(n_6194),
.B(n_41),
.Y(n_6392)
);

INVx2_ASAP7_75t_L g6393 ( 
.A(n_6180),
.Y(n_6393)
);

AND2x2_ASAP7_75t_L g6394 ( 
.A(n_6197),
.B(n_42),
.Y(n_6394)
);

INVx2_ASAP7_75t_L g6395 ( 
.A(n_6140),
.Y(n_6395)
);

INVx2_ASAP7_75t_L g6396 ( 
.A(n_6309),
.Y(n_6396)
);

INVx2_ASAP7_75t_L g6397 ( 
.A(n_6221),
.Y(n_6397)
);

INVx2_ASAP7_75t_SL g6398 ( 
.A(n_6177),
.Y(n_6398)
);

HB1xp67_ASAP7_75t_L g6399 ( 
.A(n_6216),
.Y(n_6399)
);

INVx1_ASAP7_75t_L g6400 ( 
.A(n_6230),
.Y(n_6400)
);

INVx1_ASAP7_75t_SL g6401 ( 
.A(n_6178),
.Y(n_6401)
);

AND2x2_ASAP7_75t_L g6402 ( 
.A(n_6157),
.B(n_42),
.Y(n_6402)
);

INVx2_ASAP7_75t_L g6403 ( 
.A(n_6239),
.Y(n_6403)
);

INVx1_ASAP7_75t_L g6404 ( 
.A(n_6251),
.Y(n_6404)
);

OR2x2_ASAP7_75t_L g6405 ( 
.A(n_6311),
.B(n_42),
.Y(n_6405)
);

INVx1_ASAP7_75t_L g6406 ( 
.A(n_6244),
.Y(n_6406)
);

NAND2xp5_ASAP7_75t_L g6407 ( 
.A(n_6301),
.B(n_43),
.Y(n_6407)
);

AND2x2_ASAP7_75t_L g6408 ( 
.A(n_6237),
.B(n_43),
.Y(n_6408)
);

INVx1_ASAP7_75t_L g6409 ( 
.A(n_6250),
.Y(n_6409)
);

INVx1_ASAP7_75t_L g6410 ( 
.A(n_6254),
.Y(n_6410)
);

INVx1_ASAP7_75t_L g6411 ( 
.A(n_6257),
.Y(n_6411)
);

INVx2_ASAP7_75t_L g6412 ( 
.A(n_6209),
.Y(n_6412)
);

INVx1_ASAP7_75t_L g6413 ( 
.A(n_6258),
.Y(n_6413)
);

AND2x2_ASAP7_75t_L g6414 ( 
.A(n_6237),
.B(n_43),
.Y(n_6414)
);

AND2x2_ASAP7_75t_L g6415 ( 
.A(n_6213),
.B(n_44),
.Y(n_6415)
);

INVx1_ASAP7_75t_L g6416 ( 
.A(n_6261),
.Y(n_6416)
);

AND2x2_ASAP7_75t_L g6417 ( 
.A(n_6203),
.B(n_44),
.Y(n_6417)
);

INVx1_ASAP7_75t_L g6418 ( 
.A(n_6207),
.Y(n_6418)
);

HB1xp67_ASAP7_75t_L g6419 ( 
.A(n_6216),
.Y(n_6419)
);

AND2x2_ASAP7_75t_L g6420 ( 
.A(n_6214),
.B(n_44),
.Y(n_6420)
);

INVx2_ASAP7_75t_L g6421 ( 
.A(n_6161),
.Y(n_6421)
);

INVx1_ASAP7_75t_L g6422 ( 
.A(n_6219),
.Y(n_6422)
);

INVx1_ASAP7_75t_L g6423 ( 
.A(n_6276),
.Y(n_6423)
);

INVx3_ASAP7_75t_L g6424 ( 
.A(n_6241),
.Y(n_6424)
);

AND2x2_ASAP7_75t_L g6425 ( 
.A(n_6280),
.B(n_6287),
.Y(n_6425)
);

HB1xp67_ASAP7_75t_L g6426 ( 
.A(n_6218),
.Y(n_6426)
);

OR2x2_ASAP7_75t_L g6427 ( 
.A(n_6260),
.B(n_514),
.Y(n_6427)
);

OAI21xp5_ASAP7_75t_SL g6428 ( 
.A1(n_6199),
.A2(n_515),
.B(n_516),
.Y(n_6428)
);

INVx1_ASAP7_75t_L g6429 ( 
.A(n_6218),
.Y(n_6429)
);

OR2x2_ASAP7_75t_L g6430 ( 
.A(n_6187),
.B(n_515),
.Y(n_6430)
);

AND2x2_ASAP7_75t_L g6431 ( 
.A(n_6233),
.B(n_516),
.Y(n_6431)
);

INVx1_ASAP7_75t_L g6432 ( 
.A(n_6145),
.Y(n_6432)
);

BUFx3_ASAP7_75t_L g6433 ( 
.A(n_6166),
.Y(n_6433)
);

INVx2_ASAP7_75t_L g6434 ( 
.A(n_6248),
.Y(n_6434)
);

HB1xp67_ASAP7_75t_L g6435 ( 
.A(n_6235),
.Y(n_6435)
);

INVx2_ASAP7_75t_SL g6436 ( 
.A(n_6288),
.Y(n_6436)
);

NOR2x1p5_ASAP7_75t_L g6437 ( 
.A(n_6278),
.B(n_517),
.Y(n_6437)
);

AND2x2_ASAP7_75t_L g6438 ( 
.A(n_6228),
.B(n_517),
.Y(n_6438)
);

INVx1_ASAP7_75t_SL g6439 ( 
.A(n_6170),
.Y(n_6439)
);

NOR2xp33_ASAP7_75t_L g6440 ( 
.A(n_6173),
.B(n_517),
.Y(n_6440)
);

BUFx2_ASAP7_75t_L g6441 ( 
.A(n_6231),
.Y(n_6441)
);

INVxp67_ASAP7_75t_L g6442 ( 
.A(n_6283),
.Y(n_6442)
);

INVx3_ASAP7_75t_L g6443 ( 
.A(n_6264),
.Y(n_6443)
);

BUFx3_ASAP7_75t_L g6444 ( 
.A(n_6179),
.Y(n_6444)
);

NAND2xp5_ASAP7_75t_L g6445 ( 
.A(n_6303),
.B(n_518),
.Y(n_6445)
);

INVx1_ASAP7_75t_L g6446 ( 
.A(n_6249),
.Y(n_6446)
);

AND2x4_ASAP7_75t_L g6447 ( 
.A(n_6211),
.B(n_518),
.Y(n_6447)
);

NAND2xp5_ASAP7_75t_L g6448 ( 
.A(n_6302),
.B(n_519),
.Y(n_6448)
);

NAND2xp5_ASAP7_75t_L g6449 ( 
.A(n_6232),
.B(n_519),
.Y(n_6449)
);

INVx1_ASAP7_75t_L g6450 ( 
.A(n_6277),
.Y(n_6450)
);

INVx1_ASAP7_75t_SL g6451 ( 
.A(n_6211),
.Y(n_6451)
);

INVx1_ASAP7_75t_L g6452 ( 
.A(n_6284),
.Y(n_6452)
);

INVx2_ASAP7_75t_L g6453 ( 
.A(n_6269),
.Y(n_6453)
);

INVx1_ASAP7_75t_L g6454 ( 
.A(n_6297),
.Y(n_6454)
);

INVx2_ASAP7_75t_L g6455 ( 
.A(n_6282),
.Y(n_6455)
);

INVx1_ASAP7_75t_L g6456 ( 
.A(n_6183),
.Y(n_6456)
);

OR2x2_ASAP7_75t_L g6457 ( 
.A(n_6240),
.B(n_520),
.Y(n_6457)
);

INVx2_ASAP7_75t_L g6458 ( 
.A(n_6285),
.Y(n_6458)
);

INVx1_ASAP7_75t_L g6459 ( 
.A(n_6201),
.Y(n_6459)
);

INVx2_ASAP7_75t_L g6460 ( 
.A(n_6290),
.Y(n_6460)
);

INVx4_ASAP7_75t_L g6461 ( 
.A(n_6291),
.Y(n_6461)
);

INVx2_ASAP7_75t_SL g6462 ( 
.A(n_6236),
.Y(n_6462)
);

AND2x2_ASAP7_75t_L g6463 ( 
.A(n_6202),
.B(n_520),
.Y(n_6463)
);

HB1xp67_ASAP7_75t_SL g6464 ( 
.A(n_6165),
.Y(n_6464)
);

INVx5_ASAP7_75t_L g6465 ( 
.A(n_6243),
.Y(n_6465)
);

INVx1_ASAP7_75t_L g6466 ( 
.A(n_6160),
.Y(n_6466)
);

AO21x2_ASAP7_75t_L g6467 ( 
.A1(n_6190),
.A2(n_520),
.B(n_521),
.Y(n_6467)
);

INVx1_ASAP7_75t_L g6468 ( 
.A(n_6206),
.Y(n_6468)
);

INVx2_ASAP7_75t_SL g6469 ( 
.A(n_6223),
.Y(n_6469)
);

AND2x4_ASAP7_75t_L g6470 ( 
.A(n_6165),
.B(n_521),
.Y(n_6470)
);

INVxp67_ASAP7_75t_L g6471 ( 
.A(n_6238),
.Y(n_6471)
);

INVxp67_ASAP7_75t_L g6472 ( 
.A(n_6289),
.Y(n_6472)
);

AND2x4_ASAP7_75t_L g6473 ( 
.A(n_6200),
.B(n_521),
.Y(n_6473)
);

BUFx6f_ASAP7_75t_L g6474 ( 
.A(n_6298),
.Y(n_6474)
);

AND2x4_ASAP7_75t_L g6475 ( 
.A(n_6292),
.B(n_6247),
.Y(n_6475)
);

INVx3_ASAP7_75t_L g6476 ( 
.A(n_6243),
.Y(n_6476)
);

INVx1_ASAP7_75t_L g6477 ( 
.A(n_6206),
.Y(n_6477)
);

AND2x2_ASAP7_75t_L g6478 ( 
.A(n_6220),
.B(n_522),
.Y(n_6478)
);

NOR2x1_ASAP7_75t_L g6479 ( 
.A(n_6286),
.B(n_522),
.Y(n_6479)
);

INVx2_ASAP7_75t_L g6480 ( 
.A(n_6295),
.Y(n_6480)
);

AND2x2_ASAP7_75t_L g6481 ( 
.A(n_6300),
.B(n_522),
.Y(n_6481)
);

INVx2_ASAP7_75t_L g6482 ( 
.A(n_6234),
.Y(n_6482)
);

AND2x2_ASAP7_75t_L g6483 ( 
.A(n_6268),
.B(n_523),
.Y(n_6483)
);

INVx2_ASAP7_75t_L g6484 ( 
.A(n_6256),
.Y(n_6484)
);

AND2x2_ASAP7_75t_L g6485 ( 
.A(n_6259),
.B(n_523),
.Y(n_6485)
);

INVx2_ASAP7_75t_L g6486 ( 
.A(n_6262),
.Y(n_6486)
);

OA21x2_ASAP7_75t_L g6487 ( 
.A1(n_6332),
.A2(n_6210),
.B(n_6208),
.Y(n_6487)
);

INVx1_ASAP7_75t_L g6488 ( 
.A(n_6314),
.Y(n_6488)
);

AND2x2_ASAP7_75t_L g6489 ( 
.A(n_6322),
.B(n_6274),
.Y(n_6489)
);

AOI21xp33_ASAP7_75t_L g6490 ( 
.A1(n_6314),
.A2(n_6136),
.B(n_6253),
.Y(n_6490)
);

AND2x2_ASAP7_75t_L g6491 ( 
.A(n_6321),
.B(n_6296),
.Y(n_6491)
);

INVx1_ASAP7_75t_L g6492 ( 
.A(n_6339),
.Y(n_6492)
);

INVx2_ASAP7_75t_L g6493 ( 
.A(n_6345),
.Y(n_6493)
);

INVx2_ASAP7_75t_SL g6494 ( 
.A(n_6317),
.Y(n_6494)
);

INVx1_ASAP7_75t_SL g6495 ( 
.A(n_6353),
.Y(n_6495)
);

INVx2_ASAP7_75t_L g6496 ( 
.A(n_6345),
.Y(n_6496)
);

BUFx6f_ASAP7_75t_L g6497 ( 
.A(n_6333),
.Y(n_6497)
);

INVx2_ASAP7_75t_SL g6498 ( 
.A(n_6349),
.Y(n_6498)
);

INVx2_ASAP7_75t_L g6499 ( 
.A(n_6316),
.Y(n_6499)
);

NAND2xp5_ASAP7_75t_L g6500 ( 
.A(n_6327),
.B(n_6263),
.Y(n_6500)
);

NAND2xp5_ASAP7_75t_L g6501 ( 
.A(n_6327),
.B(n_6265),
.Y(n_6501)
);

INVx2_ASAP7_75t_L g6502 ( 
.A(n_6319),
.Y(n_6502)
);

AOI221xp5_ASAP7_75t_L g6503 ( 
.A1(n_6442),
.A2(n_6139),
.B1(n_6275),
.B2(n_6255),
.C(n_6208),
.Y(n_6503)
);

INVx1_ASAP7_75t_L g6504 ( 
.A(n_6323),
.Y(n_6504)
);

INVx2_ASAP7_75t_L g6505 ( 
.A(n_6342),
.Y(n_6505)
);

INVx2_ASAP7_75t_L g6506 ( 
.A(n_6313),
.Y(n_6506)
);

INVxp67_ASAP7_75t_SL g6507 ( 
.A(n_6324),
.Y(n_6507)
);

BUFx2_ASAP7_75t_SL g6508 ( 
.A(n_6328),
.Y(n_6508)
);

AND2x2_ASAP7_75t_L g6509 ( 
.A(n_6347),
.B(n_6374),
.Y(n_6509)
);

INVx1_ASAP7_75t_L g6510 ( 
.A(n_6435),
.Y(n_6510)
);

NAND2xp5_ASAP7_75t_SL g6511 ( 
.A(n_6436),
.B(n_6243),
.Y(n_6511)
);

OA21x2_ASAP7_75t_L g6512 ( 
.A1(n_6357),
.A2(n_6212),
.B(n_6210),
.Y(n_6512)
);

AOI21xp5_ASAP7_75t_L g6513 ( 
.A1(n_6375),
.A2(n_6255),
.B(n_6212),
.Y(n_6513)
);

INVx5_ASAP7_75t_L g6514 ( 
.A(n_6315),
.Y(n_6514)
);

INVx1_ASAP7_75t_L g6515 ( 
.A(n_6352),
.Y(n_6515)
);

INVx1_ASAP7_75t_L g6516 ( 
.A(n_6481),
.Y(n_6516)
);

NOR2xp33_ASAP7_75t_L g6517 ( 
.A(n_6360),
.B(n_6281),
.Y(n_6517)
);

OAI21x1_ASAP7_75t_L g6518 ( 
.A1(n_6476),
.A2(n_6281),
.B(n_6204),
.Y(n_6518)
);

INVxp67_ASAP7_75t_SL g6519 ( 
.A(n_6354),
.Y(n_6519)
);

INVx1_ASAP7_75t_L g6520 ( 
.A(n_6315),
.Y(n_6520)
);

HB1xp67_ASAP7_75t_L g6521 ( 
.A(n_6390),
.Y(n_6521)
);

AND2x2_ASAP7_75t_L g6522 ( 
.A(n_6388),
.B(n_6281),
.Y(n_6522)
);

OA21x2_ASAP7_75t_L g6523 ( 
.A1(n_6441),
.A2(n_6205),
.B(n_6155),
.Y(n_6523)
);

INVx1_ASAP7_75t_L g6524 ( 
.A(n_6382),
.Y(n_6524)
);

OAI21x1_ASAP7_75t_L g6525 ( 
.A1(n_6383),
.A2(n_6155),
.B(n_6193),
.Y(n_6525)
);

INVx2_ASAP7_75t_L g6526 ( 
.A(n_6328),
.Y(n_6526)
);

NAND2xp5_ASAP7_75t_SL g6527 ( 
.A(n_6475),
.B(n_6155),
.Y(n_6527)
);

BUFx3_ASAP7_75t_L g6528 ( 
.A(n_6470),
.Y(n_6528)
);

AND2x6_ASAP7_75t_L g6529 ( 
.A(n_6479),
.B(n_523),
.Y(n_6529)
);

NAND4xp25_ASAP7_75t_L g6530 ( 
.A(n_6363),
.B(n_526),
.C(n_524),
.D(n_525),
.Y(n_6530)
);

NAND2xp5_ASAP7_75t_L g6531 ( 
.A(n_6385),
.B(n_524),
.Y(n_6531)
);

HB1xp67_ASAP7_75t_L g6532 ( 
.A(n_6346),
.Y(n_6532)
);

OAI21x1_ASAP7_75t_L g6533 ( 
.A1(n_6387),
.A2(n_525),
.B(n_527),
.Y(n_6533)
);

INVx1_ASAP7_75t_L g6534 ( 
.A(n_6326),
.Y(n_6534)
);

INVx1_ASAP7_75t_L g6535 ( 
.A(n_6366),
.Y(n_6535)
);

INVx3_ASAP7_75t_L g6536 ( 
.A(n_6424),
.Y(n_6536)
);

A2O1A1Ixp33_ASAP7_75t_L g6537 ( 
.A1(n_6428),
.A2(n_528),
.B(n_525),
.C(n_527),
.Y(n_6537)
);

AOI21xp5_ASAP7_75t_L g6538 ( 
.A1(n_6354),
.A2(n_527),
.B(n_528),
.Y(n_6538)
);

BUFx3_ASAP7_75t_L g6539 ( 
.A(n_6470),
.Y(n_6539)
);

A2O1A1Ixp33_ASAP7_75t_L g6540 ( 
.A1(n_6320),
.A2(n_530),
.B(n_528),
.C(n_529),
.Y(n_6540)
);

INVx1_ASAP7_75t_L g6541 ( 
.A(n_6370),
.Y(n_6541)
);

NAND3xp33_ASAP7_75t_L g6542 ( 
.A(n_6325),
.B(n_529),
.C(n_530),
.Y(n_6542)
);

INVx1_ASAP7_75t_L g6543 ( 
.A(n_6399),
.Y(n_6543)
);

INVx1_ASAP7_75t_L g6544 ( 
.A(n_6419),
.Y(n_6544)
);

OAI21xp33_ASAP7_75t_L g6545 ( 
.A1(n_6451),
.A2(n_530),
.B(n_531),
.Y(n_6545)
);

INVx1_ASAP7_75t_L g6546 ( 
.A(n_6426),
.Y(n_6546)
);

INVx2_ASAP7_75t_SL g6547 ( 
.A(n_6378),
.Y(n_6547)
);

AO21x2_ASAP7_75t_L g6548 ( 
.A1(n_6334),
.A2(n_531),
.B(n_532),
.Y(n_6548)
);

NOR2xp33_ASAP7_75t_L g6549 ( 
.A(n_6461),
.B(n_6401),
.Y(n_6549)
);

OAI21xp5_ASAP7_75t_L g6550 ( 
.A1(n_6471),
.A2(n_532),
.B(n_533),
.Y(n_6550)
);

INVx2_ASAP7_75t_L g6551 ( 
.A(n_6443),
.Y(n_6551)
);

BUFx2_ASAP7_75t_L g6552 ( 
.A(n_6337),
.Y(n_6552)
);

INVx2_ASAP7_75t_L g6553 ( 
.A(n_6447),
.Y(n_6553)
);

AND2x2_ASAP7_75t_L g6554 ( 
.A(n_6415),
.B(n_1057),
.Y(n_6554)
);

BUFx2_ASAP7_75t_L g6555 ( 
.A(n_6355),
.Y(n_6555)
);

AO22x2_ASAP7_75t_L g6556 ( 
.A1(n_6410),
.A2(n_6411),
.B1(n_6416),
.B2(n_6413),
.Y(n_6556)
);

HB1xp67_ASAP7_75t_L g6557 ( 
.A(n_6384),
.Y(n_6557)
);

INVx1_ASAP7_75t_L g6558 ( 
.A(n_6377),
.Y(n_6558)
);

INVx2_ASAP7_75t_L g6559 ( 
.A(n_6447),
.Y(n_6559)
);

INVx1_ASAP7_75t_L g6560 ( 
.A(n_6341),
.Y(n_6560)
);

INVx4_ASAP7_75t_R g6561 ( 
.A(n_6464),
.Y(n_6561)
);

INVx2_ASAP7_75t_L g6562 ( 
.A(n_6395),
.Y(n_6562)
);

INVx1_ASAP7_75t_L g6563 ( 
.A(n_6335),
.Y(n_6563)
);

INVx2_ASAP7_75t_SL g6564 ( 
.A(n_6380),
.Y(n_6564)
);

AND2x2_ASAP7_75t_L g6565 ( 
.A(n_6425),
.B(n_1058),
.Y(n_6565)
);

INVx4_ASAP7_75t_SL g6566 ( 
.A(n_6380),
.Y(n_6566)
);

AND2x4_ASAP7_75t_SL g6567 ( 
.A(n_6356),
.B(n_532),
.Y(n_6567)
);

OAI21x1_ASAP7_75t_L g6568 ( 
.A1(n_6389),
.A2(n_534),
.B(n_535),
.Y(n_6568)
);

NAND2xp5_ASAP7_75t_L g6569 ( 
.A(n_6336),
.B(n_534),
.Y(n_6569)
);

AND2x2_ASAP7_75t_L g6570 ( 
.A(n_6398),
.B(n_1066),
.Y(n_6570)
);

AOI21xp5_ASAP7_75t_L g6571 ( 
.A1(n_6359),
.A2(n_535),
.B(n_536),
.Y(n_6571)
);

OAI21x1_ASAP7_75t_L g6572 ( 
.A1(n_6361),
.A2(n_6376),
.B(n_6373),
.Y(n_6572)
);

OR2x2_ASAP7_75t_L g6573 ( 
.A(n_6372),
.B(n_535),
.Y(n_6573)
);

INVx1_ASAP7_75t_L g6574 ( 
.A(n_6391),
.Y(n_6574)
);

INVx2_ASAP7_75t_L g6575 ( 
.A(n_6396),
.Y(n_6575)
);

BUFx3_ASAP7_75t_L g6576 ( 
.A(n_6402),
.Y(n_6576)
);

INVx1_ASAP7_75t_L g6577 ( 
.A(n_6393),
.Y(n_6577)
);

INVx2_ASAP7_75t_L g6578 ( 
.A(n_6412),
.Y(n_6578)
);

INVxp67_ASAP7_75t_L g6579 ( 
.A(n_6392),
.Y(n_6579)
);

BUFx2_ASAP7_75t_L g6580 ( 
.A(n_6421),
.Y(n_6580)
);

INVxp67_ASAP7_75t_SL g6581 ( 
.A(n_6369),
.Y(n_6581)
);

INVx1_ASAP7_75t_L g6582 ( 
.A(n_6400),
.Y(n_6582)
);

AND2x2_ASAP7_75t_L g6583 ( 
.A(n_6356),
.B(n_1068),
.Y(n_6583)
);

INVx2_ASAP7_75t_L g6584 ( 
.A(n_6397),
.Y(n_6584)
);

OR2x2_ASAP7_75t_L g6585 ( 
.A(n_6430),
.B(n_536),
.Y(n_6585)
);

INVx1_ASAP7_75t_L g6586 ( 
.A(n_6404),
.Y(n_6586)
);

INVx2_ASAP7_75t_L g6587 ( 
.A(n_6403),
.Y(n_6587)
);

INVx1_ASAP7_75t_L g6588 ( 
.A(n_6423),
.Y(n_6588)
);

INVx1_ASAP7_75t_SL g6589 ( 
.A(n_6408),
.Y(n_6589)
);

AOI21xp5_ASAP7_75t_L g6590 ( 
.A1(n_6379),
.A2(n_6441),
.B(n_6351),
.Y(n_6590)
);

BUFx2_ASAP7_75t_L g6591 ( 
.A(n_6434),
.Y(n_6591)
);

INVx1_ASAP7_75t_L g6592 ( 
.A(n_6348),
.Y(n_6592)
);

NAND2xp5_ASAP7_75t_L g6593 ( 
.A(n_6422),
.B(n_537),
.Y(n_6593)
);

INVx2_ASAP7_75t_L g6594 ( 
.A(n_6453),
.Y(n_6594)
);

INVx2_ASAP7_75t_L g6595 ( 
.A(n_6455),
.Y(n_6595)
);

AO21x1_ASAP7_75t_L g6596 ( 
.A1(n_6429),
.A2(n_539),
.B(n_538),
.Y(n_6596)
);

NAND2xp5_ASAP7_75t_L g6597 ( 
.A(n_6439),
.B(n_6344),
.Y(n_6597)
);

NAND2xp5_ASAP7_75t_L g6598 ( 
.A(n_6437),
.B(n_537),
.Y(n_6598)
);

INVxp67_ASAP7_75t_L g6599 ( 
.A(n_6394),
.Y(n_6599)
);

INVx1_ASAP7_75t_L g6600 ( 
.A(n_6330),
.Y(n_6600)
);

OA21x2_ASAP7_75t_L g6601 ( 
.A1(n_6480),
.A2(n_537),
.B(n_538),
.Y(n_6601)
);

INVx2_ASAP7_75t_SL g6602 ( 
.A(n_6462),
.Y(n_6602)
);

INVx2_ASAP7_75t_L g6603 ( 
.A(n_6458),
.Y(n_6603)
);

INVx2_ASAP7_75t_L g6604 ( 
.A(n_6460),
.Y(n_6604)
);

BUFx2_ASAP7_75t_L g6605 ( 
.A(n_6367),
.Y(n_6605)
);

INVx1_ASAP7_75t_L g6606 ( 
.A(n_6371),
.Y(n_6606)
);

BUFx6f_ASAP7_75t_L g6607 ( 
.A(n_6414),
.Y(n_6607)
);

AOI21xp5_ASAP7_75t_L g6608 ( 
.A1(n_6358),
.A2(n_538),
.B(n_539),
.Y(n_6608)
);

INVx1_ASAP7_75t_L g6609 ( 
.A(n_6407),
.Y(n_6609)
);

CKINVDCx5p33_ASAP7_75t_R g6610 ( 
.A(n_6362),
.Y(n_6610)
);

OA21x2_ASAP7_75t_L g6611 ( 
.A1(n_6483),
.A2(n_539),
.B(n_540),
.Y(n_6611)
);

AND2x2_ASAP7_75t_L g6612 ( 
.A(n_6367),
.B(n_1048),
.Y(n_6612)
);

NOR2xp33_ASAP7_75t_R g6613 ( 
.A(n_6417),
.B(n_6420),
.Y(n_6613)
);

AND2x4_ASAP7_75t_L g6614 ( 
.A(n_6418),
.B(n_540),
.Y(n_6614)
);

A2O1A1Ixp33_ASAP7_75t_L g6615 ( 
.A1(n_6433),
.A2(n_542),
.B(n_540),
.C(n_541),
.Y(n_6615)
);

OR2x2_ASAP7_75t_L g6616 ( 
.A(n_6350),
.B(n_541),
.Y(n_6616)
);

OAI21xp33_ASAP7_75t_L g6617 ( 
.A1(n_6446),
.A2(n_6452),
.B(n_6450),
.Y(n_6617)
);

INVx2_ASAP7_75t_L g6618 ( 
.A(n_6469),
.Y(n_6618)
);

NAND3xp33_ASAP7_75t_L g6619 ( 
.A(n_6331),
.B(n_541),
.C(n_542),
.Y(n_6619)
);

AND2x2_ASAP7_75t_L g6620 ( 
.A(n_6431),
.B(n_6406),
.Y(n_6620)
);

INVx2_ASAP7_75t_SL g6621 ( 
.A(n_6473),
.Y(n_6621)
);

INVx3_ASAP7_75t_L g6622 ( 
.A(n_6444),
.Y(n_6622)
);

INVx2_ASAP7_75t_L g6623 ( 
.A(n_6474),
.Y(n_6623)
);

OA21x2_ASAP7_75t_L g6624 ( 
.A1(n_6472),
.A2(n_542),
.B(n_543),
.Y(n_6624)
);

INVx3_ASAP7_75t_L g6625 ( 
.A(n_6474),
.Y(n_6625)
);

INVx2_ASAP7_75t_SL g6626 ( 
.A(n_6340),
.Y(n_6626)
);

A2O1A1Ixp33_ASAP7_75t_L g6627 ( 
.A1(n_6409),
.A2(n_546),
.B(n_543),
.C(n_544),
.Y(n_6627)
);

NAND2xp5_ASAP7_75t_L g6628 ( 
.A(n_6432),
.B(n_543),
.Y(n_6628)
);

INVx1_ASAP7_75t_L g6629 ( 
.A(n_6364),
.Y(n_6629)
);

AO21x2_ASAP7_75t_L g6630 ( 
.A1(n_6454),
.A2(n_546),
.B(n_547),
.Y(n_6630)
);

INVx1_ASAP7_75t_L g6631 ( 
.A(n_6448),
.Y(n_6631)
);

O2A1O1Ixp33_ASAP7_75t_L g6632 ( 
.A1(n_6467),
.A2(n_6459),
.B(n_6445),
.C(n_6449),
.Y(n_6632)
);

AO22x2_ASAP7_75t_L g6633 ( 
.A1(n_6456),
.A2(n_549),
.B1(n_547),
.B2(n_548),
.Y(n_6633)
);

AND2x2_ASAP7_75t_L g6634 ( 
.A(n_6478),
.B(n_1056),
.Y(n_6634)
);

BUFx6f_ASAP7_75t_L g6635 ( 
.A(n_6368),
.Y(n_6635)
);

OAI211xp5_ASAP7_75t_L g6636 ( 
.A1(n_6466),
.A2(n_550),
.B(n_548),
.C(n_549),
.Y(n_6636)
);

AOI21xp5_ASAP7_75t_L g6637 ( 
.A1(n_6338),
.A2(n_6365),
.B(n_6440),
.Y(n_6637)
);

HB1xp67_ASAP7_75t_L g6638 ( 
.A(n_6463),
.Y(n_6638)
);

INVx2_ASAP7_75t_SL g6639 ( 
.A(n_6386),
.Y(n_6639)
);

INVx1_ASAP7_75t_L g6640 ( 
.A(n_6485),
.Y(n_6640)
);

AOI21xp5_ASAP7_75t_L g6641 ( 
.A1(n_6482),
.A2(n_548),
.B(n_549),
.Y(n_6641)
);

INVx2_ASAP7_75t_L g6642 ( 
.A(n_6465),
.Y(n_6642)
);

NAND3xp33_ASAP7_75t_L g6643 ( 
.A(n_6465),
.B(n_550),
.C(n_551),
.Y(n_6643)
);

INVx1_ASAP7_75t_L g6644 ( 
.A(n_6457),
.Y(n_6644)
);

INVx2_ASAP7_75t_L g6645 ( 
.A(n_6465),
.Y(n_6645)
);

INVx1_ASAP7_75t_L g6646 ( 
.A(n_6329),
.Y(n_6646)
);

INVx1_ASAP7_75t_L g6647 ( 
.A(n_6405),
.Y(n_6647)
);

INVx2_ASAP7_75t_L g6648 ( 
.A(n_6484),
.Y(n_6648)
);

NAND2xp5_ASAP7_75t_L g6649 ( 
.A(n_6486),
.B(n_550),
.Y(n_6649)
);

INVxp67_ASAP7_75t_L g6650 ( 
.A(n_6343),
.Y(n_6650)
);

OAI21xp33_ASAP7_75t_L g6651 ( 
.A1(n_6468),
.A2(n_551),
.B(n_552),
.Y(n_6651)
);

NAND2xp5_ASAP7_75t_L g6652 ( 
.A(n_6381),
.B(n_551),
.Y(n_6652)
);

INVx1_ASAP7_75t_L g6653 ( 
.A(n_6318),
.Y(n_6653)
);

AOI21xp5_ASAP7_75t_L g6654 ( 
.A1(n_6477),
.A2(n_552),
.B(n_553),
.Y(n_6654)
);

INVx1_ASAP7_75t_L g6655 ( 
.A(n_6427),
.Y(n_6655)
);

OR2x2_ASAP7_75t_L g6656 ( 
.A(n_6438),
.B(n_552),
.Y(n_6656)
);

AND2x2_ASAP7_75t_L g6657 ( 
.A(n_6322),
.B(n_553),
.Y(n_6657)
);

AND2x2_ASAP7_75t_L g6658 ( 
.A(n_6322),
.B(n_553),
.Y(n_6658)
);

OR2x2_ASAP7_75t_L g6659 ( 
.A(n_6314),
.B(n_554),
.Y(n_6659)
);

INVx1_ASAP7_75t_L g6660 ( 
.A(n_6314),
.Y(n_6660)
);

AND2x2_ASAP7_75t_L g6661 ( 
.A(n_6322),
.B(n_1045),
.Y(n_6661)
);

OA21x2_ASAP7_75t_L g6662 ( 
.A1(n_6332),
.A2(n_554),
.B(n_555),
.Y(n_6662)
);

INVx1_ASAP7_75t_L g6663 ( 
.A(n_6314),
.Y(n_6663)
);

INVx2_ASAP7_75t_L g6664 ( 
.A(n_6314),
.Y(n_6664)
);

INVx1_ASAP7_75t_L g6665 ( 
.A(n_6314),
.Y(n_6665)
);

AOI21xp5_ASAP7_75t_L g6666 ( 
.A1(n_6357),
.A2(n_554),
.B(n_555),
.Y(n_6666)
);

INVxp67_ASAP7_75t_SL g6667 ( 
.A(n_6322),
.Y(n_6667)
);

INVx1_ASAP7_75t_L g6668 ( 
.A(n_6314),
.Y(n_6668)
);

AOI21xp5_ASAP7_75t_L g6669 ( 
.A1(n_6357),
.A2(n_555),
.B(n_556),
.Y(n_6669)
);

INVx2_ASAP7_75t_L g6670 ( 
.A(n_6314),
.Y(n_6670)
);

AO21x2_ASAP7_75t_L g6671 ( 
.A1(n_6375),
.A2(n_556),
.B(n_557),
.Y(n_6671)
);

NAND2xp5_ASAP7_75t_L g6672 ( 
.A(n_6314),
.B(n_558),
.Y(n_6672)
);

AOI21x1_ASAP7_75t_L g6673 ( 
.A1(n_6441),
.A2(n_558),
.B(n_559),
.Y(n_6673)
);

INVx1_ASAP7_75t_L g6674 ( 
.A(n_6314),
.Y(n_6674)
);

OA21x2_ASAP7_75t_L g6675 ( 
.A1(n_6332),
.A2(n_558),
.B(n_559),
.Y(n_6675)
);

AND2x2_ASAP7_75t_L g6676 ( 
.A(n_6322),
.B(n_1051),
.Y(n_6676)
);

INVx2_ASAP7_75t_SL g6677 ( 
.A(n_6317),
.Y(n_6677)
);

INVx1_ASAP7_75t_L g6678 ( 
.A(n_6314),
.Y(n_6678)
);

INVx1_ASAP7_75t_L g6679 ( 
.A(n_6314),
.Y(n_6679)
);

NAND2xp5_ASAP7_75t_L g6680 ( 
.A(n_6314),
.B(n_559),
.Y(n_6680)
);

INVxp67_ASAP7_75t_L g6681 ( 
.A(n_6314),
.Y(n_6681)
);

NAND4xp25_ASAP7_75t_L g6682 ( 
.A(n_6314),
.B(n_562),
.C(n_560),
.D(n_561),
.Y(n_6682)
);

HB1xp67_ASAP7_75t_L g6683 ( 
.A(n_6323),
.Y(n_6683)
);

INVx1_ASAP7_75t_L g6684 ( 
.A(n_6314),
.Y(n_6684)
);

BUFx2_ASAP7_75t_L g6685 ( 
.A(n_6314),
.Y(n_6685)
);

AND2x4_ASAP7_75t_L g6686 ( 
.A(n_6317),
.B(n_560),
.Y(n_6686)
);

INVx1_ASAP7_75t_L g6687 ( 
.A(n_6314),
.Y(n_6687)
);

INVx4_ASAP7_75t_L g6688 ( 
.A(n_6353),
.Y(n_6688)
);

NAND3xp33_ASAP7_75t_L g6689 ( 
.A(n_6688),
.B(n_561),
.C(n_562),
.Y(n_6689)
);

AND4x1_ASAP7_75t_L g6690 ( 
.A(n_6517),
.B(n_1054),
.C(n_1055),
.D(n_1053),
.Y(n_6690)
);

AOI221xp5_ASAP7_75t_L g6691 ( 
.A1(n_6490),
.A2(n_563),
.B1(n_561),
.B2(n_562),
.C(n_564),
.Y(n_6691)
);

BUFx3_ASAP7_75t_L g6692 ( 
.A(n_6494),
.Y(n_6692)
);

INVx1_ASAP7_75t_L g6693 ( 
.A(n_6685),
.Y(n_6693)
);

AOI211xp5_ASAP7_75t_L g6694 ( 
.A1(n_6667),
.A2(n_565),
.B(n_563),
.C(n_564),
.Y(n_6694)
);

AND2x2_ASAP7_75t_L g6695 ( 
.A(n_6495),
.B(n_563),
.Y(n_6695)
);

OR2x2_ASAP7_75t_L g6696 ( 
.A(n_6664),
.B(n_564),
.Y(n_6696)
);

AND2x2_ASAP7_75t_L g6697 ( 
.A(n_6677),
.B(n_565),
.Y(n_6697)
);

NOR3xp33_ASAP7_75t_L g6698 ( 
.A(n_6625),
.B(n_567),
.C(n_566),
.Y(n_6698)
);

AOI211xp5_ASAP7_75t_L g6699 ( 
.A1(n_6549),
.A2(n_568),
.B(n_565),
.C(n_567),
.Y(n_6699)
);

OR2x2_ASAP7_75t_L g6700 ( 
.A(n_6670),
.B(n_6659),
.Y(n_6700)
);

OR2x2_ASAP7_75t_L g6701 ( 
.A(n_6488),
.B(n_567),
.Y(n_6701)
);

NAND2xp5_ASAP7_75t_SL g6702 ( 
.A(n_6514),
.B(n_568),
.Y(n_6702)
);

NAND3xp33_ASAP7_75t_SL g6703 ( 
.A(n_6590),
.B(n_568),
.C(n_569),
.Y(n_6703)
);

NOR2xp33_ASAP7_75t_L g6704 ( 
.A(n_6514),
.B(n_569),
.Y(n_6704)
);

NOR3xp33_ASAP7_75t_L g6705 ( 
.A(n_6681),
.B(n_571),
.C(n_570),
.Y(n_6705)
);

NAND3xp33_ASAP7_75t_L g6706 ( 
.A(n_6497),
.B(n_569),
.C(n_570),
.Y(n_6706)
);

NOR3xp33_ASAP7_75t_L g6707 ( 
.A(n_6672),
.B(n_574),
.C(n_573),
.Y(n_6707)
);

AOI221x1_ASAP7_75t_SL g6708 ( 
.A1(n_6660),
.A2(n_574),
.B1(n_572),
.B2(n_573),
.C(n_575),
.Y(n_6708)
);

INVx1_ASAP7_75t_L g6709 ( 
.A(n_6657),
.Y(n_6709)
);

NAND2xp5_ASAP7_75t_L g6710 ( 
.A(n_6529),
.B(n_572),
.Y(n_6710)
);

NAND4xp75_ASAP7_75t_L g6711 ( 
.A(n_6663),
.B(n_582),
.C(n_590),
.D(n_572),
.Y(n_6711)
);

BUFx2_ASAP7_75t_L g6712 ( 
.A(n_6505),
.Y(n_6712)
);

AOI22xp5_ASAP7_75t_L g6713 ( 
.A1(n_6498),
.A2(n_577),
.B1(n_573),
.B2(n_576),
.Y(n_6713)
);

NAND3xp33_ASAP7_75t_L g6714 ( 
.A(n_6497),
.B(n_576),
.C(n_577),
.Y(n_6714)
);

NAND4xp75_ASAP7_75t_L g6715 ( 
.A(n_6665),
.B(n_585),
.C(n_593),
.D(n_576),
.Y(n_6715)
);

AOI22xp33_ASAP7_75t_L g6716 ( 
.A1(n_6602),
.A2(n_580),
.B1(n_578),
.B2(n_579),
.Y(n_6716)
);

OR2x2_ASAP7_75t_L g6717 ( 
.A(n_6668),
.B(n_578),
.Y(n_6717)
);

AOI221xp5_ASAP7_75t_L g6718 ( 
.A1(n_6674),
.A2(n_581),
.B1(n_579),
.B2(n_580),
.C(n_582),
.Y(n_6718)
);

NOR2xp33_ASAP7_75t_L g6719 ( 
.A(n_6514),
.B(n_580),
.Y(n_6719)
);

NAND3xp33_ASAP7_75t_L g6720 ( 
.A(n_6678),
.B(n_581),
.C(n_582),
.Y(n_6720)
);

AND2x2_ASAP7_75t_L g6721 ( 
.A(n_6508),
.B(n_6622),
.Y(n_6721)
);

NAND3xp33_ASAP7_75t_L g6722 ( 
.A(n_6679),
.B(n_581),
.C(n_583),
.Y(n_6722)
);

NAND3xp33_ASAP7_75t_L g6723 ( 
.A(n_6684),
.B(n_583),
.C(n_584),
.Y(n_6723)
);

AOI22xp33_ASAP7_75t_L g6724 ( 
.A1(n_6536),
.A2(n_586),
.B1(n_583),
.B2(n_584),
.Y(n_6724)
);

INVx1_ASAP7_75t_L g6725 ( 
.A(n_6658),
.Y(n_6725)
);

NAND2xp5_ASAP7_75t_L g6726 ( 
.A(n_6529),
.B(n_586),
.Y(n_6726)
);

NAND3xp33_ASAP7_75t_L g6727 ( 
.A(n_6687),
.B(n_586),
.C(n_587),
.Y(n_6727)
);

NAND2xp5_ASAP7_75t_L g6728 ( 
.A(n_6529),
.B(n_587),
.Y(n_6728)
);

AND2x4_ASAP7_75t_L g6729 ( 
.A(n_6566),
.B(n_587),
.Y(n_6729)
);

AND2x2_ASAP7_75t_SL g6730 ( 
.A(n_6662),
.B(n_588),
.Y(n_6730)
);

NAND2xp5_ASAP7_75t_L g6731 ( 
.A(n_6610),
.B(n_588),
.Y(n_6731)
);

NAND4xp75_ASAP7_75t_L g6732 ( 
.A(n_6504),
.B(n_597),
.C(n_605),
.D(n_589),
.Y(n_6732)
);

INVx2_ASAP7_75t_L g6733 ( 
.A(n_6661),
.Y(n_6733)
);

OA211x2_ASAP7_75t_L g6734 ( 
.A1(n_6503),
.A2(n_591),
.B(n_589),
.C(n_590),
.Y(n_6734)
);

NOR3xp33_ASAP7_75t_L g6735 ( 
.A(n_6680),
.B(n_591),
.C(n_590),
.Y(n_6735)
);

OAI211xp5_ASAP7_75t_SL g6736 ( 
.A1(n_6617),
.A2(n_592),
.B(n_589),
.C(n_591),
.Y(n_6736)
);

AO21x2_ASAP7_75t_L g6737 ( 
.A1(n_6519),
.A2(n_592),
.B(n_593),
.Y(n_6737)
);

OAI211xp5_ASAP7_75t_SL g6738 ( 
.A1(n_6510),
.A2(n_595),
.B(n_592),
.C(n_594),
.Y(n_6738)
);

NOR2xp33_ASAP7_75t_L g6739 ( 
.A(n_6547),
.B(n_6635),
.Y(n_6739)
);

INVxp67_ASAP7_75t_L g6740 ( 
.A(n_6676),
.Y(n_6740)
);

AND2x2_ASAP7_75t_L g6741 ( 
.A(n_6491),
.B(n_594),
.Y(n_6741)
);

OAI221xp5_ASAP7_75t_L g6742 ( 
.A1(n_6537),
.A2(n_597),
.B1(n_594),
.B2(n_596),
.C(n_598),
.Y(n_6742)
);

AND2x2_ASAP7_75t_L g6743 ( 
.A(n_6509),
.B(n_596),
.Y(n_6743)
);

NOR3xp33_ASAP7_75t_SL g6744 ( 
.A(n_6511),
.B(n_6682),
.C(n_6501),
.Y(n_6744)
);

NAND2xp5_ASAP7_75t_L g6745 ( 
.A(n_6507),
.B(n_597),
.Y(n_6745)
);

NAND2xp5_ASAP7_75t_L g6746 ( 
.A(n_6666),
.B(n_598),
.Y(n_6746)
);

OAI211xp5_ASAP7_75t_SL g6747 ( 
.A1(n_6535),
.A2(n_601),
.B(n_599),
.C(n_600),
.Y(n_6747)
);

AOI22xp33_ASAP7_75t_L g6748 ( 
.A1(n_6551),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.Y(n_6748)
);

AND2x2_ASAP7_75t_L g6749 ( 
.A(n_6526),
.B(n_6565),
.Y(n_6749)
);

AOI221xp5_ASAP7_75t_L g6750 ( 
.A1(n_6632),
.A2(n_601),
.B1(n_599),
.B2(n_600),
.C(n_602),
.Y(n_6750)
);

NOR3xp33_ASAP7_75t_L g6751 ( 
.A(n_6623),
.B(n_604),
.C(n_603),
.Y(n_6751)
);

NAND3xp33_ASAP7_75t_L g6752 ( 
.A(n_6642),
.B(n_602),
.C(n_604),
.Y(n_6752)
);

AND2x2_ASAP7_75t_L g6753 ( 
.A(n_6493),
.B(n_602),
.Y(n_6753)
);

AND2x2_ASAP7_75t_L g6754 ( 
.A(n_6496),
.B(n_605),
.Y(n_6754)
);

AND2x2_ASAP7_75t_L g6755 ( 
.A(n_6555),
.B(n_605),
.Y(n_6755)
);

AND2x2_ASAP7_75t_L g6756 ( 
.A(n_6620),
.B(n_606),
.Y(n_6756)
);

AOI22xp5_ASAP7_75t_L g6757 ( 
.A1(n_6564),
.A2(n_609),
.B1(n_607),
.B2(n_608),
.Y(n_6757)
);

OR2x2_ASAP7_75t_L g6758 ( 
.A(n_6578),
.B(n_607),
.Y(n_6758)
);

NOR3xp33_ASAP7_75t_L g6759 ( 
.A(n_6643),
.B(n_609),
.C(n_608),
.Y(n_6759)
);

NAND3xp33_ASAP7_75t_L g6760 ( 
.A(n_6645),
.B(n_607),
.C(n_608),
.Y(n_6760)
);

AOI211xp5_ASAP7_75t_L g6761 ( 
.A1(n_6522),
.A2(n_611),
.B(n_609),
.C(n_610),
.Y(n_6761)
);

NAND3xp33_ASAP7_75t_L g6762 ( 
.A(n_6683),
.B(n_6520),
.C(n_6675),
.Y(n_6762)
);

NAND2xp5_ASAP7_75t_SL g6763 ( 
.A(n_6635),
.B(n_610),
.Y(n_6763)
);

NAND3xp33_ASAP7_75t_L g6764 ( 
.A(n_6532),
.B(n_610),
.C(n_611),
.Y(n_6764)
);

NAND3xp33_ASAP7_75t_L g6765 ( 
.A(n_6521),
.B(n_611),
.C(n_612),
.Y(n_6765)
);

NOR3xp33_ASAP7_75t_SL g6766 ( 
.A(n_6500),
.B(n_613),
.C(n_614),
.Y(n_6766)
);

INVx2_ASAP7_75t_L g6767 ( 
.A(n_6528),
.Y(n_6767)
);

AND2x4_ASAP7_75t_L g6768 ( 
.A(n_6566),
.B(n_6489),
.Y(n_6768)
);

NOR3xp33_ASAP7_75t_L g6769 ( 
.A(n_6619),
.B(n_617),
.C(n_616),
.Y(n_6769)
);

INVx1_ASAP7_75t_L g6770 ( 
.A(n_6512),
.Y(n_6770)
);

INVx3_ASAP7_75t_L g6771 ( 
.A(n_6686),
.Y(n_6771)
);

AND2x2_ASAP7_75t_L g6772 ( 
.A(n_6576),
.B(n_615),
.Y(n_6772)
);

INVx1_ASAP7_75t_L g6773 ( 
.A(n_6512),
.Y(n_6773)
);

AND2x2_ASAP7_75t_L g6774 ( 
.A(n_6552),
.B(n_615),
.Y(n_6774)
);

NAND3xp33_ASAP7_75t_L g6775 ( 
.A(n_6541),
.B(n_616),
.C(n_618),
.Y(n_6775)
);

AND2x2_ASAP7_75t_L g6776 ( 
.A(n_6618),
.B(n_616),
.Y(n_6776)
);

INVx1_ASAP7_75t_L g6777 ( 
.A(n_6557),
.Y(n_6777)
);

NOR3xp33_ASAP7_75t_L g6778 ( 
.A(n_6545),
.B(n_620),
.C(n_619),
.Y(n_6778)
);

AO21x2_ASAP7_75t_L g6779 ( 
.A1(n_6673),
.A2(n_618),
.B(n_619),
.Y(n_6779)
);

NAND3xp33_ASAP7_75t_L g6780 ( 
.A(n_6543),
.B(n_618),
.C(n_619),
.Y(n_6780)
);

OR2x2_ASAP7_75t_L g6781 ( 
.A(n_6506),
.B(n_620),
.Y(n_6781)
);

NAND3xp33_ASAP7_75t_L g6782 ( 
.A(n_6544),
.B(n_621),
.C(n_622),
.Y(n_6782)
);

BUFx2_ASAP7_75t_L g6783 ( 
.A(n_6591),
.Y(n_6783)
);

AND2x2_ASAP7_75t_L g6784 ( 
.A(n_6499),
.B(n_621),
.Y(n_6784)
);

NOR3xp33_ASAP7_75t_L g6785 ( 
.A(n_6636),
.B(n_625),
.C(n_624),
.Y(n_6785)
);

NAND2xp5_ASAP7_75t_L g6786 ( 
.A(n_6669),
.B(n_623),
.Y(n_6786)
);

NAND2xp5_ASAP7_75t_L g6787 ( 
.A(n_6639),
.B(n_623),
.Y(n_6787)
);

NAND3xp33_ASAP7_75t_L g6788 ( 
.A(n_6546),
.B(n_6624),
.C(n_6542),
.Y(n_6788)
);

AND2x4_ASAP7_75t_L g6789 ( 
.A(n_6539),
.B(n_623),
.Y(n_6789)
);

NAND2xp5_ASAP7_75t_L g6790 ( 
.A(n_6626),
.B(n_624),
.Y(n_6790)
);

AND2x2_ASAP7_75t_L g6791 ( 
.A(n_6502),
.B(n_624),
.Y(n_6791)
);

NAND3xp33_ASAP7_75t_L g6792 ( 
.A(n_6524),
.B(n_625),
.C(n_626),
.Y(n_6792)
);

NAND2xp5_ASAP7_75t_L g6793 ( 
.A(n_6589),
.B(n_626),
.Y(n_6793)
);

AO21x2_ASAP7_75t_L g6794 ( 
.A1(n_6572),
.A2(n_627),
.B(n_628),
.Y(n_6794)
);

OR2x2_ASAP7_75t_L g6795 ( 
.A(n_6531),
.B(n_627),
.Y(n_6795)
);

HB1xp67_ASAP7_75t_L g6796 ( 
.A(n_6570),
.Y(n_6796)
);

INVx2_ASAP7_75t_L g6797 ( 
.A(n_6562),
.Y(n_6797)
);

NAND2xp5_ASAP7_75t_SL g6798 ( 
.A(n_6607),
.B(n_627),
.Y(n_6798)
);

INVx2_ASAP7_75t_L g6799 ( 
.A(n_6575),
.Y(n_6799)
);

OR2x2_ASAP7_75t_L g6800 ( 
.A(n_6597),
.B(n_6534),
.Y(n_6800)
);

AND2x2_ASAP7_75t_L g6801 ( 
.A(n_6580),
.B(n_628),
.Y(n_6801)
);

NAND2xp5_ASAP7_75t_L g6802 ( 
.A(n_6538),
.B(n_628),
.Y(n_6802)
);

AND2x2_ASAP7_75t_L g6803 ( 
.A(n_6605),
.B(n_629),
.Y(n_6803)
);

NAND2xp5_ASAP7_75t_L g6804 ( 
.A(n_6637),
.B(n_629),
.Y(n_6804)
);

NAND2xp5_ASAP7_75t_L g6805 ( 
.A(n_6579),
.B(n_629),
.Y(n_6805)
);

NAND2xp5_ASAP7_75t_SL g6806 ( 
.A(n_6607),
.B(n_630),
.Y(n_6806)
);

INVx2_ASAP7_75t_L g6807 ( 
.A(n_6584),
.Y(n_6807)
);

AND2x4_ASAP7_75t_L g6808 ( 
.A(n_6621),
.B(n_631),
.Y(n_6808)
);

NOR3xp33_ASAP7_75t_L g6809 ( 
.A(n_6530),
.B(n_633),
.C(n_632),
.Y(n_6809)
);

NOR2x1_ASAP7_75t_SL g6810 ( 
.A(n_6553),
.B(n_631),
.Y(n_6810)
);

AOI221xp5_ASAP7_75t_L g6811 ( 
.A1(n_6556),
.A2(n_634),
.B1(n_631),
.B2(n_632),
.C(n_635),
.Y(n_6811)
);

AND2x2_ASAP7_75t_L g6812 ( 
.A(n_6638),
.B(n_632),
.Y(n_6812)
);

AND2x2_ASAP7_75t_L g6813 ( 
.A(n_6559),
.B(n_634),
.Y(n_6813)
);

NOR3xp33_ASAP7_75t_L g6814 ( 
.A(n_6651),
.B(n_637),
.C(n_636),
.Y(n_6814)
);

NOR3xp33_ASAP7_75t_L g6815 ( 
.A(n_6550),
.B(n_638),
.C(n_636),
.Y(n_6815)
);

AND2x2_ASAP7_75t_L g6816 ( 
.A(n_6558),
.B(n_635),
.Y(n_6816)
);

NAND2xp5_ASAP7_75t_L g6817 ( 
.A(n_6599),
.B(n_636),
.Y(n_6817)
);

INVx1_ASAP7_75t_L g6818 ( 
.A(n_6487),
.Y(n_6818)
);

NOR3xp33_ASAP7_75t_L g6819 ( 
.A(n_6615),
.B(n_640),
.C(n_639),
.Y(n_6819)
);

BUFx3_ASAP7_75t_L g6820 ( 
.A(n_6587),
.Y(n_6820)
);

AOI221xp5_ASAP7_75t_L g6821 ( 
.A1(n_6556),
.A2(n_640),
.B1(n_638),
.B2(n_639),
.C(n_641),
.Y(n_6821)
);

BUFx2_ASAP7_75t_L g6822 ( 
.A(n_6594),
.Y(n_6822)
);

OR2x2_ASAP7_75t_L g6823 ( 
.A(n_6595),
.B(n_6603),
.Y(n_6823)
);

OR2x2_ASAP7_75t_L g6824 ( 
.A(n_6604),
.B(n_638),
.Y(n_6824)
);

NAND4xp25_ASAP7_75t_L g6825 ( 
.A(n_6560),
.B(n_642),
.C(n_640),
.D(n_641),
.Y(n_6825)
);

AOI22xp33_ASAP7_75t_L g6826 ( 
.A1(n_6631),
.A2(n_6609),
.B1(n_6606),
.B2(n_6644),
.Y(n_6826)
);

AND2x2_ASAP7_75t_L g6827 ( 
.A(n_6492),
.B(n_641),
.Y(n_6827)
);

NAND3xp33_ASAP7_75t_L g6828 ( 
.A(n_6574),
.B(n_642),
.C(n_643),
.Y(n_6828)
);

NAND2xp5_ASAP7_75t_L g6829 ( 
.A(n_6650),
.B(n_642),
.Y(n_6829)
);

OR2x2_ASAP7_75t_SL g6830 ( 
.A(n_6611),
.B(n_644),
.Y(n_6830)
);

NAND3xp33_ASAP7_75t_L g6831 ( 
.A(n_6577),
.B(n_644),
.C(n_645),
.Y(n_6831)
);

INVx2_ASAP7_75t_L g6832 ( 
.A(n_6567),
.Y(n_6832)
);

AND2x2_ASAP7_75t_L g6833 ( 
.A(n_6515),
.B(n_644),
.Y(n_6833)
);

AOI22xp33_ASAP7_75t_L g6834 ( 
.A1(n_6582),
.A2(n_647),
.B1(n_645),
.B2(n_646),
.Y(n_6834)
);

AND2x2_ASAP7_75t_L g6835 ( 
.A(n_6646),
.B(n_645),
.Y(n_6835)
);

XOR2x2_ASAP7_75t_L g6836 ( 
.A(n_6571),
.B(n_646),
.Y(n_6836)
);

OAI21xp5_ASAP7_75t_L g6837 ( 
.A1(n_6518),
.A2(n_647),
.B(n_648),
.Y(n_6837)
);

NAND3xp33_ASAP7_75t_L g6838 ( 
.A(n_6540),
.B(n_6601),
.C(n_6513),
.Y(n_6838)
);

BUFx2_ASAP7_75t_L g6839 ( 
.A(n_6613),
.Y(n_6839)
);

AND2x2_ASAP7_75t_L g6840 ( 
.A(n_6516),
.B(n_647),
.Y(n_6840)
);

NOR3xp33_ASAP7_75t_L g6841 ( 
.A(n_6649),
.B(n_651),
.C(n_650),
.Y(n_6841)
);

NAND2xp5_ASAP7_75t_L g6842 ( 
.A(n_6581),
.B(n_649),
.Y(n_6842)
);

NAND3xp33_ASAP7_75t_L g6843 ( 
.A(n_6627),
.B(n_649),
.C(n_651),
.Y(n_6843)
);

NOR2xp33_ASAP7_75t_L g6844 ( 
.A(n_6600),
.B(n_649),
.Y(n_6844)
);

AND2x2_ASAP7_75t_L g6845 ( 
.A(n_6640),
.B(n_652),
.Y(n_6845)
);

INVx1_ASAP7_75t_L g6846 ( 
.A(n_6554),
.Y(n_6846)
);

OR2x2_ASAP7_75t_L g6847 ( 
.A(n_6569),
.B(n_6628),
.Y(n_6847)
);

OR2x2_ASAP7_75t_L g6848 ( 
.A(n_6593),
.B(n_6629),
.Y(n_6848)
);

AOI22xp5_ASAP7_75t_L g6849 ( 
.A1(n_6647),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.Y(n_6849)
);

AOI221xp5_ASAP7_75t_L g6850 ( 
.A1(n_6563),
.A2(n_654),
.B1(n_652),
.B2(n_653),
.C(n_655),
.Y(n_6850)
);

INVx2_ASAP7_75t_SL g6851 ( 
.A(n_6561),
.Y(n_6851)
);

AOI221xp5_ASAP7_75t_L g6852 ( 
.A1(n_6592),
.A2(n_6588),
.B1(n_6586),
.B2(n_6527),
.C(n_6648),
.Y(n_6852)
);

NOR3xp33_ASAP7_75t_L g6853 ( 
.A(n_6598),
.B(n_656),
.C(n_655),
.Y(n_6853)
);

OR2x2_ASAP7_75t_L g6854 ( 
.A(n_6671),
.B(n_653),
.Y(n_6854)
);

HB1xp67_ASAP7_75t_L g6855 ( 
.A(n_6533),
.Y(n_6855)
);

INVx1_ASAP7_75t_SL g6856 ( 
.A(n_6692),
.Y(n_6856)
);

AND2x2_ASAP7_75t_L g6857 ( 
.A(n_6851),
.B(n_6653),
.Y(n_6857)
);

BUFx2_ASAP7_75t_L g6858 ( 
.A(n_6721),
.Y(n_6858)
);

NAND2xp5_ASAP7_75t_L g6859 ( 
.A(n_6729),
.B(n_6633),
.Y(n_6859)
);

INVx2_ASAP7_75t_L g6860 ( 
.A(n_6820),
.Y(n_6860)
);

INVx1_ASAP7_75t_SL g6861 ( 
.A(n_6697),
.Y(n_6861)
);

OR2x2_ASAP7_75t_L g6862 ( 
.A(n_6823),
.B(n_6573),
.Y(n_6862)
);

INVx1_ASAP7_75t_L g6863 ( 
.A(n_6770),
.Y(n_6863)
);

NAND2xp5_ASAP7_75t_L g6864 ( 
.A(n_6729),
.B(n_6633),
.Y(n_6864)
);

NOR3xp33_ASAP7_75t_SL g6865 ( 
.A(n_6703),
.B(n_6739),
.C(n_6762),
.Y(n_6865)
);

INVx1_ASAP7_75t_L g6866 ( 
.A(n_6773),
.Y(n_6866)
);

OR2x2_ASAP7_75t_L g6867 ( 
.A(n_6710),
.B(n_6655),
.Y(n_6867)
);

AND2x4_ASAP7_75t_L g6868 ( 
.A(n_6767),
.B(n_6614),
.Y(n_6868)
);

AND2x2_ASAP7_75t_L g6869 ( 
.A(n_6839),
.B(n_6634),
.Y(n_6869)
);

NAND2xp5_ASAP7_75t_L g6870 ( 
.A(n_6730),
.B(n_6548),
.Y(n_6870)
);

OAI211xp5_ASAP7_75t_SL g6871 ( 
.A1(n_6693),
.A2(n_6608),
.B(n_6654),
.C(n_6641),
.Y(n_6871)
);

NOR2x1_ASAP7_75t_R g6872 ( 
.A(n_6731),
.B(n_6652),
.Y(n_6872)
);

NOR2xp33_ASAP7_75t_L g6873 ( 
.A(n_6783),
.B(n_6596),
.Y(n_6873)
);

INVx1_ASAP7_75t_L g6874 ( 
.A(n_6695),
.Y(n_6874)
);

INVx2_ASAP7_75t_L g6875 ( 
.A(n_6712),
.Y(n_6875)
);

OAI31xp33_ASAP7_75t_L g6876 ( 
.A1(n_6838),
.A2(n_6818),
.A3(n_6736),
.B(n_6768),
.Y(n_6876)
);

NAND2xp5_ASAP7_75t_L g6877 ( 
.A(n_6808),
.B(n_6755),
.Y(n_6877)
);

NOR3xp33_ASAP7_75t_L g6878 ( 
.A(n_6702),
.B(n_6568),
.C(n_6585),
.Y(n_6878)
);

INVx1_ASAP7_75t_L g6879 ( 
.A(n_6774),
.Y(n_6879)
);

AND2x2_ASAP7_75t_L g6880 ( 
.A(n_6741),
.B(n_6656),
.Y(n_6880)
);

INVx1_ASAP7_75t_L g6881 ( 
.A(n_6801),
.Y(n_6881)
);

OAI33xp33_ASAP7_75t_L g6882 ( 
.A1(n_6777),
.A2(n_6616),
.A3(n_6525),
.B1(n_6630),
.B2(n_6523),
.B3(n_6612),
.Y(n_6882)
);

AND2x2_ASAP7_75t_L g6883 ( 
.A(n_6768),
.B(n_6583),
.Y(n_6883)
);

OR2x2_ASAP7_75t_L g6884 ( 
.A(n_6726),
.B(n_655),
.Y(n_6884)
);

AND2x2_ASAP7_75t_L g6885 ( 
.A(n_6756),
.B(n_6772),
.Y(n_6885)
);

INVx2_ASAP7_75t_SL g6886 ( 
.A(n_6797),
.Y(n_6886)
);

NAND2xp5_ASAP7_75t_L g6887 ( 
.A(n_6808),
.B(n_656),
.Y(n_6887)
);

OAI221xp5_ASAP7_75t_L g6888 ( 
.A1(n_6837),
.A2(n_658),
.B1(n_656),
.B2(n_657),
.C(n_659),
.Y(n_6888)
);

OAI31xp33_ASAP7_75t_L g6889 ( 
.A1(n_6788),
.A2(n_6855),
.A3(n_6719),
.B(n_6704),
.Y(n_6889)
);

NOR2x1_ASAP7_75t_L g6890 ( 
.A(n_6737),
.B(n_657),
.Y(n_6890)
);

INVx3_ASAP7_75t_L g6891 ( 
.A(n_6789),
.Y(n_6891)
);

INVx2_ASAP7_75t_L g6892 ( 
.A(n_6789),
.Y(n_6892)
);

OAI22xp33_ASAP7_75t_L g6893 ( 
.A1(n_6804),
.A2(n_660),
.B1(n_658),
.B2(n_659),
.Y(n_6893)
);

NOR4xp25_ASAP7_75t_L g6894 ( 
.A(n_6852),
.B(n_662),
.C(n_658),
.D(n_661),
.Y(n_6894)
);

NAND2xp5_ASAP7_75t_L g6895 ( 
.A(n_6803),
.B(n_661),
.Y(n_6895)
);

INVx1_ASAP7_75t_L g6896 ( 
.A(n_6822),
.Y(n_6896)
);

AND2x4_ASAP7_75t_L g6897 ( 
.A(n_6832),
.B(n_662),
.Y(n_6897)
);

AOI221xp5_ASAP7_75t_L g6898 ( 
.A1(n_6750),
.A2(n_665),
.B1(n_662),
.B2(n_664),
.C(n_666),
.Y(n_6898)
);

INVx2_ASAP7_75t_L g6899 ( 
.A(n_6771),
.Y(n_6899)
);

OAI31xp33_ASAP7_75t_L g6900 ( 
.A1(n_6843),
.A2(n_666),
.A3(n_664),
.B(n_665),
.Y(n_6900)
);

AND2x2_ASAP7_75t_L g6901 ( 
.A(n_6753),
.B(n_664),
.Y(n_6901)
);

NAND2xp5_ASAP7_75t_SL g6902 ( 
.A(n_6811),
.B(n_666),
.Y(n_6902)
);

BUFx3_ASAP7_75t_L g6903 ( 
.A(n_6799),
.Y(n_6903)
);

HB1xp67_ASAP7_75t_L g6904 ( 
.A(n_6807),
.Y(n_6904)
);

INVx1_ASAP7_75t_L g6905 ( 
.A(n_6754),
.Y(n_6905)
);

INVx4_ASAP7_75t_L g6906 ( 
.A(n_6795),
.Y(n_6906)
);

NAND2x1_ASAP7_75t_SL g6907 ( 
.A(n_6743),
.B(n_667),
.Y(n_6907)
);

OAI31xp33_ASAP7_75t_L g6908 ( 
.A1(n_6785),
.A2(n_669),
.A3(n_667),
.B(n_668),
.Y(n_6908)
);

OA332x1_ASAP7_75t_L g6909 ( 
.A1(n_6744),
.A2(n_1076),
.A3(n_673),
.B1(n_670),
.B2(n_674),
.B3(n_672),
.C1(n_667),
.C2(n_668),
.Y(n_6909)
);

INVx2_ASAP7_75t_L g6910 ( 
.A(n_6810),
.Y(n_6910)
);

INVx1_ASAP7_75t_L g6911 ( 
.A(n_6700),
.Y(n_6911)
);

AND2x2_ASAP7_75t_L g6912 ( 
.A(n_6813),
.B(n_668),
.Y(n_6912)
);

OR2x2_ASAP7_75t_L g6913 ( 
.A(n_6728),
.B(n_670),
.Y(n_6913)
);

OAI31xp33_ASAP7_75t_L g6914 ( 
.A1(n_6747),
.A2(n_672),
.A3(n_670),
.B(n_671),
.Y(n_6914)
);

INVx1_ASAP7_75t_L g6915 ( 
.A(n_6854),
.Y(n_6915)
);

NOR2xp33_ASAP7_75t_L g6916 ( 
.A(n_6740),
.B(n_6830),
.Y(n_6916)
);

AND2x4_ASAP7_75t_SL g6917 ( 
.A(n_6749),
.B(n_671),
.Y(n_6917)
);

INVx2_ASAP7_75t_L g6918 ( 
.A(n_6758),
.Y(n_6918)
);

HB1xp67_ASAP7_75t_L g6919 ( 
.A(n_6711),
.Y(n_6919)
);

INVx2_ASAP7_75t_L g6920 ( 
.A(n_6781),
.Y(n_6920)
);

BUFx2_ASAP7_75t_L g6921 ( 
.A(n_6776),
.Y(n_6921)
);

INVx1_ASAP7_75t_L g6922 ( 
.A(n_6800),
.Y(n_6922)
);

OAI32xp33_ASAP7_75t_L g6923 ( 
.A1(n_6848),
.A2(n_673),
.A3(n_671),
.B1(n_672),
.B2(n_674),
.Y(n_6923)
);

OAI221xp5_ASAP7_75t_L g6924 ( 
.A1(n_6821),
.A2(n_676),
.B1(n_673),
.B2(n_675),
.C(n_677),
.Y(n_6924)
);

INVx1_ASAP7_75t_L g6925 ( 
.A(n_6784),
.Y(n_6925)
);

AOI322xp5_ASAP7_75t_L g6926 ( 
.A1(n_6826),
.A2(n_680),
.A3(n_679),
.B1(n_677),
.B2(n_675),
.C1(n_676),
.C2(n_678),
.Y(n_6926)
);

AND2x2_ASAP7_75t_L g6927 ( 
.A(n_6827),
.B(n_675),
.Y(n_6927)
);

AND2x2_ASAP7_75t_L g6928 ( 
.A(n_6833),
.B(n_6816),
.Y(n_6928)
);

INVx1_ASAP7_75t_L g6929 ( 
.A(n_6791),
.Y(n_6929)
);

INVx1_ASAP7_75t_L g6930 ( 
.A(n_6696),
.Y(n_6930)
);

INVx1_ASAP7_75t_L g6931 ( 
.A(n_6787),
.Y(n_6931)
);

INVx1_ASAP7_75t_L g6932 ( 
.A(n_6790),
.Y(n_6932)
);

HB1xp67_ASAP7_75t_L g6933 ( 
.A(n_6715),
.Y(n_6933)
);

AND2x2_ASAP7_75t_L g6934 ( 
.A(n_6835),
.B(n_676),
.Y(n_6934)
);

HB1xp67_ASAP7_75t_L g6935 ( 
.A(n_6732),
.Y(n_6935)
);

INVx1_ASAP7_75t_L g6936 ( 
.A(n_6812),
.Y(n_6936)
);

NAND2xp5_ASAP7_75t_L g6937 ( 
.A(n_6708),
.B(n_677),
.Y(n_6937)
);

NAND2xp5_ASAP7_75t_L g6938 ( 
.A(n_6809),
.B(n_6691),
.Y(n_6938)
);

AOI211xp5_ASAP7_75t_L g6939 ( 
.A1(n_6769),
.A2(n_680),
.B(n_678),
.C(n_679),
.Y(n_6939)
);

INVx1_ASAP7_75t_L g6940 ( 
.A(n_6701),
.Y(n_6940)
);

INVx1_ASAP7_75t_L g6941 ( 
.A(n_6717),
.Y(n_6941)
);

INVx2_ASAP7_75t_L g6942 ( 
.A(n_6824),
.Y(n_6942)
);

AND2x4_ASAP7_75t_L g6943 ( 
.A(n_6733),
.B(n_678),
.Y(n_6943)
);

OAI22xp33_ASAP7_75t_L g6944 ( 
.A1(n_6793),
.A2(n_681),
.B1(n_679),
.B2(n_680),
.Y(n_6944)
);

OAI21xp33_ASAP7_75t_L g6945 ( 
.A1(n_6709),
.A2(n_681),
.B(n_682),
.Y(n_6945)
);

AND2x2_ASAP7_75t_L g6946 ( 
.A(n_6840),
.B(n_682),
.Y(n_6946)
);

INVx3_ASAP7_75t_L g6947 ( 
.A(n_6690),
.Y(n_6947)
);

NAND2xp5_ASAP7_75t_L g6948 ( 
.A(n_6694),
.B(n_6779),
.Y(n_6948)
);

BUFx3_ASAP7_75t_L g6949 ( 
.A(n_6745),
.Y(n_6949)
);

AND2x2_ASAP7_75t_L g6950 ( 
.A(n_6845),
.B(n_682),
.Y(n_6950)
);

NAND3xp33_ASAP7_75t_L g6951 ( 
.A(n_6699),
.B(n_683),
.C(n_684),
.Y(n_6951)
);

AND2x2_ASAP7_75t_L g6952 ( 
.A(n_6796),
.B(n_683),
.Y(n_6952)
);

CKINVDCx16_ASAP7_75t_R g6953 ( 
.A(n_6757),
.Y(n_6953)
);

OAI33xp33_ASAP7_75t_L g6954 ( 
.A1(n_6725),
.A2(n_686),
.A3(n_688),
.B1(n_684),
.B2(n_685),
.B3(n_687),
.Y(n_6954)
);

INVx1_ASAP7_75t_L g6955 ( 
.A(n_6752),
.Y(n_6955)
);

NOR3xp33_ASAP7_75t_SL g6956 ( 
.A(n_6689),
.B(n_1068),
.C(n_685),
.Y(n_6956)
);

INVx2_ASAP7_75t_SL g6957 ( 
.A(n_6836),
.Y(n_6957)
);

AOI22xp5_ASAP7_75t_L g6958 ( 
.A1(n_6759),
.A2(n_687),
.B1(n_685),
.B2(n_686),
.Y(n_6958)
);

INVx1_ASAP7_75t_SL g6959 ( 
.A(n_6805),
.Y(n_6959)
);

HB1xp67_ASAP7_75t_L g6960 ( 
.A(n_6817),
.Y(n_6960)
);

INVx1_ASAP7_75t_SL g6961 ( 
.A(n_6829),
.Y(n_6961)
);

INVx1_ASAP7_75t_SL g6962 ( 
.A(n_6763),
.Y(n_6962)
);

AOI211xp5_ASAP7_75t_L g6963 ( 
.A1(n_6844),
.A2(n_690),
.B(n_688),
.C(n_689),
.Y(n_6963)
);

AND2x2_ASAP7_75t_L g6964 ( 
.A(n_6846),
.B(n_689),
.Y(n_6964)
);

OR2x2_ASAP7_75t_L g6965 ( 
.A(n_6746),
.B(n_689),
.Y(n_6965)
);

INVx1_ASAP7_75t_L g6966 ( 
.A(n_6760),
.Y(n_6966)
);

NAND2xp5_ASAP7_75t_L g6967 ( 
.A(n_6698),
.B(n_690),
.Y(n_6967)
);

INVx1_ASAP7_75t_L g6968 ( 
.A(n_6794),
.Y(n_6968)
);

INVx1_ASAP7_75t_L g6969 ( 
.A(n_6842),
.Y(n_6969)
);

OAI31xp33_ASAP7_75t_SL g6970 ( 
.A1(n_6765),
.A2(n_693),
.A3(n_691),
.B(n_692),
.Y(n_6970)
);

AND2x4_ASAP7_75t_L g6971 ( 
.A(n_6706),
.B(n_691),
.Y(n_6971)
);

AOI22xp33_ASAP7_75t_L g6972 ( 
.A1(n_6734),
.A2(n_693),
.B1(n_691),
.B2(n_692),
.Y(n_6972)
);

INVx3_ASAP7_75t_L g6973 ( 
.A(n_6847),
.Y(n_6973)
);

NAND4xp25_ASAP7_75t_L g6974 ( 
.A(n_6761),
.B(n_694),
.C(n_692),
.D(n_693),
.Y(n_6974)
);

NOR3xp33_ASAP7_75t_L g6975 ( 
.A(n_6764),
.B(n_694),
.C(n_695),
.Y(n_6975)
);

AND2x2_ASAP7_75t_L g6976 ( 
.A(n_6766),
.B(n_694),
.Y(n_6976)
);

INVx1_ASAP7_75t_L g6977 ( 
.A(n_6714),
.Y(n_6977)
);

OR2x2_ASAP7_75t_L g6978 ( 
.A(n_6786),
.B(n_6802),
.Y(n_6978)
);

BUFx3_ASAP7_75t_L g6979 ( 
.A(n_6828),
.Y(n_6979)
);

OAI31xp33_ASAP7_75t_L g6980 ( 
.A1(n_6738),
.A2(n_6831),
.A3(n_6720),
.B(n_6723),
.Y(n_6980)
);

NAND3xp33_ASAP7_75t_L g6981 ( 
.A(n_6705),
.B(n_695),
.C(n_696),
.Y(n_6981)
);

AOI33xp33_ASAP7_75t_L g6982 ( 
.A1(n_6716),
.A2(n_6748),
.A3(n_6724),
.B1(n_6834),
.B2(n_6718),
.B3(n_6850),
.Y(n_6982)
);

INVx2_ASAP7_75t_L g6983 ( 
.A(n_6798),
.Y(n_6983)
);

INVx1_ASAP7_75t_L g6984 ( 
.A(n_6713),
.Y(n_6984)
);

BUFx2_ASAP7_75t_L g6985 ( 
.A(n_6849),
.Y(n_6985)
);

INVx1_ASAP7_75t_L g6986 ( 
.A(n_6806),
.Y(n_6986)
);

OR2x2_ASAP7_75t_L g6987 ( 
.A(n_6722),
.B(n_696),
.Y(n_6987)
);

AND2x2_ASAP7_75t_L g6988 ( 
.A(n_6853),
.B(n_696),
.Y(n_6988)
);

AND2x2_ASAP7_75t_L g6989 ( 
.A(n_6841),
.B(n_697),
.Y(n_6989)
);

INVx1_ASAP7_75t_SL g6990 ( 
.A(n_6727),
.Y(n_6990)
);

AOI221xp5_ASAP7_75t_L g6991 ( 
.A1(n_6819),
.A2(n_699),
.B1(n_697),
.B2(n_698),
.C(n_700),
.Y(n_6991)
);

OAI33xp33_ASAP7_75t_L g6992 ( 
.A1(n_6825),
.A2(n_700),
.A3(n_702),
.B1(n_698),
.B2(n_699),
.B3(n_701),
.Y(n_6992)
);

AND2x2_ASAP7_75t_L g6993 ( 
.A(n_6707),
.B(n_698),
.Y(n_6993)
);

INVx2_ASAP7_75t_L g6994 ( 
.A(n_6775),
.Y(n_6994)
);

AND2x2_ASAP7_75t_L g6995 ( 
.A(n_6735),
.B(n_6778),
.Y(n_6995)
);

NAND2xp5_ASAP7_75t_L g6996 ( 
.A(n_6751),
.B(n_699),
.Y(n_6996)
);

AND2x2_ASAP7_75t_L g6997 ( 
.A(n_6814),
.B(n_700),
.Y(n_6997)
);

HB1xp67_ASAP7_75t_L g6998 ( 
.A(n_6780),
.Y(n_6998)
);

NAND2xp5_ASAP7_75t_L g6999 ( 
.A(n_6815),
.B(n_701),
.Y(n_6999)
);

AND2x2_ASAP7_75t_L g7000 ( 
.A(n_6782),
.B(n_701),
.Y(n_7000)
);

INVx1_ASAP7_75t_L g7001 ( 
.A(n_6792),
.Y(n_7001)
);

AOI22xp5_ASAP7_75t_L g7002 ( 
.A1(n_6742),
.A2(n_1067),
.B1(n_704),
.B2(n_702),
.Y(n_7002)
);

NAND2xp5_ASAP7_75t_L g7003 ( 
.A(n_6692),
.B(n_702),
.Y(n_7003)
);

AND2x2_ASAP7_75t_L g7004 ( 
.A(n_6851),
.B(n_703),
.Y(n_7004)
);

OAI33xp33_ASAP7_75t_L g7005 ( 
.A1(n_6693),
.A2(n_705),
.A3(n_707),
.B1(n_703),
.B2(n_704),
.B3(n_706),
.Y(n_7005)
);

INVx2_ASAP7_75t_L g7006 ( 
.A(n_6692),
.Y(n_7006)
);

BUFx3_ASAP7_75t_L g7007 ( 
.A(n_6692),
.Y(n_7007)
);

NAND2x1_ASAP7_75t_SL g7008 ( 
.A(n_6721),
.B(n_703),
.Y(n_7008)
);

INVx1_ASAP7_75t_L g7009 ( 
.A(n_6770),
.Y(n_7009)
);

NOR2xp33_ASAP7_75t_L g7010 ( 
.A(n_6851),
.B(n_705),
.Y(n_7010)
);

INVx1_ASAP7_75t_L g7011 ( 
.A(n_6770),
.Y(n_7011)
);

INVx1_ASAP7_75t_SL g7012 ( 
.A(n_6692),
.Y(n_7012)
);

INVx1_ASAP7_75t_L g7013 ( 
.A(n_6770),
.Y(n_7013)
);

AND2x2_ASAP7_75t_L g7014 ( 
.A(n_6851),
.B(n_706),
.Y(n_7014)
);

INVx2_ASAP7_75t_SL g7015 ( 
.A(n_6692),
.Y(n_7015)
);

INVx1_ASAP7_75t_L g7016 ( 
.A(n_6770),
.Y(n_7016)
);

INVx1_ASAP7_75t_L g7017 ( 
.A(n_6770),
.Y(n_7017)
);

NAND3xp33_ASAP7_75t_L g7018 ( 
.A(n_6851),
.B(n_706),
.C(n_707),
.Y(n_7018)
);

INVx4_ASAP7_75t_L g7019 ( 
.A(n_6692),
.Y(n_7019)
);

INVx1_ASAP7_75t_L g7020 ( 
.A(n_6770),
.Y(n_7020)
);

OAI22xp5_ASAP7_75t_L g7021 ( 
.A1(n_6851),
.A2(n_710),
.B1(n_708),
.B2(n_709),
.Y(n_7021)
);

INVx1_ASAP7_75t_L g7022 ( 
.A(n_6770),
.Y(n_7022)
);

AND2x2_ASAP7_75t_L g7023 ( 
.A(n_6851),
.B(n_708),
.Y(n_7023)
);

INVx1_ASAP7_75t_L g7024 ( 
.A(n_6770),
.Y(n_7024)
);

OR2x2_ASAP7_75t_L g7025 ( 
.A(n_6692),
.B(n_708),
.Y(n_7025)
);

OAI32xp33_ASAP7_75t_L g7026 ( 
.A1(n_6770),
.A2(n_712),
.A3(n_710),
.B1(n_711),
.B2(n_713),
.Y(n_7026)
);

INVx1_ASAP7_75t_L g7027 ( 
.A(n_6770),
.Y(n_7027)
);

INVx2_ASAP7_75t_L g7028 ( 
.A(n_7007),
.Y(n_7028)
);

INVx1_ASAP7_75t_L g7029 ( 
.A(n_6863),
.Y(n_7029)
);

INVx1_ASAP7_75t_L g7030 ( 
.A(n_6866),
.Y(n_7030)
);

NAND2xp5_ASAP7_75t_L g7031 ( 
.A(n_6856),
.B(n_710),
.Y(n_7031)
);

NAND2xp5_ASAP7_75t_L g7032 ( 
.A(n_7012),
.B(n_711),
.Y(n_7032)
);

AND2x2_ASAP7_75t_L g7033 ( 
.A(n_7019),
.B(n_712),
.Y(n_7033)
);

INVx1_ASAP7_75t_L g7034 ( 
.A(n_7009),
.Y(n_7034)
);

INVx3_ASAP7_75t_L g7035 ( 
.A(n_7006),
.Y(n_7035)
);

AND2x2_ASAP7_75t_L g7036 ( 
.A(n_6858),
.B(n_712),
.Y(n_7036)
);

OR2x2_ASAP7_75t_L g7037 ( 
.A(n_7015),
.B(n_7003),
.Y(n_7037)
);

AND2x2_ASAP7_75t_L g7038 ( 
.A(n_6869),
.B(n_713),
.Y(n_7038)
);

OAI33xp33_ASAP7_75t_L g7039 ( 
.A1(n_7011),
.A2(n_715),
.A3(n_717),
.B1(n_713),
.B2(n_714),
.B3(n_716),
.Y(n_7039)
);

AND2x2_ASAP7_75t_L g7040 ( 
.A(n_7004),
.B(n_714),
.Y(n_7040)
);

OR2x2_ASAP7_75t_L g7041 ( 
.A(n_6860),
.B(n_715),
.Y(n_7041)
);

INVx2_ASAP7_75t_SL g7042 ( 
.A(n_6903),
.Y(n_7042)
);

INVx2_ASAP7_75t_L g7043 ( 
.A(n_6897),
.Y(n_7043)
);

INVx1_ASAP7_75t_L g7044 ( 
.A(n_7013),
.Y(n_7044)
);

INVx1_ASAP7_75t_L g7045 ( 
.A(n_7016),
.Y(n_7045)
);

AND2x2_ASAP7_75t_L g7046 ( 
.A(n_7014),
.B(n_716),
.Y(n_7046)
);

INVx1_ASAP7_75t_L g7047 ( 
.A(n_7017),
.Y(n_7047)
);

NOR2xp33_ASAP7_75t_L g7048 ( 
.A(n_6910),
.B(n_716),
.Y(n_7048)
);

AND2x2_ASAP7_75t_L g7049 ( 
.A(n_7023),
.B(n_717),
.Y(n_7049)
);

INVx1_ASAP7_75t_L g7050 ( 
.A(n_7020),
.Y(n_7050)
);

INVx2_ASAP7_75t_SL g7051 ( 
.A(n_6868),
.Y(n_7051)
);

OR2x2_ASAP7_75t_L g7052 ( 
.A(n_7025),
.B(n_717),
.Y(n_7052)
);

NAND2xp5_ASAP7_75t_SL g7053 ( 
.A(n_6876),
.B(n_718),
.Y(n_7053)
);

INVx2_ASAP7_75t_SL g7054 ( 
.A(n_6868),
.Y(n_7054)
);

INVx1_ASAP7_75t_L g7055 ( 
.A(n_7022),
.Y(n_7055)
);

AND2x2_ASAP7_75t_L g7056 ( 
.A(n_6857),
.B(n_718),
.Y(n_7056)
);

NAND2xp5_ASAP7_75t_L g7057 ( 
.A(n_6897),
.B(n_6972),
.Y(n_7057)
);

BUFx2_ASAP7_75t_L g7058 ( 
.A(n_7008),
.Y(n_7058)
);

INVx1_ASAP7_75t_L g7059 ( 
.A(n_7024),
.Y(n_7059)
);

AND2x2_ASAP7_75t_L g7060 ( 
.A(n_6976),
.B(n_719),
.Y(n_7060)
);

NAND2xp5_ASAP7_75t_L g7061 ( 
.A(n_6926),
.B(n_719),
.Y(n_7061)
);

OAI22xp5_ASAP7_75t_L g7062 ( 
.A1(n_7018),
.A2(n_722),
.B1(n_720),
.B2(n_721),
.Y(n_7062)
);

AND2x2_ASAP7_75t_L g7063 ( 
.A(n_6883),
.B(n_6885),
.Y(n_7063)
);

INVxp67_ASAP7_75t_L g7064 ( 
.A(n_7010),
.Y(n_7064)
);

AND2x2_ASAP7_75t_L g7065 ( 
.A(n_6901),
.B(n_720),
.Y(n_7065)
);

NAND2xp5_ASAP7_75t_L g7066 ( 
.A(n_6886),
.B(n_721),
.Y(n_7066)
);

NOR2xp33_ASAP7_75t_L g7067 ( 
.A(n_6882),
.B(n_721),
.Y(n_7067)
);

OAI22xp5_ASAP7_75t_L g7068 ( 
.A1(n_6875),
.A2(n_724),
.B1(n_722),
.B2(n_723),
.Y(n_7068)
);

HB1xp67_ASAP7_75t_L g7069 ( 
.A(n_6904),
.Y(n_7069)
);

INVx1_ASAP7_75t_L g7070 ( 
.A(n_7027),
.Y(n_7070)
);

AND2x2_ASAP7_75t_L g7071 ( 
.A(n_6912),
.B(n_722),
.Y(n_7071)
);

NAND2xp5_ASAP7_75t_L g7072 ( 
.A(n_6947),
.B(n_723),
.Y(n_7072)
);

INVx2_ASAP7_75t_L g7073 ( 
.A(n_6899),
.Y(n_7073)
);

HB1xp67_ASAP7_75t_L g7074 ( 
.A(n_7021),
.Y(n_7074)
);

INVx1_ASAP7_75t_L g7075 ( 
.A(n_6887),
.Y(n_7075)
);

OR2x2_ASAP7_75t_L g7076 ( 
.A(n_6877),
.B(n_724),
.Y(n_7076)
);

INVx1_ASAP7_75t_L g7077 ( 
.A(n_6862),
.Y(n_7077)
);

INVx1_ASAP7_75t_L g7078 ( 
.A(n_6987),
.Y(n_7078)
);

AND2x4_ASAP7_75t_L g7079 ( 
.A(n_6896),
.B(n_724),
.Y(n_7079)
);

INVx1_ASAP7_75t_SL g7080 ( 
.A(n_6917),
.Y(n_7080)
);

INVx2_ASAP7_75t_L g7081 ( 
.A(n_6891),
.Y(n_7081)
);

AND2x2_ASAP7_75t_L g7082 ( 
.A(n_6928),
.B(n_725),
.Y(n_7082)
);

INVx1_ASAP7_75t_L g7083 ( 
.A(n_6943),
.Y(n_7083)
);

NOR2xp33_ASAP7_75t_L g7084 ( 
.A(n_6954),
.B(n_7005),
.Y(n_7084)
);

INVxp67_ASAP7_75t_SL g7085 ( 
.A(n_6895),
.Y(n_7085)
);

INVx2_ASAP7_75t_L g7086 ( 
.A(n_6892),
.Y(n_7086)
);

OR2x2_ASAP7_75t_L g7087 ( 
.A(n_6859),
.B(n_725),
.Y(n_7087)
);

AND2x2_ASAP7_75t_L g7088 ( 
.A(n_6880),
.B(n_6927),
.Y(n_7088)
);

NAND2xp5_ASAP7_75t_L g7089 ( 
.A(n_6934),
.B(n_725),
.Y(n_7089)
);

AND2x2_ASAP7_75t_L g7090 ( 
.A(n_6946),
.B(n_726),
.Y(n_7090)
);

INVx1_ASAP7_75t_SL g7091 ( 
.A(n_6943),
.Y(n_7091)
);

OR2x2_ASAP7_75t_L g7092 ( 
.A(n_6864),
.B(n_726),
.Y(n_7092)
);

OAI21xp33_ASAP7_75t_L g7093 ( 
.A1(n_6982),
.A2(n_726),
.B(n_727),
.Y(n_7093)
);

AND2x2_ASAP7_75t_L g7094 ( 
.A(n_6950),
.B(n_727),
.Y(n_7094)
);

INVx2_ASAP7_75t_L g7095 ( 
.A(n_6911),
.Y(n_7095)
);

NAND2xp5_ASAP7_75t_L g7096 ( 
.A(n_6894),
.B(n_727),
.Y(n_7096)
);

AND2x2_ASAP7_75t_L g7097 ( 
.A(n_6952),
.B(n_728),
.Y(n_7097)
);

INVx2_ASAP7_75t_L g7098 ( 
.A(n_6971),
.Y(n_7098)
);

AND2x2_ASAP7_75t_L g7099 ( 
.A(n_6964),
.B(n_728),
.Y(n_7099)
);

NOR2xp33_ASAP7_75t_L g7100 ( 
.A(n_6871),
.B(n_7026),
.Y(n_7100)
);

INVx2_ASAP7_75t_L g7101 ( 
.A(n_6971),
.Y(n_7101)
);

AND2x2_ASAP7_75t_L g7102 ( 
.A(n_6865),
.B(n_729),
.Y(n_7102)
);

INVxp33_ASAP7_75t_SL g7103 ( 
.A(n_6919),
.Y(n_7103)
);

INVx2_ASAP7_75t_L g7104 ( 
.A(n_6918),
.Y(n_7104)
);

INVx2_ASAP7_75t_L g7105 ( 
.A(n_6920),
.Y(n_7105)
);

AND3x1_ASAP7_75t_L g7106 ( 
.A(n_6956),
.B(n_729),
.C(n_730),
.Y(n_7106)
);

INVx1_ASAP7_75t_L g7107 ( 
.A(n_6965),
.Y(n_7107)
);

AND2x2_ASAP7_75t_SL g7108 ( 
.A(n_6933),
.B(n_6935),
.Y(n_7108)
);

INVx1_ASAP7_75t_L g7109 ( 
.A(n_6922),
.Y(n_7109)
);

INVx1_ASAP7_75t_L g7110 ( 
.A(n_7000),
.Y(n_7110)
);

INVx1_ASAP7_75t_L g7111 ( 
.A(n_6921),
.Y(n_7111)
);

AND2x2_ASAP7_75t_L g7112 ( 
.A(n_6997),
.B(n_729),
.Y(n_7112)
);

OR2x2_ASAP7_75t_L g7113 ( 
.A(n_6996),
.B(n_730),
.Y(n_7113)
);

AND2x2_ASAP7_75t_L g7114 ( 
.A(n_6957),
.B(n_730),
.Y(n_7114)
);

OR2x2_ASAP7_75t_L g7115 ( 
.A(n_6861),
.B(n_731),
.Y(n_7115)
);

OR2x2_ASAP7_75t_L g7116 ( 
.A(n_6999),
.B(n_731),
.Y(n_7116)
);

INVx1_ASAP7_75t_L g7117 ( 
.A(n_6884),
.Y(n_7117)
);

OR2x2_ASAP7_75t_L g7118 ( 
.A(n_6915),
.B(n_731),
.Y(n_7118)
);

INVx1_ASAP7_75t_L g7119 ( 
.A(n_6913),
.Y(n_7119)
);

AOI22xp5_ASAP7_75t_L g7120 ( 
.A1(n_6992),
.A2(n_734),
.B1(n_732),
.B2(n_733),
.Y(n_7120)
);

OR2x2_ASAP7_75t_L g7121 ( 
.A(n_6902),
.B(n_732),
.Y(n_7121)
);

INVx1_ASAP7_75t_L g7122 ( 
.A(n_6905),
.Y(n_7122)
);

AND2x2_ASAP7_75t_L g7123 ( 
.A(n_6988),
.B(n_733),
.Y(n_7123)
);

OAI21xp33_ASAP7_75t_L g7124 ( 
.A1(n_6938),
.A2(n_733),
.B(n_735),
.Y(n_7124)
);

INVx1_ASAP7_75t_L g7125 ( 
.A(n_6874),
.Y(n_7125)
);

NAND2xp5_ASAP7_75t_L g7126 ( 
.A(n_6908),
.B(n_735),
.Y(n_7126)
);

NOR2xp33_ASAP7_75t_L g7127 ( 
.A(n_6937),
.B(n_6953),
.Y(n_7127)
);

AND2x4_ASAP7_75t_L g7128 ( 
.A(n_6977),
.B(n_735),
.Y(n_7128)
);

INVx3_ASAP7_75t_L g7129 ( 
.A(n_6906),
.Y(n_7129)
);

INVx2_ASAP7_75t_L g7130 ( 
.A(n_6942),
.Y(n_7130)
);

OR2x2_ASAP7_75t_L g7131 ( 
.A(n_6967),
.B(n_736),
.Y(n_7131)
);

NAND2xp5_ASAP7_75t_L g7132 ( 
.A(n_6970),
.B(n_736),
.Y(n_7132)
);

AND2x2_ASAP7_75t_L g7133 ( 
.A(n_6993),
.B(n_736),
.Y(n_7133)
);

NAND2xp5_ASAP7_75t_L g7134 ( 
.A(n_6873),
.B(n_737),
.Y(n_7134)
);

AND2x2_ASAP7_75t_L g7135 ( 
.A(n_6989),
.B(n_737),
.Y(n_7135)
);

NAND2xp5_ASAP7_75t_L g7136 ( 
.A(n_6914),
.B(n_737),
.Y(n_7136)
);

INVx1_ASAP7_75t_L g7137 ( 
.A(n_6955),
.Y(n_7137)
);

INVx2_ASAP7_75t_L g7138 ( 
.A(n_6930),
.Y(n_7138)
);

AOI22xp33_ASAP7_75t_L g7139 ( 
.A1(n_6979),
.A2(n_6878),
.B1(n_6966),
.B2(n_6984),
.Y(n_7139)
);

INVx3_ASAP7_75t_L g7140 ( 
.A(n_6906),
.Y(n_7140)
);

AND2x2_ASAP7_75t_L g7141 ( 
.A(n_6995),
.B(n_738),
.Y(n_7141)
);

AND2x2_ASAP7_75t_L g7142 ( 
.A(n_6879),
.B(n_738),
.Y(n_7142)
);

AND2x2_ASAP7_75t_L g7143 ( 
.A(n_6881),
.B(n_738),
.Y(n_7143)
);

INVxp67_ASAP7_75t_SL g7144 ( 
.A(n_6944),
.Y(n_7144)
);

NAND2xp5_ASAP7_75t_SL g7145 ( 
.A(n_6889),
.B(n_739),
.Y(n_7145)
);

AND2x2_ASAP7_75t_L g7146 ( 
.A(n_6936),
.B(n_740),
.Y(n_7146)
);

INVx1_ASAP7_75t_L g7147 ( 
.A(n_6925),
.Y(n_7147)
);

INVxp33_ASAP7_75t_L g7148 ( 
.A(n_6872),
.Y(n_7148)
);

AOI21xp5_ASAP7_75t_L g7149 ( 
.A1(n_6870),
.A2(n_740),
.B(n_741),
.Y(n_7149)
);

AND2x2_ASAP7_75t_L g7150 ( 
.A(n_6962),
.B(n_740),
.Y(n_7150)
);

NAND2xp5_ASAP7_75t_L g7151 ( 
.A(n_6907),
.B(n_741),
.Y(n_7151)
);

NAND2xp5_ASAP7_75t_L g7152 ( 
.A(n_6939),
.B(n_741),
.Y(n_7152)
);

OR2x2_ASAP7_75t_L g7153 ( 
.A(n_6974),
.B(n_742),
.Y(n_7153)
);

NOR2xp33_ASAP7_75t_L g7154 ( 
.A(n_6945),
.B(n_742),
.Y(n_7154)
);

OR2x2_ASAP7_75t_L g7155 ( 
.A(n_6990),
.B(n_743),
.Y(n_7155)
);

INVx1_ASAP7_75t_L g7156 ( 
.A(n_6929),
.Y(n_7156)
);

NAND2xp5_ASAP7_75t_SL g7157 ( 
.A(n_6980),
.B(n_743),
.Y(n_7157)
);

OR2x2_ASAP7_75t_L g7158 ( 
.A(n_6994),
.B(n_743),
.Y(n_7158)
);

AND2x2_ASAP7_75t_L g7159 ( 
.A(n_6983),
.B(n_744),
.Y(n_7159)
);

INVx2_ASAP7_75t_L g7160 ( 
.A(n_6973),
.Y(n_7160)
);

NAND2xp5_ASAP7_75t_L g7161 ( 
.A(n_6890),
.B(n_744),
.Y(n_7161)
);

AOI22xp5_ASAP7_75t_L g7162 ( 
.A1(n_7106),
.A2(n_6916),
.B1(n_6975),
.B2(n_6951),
.Y(n_7162)
);

NAND2xp5_ASAP7_75t_L g7163 ( 
.A(n_7051),
.B(n_6900),
.Y(n_7163)
);

NAND2xp5_ASAP7_75t_L g7164 ( 
.A(n_7054),
.B(n_6898),
.Y(n_7164)
);

INVx2_ASAP7_75t_SL g7165 ( 
.A(n_7028),
.Y(n_7165)
);

AND2x2_ASAP7_75t_L g7166 ( 
.A(n_7063),
.B(n_6985),
.Y(n_7166)
);

INVx1_ASAP7_75t_L g7167 ( 
.A(n_7035),
.Y(n_7167)
);

AOI22xp5_ASAP7_75t_L g7168 ( 
.A1(n_7042),
.A2(n_6986),
.B1(n_7001),
.B2(n_6998),
.Y(n_7168)
);

OR2x2_ASAP7_75t_L g7169 ( 
.A(n_7035),
.B(n_6867),
.Y(n_7169)
);

INVxp67_ASAP7_75t_L g7170 ( 
.A(n_7048),
.Y(n_7170)
);

NOR2xp33_ASAP7_75t_L g7171 ( 
.A(n_7103),
.B(n_6948),
.Y(n_7171)
);

INVx1_ASAP7_75t_L g7172 ( 
.A(n_7033),
.Y(n_7172)
);

AOI32xp33_ASAP7_75t_L g7173 ( 
.A1(n_7084),
.A2(n_6959),
.A3(n_6961),
.B1(n_6941),
.B2(n_6940),
.Y(n_7173)
);

INVx1_ASAP7_75t_L g7174 ( 
.A(n_7069),
.Y(n_7174)
);

INVx1_ASAP7_75t_L g7175 ( 
.A(n_7056),
.Y(n_7175)
);

AND2x2_ASAP7_75t_L g7176 ( 
.A(n_7038),
.B(n_6949),
.Y(n_7176)
);

NAND2xp5_ASAP7_75t_SL g7177 ( 
.A(n_7073),
.B(n_6893),
.Y(n_7177)
);

AOI21xp5_ASAP7_75t_L g7178 ( 
.A1(n_7053),
.A2(n_6923),
.B(n_6968),
.Y(n_7178)
);

AOI22xp5_ASAP7_75t_L g7179 ( 
.A1(n_7102),
.A2(n_6981),
.B1(n_6931),
.B2(n_6932),
.Y(n_7179)
);

AOI22xp5_ASAP7_75t_L g7180 ( 
.A1(n_7093),
.A2(n_6969),
.B1(n_6958),
.B2(n_6888),
.Y(n_7180)
);

INVx1_ASAP7_75t_L g7181 ( 
.A(n_7159),
.Y(n_7181)
);

NAND2xp5_ASAP7_75t_L g7182 ( 
.A(n_7120),
.B(n_6963),
.Y(n_7182)
);

OAI22xp5_ASAP7_75t_L g7183 ( 
.A1(n_7139),
.A2(n_6978),
.B1(n_6960),
.B2(n_7002),
.Y(n_7183)
);

NAND3xp33_ASAP7_75t_L g7184 ( 
.A(n_7067),
.B(n_6991),
.C(n_6924),
.Y(n_7184)
);

OR2x2_ASAP7_75t_L g7185 ( 
.A(n_7091),
.B(n_6909),
.Y(n_7185)
);

NOR2xp33_ASAP7_75t_SL g7186 ( 
.A(n_7080),
.B(n_744),
.Y(n_7186)
);

INVx1_ASAP7_75t_L g7187 ( 
.A(n_7031),
.Y(n_7187)
);

OAI21xp33_ASAP7_75t_L g7188 ( 
.A1(n_7148),
.A2(n_745),
.B(n_746),
.Y(n_7188)
);

NAND2xp5_ASAP7_75t_L g7189 ( 
.A(n_7036),
.B(n_745),
.Y(n_7189)
);

INVx1_ASAP7_75t_L g7190 ( 
.A(n_7032),
.Y(n_7190)
);

INVxp67_ASAP7_75t_L g7191 ( 
.A(n_7057),
.Y(n_7191)
);

AOI32xp33_ASAP7_75t_L g7192 ( 
.A1(n_7058),
.A2(n_748),
.A3(n_746),
.B1(n_747),
.B2(n_749),
.Y(n_7192)
);

OAI211xp5_ASAP7_75t_L g7193 ( 
.A1(n_7145),
.A2(n_750),
.B(n_746),
.C(n_748),
.Y(n_7193)
);

OAI21xp33_ASAP7_75t_SL g7194 ( 
.A1(n_7157),
.A2(n_748),
.B(n_750),
.Y(n_7194)
);

BUFx2_ASAP7_75t_L g7195 ( 
.A(n_7079),
.Y(n_7195)
);

AOI22xp33_ASAP7_75t_L g7196 ( 
.A1(n_7160),
.A2(n_7086),
.B1(n_7081),
.B2(n_7074),
.Y(n_7196)
);

AOI21xp33_ASAP7_75t_SL g7197 ( 
.A1(n_7153),
.A2(n_750),
.B(n_751),
.Y(n_7197)
);

INVx1_ASAP7_75t_L g7198 ( 
.A(n_7060),
.Y(n_7198)
);

OAI22xp33_ASAP7_75t_L g7199 ( 
.A1(n_7096),
.A2(n_1067),
.B1(n_754),
.B2(n_752),
.Y(n_7199)
);

AOI22xp5_ASAP7_75t_L g7200 ( 
.A1(n_7144),
.A2(n_754),
.B1(n_752),
.B2(n_753),
.Y(n_7200)
);

OAI21xp33_ASAP7_75t_L g7201 ( 
.A1(n_7127),
.A2(n_753),
.B(n_754),
.Y(n_7201)
);

INVx2_ASAP7_75t_SL g7202 ( 
.A(n_7043),
.Y(n_7202)
);

OAI31xp33_ASAP7_75t_L g7203 ( 
.A1(n_7124),
.A2(n_756),
.A3(n_753),
.B(n_755),
.Y(n_7203)
);

OR2x2_ASAP7_75t_L g7204 ( 
.A(n_7151),
.B(n_756),
.Y(n_7204)
);

INVx2_ASAP7_75t_L g7205 ( 
.A(n_7129),
.Y(n_7205)
);

INVx1_ASAP7_75t_L g7206 ( 
.A(n_7150),
.Y(n_7206)
);

OR2x2_ASAP7_75t_L g7207 ( 
.A(n_7129),
.B(n_757),
.Y(n_7207)
);

AND2x2_ASAP7_75t_L g7208 ( 
.A(n_7040),
.B(n_7046),
.Y(n_7208)
);

AOI22xp5_ASAP7_75t_L g7209 ( 
.A1(n_7100),
.A2(n_759),
.B1(n_757),
.B2(n_758),
.Y(n_7209)
);

AND2x2_ASAP7_75t_L g7210 ( 
.A(n_7049),
.B(n_758),
.Y(n_7210)
);

INVx1_ASAP7_75t_SL g7211 ( 
.A(n_7037),
.Y(n_7211)
);

INVx1_ASAP7_75t_SL g7212 ( 
.A(n_7041),
.Y(n_7212)
);

AND2x2_ASAP7_75t_L g7213 ( 
.A(n_7097),
.B(n_758),
.Y(n_7213)
);

AOI22xp33_ASAP7_75t_L g7214 ( 
.A1(n_7095),
.A2(n_7108),
.B1(n_7077),
.B2(n_7140),
.Y(n_7214)
);

OAI22xp33_ASAP7_75t_L g7215 ( 
.A1(n_7061),
.A2(n_1065),
.B1(n_761),
.B2(n_759),
.Y(n_7215)
);

OAI33xp33_ASAP7_75t_L g7216 ( 
.A1(n_7109),
.A2(n_761),
.A3(n_763),
.B1(n_759),
.B2(n_760),
.B3(n_762),
.Y(n_7216)
);

NAND2xp5_ASAP7_75t_L g7217 ( 
.A(n_7140),
.B(n_760),
.Y(n_7217)
);

NOR2xp33_ASAP7_75t_L g7218 ( 
.A(n_7039),
.B(n_760),
.Y(n_7218)
);

INVx1_ASAP7_75t_L g7219 ( 
.A(n_7114),
.Y(n_7219)
);

NOR2xp67_ASAP7_75t_SL g7220 ( 
.A(n_7137),
.B(n_761),
.Y(n_7220)
);

NOR2xp33_ASAP7_75t_L g7221 ( 
.A(n_7132),
.B(n_7083),
.Y(n_7221)
);

INVx1_ASAP7_75t_L g7222 ( 
.A(n_7079),
.Y(n_7222)
);

AOI32xp33_ASAP7_75t_L g7223 ( 
.A1(n_7128),
.A2(n_764),
.A3(n_762),
.B1(n_763),
.B2(n_765),
.Y(n_7223)
);

AND3x1_ASAP7_75t_L g7224 ( 
.A(n_7141),
.B(n_762),
.C(n_763),
.Y(n_7224)
);

CKINVDCx16_ASAP7_75t_R g7225 ( 
.A(n_7076),
.Y(n_7225)
);

INVx2_ASAP7_75t_SL g7226 ( 
.A(n_7104),
.Y(n_7226)
);

OAI22xp5_ASAP7_75t_L g7227 ( 
.A1(n_7134),
.A2(n_766),
.B1(n_764),
.B2(n_765),
.Y(n_7227)
);

INVx1_ASAP7_75t_L g7228 ( 
.A(n_7066),
.Y(n_7228)
);

INVx2_ASAP7_75t_L g7229 ( 
.A(n_7098),
.Y(n_7229)
);

OAI21xp5_ASAP7_75t_L g7230 ( 
.A1(n_7149),
.A2(n_764),
.B(n_765),
.Y(n_7230)
);

INVx2_ASAP7_75t_L g7231 ( 
.A(n_7101),
.Y(n_7231)
);

INVx1_ASAP7_75t_L g7232 ( 
.A(n_7052),
.Y(n_7232)
);

INVx1_ASAP7_75t_L g7233 ( 
.A(n_7072),
.Y(n_7233)
);

OA222x2_ASAP7_75t_L g7234 ( 
.A1(n_7121),
.A2(n_768),
.B1(n_770),
.B2(n_766),
.C1(n_767),
.C2(n_769),
.Y(n_7234)
);

INVx1_ASAP7_75t_SL g7235 ( 
.A(n_7128),
.Y(n_7235)
);

INVxp67_ASAP7_75t_L g7236 ( 
.A(n_7154),
.Y(n_7236)
);

NAND3xp33_ASAP7_75t_L g7237 ( 
.A(n_7068),
.B(n_766),
.C(n_767),
.Y(n_7237)
);

HB1xp67_ASAP7_75t_L g7238 ( 
.A(n_7105),
.Y(n_7238)
);

NAND2x1_ASAP7_75t_L g7239 ( 
.A(n_7130),
.B(n_767),
.Y(n_7239)
);

OR2x2_ASAP7_75t_L g7240 ( 
.A(n_7118),
.B(n_768),
.Y(n_7240)
);

AO22x1_ASAP7_75t_L g7241 ( 
.A1(n_7123),
.A2(n_771),
.B1(n_769),
.B2(n_770),
.Y(n_7241)
);

INVx1_ASAP7_75t_L g7242 ( 
.A(n_7115),
.Y(n_7242)
);

INVx1_ASAP7_75t_L g7243 ( 
.A(n_7082),
.Y(n_7243)
);

NAND2xp5_ASAP7_75t_L g7244 ( 
.A(n_7099),
.B(n_771),
.Y(n_7244)
);

AND2x2_ASAP7_75t_L g7245 ( 
.A(n_7088),
.B(n_771),
.Y(n_7245)
);

AND2x2_ASAP7_75t_L g7246 ( 
.A(n_7090),
.B(n_772),
.Y(n_7246)
);

INVx1_ASAP7_75t_L g7247 ( 
.A(n_7133),
.Y(n_7247)
);

NAND2xp5_ASAP7_75t_L g7248 ( 
.A(n_7112),
.B(n_773),
.Y(n_7248)
);

INVx1_ASAP7_75t_L g7249 ( 
.A(n_7135),
.Y(n_7249)
);

INVx2_ASAP7_75t_L g7250 ( 
.A(n_7138),
.Y(n_7250)
);

INVx1_ASAP7_75t_L g7251 ( 
.A(n_7155),
.Y(n_7251)
);

INVx1_ASAP7_75t_SL g7252 ( 
.A(n_7158),
.Y(n_7252)
);

OAI21xp33_ASAP7_75t_L g7253 ( 
.A1(n_7111),
.A2(n_773),
.B(n_774),
.Y(n_7253)
);

INVx1_ASAP7_75t_L g7254 ( 
.A(n_7089),
.Y(n_7254)
);

AND2x2_ASAP7_75t_L g7255 ( 
.A(n_7094),
.B(n_774),
.Y(n_7255)
);

INVx2_ASAP7_75t_SL g7256 ( 
.A(n_7146),
.Y(n_7256)
);

OR2x6_ASAP7_75t_L g7257 ( 
.A(n_7161),
.B(n_775),
.Y(n_7257)
);

INVx1_ASAP7_75t_L g7258 ( 
.A(n_7142),
.Y(n_7258)
);

HB1xp67_ASAP7_75t_L g7259 ( 
.A(n_7078),
.Y(n_7259)
);

INVx2_ASAP7_75t_L g7260 ( 
.A(n_7107),
.Y(n_7260)
);

INVxp67_ASAP7_75t_SL g7261 ( 
.A(n_7136),
.Y(n_7261)
);

INVx1_ASAP7_75t_L g7262 ( 
.A(n_7143),
.Y(n_7262)
);

AND2x2_ASAP7_75t_L g7263 ( 
.A(n_7065),
.B(n_775),
.Y(n_7263)
);

INVx1_ASAP7_75t_L g7264 ( 
.A(n_7071),
.Y(n_7264)
);

OR2x2_ASAP7_75t_L g7265 ( 
.A(n_7126),
.B(n_775),
.Y(n_7265)
);

INVx1_ASAP7_75t_L g7266 ( 
.A(n_7087),
.Y(n_7266)
);

INVx3_ASAP7_75t_L g7267 ( 
.A(n_7116),
.Y(n_7267)
);

NAND2x1_ASAP7_75t_L g7268 ( 
.A(n_7117),
.B(n_776),
.Y(n_7268)
);

INVx1_ASAP7_75t_L g7269 ( 
.A(n_7092),
.Y(n_7269)
);

INVx2_ASAP7_75t_L g7270 ( 
.A(n_7119),
.Y(n_7270)
);

INVx3_ASAP7_75t_L g7271 ( 
.A(n_7131),
.Y(n_7271)
);

AOI211xp5_ASAP7_75t_SL g7272 ( 
.A1(n_7064),
.A2(n_778),
.B(n_776),
.C(n_777),
.Y(n_7272)
);

INVx2_ASAP7_75t_L g7273 ( 
.A(n_7029),
.Y(n_7273)
);

AND2x2_ASAP7_75t_L g7274 ( 
.A(n_7110),
.B(n_777),
.Y(n_7274)
);

NOR2xp33_ASAP7_75t_L g7275 ( 
.A(n_7152),
.B(n_777),
.Y(n_7275)
);

NOR2xp33_ASAP7_75t_L g7276 ( 
.A(n_7030),
.B(n_779),
.Y(n_7276)
);

INVx1_ASAP7_75t_L g7277 ( 
.A(n_7062),
.Y(n_7277)
);

OR2x2_ASAP7_75t_L g7278 ( 
.A(n_7113),
.B(n_779),
.Y(n_7278)
);

INVx1_ASAP7_75t_L g7279 ( 
.A(n_7034),
.Y(n_7279)
);

INVx1_ASAP7_75t_L g7280 ( 
.A(n_7044),
.Y(n_7280)
);

OA222x2_ASAP7_75t_L g7281 ( 
.A1(n_7045),
.A2(n_781),
.B1(n_783),
.B2(n_779),
.C1(n_780),
.C2(n_782),
.Y(n_7281)
);

INVx1_ASAP7_75t_L g7282 ( 
.A(n_7047),
.Y(n_7282)
);

OAI22xp33_ASAP7_75t_L g7283 ( 
.A1(n_7125),
.A2(n_1063),
.B1(n_782),
.B2(n_780),
.Y(n_7283)
);

INVx1_ASAP7_75t_L g7284 ( 
.A(n_7050),
.Y(n_7284)
);

OAI22xp33_ASAP7_75t_L g7285 ( 
.A1(n_7122),
.A2(n_783),
.B1(n_781),
.B2(n_782),
.Y(n_7285)
);

AOI22xp5_ASAP7_75t_L g7286 ( 
.A1(n_7147),
.A2(n_785),
.B1(n_781),
.B2(n_784),
.Y(n_7286)
);

AND2x2_ASAP7_75t_L g7287 ( 
.A(n_7156),
.B(n_784),
.Y(n_7287)
);

OAI322xp33_ASAP7_75t_L g7288 ( 
.A1(n_7055),
.A2(n_790),
.A3(n_789),
.B1(n_787),
.B2(n_785),
.C1(n_786),
.C2(n_788),
.Y(n_7288)
);

AND2x4_ASAP7_75t_L g7289 ( 
.A(n_7059),
.B(n_786),
.Y(n_7289)
);

INVx2_ASAP7_75t_L g7290 ( 
.A(n_7070),
.Y(n_7290)
);

INVx2_ASAP7_75t_L g7291 ( 
.A(n_7075),
.Y(n_7291)
);

OAI22xp5_ASAP7_75t_L g7292 ( 
.A1(n_7085),
.A2(n_789),
.B1(n_786),
.B2(n_788),
.Y(n_7292)
);

NAND3xp33_ASAP7_75t_L g7293 ( 
.A(n_7067),
.B(n_788),
.C(n_789),
.Y(n_7293)
);

NAND2x1_ASAP7_75t_L g7294 ( 
.A(n_7035),
.B(n_790),
.Y(n_7294)
);

OR2x2_ASAP7_75t_L g7295 ( 
.A(n_7028),
.B(n_790),
.Y(n_7295)
);

HB1xp67_ASAP7_75t_L g7296 ( 
.A(n_7035),
.Y(n_7296)
);

INVx1_ASAP7_75t_L g7297 ( 
.A(n_7035),
.Y(n_7297)
);

INVx1_ASAP7_75t_L g7298 ( 
.A(n_7035),
.Y(n_7298)
);

INVx1_ASAP7_75t_L g7299 ( 
.A(n_7035),
.Y(n_7299)
);

INVx2_ASAP7_75t_L g7300 ( 
.A(n_7028),
.Y(n_7300)
);

OAI21xp33_ASAP7_75t_L g7301 ( 
.A1(n_7093),
.A2(n_791),
.B(n_792),
.Y(n_7301)
);

NOR2xp33_ASAP7_75t_SL g7302 ( 
.A(n_7300),
.B(n_791),
.Y(n_7302)
);

INVx1_ASAP7_75t_L g7303 ( 
.A(n_7296),
.Y(n_7303)
);

INVx1_ASAP7_75t_L g7304 ( 
.A(n_7238),
.Y(n_7304)
);

INVx1_ASAP7_75t_L g7305 ( 
.A(n_7165),
.Y(n_7305)
);

OR2x2_ASAP7_75t_L g7306 ( 
.A(n_7205),
.B(n_792),
.Y(n_7306)
);

INVx1_ASAP7_75t_L g7307 ( 
.A(n_7169),
.Y(n_7307)
);

OR2x2_ASAP7_75t_L g7308 ( 
.A(n_7226),
.B(n_793),
.Y(n_7308)
);

AND2x2_ASAP7_75t_L g7309 ( 
.A(n_7166),
.B(n_793),
.Y(n_7309)
);

AND2x2_ASAP7_75t_L g7310 ( 
.A(n_7245),
.B(n_1063),
.Y(n_7310)
);

AND2x2_ASAP7_75t_SL g7311 ( 
.A(n_7224),
.B(n_794),
.Y(n_7311)
);

INVx2_ASAP7_75t_L g7312 ( 
.A(n_7202),
.Y(n_7312)
);

HB1xp67_ASAP7_75t_L g7313 ( 
.A(n_7294),
.Y(n_7313)
);

AND2x2_ASAP7_75t_L g7314 ( 
.A(n_7210),
.B(n_794),
.Y(n_7314)
);

INVx1_ASAP7_75t_L g7315 ( 
.A(n_7207),
.Y(n_7315)
);

AOI22xp33_ASAP7_75t_L g7316 ( 
.A1(n_7250),
.A2(n_796),
.B1(n_794),
.B2(n_795),
.Y(n_7316)
);

NAND2xp5_ASAP7_75t_L g7317 ( 
.A(n_7241),
.B(n_7196),
.Y(n_7317)
);

INVx3_ASAP7_75t_L g7318 ( 
.A(n_7229),
.Y(n_7318)
);

NAND2x1_ASAP7_75t_L g7319 ( 
.A(n_7167),
.B(n_1054),
.Y(n_7319)
);

NAND2xp5_ASAP7_75t_L g7320 ( 
.A(n_7297),
.B(n_795),
.Y(n_7320)
);

NAND2xp5_ASAP7_75t_L g7321 ( 
.A(n_7298),
.B(n_795),
.Y(n_7321)
);

INVx1_ASAP7_75t_L g7322 ( 
.A(n_7217),
.Y(n_7322)
);

AND2x2_ASAP7_75t_L g7323 ( 
.A(n_7246),
.B(n_1053),
.Y(n_7323)
);

INVx1_ASAP7_75t_L g7324 ( 
.A(n_7239),
.Y(n_7324)
);

INVx1_ASAP7_75t_L g7325 ( 
.A(n_7299),
.Y(n_7325)
);

INVx2_ASAP7_75t_L g7326 ( 
.A(n_7231),
.Y(n_7326)
);

NOR2x1_ASAP7_75t_L g7327 ( 
.A(n_7174),
.B(n_796),
.Y(n_7327)
);

NOR2x1_ASAP7_75t_L g7328 ( 
.A(n_7193),
.B(n_7293),
.Y(n_7328)
);

INVx2_ASAP7_75t_L g7329 ( 
.A(n_7211),
.Y(n_7329)
);

INVx1_ASAP7_75t_L g7330 ( 
.A(n_7195),
.Y(n_7330)
);

NAND2xp5_ASAP7_75t_L g7331 ( 
.A(n_7218),
.B(n_796),
.Y(n_7331)
);

AND2x2_ASAP7_75t_L g7332 ( 
.A(n_7255),
.B(n_1052),
.Y(n_7332)
);

INVx1_ASAP7_75t_SL g7333 ( 
.A(n_7235),
.Y(n_7333)
);

INVx2_ASAP7_75t_L g7334 ( 
.A(n_7295),
.Y(n_7334)
);

AND2x4_ASAP7_75t_L g7335 ( 
.A(n_7222),
.B(n_797),
.Y(n_7335)
);

CKINVDCx5p33_ASAP7_75t_R g7336 ( 
.A(n_7200),
.Y(n_7336)
);

AND2x2_ASAP7_75t_L g7337 ( 
.A(n_7263),
.B(n_7213),
.Y(n_7337)
);

INVx1_ASAP7_75t_L g7338 ( 
.A(n_7163),
.Y(n_7338)
);

HB1xp67_ASAP7_75t_L g7339 ( 
.A(n_7289),
.Y(n_7339)
);

AND2x2_ASAP7_75t_L g7340 ( 
.A(n_7208),
.B(n_1052),
.Y(n_7340)
);

INVx2_ASAP7_75t_L g7341 ( 
.A(n_7260),
.Y(n_7341)
);

INVx1_ASAP7_75t_SL g7342 ( 
.A(n_7212),
.Y(n_7342)
);

INVx1_ASAP7_75t_SL g7343 ( 
.A(n_7252),
.Y(n_7343)
);

INVx1_ASAP7_75t_L g7344 ( 
.A(n_7176),
.Y(n_7344)
);

INVx1_ASAP7_75t_L g7345 ( 
.A(n_7268),
.Y(n_7345)
);

NAND2xp5_ASAP7_75t_L g7346 ( 
.A(n_7272),
.B(n_797),
.Y(n_7346)
);

INVx1_ASAP7_75t_L g7347 ( 
.A(n_7289),
.Y(n_7347)
);

INVx2_ASAP7_75t_SL g7348 ( 
.A(n_7270),
.Y(n_7348)
);

NAND2xp5_ASAP7_75t_L g7349 ( 
.A(n_7287),
.B(n_797),
.Y(n_7349)
);

INVx1_ASAP7_75t_SL g7350 ( 
.A(n_7278),
.Y(n_7350)
);

AOI22xp33_ASAP7_75t_L g7351 ( 
.A1(n_7301),
.A2(n_7184),
.B1(n_7216),
.B2(n_7277),
.Y(n_7351)
);

NAND2x1_ASAP7_75t_SL g7352 ( 
.A(n_7274),
.B(n_7168),
.Y(n_7352)
);

AOI22xp33_ASAP7_75t_L g7353 ( 
.A1(n_7171),
.A2(n_800),
.B1(n_798),
.B2(n_799),
.Y(n_7353)
);

NOR2xp33_ASAP7_75t_L g7354 ( 
.A(n_7186),
.B(n_798),
.Y(n_7354)
);

INVx2_ASAP7_75t_L g7355 ( 
.A(n_7291),
.Y(n_7355)
);

INVx2_ASAP7_75t_L g7356 ( 
.A(n_7273),
.Y(n_7356)
);

NAND2xp5_ASAP7_75t_L g7357 ( 
.A(n_7214),
.B(n_798),
.Y(n_7357)
);

NAND2xp5_ASAP7_75t_L g7358 ( 
.A(n_7225),
.B(n_800),
.Y(n_7358)
);

NOR2x1_ASAP7_75t_L g7359 ( 
.A(n_7199),
.B(n_7215),
.Y(n_7359)
);

INVx1_ASAP7_75t_L g7360 ( 
.A(n_7220),
.Y(n_7360)
);

INVx1_ASAP7_75t_L g7361 ( 
.A(n_7244),
.Y(n_7361)
);

AND2x4_ASAP7_75t_L g7362 ( 
.A(n_7290),
.B(n_800),
.Y(n_7362)
);

HB1xp67_ASAP7_75t_L g7363 ( 
.A(n_7259),
.Y(n_7363)
);

NAND2xp5_ASAP7_75t_L g7364 ( 
.A(n_7173),
.B(n_801),
.Y(n_7364)
);

OR2x2_ASAP7_75t_L g7365 ( 
.A(n_7248),
.B(n_801),
.Y(n_7365)
);

OR2x2_ASAP7_75t_L g7366 ( 
.A(n_7189),
.B(n_801),
.Y(n_7366)
);

INVxp67_ASAP7_75t_SL g7367 ( 
.A(n_7283),
.Y(n_7367)
);

INVxp67_ASAP7_75t_SL g7368 ( 
.A(n_7285),
.Y(n_7368)
);

NAND2xp5_ASAP7_75t_L g7369 ( 
.A(n_7223),
.B(n_802),
.Y(n_7369)
);

INVx1_ASAP7_75t_L g7370 ( 
.A(n_7204),
.Y(n_7370)
);

NAND3xp33_ASAP7_75t_L g7371 ( 
.A(n_7192),
.B(n_802),
.C(n_803),
.Y(n_7371)
);

AND2x2_ASAP7_75t_L g7372 ( 
.A(n_7234),
.B(n_802),
.Y(n_7372)
);

AND2x2_ASAP7_75t_L g7373 ( 
.A(n_7243),
.B(n_7281),
.Y(n_7373)
);

INVx2_ASAP7_75t_L g7374 ( 
.A(n_7267),
.Y(n_7374)
);

AND2x4_ASAP7_75t_L g7375 ( 
.A(n_7237),
.B(n_7251),
.Y(n_7375)
);

INVx2_ASAP7_75t_L g7376 ( 
.A(n_7267),
.Y(n_7376)
);

INVx1_ASAP7_75t_L g7377 ( 
.A(n_7265),
.Y(n_7377)
);

INVx1_ASAP7_75t_L g7378 ( 
.A(n_7240),
.Y(n_7378)
);

INVx1_ASAP7_75t_SL g7379 ( 
.A(n_7177),
.Y(n_7379)
);

BUFx3_ASAP7_75t_L g7380 ( 
.A(n_7242),
.Y(n_7380)
);

INVx1_ASAP7_75t_L g7381 ( 
.A(n_7164),
.Y(n_7381)
);

AND2x2_ASAP7_75t_L g7382 ( 
.A(n_7175),
.B(n_1052),
.Y(n_7382)
);

INVx2_ASAP7_75t_L g7383 ( 
.A(n_7271),
.Y(n_7383)
);

NOR2xp67_ASAP7_75t_L g7384 ( 
.A(n_7194),
.B(n_803),
.Y(n_7384)
);

OR2x2_ASAP7_75t_L g7385 ( 
.A(n_7256),
.B(n_804),
.Y(n_7385)
);

NAND2xp5_ASAP7_75t_SL g7386 ( 
.A(n_7326),
.B(n_7312),
.Y(n_7386)
);

OAI222xp33_ASAP7_75t_L g7387 ( 
.A1(n_7333),
.A2(n_7162),
.B1(n_7191),
.B2(n_7185),
.C1(n_7180),
.C2(n_7182),
.Y(n_7387)
);

OAI22xp5_ASAP7_75t_L g7388 ( 
.A1(n_7305),
.A2(n_7179),
.B1(n_7170),
.B2(n_7236),
.Y(n_7388)
);

NAND2xp5_ASAP7_75t_L g7389 ( 
.A(n_7309),
.B(n_7197),
.Y(n_7389)
);

INVx1_ASAP7_75t_L g7390 ( 
.A(n_7319),
.Y(n_7390)
);

HB1xp67_ASAP7_75t_L g7391 ( 
.A(n_7307),
.Y(n_7391)
);

NOR2x1_ASAP7_75t_L g7392 ( 
.A(n_7357),
.B(n_7279),
.Y(n_7392)
);

AND2x4_ASAP7_75t_L g7393 ( 
.A(n_7318),
.B(n_7181),
.Y(n_7393)
);

INVx1_ASAP7_75t_L g7394 ( 
.A(n_7319),
.Y(n_7394)
);

AOI21xp5_ASAP7_75t_L g7395 ( 
.A1(n_7364),
.A2(n_7178),
.B(n_7230),
.Y(n_7395)
);

INVx1_ASAP7_75t_L g7396 ( 
.A(n_7335),
.Y(n_7396)
);

NOR2xp33_ASAP7_75t_L g7397 ( 
.A(n_7329),
.B(n_7253),
.Y(n_7397)
);

INVx1_ASAP7_75t_SL g7398 ( 
.A(n_7342),
.Y(n_7398)
);

INVx1_ASAP7_75t_L g7399 ( 
.A(n_7335),
.Y(n_7399)
);

AND2x2_ASAP7_75t_L g7400 ( 
.A(n_7340),
.B(n_7172),
.Y(n_7400)
);

NAND2x1_ASAP7_75t_L g7401 ( 
.A(n_7304),
.B(n_7271),
.Y(n_7401)
);

AOI222xp33_ASAP7_75t_L g7402 ( 
.A1(n_7379),
.A2(n_7201),
.B1(n_7183),
.B2(n_7276),
.C1(n_7261),
.C2(n_7206),
.Y(n_7402)
);

AOI221xp5_ASAP7_75t_L g7403 ( 
.A1(n_7344),
.A2(n_7188),
.B1(n_7292),
.B2(n_7227),
.C(n_7288),
.Y(n_7403)
);

OAI22xp5_ASAP7_75t_L g7404 ( 
.A1(n_7351),
.A2(n_7219),
.B1(n_7269),
.B2(n_7266),
.Y(n_7404)
);

NAND2xp5_ASAP7_75t_L g7405 ( 
.A(n_7311),
.B(n_7372),
.Y(n_7405)
);

INVx2_ASAP7_75t_L g7406 ( 
.A(n_7341),
.Y(n_7406)
);

INVx1_ASAP7_75t_L g7407 ( 
.A(n_7362),
.Y(n_7407)
);

AOI22xp5_ASAP7_75t_L g7408 ( 
.A1(n_7367),
.A2(n_7275),
.B1(n_7221),
.B2(n_7198),
.Y(n_7408)
);

INVx1_ASAP7_75t_L g7409 ( 
.A(n_7362),
.Y(n_7409)
);

INVxp67_ASAP7_75t_L g7410 ( 
.A(n_7302),
.Y(n_7410)
);

OAI22xp33_ASAP7_75t_L g7411 ( 
.A1(n_7346),
.A2(n_7257),
.B1(n_7264),
.B2(n_7262),
.Y(n_7411)
);

OAI222xp33_ASAP7_75t_L g7412 ( 
.A1(n_7343),
.A2(n_7303),
.B1(n_7348),
.B2(n_7308),
.C1(n_7330),
.C2(n_7331),
.Y(n_7412)
);

NAND2xp5_ASAP7_75t_L g7413 ( 
.A(n_7384),
.B(n_7286),
.Y(n_7413)
);

AOI221xp5_ASAP7_75t_L g7414 ( 
.A1(n_7354),
.A2(n_7280),
.B1(n_7284),
.B2(n_7282),
.C(n_7258),
.Y(n_7414)
);

INVx1_ASAP7_75t_L g7415 ( 
.A(n_7363),
.Y(n_7415)
);

AOI22xp33_ASAP7_75t_L g7416 ( 
.A1(n_7355),
.A2(n_7232),
.B1(n_7249),
.B2(n_7247),
.Y(n_7416)
);

AOI22xp5_ASAP7_75t_L g7417 ( 
.A1(n_7368),
.A2(n_7190),
.B1(n_7187),
.B2(n_7233),
.Y(n_7417)
);

OAI22xp33_ASAP7_75t_L g7418 ( 
.A1(n_7317),
.A2(n_7257),
.B1(n_7209),
.B2(n_7228),
.Y(n_7418)
);

OAI21xp33_ASAP7_75t_L g7419 ( 
.A1(n_7352),
.A2(n_7254),
.B(n_7203),
.Y(n_7419)
);

NOR2xp33_ASAP7_75t_L g7420 ( 
.A(n_7349),
.B(n_804),
.Y(n_7420)
);

INVx1_ASAP7_75t_L g7421 ( 
.A(n_7339),
.Y(n_7421)
);

AOI211xp5_ASAP7_75t_SL g7422 ( 
.A1(n_7369),
.A2(n_806),
.B(n_804),
.C(n_805),
.Y(n_7422)
);

NAND2xp5_ASAP7_75t_L g7423 ( 
.A(n_7310),
.B(n_805),
.Y(n_7423)
);

INVx1_ASAP7_75t_L g7424 ( 
.A(n_7313),
.Y(n_7424)
);

INVxp67_ASAP7_75t_L g7425 ( 
.A(n_7327),
.Y(n_7425)
);

OAI221xp5_ASAP7_75t_SL g7426 ( 
.A1(n_7306),
.A2(n_808),
.B1(n_806),
.B2(n_807),
.C(n_809),
.Y(n_7426)
);

INVx1_ASAP7_75t_L g7427 ( 
.A(n_7320),
.Y(n_7427)
);

AOI221xp5_ASAP7_75t_L g7428 ( 
.A1(n_7371),
.A2(n_810),
.B1(n_808),
.B2(n_809),
.C(n_811),
.Y(n_7428)
);

NAND2x1_ASAP7_75t_SL g7429 ( 
.A(n_7382),
.B(n_1051),
.Y(n_7429)
);

NOR2xp33_ASAP7_75t_L g7430 ( 
.A(n_7356),
.B(n_808),
.Y(n_7430)
);

AND2x2_ASAP7_75t_L g7431 ( 
.A(n_7314),
.B(n_809),
.Y(n_7431)
);

OR2x2_ASAP7_75t_L g7432 ( 
.A(n_7385),
.B(n_810),
.Y(n_7432)
);

INVx1_ASAP7_75t_L g7433 ( 
.A(n_7321),
.Y(n_7433)
);

INVx3_ASAP7_75t_L g7434 ( 
.A(n_7380),
.Y(n_7434)
);

INVx1_ASAP7_75t_L g7435 ( 
.A(n_7358),
.Y(n_7435)
);

INVx1_ASAP7_75t_SL g7436 ( 
.A(n_7325),
.Y(n_7436)
);

NOR2xp33_ASAP7_75t_L g7437 ( 
.A(n_7347),
.B(n_811),
.Y(n_7437)
);

OR2x2_ASAP7_75t_L g7438 ( 
.A(n_7374),
.B(n_811),
.Y(n_7438)
);

AOI21xp33_ASAP7_75t_SL g7439 ( 
.A1(n_7338),
.A2(n_812),
.B(n_813),
.Y(n_7439)
);

OAI21xp33_ASAP7_75t_L g7440 ( 
.A1(n_7381),
.A2(n_812),
.B(n_813),
.Y(n_7440)
);

INVx1_ASAP7_75t_L g7441 ( 
.A(n_7323),
.Y(n_7441)
);

INVx1_ASAP7_75t_SL g7442 ( 
.A(n_7376),
.Y(n_7442)
);

AND2x2_ASAP7_75t_L g7443 ( 
.A(n_7332),
.B(n_813),
.Y(n_7443)
);

OAI31xp33_ASAP7_75t_L g7444 ( 
.A1(n_7360),
.A2(n_816),
.A3(n_814),
.B(n_815),
.Y(n_7444)
);

INVx2_ASAP7_75t_L g7445 ( 
.A(n_7383),
.Y(n_7445)
);

OR2x2_ASAP7_75t_L g7446 ( 
.A(n_7365),
.B(n_814),
.Y(n_7446)
);

OR2x2_ASAP7_75t_L g7447 ( 
.A(n_7366),
.B(n_814),
.Y(n_7447)
);

OAI21xp5_ASAP7_75t_L g7448 ( 
.A1(n_7328),
.A2(n_815),
.B(n_816),
.Y(n_7448)
);

OAI21xp5_ASAP7_75t_L g7449 ( 
.A1(n_7359),
.A2(n_816),
.B(n_817),
.Y(n_7449)
);

INVx1_ASAP7_75t_L g7450 ( 
.A(n_7345),
.Y(n_7450)
);

AOI22xp5_ASAP7_75t_L g7451 ( 
.A1(n_7375),
.A2(n_819),
.B1(n_817),
.B2(n_818),
.Y(n_7451)
);

NOR2xp33_ASAP7_75t_L g7452 ( 
.A(n_7324),
.B(n_817),
.Y(n_7452)
);

NOR2xp33_ASAP7_75t_L g7453 ( 
.A(n_7350),
.B(n_818),
.Y(n_7453)
);

INVx1_ASAP7_75t_L g7454 ( 
.A(n_7315),
.Y(n_7454)
);

NAND2xp5_ASAP7_75t_L g7455 ( 
.A(n_7316),
.B(n_7337),
.Y(n_7455)
);

NAND2xp5_ASAP7_75t_L g7456 ( 
.A(n_7353),
.B(n_818),
.Y(n_7456)
);

INVx1_ASAP7_75t_L g7457 ( 
.A(n_7334),
.Y(n_7457)
);

NAND2xp5_ASAP7_75t_L g7458 ( 
.A(n_7373),
.B(n_819),
.Y(n_7458)
);

OAI21xp33_ASAP7_75t_L g7459 ( 
.A1(n_7336),
.A2(n_819),
.B(n_820),
.Y(n_7459)
);

INVx1_ASAP7_75t_L g7460 ( 
.A(n_7375),
.Y(n_7460)
);

AOI211xp5_ASAP7_75t_L g7461 ( 
.A1(n_7378),
.A2(n_822),
.B(n_820),
.C(n_821),
.Y(n_7461)
);

INVx1_ASAP7_75t_L g7462 ( 
.A(n_7370),
.Y(n_7462)
);

O2A1O1Ixp33_ASAP7_75t_L g7463 ( 
.A1(n_7377),
.A2(n_824),
.B(n_822),
.C(n_823),
.Y(n_7463)
);

INVx1_ASAP7_75t_SL g7464 ( 
.A(n_7322),
.Y(n_7464)
);

OAI21xp33_ASAP7_75t_L g7465 ( 
.A1(n_7361),
.A2(n_823),
.B(n_824),
.Y(n_7465)
);

NAND4xp25_ASAP7_75t_SL g7466 ( 
.A(n_7333),
.B(n_827),
.C(n_825),
.D(n_826),
.Y(n_7466)
);

OAI322xp33_ASAP7_75t_L g7467 ( 
.A1(n_7333),
.A2(n_825),
.A3(n_826),
.B1(n_827),
.B2(n_828),
.C1(n_829),
.C2(n_830),
.Y(n_7467)
);

NAND2xp5_ASAP7_75t_L g7468 ( 
.A(n_7326),
.B(n_825),
.Y(n_7468)
);

AOI22xp5_ASAP7_75t_L g7469 ( 
.A1(n_7305),
.A2(n_828),
.B1(n_826),
.B2(n_827),
.Y(n_7469)
);

AOI22xp5_ASAP7_75t_L g7470 ( 
.A1(n_7305),
.A2(n_830),
.B1(n_828),
.B2(n_829),
.Y(n_7470)
);

INVx2_ASAP7_75t_L g7471 ( 
.A(n_7326),
.Y(n_7471)
);

AOI22xp33_ASAP7_75t_L g7472 ( 
.A1(n_7326),
.A2(n_831),
.B1(n_829),
.B2(n_830),
.Y(n_7472)
);

OR2x2_ASAP7_75t_L g7473 ( 
.A(n_7326),
.B(n_831),
.Y(n_7473)
);

NAND2xp5_ASAP7_75t_L g7474 ( 
.A(n_7326),
.B(n_831),
.Y(n_7474)
);

OR2x2_ASAP7_75t_L g7475 ( 
.A(n_7326),
.B(n_832),
.Y(n_7475)
);

OAI32xp33_ASAP7_75t_L g7476 ( 
.A1(n_7333),
.A2(n_834),
.A3(n_832),
.B1(n_833),
.B2(n_835),
.Y(n_7476)
);

INVx1_ASAP7_75t_L g7477 ( 
.A(n_7326),
.Y(n_7477)
);

INVxp67_ASAP7_75t_L g7478 ( 
.A(n_7302),
.Y(n_7478)
);

AOI22xp33_ASAP7_75t_L g7479 ( 
.A1(n_7326),
.A2(n_834),
.B1(n_832),
.B2(n_833),
.Y(n_7479)
);

OR2x2_ASAP7_75t_L g7480 ( 
.A(n_7326),
.B(n_833),
.Y(n_7480)
);

AO221x1_ASAP7_75t_L g7481 ( 
.A1(n_7387),
.A2(n_838),
.B1(n_835),
.B2(n_837),
.C(n_839),
.Y(n_7481)
);

INVxp67_ASAP7_75t_L g7482 ( 
.A(n_7391),
.Y(n_7482)
);

AND2x2_ASAP7_75t_L g7483 ( 
.A(n_7398),
.B(n_835),
.Y(n_7483)
);

OAI22xp33_ASAP7_75t_L g7484 ( 
.A1(n_7442),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_7484)
);

OAI22xp33_ASAP7_75t_L g7485 ( 
.A1(n_7471),
.A2(n_839),
.B1(n_837),
.B2(n_838),
.Y(n_7485)
);

OAI22xp33_ASAP7_75t_L g7486 ( 
.A1(n_7477),
.A2(n_842),
.B1(n_840),
.B2(n_841),
.Y(n_7486)
);

AOI22x1_ASAP7_75t_L g7487 ( 
.A1(n_7406),
.A2(n_842),
.B1(n_840),
.B2(n_841),
.Y(n_7487)
);

INVxp67_ASAP7_75t_L g7488 ( 
.A(n_7386),
.Y(n_7488)
);

OR2x2_ASAP7_75t_L g7489 ( 
.A(n_7445),
.B(n_840),
.Y(n_7489)
);

INVx1_ASAP7_75t_L g7490 ( 
.A(n_7468),
.Y(n_7490)
);

AOI21xp5_ASAP7_75t_L g7491 ( 
.A1(n_7458),
.A2(n_843),
.B(n_844),
.Y(n_7491)
);

AOI22xp5_ASAP7_75t_L g7492 ( 
.A1(n_7460),
.A2(n_1051),
.B1(n_845),
.B2(n_843),
.Y(n_7492)
);

INVx1_ASAP7_75t_L g7493 ( 
.A(n_7474),
.Y(n_7493)
);

INVx1_ASAP7_75t_L g7494 ( 
.A(n_7438),
.Y(n_7494)
);

NAND2xp5_ASAP7_75t_L g7495 ( 
.A(n_7421),
.B(n_843),
.Y(n_7495)
);

OAI21xp5_ASAP7_75t_SL g7496 ( 
.A1(n_7408),
.A2(n_844),
.B(n_845),
.Y(n_7496)
);

OA21x2_ASAP7_75t_L g7497 ( 
.A1(n_7405),
.A2(n_1050),
.B(n_844),
.Y(n_7497)
);

NAND3xp33_ASAP7_75t_L g7498 ( 
.A(n_7461),
.B(n_845),
.C(n_846),
.Y(n_7498)
);

AOI22xp5_ASAP7_75t_L g7499 ( 
.A1(n_7397),
.A2(n_1050),
.B1(n_848),
.B2(n_846),
.Y(n_7499)
);

OAI21xp33_ASAP7_75t_L g7500 ( 
.A1(n_7416),
.A2(n_7419),
.B(n_7457),
.Y(n_7500)
);

AOI22xp33_ASAP7_75t_SL g7501 ( 
.A1(n_7434),
.A2(n_849),
.B1(n_847),
.B2(n_848),
.Y(n_7501)
);

NAND2xp5_ASAP7_75t_L g7502 ( 
.A(n_7431),
.B(n_847),
.Y(n_7502)
);

INVx1_ASAP7_75t_L g7503 ( 
.A(n_7432),
.Y(n_7503)
);

OAI21xp5_ASAP7_75t_L g7504 ( 
.A1(n_7395),
.A2(n_847),
.B(n_848),
.Y(n_7504)
);

AND2x2_ASAP7_75t_L g7505 ( 
.A(n_7443),
.B(n_850),
.Y(n_7505)
);

OAI21xp5_ASAP7_75t_L g7506 ( 
.A1(n_7452),
.A2(n_7437),
.B(n_7422),
.Y(n_7506)
);

NAND2xp5_ASAP7_75t_L g7507 ( 
.A(n_7434),
.B(n_850),
.Y(n_7507)
);

INVx2_ASAP7_75t_L g7508 ( 
.A(n_7393),
.Y(n_7508)
);

OAI22xp5_ASAP7_75t_L g7509 ( 
.A1(n_7424),
.A2(n_852),
.B1(n_850),
.B2(n_851),
.Y(n_7509)
);

INVx2_ASAP7_75t_L g7510 ( 
.A(n_7393),
.Y(n_7510)
);

INVx1_ASAP7_75t_L g7511 ( 
.A(n_7473),
.Y(n_7511)
);

OAI222xp33_ASAP7_75t_L g7512 ( 
.A1(n_7436),
.A2(n_851),
.B1(n_852),
.B2(n_853),
.C1(n_854),
.C2(n_855),
.Y(n_7512)
);

OAI22xp5_ASAP7_75t_L g7513 ( 
.A1(n_7417),
.A2(n_855),
.B1(n_851),
.B2(n_854),
.Y(n_7513)
);

INVx1_ASAP7_75t_L g7514 ( 
.A(n_7475),
.Y(n_7514)
);

INVx1_ASAP7_75t_L g7515 ( 
.A(n_7480),
.Y(n_7515)
);

NOR2xp33_ASAP7_75t_L g7516 ( 
.A(n_7459),
.B(n_854),
.Y(n_7516)
);

AND2x2_ASAP7_75t_L g7517 ( 
.A(n_7400),
.B(n_856),
.Y(n_7517)
);

OAI21xp5_ASAP7_75t_L g7518 ( 
.A1(n_7449),
.A2(n_856),
.B(n_857),
.Y(n_7518)
);

INVx1_ASAP7_75t_L g7519 ( 
.A(n_7396),
.Y(n_7519)
);

OAI221xp5_ASAP7_75t_SL g7520 ( 
.A1(n_7444),
.A2(n_858),
.B1(n_856),
.B2(n_857),
.C(n_859),
.Y(n_7520)
);

AOI222xp33_ASAP7_75t_L g7521 ( 
.A1(n_7428),
.A2(n_857),
.B1(n_858),
.B2(n_859),
.C1(n_860),
.C2(n_861),
.Y(n_7521)
);

INVxp67_ASAP7_75t_L g7522 ( 
.A(n_7430),
.Y(n_7522)
);

INVx1_ASAP7_75t_L g7523 ( 
.A(n_7399),
.Y(n_7523)
);

AND2x2_ASAP7_75t_L g7524 ( 
.A(n_7415),
.B(n_858),
.Y(n_7524)
);

OAI21xp5_ASAP7_75t_L g7525 ( 
.A1(n_7453),
.A2(n_859),
.B(n_860),
.Y(n_7525)
);

HB1xp67_ASAP7_75t_L g7526 ( 
.A(n_7401),
.Y(n_7526)
);

INVx1_ASAP7_75t_L g7527 ( 
.A(n_7423),
.Y(n_7527)
);

INVx1_ASAP7_75t_L g7528 ( 
.A(n_7526),
.Y(n_7528)
);

NAND2xp5_ASAP7_75t_L g7529 ( 
.A(n_7508),
.B(n_7472),
.Y(n_7529)
);

NOR2xp33_ASAP7_75t_SL g7530 ( 
.A(n_7500),
.B(n_7450),
.Y(n_7530)
);

HB1xp67_ASAP7_75t_L g7531 ( 
.A(n_7510),
.Y(n_7531)
);

AND2x2_ASAP7_75t_L g7532 ( 
.A(n_7517),
.B(n_7441),
.Y(n_7532)
);

NAND2xp5_ASAP7_75t_L g7533 ( 
.A(n_7481),
.B(n_7524),
.Y(n_7533)
);

NAND2xp5_ASAP7_75t_SL g7534 ( 
.A(n_7488),
.B(n_7403),
.Y(n_7534)
);

NAND2xp5_ASAP7_75t_L g7535 ( 
.A(n_7483),
.B(n_7479),
.Y(n_7535)
);

INVx1_ASAP7_75t_L g7536 ( 
.A(n_7497),
.Y(n_7536)
);

NOR2xp33_ASAP7_75t_L g7537 ( 
.A(n_7482),
.B(n_7412),
.Y(n_7537)
);

NAND2xp5_ASAP7_75t_L g7538 ( 
.A(n_7501),
.B(n_7407),
.Y(n_7538)
);

HB1xp67_ASAP7_75t_L g7539 ( 
.A(n_7497),
.Y(n_7539)
);

AOI22xp33_ASAP7_75t_SL g7540 ( 
.A1(n_7487),
.A2(n_7420),
.B1(n_7454),
.B2(n_7462),
.Y(n_7540)
);

INVx2_ASAP7_75t_SL g7541 ( 
.A(n_7519),
.Y(n_7541)
);

INVx2_ASAP7_75t_L g7542 ( 
.A(n_7523),
.Y(n_7542)
);

NAND2xp5_ASAP7_75t_L g7543 ( 
.A(n_7505),
.B(n_7409),
.Y(n_7543)
);

AOI22xp33_ASAP7_75t_L g7544 ( 
.A1(n_7516),
.A2(n_7466),
.B1(n_7440),
.B2(n_7465),
.Y(n_7544)
);

AND2x2_ASAP7_75t_L g7545 ( 
.A(n_7503),
.B(n_7464),
.Y(n_7545)
);

NAND3xp33_ASAP7_75t_SL g7546 ( 
.A(n_7521),
.B(n_7414),
.C(n_7402),
.Y(n_7546)
);

INVx1_ASAP7_75t_L g7547 ( 
.A(n_7507),
.Y(n_7547)
);

NOR2xp33_ASAP7_75t_L g7548 ( 
.A(n_7502),
.B(n_7390),
.Y(n_7548)
);

INVx1_ASAP7_75t_L g7549 ( 
.A(n_7495),
.Y(n_7549)
);

NAND2xp5_ASAP7_75t_L g7550 ( 
.A(n_7484),
.B(n_7394),
.Y(n_7550)
);

INVx1_ASAP7_75t_L g7551 ( 
.A(n_7489),
.Y(n_7551)
);

INVxp67_ASAP7_75t_L g7552 ( 
.A(n_7509),
.Y(n_7552)
);

NAND2xp5_ASAP7_75t_L g7553 ( 
.A(n_7486),
.B(n_7451),
.Y(n_7553)
);

OR2x2_ASAP7_75t_L g7554 ( 
.A(n_7513),
.B(n_7446),
.Y(n_7554)
);

NAND2xp5_ASAP7_75t_L g7555 ( 
.A(n_7492),
.B(n_7439),
.Y(n_7555)
);

AND2x2_ASAP7_75t_L g7556 ( 
.A(n_7494),
.B(n_7392),
.Y(n_7556)
);

OR2x2_ASAP7_75t_L g7557 ( 
.A(n_7520),
.B(n_7447),
.Y(n_7557)
);

INVx1_ASAP7_75t_SL g7558 ( 
.A(n_7511),
.Y(n_7558)
);

AOI22xp33_ASAP7_75t_L g7559 ( 
.A1(n_7498),
.A2(n_7456),
.B1(n_7404),
.B2(n_7435),
.Y(n_7559)
);

NAND2xp5_ASAP7_75t_L g7560 ( 
.A(n_7485),
.B(n_7469),
.Y(n_7560)
);

INVx1_ASAP7_75t_L g7561 ( 
.A(n_7499),
.Y(n_7561)
);

NAND2xp5_ASAP7_75t_L g7562 ( 
.A(n_7491),
.B(n_7470),
.Y(n_7562)
);

INVx1_ASAP7_75t_L g7563 ( 
.A(n_7514),
.Y(n_7563)
);

INVx1_ASAP7_75t_L g7564 ( 
.A(n_7515),
.Y(n_7564)
);

NOR2x1p5_ASAP7_75t_L g7565 ( 
.A(n_7490),
.B(n_7455),
.Y(n_7565)
);

AND2x2_ASAP7_75t_L g7566 ( 
.A(n_7506),
.B(n_7410),
.Y(n_7566)
);

INVx1_ASAP7_75t_L g7567 ( 
.A(n_7504),
.Y(n_7567)
);

INVx1_ASAP7_75t_L g7568 ( 
.A(n_7496),
.Y(n_7568)
);

OR2x2_ASAP7_75t_L g7569 ( 
.A(n_7527),
.B(n_7426),
.Y(n_7569)
);

NAND2xp5_ASAP7_75t_L g7570 ( 
.A(n_7493),
.B(n_7429),
.Y(n_7570)
);

INVx1_ASAP7_75t_L g7571 ( 
.A(n_7525),
.Y(n_7571)
);

NAND2xp33_ASAP7_75t_L g7572 ( 
.A(n_7518),
.B(n_7388),
.Y(n_7572)
);

AND2x2_ASAP7_75t_L g7573 ( 
.A(n_7522),
.B(n_7478),
.Y(n_7573)
);

INVx1_ASAP7_75t_L g7574 ( 
.A(n_7512),
.Y(n_7574)
);

INVx1_ASAP7_75t_L g7575 ( 
.A(n_7526),
.Y(n_7575)
);

NAND2xp5_ASAP7_75t_L g7576 ( 
.A(n_7526),
.B(n_7411),
.Y(n_7576)
);

INVx2_ASAP7_75t_SL g7577 ( 
.A(n_7508),
.Y(n_7577)
);

OAI221xp5_ASAP7_75t_SL g7578 ( 
.A1(n_7500),
.A2(n_7463),
.B1(n_7389),
.B2(n_7418),
.C(n_7413),
.Y(n_7578)
);

INVx1_ASAP7_75t_L g7579 ( 
.A(n_7526),
.Y(n_7579)
);

INVx1_ASAP7_75t_L g7580 ( 
.A(n_7526),
.Y(n_7580)
);

OAI221xp5_ASAP7_75t_L g7581 ( 
.A1(n_7530),
.A2(n_7448),
.B1(n_7425),
.B2(n_7433),
.C(n_7427),
.Y(n_7581)
);

NAND2xp5_ASAP7_75t_L g7582 ( 
.A(n_7531),
.B(n_7476),
.Y(n_7582)
);

AOI21xp33_ASAP7_75t_L g7583 ( 
.A1(n_7528),
.A2(n_7467),
.B(n_860),
.Y(n_7583)
);

NAND2xp5_ASAP7_75t_L g7584 ( 
.A(n_7577),
.B(n_861),
.Y(n_7584)
);

INVx1_ASAP7_75t_L g7585 ( 
.A(n_7575),
.Y(n_7585)
);

HB1xp67_ASAP7_75t_L g7586 ( 
.A(n_7579),
.Y(n_7586)
);

NAND2xp5_ASAP7_75t_L g7587 ( 
.A(n_7536),
.B(n_861),
.Y(n_7587)
);

INVx1_ASAP7_75t_L g7588 ( 
.A(n_7580),
.Y(n_7588)
);

NAND2xp5_ASAP7_75t_L g7589 ( 
.A(n_7539),
.B(n_862),
.Y(n_7589)
);

INVx1_ASAP7_75t_SL g7590 ( 
.A(n_7545),
.Y(n_7590)
);

AOI211xp5_ASAP7_75t_L g7591 ( 
.A1(n_7578),
.A2(n_864),
.B(n_862),
.C(n_863),
.Y(n_7591)
);

NAND3xp33_ASAP7_75t_L g7592 ( 
.A(n_7530),
.B(n_862),
.C(n_863),
.Y(n_7592)
);

NOR2xp33_ASAP7_75t_L g7593 ( 
.A(n_7534),
.B(n_864),
.Y(n_7593)
);

AOI22xp5_ASAP7_75t_L g7594 ( 
.A1(n_7537),
.A2(n_866),
.B1(n_864),
.B2(n_865),
.Y(n_7594)
);

AND3x2_ASAP7_75t_L g7595 ( 
.A(n_7552),
.B(n_1049),
.C(n_865),
.Y(n_7595)
);

AO221x1_ASAP7_75t_L g7596 ( 
.A1(n_7551),
.A2(n_868),
.B1(n_866),
.B2(n_867),
.C(n_869),
.Y(n_7596)
);

NAND2xp5_ASAP7_75t_SL g7597 ( 
.A(n_7576),
.B(n_867),
.Y(n_7597)
);

OA22x2_ASAP7_75t_L g7598 ( 
.A1(n_7541),
.A2(n_870),
.B1(n_867),
.B2(n_869),
.Y(n_7598)
);

INVxp67_ASAP7_75t_L g7599 ( 
.A(n_7533),
.Y(n_7599)
);

NAND5xp2_ASAP7_75t_L g7600 ( 
.A(n_7544),
.B(n_872),
.C(n_870),
.D(n_871),
.E(n_873),
.Y(n_7600)
);

NAND2xp5_ASAP7_75t_SL g7601 ( 
.A(n_7542),
.B(n_870),
.Y(n_7601)
);

NAND5xp2_ASAP7_75t_L g7602 ( 
.A(n_7559),
.B(n_873),
.C(n_871),
.D(n_872),
.E(n_874),
.Y(n_7602)
);

NAND2xp5_ASAP7_75t_L g7603 ( 
.A(n_7532),
.B(n_871),
.Y(n_7603)
);

NOR2x1_ASAP7_75t_L g7604 ( 
.A(n_7546),
.B(n_872),
.Y(n_7604)
);

OAI21xp33_ASAP7_75t_SL g7605 ( 
.A1(n_7529),
.A2(n_874),
.B(n_875),
.Y(n_7605)
);

INVx2_ASAP7_75t_L g7606 ( 
.A(n_7565),
.Y(n_7606)
);

INVxp67_ASAP7_75t_L g7607 ( 
.A(n_7548),
.Y(n_7607)
);

NAND3xp33_ASAP7_75t_L g7608 ( 
.A(n_7572),
.B(n_874),
.C(n_875),
.Y(n_7608)
);

NAND3xp33_ASAP7_75t_SL g7609 ( 
.A(n_7558),
.B(n_875),
.C(n_876),
.Y(n_7609)
);

OAI21xp33_ASAP7_75t_SL g7610 ( 
.A1(n_7550),
.A2(n_876),
.B(n_877),
.Y(n_7610)
);

NAND5xp2_ASAP7_75t_L g7611 ( 
.A(n_7540),
.B(n_879),
.C(n_877),
.D(n_878),
.E(n_880),
.Y(n_7611)
);

NOR2xp33_ASAP7_75t_L g7612 ( 
.A(n_7574),
.B(n_878),
.Y(n_7612)
);

INVx1_ASAP7_75t_L g7613 ( 
.A(n_7557),
.Y(n_7613)
);

NAND3xp33_ASAP7_75t_L g7614 ( 
.A(n_7568),
.B(n_878),
.C(n_879),
.Y(n_7614)
);

AOI21xp5_ASAP7_75t_L g7615 ( 
.A1(n_7538),
.A2(n_879),
.B(n_880),
.Y(n_7615)
);

AND2x2_ASAP7_75t_L g7616 ( 
.A(n_7590),
.B(n_7556),
.Y(n_7616)
);

INVxp67_ASAP7_75t_L g7617 ( 
.A(n_7612),
.Y(n_7617)
);

INVxp67_ASAP7_75t_L g7618 ( 
.A(n_7593),
.Y(n_7618)
);

INVx1_ASAP7_75t_L g7619 ( 
.A(n_7587),
.Y(n_7619)
);

INVx2_ASAP7_75t_L g7620 ( 
.A(n_7613),
.Y(n_7620)
);

XNOR2xp5_ASAP7_75t_L g7621 ( 
.A(n_7586),
.B(n_7563),
.Y(n_7621)
);

INVx2_ASAP7_75t_L g7622 ( 
.A(n_7585),
.Y(n_7622)
);

NAND3xp33_ASAP7_75t_L g7623 ( 
.A(n_7591),
.B(n_7564),
.C(n_7569),
.Y(n_7623)
);

OR2x2_ASAP7_75t_L g7624 ( 
.A(n_7603),
.B(n_7543),
.Y(n_7624)
);

INVx1_ASAP7_75t_L g7625 ( 
.A(n_7598),
.Y(n_7625)
);

NOR3x1_ASAP7_75t_L g7626 ( 
.A(n_7596),
.B(n_7535),
.C(n_7553),
.Y(n_7626)
);

INVx1_ASAP7_75t_L g7627 ( 
.A(n_7589),
.Y(n_7627)
);

NAND2xp5_ASAP7_75t_L g7628 ( 
.A(n_7595),
.B(n_7566),
.Y(n_7628)
);

NAND4xp25_ASAP7_75t_L g7629 ( 
.A(n_7600),
.B(n_7573),
.C(n_7560),
.D(n_7562),
.Y(n_7629)
);

AOI21xp5_ASAP7_75t_L g7630 ( 
.A1(n_7615),
.A2(n_7555),
.B(n_7570),
.Y(n_7630)
);

INVx1_ASAP7_75t_L g7631 ( 
.A(n_7584),
.Y(n_7631)
);

NAND3xp33_ASAP7_75t_L g7632 ( 
.A(n_7594),
.B(n_7561),
.C(n_7567),
.Y(n_7632)
);

NOR2xp33_ASAP7_75t_L g7633 ( 
.A(n_7583),
.B(n_7554),
.Y(n_7633)
);

NOR3xp33_ASAP7_75t_L g7634 ( 
.A(n_7581),
.B(n_7547),
.C(n_7549),
.Y(n_7634)
);

OAI22xp5_ASAP7_75t_L g7635 ( 
.A1(n_7599),
.A2(n_7571),
.B1(n_882),
.B2(n_880),
.Y(n_7635)
);

NAND3xp33_ASAP7_75t_L g7636 ( 
.A(n_7614),
.B(n_881),
.C(n_882),
.Y(n_7636)
);

NAND2xp5_ASAP7_75t_SL g7637 ( 
.A(n_7588),
.B(n_881),
.Y(n_7637)
);

NAND2xp5_ASAP7_75t_L g7638 ( 
.A(n_7604),
.B(n_881),
.Y(n_7638)
);

NAND4xp25_ASAP7_75t_L g7639 ( 
.A(n_7602),
.B(n_885),
.C(n_883),
.D(n_884),
.Y(n_7639)
);

NAND2xp5_ASAP7_75t_SL g7640 ( 
.A(n_7610),
.B(n_883),
.Y(n_7640)
);

INVx1_ASAP7_75t_SL g7641 ( 
.A(n_7582),
.Y(n_7641)
);

NAND2xp5_ASAP7_75t_SL g7642 ( 
.A(n_7605),
.B(n_884),
.Y(n_7642)
);

AND2x2_ASAP7_75t_L g7643 ( 
.A(n_7606),
.B(n_885),
.Y(n_7643)
);

BUFx2_ASAP7_75t_L g7644 ( 
.A(n_7607),
.Y(n_7644)
);

O2A1O1Ixp5_ASAP7_75t_SL g7645 ( 
.A1(n_7597),
.A2(n_887),
.B(n_885),
.C(n_886),
.Y(n_7645)
);

NAND2xp5_ASAP7_75t_L g7646 ( 
.A(n_7608),
.B(n_888),
.Y(n_7646)
);

NOR2x1_ASAP7_75t_L g7647 ( 
.A(n_7609),
.B(n_888),
.Y(n_7647)
);

NAND4xp25_ASAP7_75t_L g7648 ( 
.A(n_7611),
.B(n_891),
.C(n_889),
.D(n_890),
.Y(n_7648)
);

NAND2xp5_ASAP7_75t_L g7649 ( 
.A(n_7592),
.B(n_1049),
.Y(n_7649)
);

NAND3xp33_ASAP7_75t_L g7650 ( 
.A(n_7601),
.B(n_889),
.C(n_890),
.Y(n_7650)
);

NAND2xp5_ASAP7_75t_L g7651 ( 
.A(n_7590),
.B(n_891),
.Y(n_7651)
);

INVx1_ASAP7_75t_L g7652 ( 
.A(n_7587),
.Y(n_7652)
);

INVx2_ASAP7_75t_L g7653 ( 
.A(n_7613),
.Y(n_7653)
);

OAI221xp5_ASAP7_75t_L g7654 ( 
.A1(n_7591),
.A2(n_893),
.B1(n_891),
.B2(n_892),
.C(n_894),
.Y(n_7654)
);

OAI21xp33_ASAP7_75t_L g7655 ( 
.A1(n_7613),
.A2(n_892),
.B(n_893),
.Y(n_7655)
);

INVx1_ASAP7_75t_L g7656 ( 
.A(n_7587),
.Y(n_7656)
);

AOI22xp5_ASAP7_75t_L g7657 ( 
.A1(n_7613),
.A2(n_895),
.B1(n_892),
.B2(n_894),
.Y(n_7657)
);

OAI22xp5_ASAP7_75t_L g7658 ( 
.A1(n_7613),
.A2(n_896),
.B1(n_894),
.B2(n_895),
.Y(n_7658)
);

AOI211xp5_ASAP7_75t_SL g7659 ( 
.A1(n_7583),
.A2(n_897),
.B(n_895),
.C(n_896),
.Y(n_7659)
);

NAND2xp5_ASAP7_75t_L g7660 ( 
.A(n_7590),
.B(n_1047),
.Y(n_7660)
);

INVx1_ASAP7_75t_L g7661 ( 
.A(n_7616),
.Y(n_7661)
);

AND2x2_ASAP7_75t_L g7662 ( 
.A(n_7643),
.B(n_896),
.Y(n_7662)
);

NAND4xp25_ASAP7_75t_L g7663 ( 
.A(n_7626),
.B(n_899),
.C(n_897),
.D(n_898),
.Y(n_7663)
);

INVx1_ASAP7_75t_L g7664 ( 
.A(n_7651),
.Y(n_7664)
);

AOI21xp5_ASAP7_75t_L g7665 ( 
.A1(n_7637),
.A2(n_898),
.B(n_899),
.Y(n_7665)
);

XOR2x2_ASAP7_75t_L g7666 ( 
.A(n_7621),
.B(n_7623),
.Y(n_7666)
);

OAI22xp5_ASAP7_75t_L g7667 ( 
.A1(n_7641),
.A2(n_901),
.B1(n_899),
.B2(n_900),
.Y(n_7667)
);

XOR2xp5_ASAP7_75t_L g7668 ( 
.A(n_7629),
.B(n_900),
.Y(n_7668)
);

AOI21xp5_ASAP7_75t_L g7669 ( 
.A1(n_7660),
.A2(n_901),
.B(n_902),
.Y(n_7669)
);

OAI22xp5_ASAP7_75t_L g7670 ( 
.A1(n_7620),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_7670)
);

AOI22xp5_ASAP7_75t_L g7671 ( 
.A1(n_7653),
.A2(n_905),
.B1(n_903),
.B2(n_904),
.Y(n_7671)
);

NAND2xp5_ASAP7_75t_SL g7672 ( 
.A(n_7622),
.B(n_903),
.Y(n_7672)
);

NAND2xp5_ASAP7_75t_L g7673 ( 
.A(n_7657),
.B(n_904),
.Y(n_7673)
);

HB1xp67_ASAP7_75t_L g7674 ( 
.A(n_7635),
.Y(n_7674)
);

XNOR2x2_ASAP7_75t_SL g7675 ( 
.A(n_7636),
.B(n_905),
.Y(n_7675)
);

NAND4xp25_ASAP7_75t_L g7676 ( 
.A(n_7633),
.B(n_908),
.C(n_906),
.D(n_907),
.Y(n_7676)
);

OAI22xp5_ASAP7_75t_L g7677 ( 
.A1(n_7632),
.A2(n_908),
.B1(n_906),
.B2(n_907),
.Y(n_7677)
);

AOI22xp5_ASAP7_75t_L g7678 ( 
.A1(n_7634),
.A2(n_909),
.B1(n_907),
.B2(n_908),
.Y(n_7678)
);

INVxp67_ASAP7_75t_L g7679 ( 
.A(n_7649),
.Y(n_7679)
);

INVx1_ASAP7_75t_L g7680 ( 
.A(n_7658),
.Y(n_7680)
);

NAND3xp33_ASAP7_75t_L g7681 ( 
.A(n_7659),
.B(n_909),
.C(n_910),
.Y(n_7681)
);

NOR2xp33_ASAP7_75t_L g7682 ( 
.A(n_7639),
.B(n_910),
.Y(n_7682)
);

NAND3xp33_ASAP7_75t_L g7683 ( 
.A(n_7654),
.B(n_911),
.C(n_912),
.Y(n_7683)
);

NAND3xp33_ASAP7_75t_L g7684 ( 
.A(n_7650),
.B(n_911),
.C(n_912),
.Y(n_7684)
);

INVx1_ASAP7_75t_L g7685 ( 
.A(n_7646),
.Y(n_7685)
);

NAND2xp5_ASAP7_75t_L g7686 ( 
.A(n_7655),
.B(n_912),
.Y(n_7686)
);

INVxp67_ASAP7_75t_L g7687 ( 
.A(n_7647),
.Y(n_7687)
);

INVx1_ASAP7_75t_L g7688 ( 
.A(n_7638),
.Y(n_7688)
);

OAI21xp5_ASAP7_75t_L g7689 ( 
.A1(n_7630),
.A2(n_913),
.B(n_914),
.Y(n_7689)
);

AOI22xp5_ASAP7_75t_L g7690 ( 
.A1(n_7648),
.A2(n_915),
.B1(n_913),
.B2(n_914),
.Y(n_7690)
);

AOI22xp33_ASAP7_75t_L g7691 ( 
.A1(n_7625),
.A2(n_7644),
.B1(n_7652),
.B2(n_7619),
.Y(n_7691)
);

XOR2x2_ASAP7_75t_L g7692 ( 
.A(n_7640),
.B(n_913),
.Y(n_7692)
);

NAND2xp5_ASAP7_75t_L g7693 ( 
.A(n_7656),
.B(n_914),
.Y(n_7693)
);

NAND2xp5_ASAP7_75t_L g7694 ( 
.A(n_7624),
.B(n_915),
.Y(n_7694)
);

OAI21xp5_ASAP7_75t_SL g7695 ( 
.A1(n_7628),
.A2(n_915),
.B(n_916),
.Y(n_7695)
);

OAI22xp33_ASAP7_75t_L g7696 ( 
.A1(n_7627),
.A2(n_918),
.B1(n_916),
.B2(n_917),
.Y(n_7696)
);

AND2x4_ASAP7_75t_L g7697 ( 
.A(n_7631),
.B(n_918),
.Y(n_7697)
);

AOI22xp5_ASAP7_75t_L g7698 ( 
.A1(n_7617),
.A2(n_920),
.B1(n_918),
.B2(n_919),
.Y(n_7698)
);

INVx1_ASAP7_75t_L g7699 ( 
.A(n_7642),
.Y(n_7699)
);

NAND2xp5_ASAP7_75t_SL g7700 ( 
.A(n_7618),
.B(n_919),
.Y(n_7700)
);

HB1xp67_ASAP7_75t_L g7701 ( 
.A(n_7645),
.Y(n_7701)
);

AOI22xp5_ASAP7_75t_L g7702 ( 
.A1(n_7661),
.A2(n_7668),
.B1(n_7682),
.B2(n_7662),
.Y(n_7702)
);

INVx1_ASAP7_75t_L g7703 ( 
.A(n_7677),
.Y(n_7703)
);

INVx1_ASAP7_75t_L g7704 ( 
.A(n_7678),
.Y(n_7704)
);

INVx1_ASAP7_75t_L g7705 ( 
.A(n_7698),
.Y(n_7705)
);

OAI22xp33_ASAP7_75t_L g7706 ( 
.A1(n_7690),
.A2(n_7693),
.B1(n_7663),
.B2(n_7694),
.Y(n_7706)
);

AO22x2_ASAP7_75t_L g7707 ( 
.A1(n_7680),
.A2(n_921),
.B1(n_919),
.B2(n_920),
.Y(n_7707)
);

INVx1_ASAP7_75t_SL g7708 ( 
.A(n_7697),
.Y(n_7708)
);

AOI22xp5_ASAP7_75t_L g7709 ( 
.A1(n_7666),
.A2(n_922),
.B1(n_920),
.B2(n_921),
.Y(n_7709)
);

AOI22xp5_ASAP7_75t_L g7710 ( 
.A1(n_7674),
.A2(n_923),
.B1(n_921),
.B2(n_922),
.Y(n_7710)
);

INVxp67_ASAP7_75t_SL g7711 ( 
.A(n_7696),
.Y(n_7711)
);

INVx1_ASAP7_75t_L g7712 ( 
.A(n_7697),
.Y(n_7712)
);

AOI22xp5_ASAP7_75t_L g7713 ( 
.A1(n_7664),
.A2(n_924),
.B1(n_922),
.B2(n_923),
.Y(n_7713)
);

NOR2x1_ASAP7_75t_L g7714 ( 
.A(n_7681),
.B(n_923),
.Y(n_7714)
);

AOI22xp5_ASAP7_75t_L g7715 ( 
.A1(n_7691),
.A2(n_926),
.B1(n_924),
.B2(n_925),
.Y(n_7715)
);

NOR2xp33_ASAP7_75t_L g7716 ( 
.A(n_7695),
.B(n_924),
.Y(n_7716)
);

AO22x2_ASAP7_75t_L g7717 ( 
.A1(n_7683),
.A2(n_927),
.B1(n_925),
.B2(n_926),
.Y(n_7717)
);

AOI22xp5_ASAP7_75t_L g7718 ( 
.A1(n_7685),
.A2(n_928),
.B1(n_926),
.B2(n_927),
.Y(n_7718)
);

NOR2xp33_ASAP7_75t_L g7719 ( 
.A(n_7686),
.B(n_927),
.Y(n_7719)
);

OAI22xp5_ASAP7_75t_SL g7720 ( 
.A1(n_7684),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.Y(n_7720)
);

OAI22xp5_ASAP7_75t_L g7721 ( 
.A1(n_7687),
.A2(n_930),
.B1(n_928),
.B2(n_929),
.Y(n_7721)
);

AOI22xp5_ASAP7_75t_L g7722 ( 
.A1(n_7699),
.A2(n_931),
.B1(n_929),
.B2(n_930),
.Y(n_7722)
);

INVx2_ASAP7_75t_L g7723 ( 
.A(n_7675),
.Y(n_7723)
);

NOR3xp33_ASAP7_75t_SL g7724 ( 
.A(n_7676),
.B(n_931),
.C(n_932),
.Y(n_7724)
);

NOR4xp25_ASAP7_75t_L g7725 ( 
.A(n_7700),
.B(n_933),
.C(n_931),
.D(n_932),
.Y(n_7725)
);

AOI22xp5_ASAP7_75t_L g7726 ( 
.A1(n_7688),
.A2(n_934),
.B1(n_932),
.B2(n_933),
.Y(n_7726)
);

NOR2x1_ASAP7_75t_L g7727 ( 
.A(n_7673),
.B(n_934),
.Y(n_7727)
);

NAND2xp5_ASAP7_75t_L g7728 ( 
.A(n_7671),
.B(n_935),
.Y(n_7728)
);

NOR2x1_ASAP7_75t_L g7729 ( 
.A(n_7672),
.B(n_935),
.Y(n_7729)
);

NOR4xp25_ASAP7_75t_L g7730 ( 
.A(n_7689),
.B(n_937),
.C(n_935),
.D(n_936),
.Y(n_7730)
);

INVx1_ASAP7_75t_L g7731 ( 
.A(n_7707),
.Y(n_7731)
);

INVx1_ASAP7_75t_L g7732 ( 
.A(n_7707),
.Y(n_7732)
);

OAI31xp33_ASAP7_75t_L g7733 ( 
.A1(n_7719),
.A2(n_7706),
.A3(n_7716),
.B(n_7703),
.Y(n_7733)
);

XOR2x2_ASAP7_75t_L g7734 ( 
.A(n_7702),
.B(n_7692),
.Y(n_7734)
);

INVx1_ASAP7_75t_L g7735 ( 
.A(n_7710),
.Y(n_7735)
);

NOR3xp33_ASAP7_75t_L g7736 ( 
.A(n_7711),
.B(n_7679),
.C(n_7667),
.Y(n_7736)
);

NAND2xp5_ASAP7_75t_L g7737 ( 
.A(n_7715),
.B(n_7669),
.Y(n_7737)
);

NAND2xp5_ASAP7_75t_L g7738 ( 
.A(n_7709),
.B(n_7665),
.Y(n_7738)
);

NAND2xp5_ASAP7_75t_L g7739 ( 
.A(n_7722),
.B(n_7670),
.Y(n_7739)
);

NOR2x1p5_ASAP7_75t_L g7740 ( 
.A(n_7723),
.B(n_7701),
.Y(n_7740)
);

NOR2x1_ASAP7_75t_L g7741 ( 
.A(n_7714),
.B(n_936),
.Y(n_7741)
);

NAND2xp5_ASAP7_75t_L g7742 ( 
.A(n_7718),
.B(n_937),
.Y(n_7742)
);

NAND2xp5_ASAP7_75t_L g7743 ( 
.A(n_7726),
.B(n_937),
.Y(n_7743)
);

NAND2x2_ASAP7_75t_L g7744 ( 
.A(n_7728),
.B(n_938),
.Y(n_7744)
);

INVx1_ASAP7_75t_L g7745 ( 
.A(n_7713),
.Y(n_7745)
);

OR2x2_ASAP7_75t_L g7746 ( 
.A(n_7708),
.B(n_938),
.Y(n_7746)
);

NAND2xp5_ASAP7_75t_L g7747 ( 
.A(n_7721),
.B(n_939),
.Y(n_7747)
);

INVxp67_ASAP7_75t_L g7748 ( 
.A(n_7727),
.Y(n_7748)
);

INVx1_ASAP7_75t_L g7749 ( 
.A(n_7720),
.Y(n_7749)
);

NAND4xp25_ASAP7_75t_L g7750 ( 
.A(n_7704),
.B(n_941),
.C(n_939),
.D(n_940),
.Y(n_7750)
);

NAND2xp5_ASAP7_75t_L g7751 ( 
.A(n_7712),
.B(n_939),
.Y(n_7751)
);

NAND2xp5_ASAP7_75t_SL g7752 ( 
.A(n_7733),
.B(n_7705),
.Y(n_7752)
);

INVx1_ASAP7_75t_L g7753 ( 
.A(n_7751),
.Y(n_7753)
);

NOR2xp67_ASAP7_75t_L g7754 ( 
.A(n_7746),
.B(n_7724),
.Y(n_7754)
);

NAND4xp25_ASAP7_75t_L g7755 ( 
.A(n_7736),
.B(n_7729),
.C(n_7717),
.D(n_7730),
.Y(n_7755)
);

NOR2x1_ASAP7_75t_L g7756 ( 
.A(n_7740),
.B(n_7725),
.Y(n_7756)
);

AOI31xp33_ASAP7_75t_L g7757 ( 
.A1(n_7749),
.A2(n_7739),
.A3(n_7737),
.B(n_7735),
.Y(n_7757)
);

NOR2xp33_ASAP7_75t_L g7758 ( 
.A(n_7748),
.B(n_940),
.Y(n_7758)
);

NAND4xp75_ASAP7_75t_L g7759 ( 
.A(n_7741),
.B(n_942),
.C(n_940),
.D(n_941),
.Y(n_7759)
);

NAND3xp33_ASAP7_75t_SL g7760 ( 
.A(n_7738),
.B(n_941),
.C(n_942),
.Y(n_7760)
);

INVx1_ASAP7_75t_L g7761 ( 
.A(n_7750),
.Y(n_7761)
);

AND2x4_ASAP7_75t_L g7762 ( 
.A(n_7745),
.B(n_943),
.Y(n_7762)
);

OR2x2_ASAP7_75t_L g7763 ( 
.A(n_7734),
.B(n_943),
.Y(n_7763)
);

NAND4xp25_ASAP7_75t_SL g7764 ( 
.A(n_7747),
.B(n_946),
.C(n_944),
.D(n_945),
.Y(n_7764)
);

AND2x4_ASAP7_75t_L g7765 ( 
.A(n_7731),
.B(n_945),
.Y(n_7765)
);

NAND4xp25_ASAP7_75t_SL g7766 ( 
.A(n_7756),
.B(n_7732),
.C(n_7743),
.D(n_7742),
.Y(n_7766)
);

NAND4xp75_ASAP7_75t_L g7767 ( 
.A(n_7752),
.B(n_7744),
.C(n_947),
.D(n_945),
.Y(n_7767)
);

NOR2xp33_ASAP7_75t_L g7768 ( 
.A(n_7757),
.B(n_1047),
.Y(n_7768)
);

NOR2x1_ASAP7_75t_L g7769 ( 
.A(n_7755),
.B(n_946),
.Y(n_7769)
);

INVx2_ASAP7_75t_L g7770 ( 
.A(n_7765),
.Y(n_7770)
);

NAND3x1_ASAP7_75t_L g7771 ( 
.A(n_7768),
.B(n_7761),
.C(n_7769),
.Y(n_7771)
);

HB1xp67_ASAP7_75t_L g7772 ( 
.A(n_7771),
.Y(n_7772)
);

AOI221xp5_ASAP7_75t_L g7773 ( 
.A1(n_7771),
.A2(n_7766),
.B1(n_7753),
.B2(n_7770),
.C(n_7754),
.Y(n_7773)
);

OR3x1_ASAP7_75t_L g7774 ( 
.A(n_7772),
.B(n_7763),
.C(n_7758),
.Y(n_7774)
);

INVx1_ASAP7_75t_L g7775 ( 
.A(n_7773),
.Y(n_7775)
);

INVx1_ASAP7_75t_L g7776 ( 
.A(n_7774),
.Y(n_7776)
);

XNOR2xp5_ASAP7_75t_L g7777 ( 
.A(n_7775),
.B(n_7762),
.Y(n_7777)
);

INVx1_ASAP7_75t_L g7778 ( 
.A(n_7777),
.Y(n_7778)
);

INVx1_ASAP7_75t_L g7779 ( 
.A(n_7778),
.Y(n_7779)
);

AOI22xp5_ASAP7_75t_L g7780 ( 
.A1(n_7779),
.A2(n_7776),
.B1(n_7767),
.B2(n_7760),
.Y(n_7780)
);

NAND2xp5_ASAP7_75t_L g7781 ( 
.A(n_7780),
.B(n_7759),
.Y(n_7781)
);

NAND2xp5_ASAP7_75t_L g7782 ( 
.A(n_7781),
.B(n_7764),
.Y(n_7782)
);

AOI21xp5_ASAP7_75t_L g7783 ( 
.A1(n_7782),
.A2(n_946),
.B(n_947),
.Y(n_7783)
);

NAND2xp5_ASAP7_75t_L g7784 ( 
.A(n_7783),
.B(n_948),
.Y(n_7784)
);

OA331x2_ASAP7_75t_L g7785 ( 
.A1(n_7784),
.A2(n_948),
.A3(n_949),
.B1(n_950),
.B2(n_951),
.B3(n_952),
.C1(n_953),
.Y(n_7785)
);

OAI221xp5_ASAP7_75t_R g7786 ( 
.A1(n_7785),
.A2(n_948),
.B1(n_949),
.B2(n_950),
.C(n_951),
.Y(n_7786)
);

AOI21xp33_ASAP7_75t_L g7787 ( 
.A1(n_7786),
.A2(n_950),
.B(n_951),
.Y(n_7787)
);

AOI211xp5_ASAP7_75t_L g7788 ( 
.A1(n_7787),
.A2(n_955),
.B(n_952),
.C(n_954),
.Y(n_7788)
);


endmodule