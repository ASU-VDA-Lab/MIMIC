module fake_jpeg_28269_n_336 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_336);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_336;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_42),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

AND2x4_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_17),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_48),
.A2(n_60),
.B1(n_17),
.B2(n_18),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_30),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_55),
.B(n_19),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_38),
.A2(n_20),
.B1(n_24),
.B2(n_25),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_18),
.B1(n_34),
.B2(n_35),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_38),
.A2(n_24),
.B1(n_20),
.B2(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g72 ( 
.A(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_66),
.B(n_71),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_47),
.A2(n_46),
.B1(n_39),
.B2(n_44),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_76),
.B1(n_88),
.B2(n_104),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_68),
.B(n_69),
.Y(n_117)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

NOR2x1_ASAP7_75t_R g136 ( 
.A(n_70),
.B(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_27),
.Y(n_71)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_77),
.Y(n_121)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_62),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_79),
.Y(n_127)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_80),
.B(n_82),
.Y(n_128)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_81),
.Y(n_108)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_47),
.B(n_17),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_84),
.A2(n_88),
.B1(n_90),
.B2(n_94),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_47),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_85),
.B(n_91),
.Y(n_135)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_64),
.Y(n_87)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_64),
.A2(n_28),
.B1(n_33),
.B2(n_29),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_32),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_32),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_92),
.B(n_99),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_22),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_53),
.A2(n_28),
.B1(n_33),
.B2(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

AOI32xp33_ASAP7_75t_L g96 ( 
.A1(n_50),
.A2(n_31),
.A3(n_45),
.B1(n_37),
.B2(n_41),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_105),
.C(n_21),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_97),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_98),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_59),
.B(n_29),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_49),
.B(n_29),
.Y(n_102)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_103),
.Y(n_120)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_22),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_106),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_83),
.B1(n_87),
.B2(n_100),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_37),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_70),
.B(n_41),
.C(n_37),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_41),
.C(n_40),
.Y(n_150)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_65),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_134),
.B(n_106),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_139),
.A2(n_151),
.B1(n_114),
.B2(n_18),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_107),
.A2(n_84),
.B1(n_67),
.B2(n_94),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_140),
.A2(n_148),
.B1(n_156),
.B2(n_165),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_118),
.A2(n_72),
.B(n_105),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_141),
.A2(n_143),
.B(n_145),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_107),
.A2(n_78),
.B1(n_100),
.B2(n_30),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_142),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_37),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_144),
.B(n_149),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_131),
.B(n_129),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_146),
.Y(n_191)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_124),
.A2(n_90),
.B1(n_77),
.B2(n_79),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_127),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_111),
.C(n_43),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_120),
.A2(n_23),
.B1(n_35),
.B2(n_34),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g152 ( 
.A(n_133),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_152),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_98),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_155),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_125),
.B(n_135),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_165),
.B(n_136),
.Y(n_168)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_137),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_135),
.A2(n_81),
.B1(n_73),
.B2(n_72),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_160),
.B1(n_166),
.B2(n_130),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_128),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_158),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_108),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_159),
.Y(n_172)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_121),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_110),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_161),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_110),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_162),
.Y(n_179)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_108),
.Y(n_163)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_122),
.B(n_41),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_167),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_136),
.B(n_39),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_168),
.A2(n_192),
.B(n_146),
.Y(n_211)
);

AO21x1_ASAP7_75t_L g173 ( 
.A1(n_165),
.A2(n_143),
.B(n_138),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_173),
.B(n_200),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_141),
.B(n_116),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_174),
.B(n_180),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_175),
.B(n_185),
.C(n_44),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_177),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_116),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_140),
.A2(n_120),
.B1(n_111),
.B2(n_133),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_195),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_134),
.C(n_132),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_109),
.B1(n_126),
.B2(n_123),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_126),
.B1(n_123),
.B2(n_113),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_119),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_188),
.B(n_190),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_189),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_164),
.B(n_149),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_138),
.A2(n_112),
.B(n_113),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_112),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_45),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_119),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_198),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_130),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_144),
.B(n_114),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_198),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_201),
.B(n_208),
.Y(n_236)
);

OAI21xp33_ASAP7_75t_SL g204 ( 
.A1(n_190),
.A2(n_143),
.B(n_19),
.Y(n_204)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_204),
.B(n_205),
.Y(n_251)
);

OAI21xp33_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_23),
.B(n_34),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_176),
.A2(n_167),
.B1(n_163),
.B2(n_23),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_225),
.B1(n_181),
.B2(n_183),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_207),
.Y(n_242)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_188),
.B(n_35),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_210),
.B(n_214),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_211),
.B(n_168),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_213),
.B(n_196),
.Y(n_232)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_170),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_179),
.B(n_159),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_215),
.B(n_216),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_184),
.B(n_159),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_226),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_221),
.B(n_175),
.C(n_194),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_182),
.B(n_159),
.Y(n_222)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_228),
.Y(n_238)
);

NAND2x1_ASAP7_75t_SL g225 ( 
.A(n_176),
.B(n_44),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_197),
.B(n_9),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_227),
.B(n_229),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_181),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_169),
.B(n_21),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_230),
.B(n_217),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_235),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_233),
.B(n_254),
.C(n_219),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_221),
.Y(n_234)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_234),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_241),
.B(n_39),
.Y(n_275)
);

NOR2x1p5_ASAP7_75t_L g244 ( 
.A(n_228),
.B(n_171),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_245),
.B(n_248),
.Y(n_274)
);

INVxp33_ASAP7_75t_SL g246 ( 
.A(n_225),
.Y(n_246)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_220),
.A2(n_171),
.B1(n_177),
.B2(n_196),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_247),
.A2(n_227),
.B1(n_225),
.B2(n_211),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g248 ( 
.A(n_206),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_180),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_219),
.Y(n_267)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_209),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_202),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_220),
.A2(n_185),
.B1(n_173),
.B2(n_174),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_252),
.A2(n_248),
.B1(n_203),
.B2(n_251),
.Y(n_258)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_213),
.B(n_212),
.C(n_202),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_262),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_231),
.A2(n_217),
.B1(n_223),
.B2(n_230),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_260),
.B(n_268),
.Y(n_288)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_261),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_233),
.B(n_214),
.C(n_208),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_264),
.B(n_269),
.C(n_271),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_239),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_265),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_270),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_235),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_247),
.A2(n_224),
.B1(n_200),
.B2(n_193),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_254),
.B(n_193),
.C(n_191),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_21),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_249),
.B(n_43),
.C(n_101),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_246),
.A2(n_39),
.B1(n_43),
.B2(n_2),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_237),
.B1(n_244),
.B2(n_240),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_251),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_243),
.Y(n_276)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_277),
.A2(n_292),
.B1(n_7),
.B2(n_14),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_238),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_293),
.Y(n_306)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_282),
.Y(n_302)
);

XNOR2x1_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_232),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_283),
.A2(n_7),
.B1(n_13),
.B2(n_12),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_274),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_286),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_238),
.B(n_244),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_285),
.Y(n_301)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_275),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_257),
.B(n_0),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_255),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_297),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_291),
.B(n_262),
.C(n_269),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_295),
.B(n_296),
.C(n_305),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_271),
.C(n_267),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_280),
.B(n_260),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_290),
.B(n_273),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_300),
.B(n_303),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_280),
.B(n_7),
.C(n_14),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_11),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_310),
.A2(n_313),
.B1(n_5),
.B2(n_15),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_298),
.B(n_299),
.Y(n_311)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_311),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_281),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_312),
.B(n_315),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_289),
.B1(n_288),
.B2(n_286),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_287),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_285),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_304),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_305),
.A2(n_293),
.B1(n_278),
.B2(n_6),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_5),
.B1(n_15),
.B2(n_9),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_295),
.C(n_296),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_308),
.B(n_294),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_323),
.A2(n_309),
.B(n_314),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_325),
.B(n_326),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_310),
.B(n_316),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_327),
.Y(n_330)
);

OAI321xp33_ASAP7_75t_L g331 ( 
.A1(n_330),
.A2(n_328),
.A3(n_318),
.B1(n_319),
.B2(n_309),
.C(n_324),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_331),
.A2(n_329),
.B(n_4),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_4),
.C(n_8),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_4),
.B(n_8),
.C(n_6),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_3),
.B(n_8),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_15),
.Y(n_336)
);


endmodule