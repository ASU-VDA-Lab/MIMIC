module fake_netlist_6_2404_n_2328 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2328);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2328;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_726;
wire n_2157;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2179;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_2291;
wire n_415;
wire n_830;
wire n_2299;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_1985;
wire n_447;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_2074;
wire n_522;
wire n_2129;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2018;
wire n_2094;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_2058;
wire n_2090;
wire n_405;
wire n_538;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_2108;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_2085;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_407;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_2300;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_577;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_2093;
wire n_483;
wire n_2207;
wire n_1970;
wire n_608;
wire n_261;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_541;
wire n_512;
wire n_2073;
wire n_2273;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_2031;
wire n_354;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_487;
wire n_241;
wire n_2068;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_2193;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2206;
wire n_604;
wire n_2319;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_2096;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_2178;
wire n_950;
wire n_388;
wire n_484;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_2075;
wire n_2194;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_2279;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_673;
wire n_382;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_2148;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_2060;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_2138;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2057;
wire n_2103;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_2231;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2238;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_399;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_2292;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2209;
wire n_2301;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_2025;
wire n_1125;
wire n_970;
wire n_2224;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_2237;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_2115;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_1093;
wire n_418;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_732;
wire n_974;
wire n_2240;
wire n_392;
wire n_2278;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_238;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_1847;
wire n_2052;
wire n_248;
wire n_2302;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_2177;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_2264;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_2220;
wire n_1262;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2164;
wire n_2225;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_2169;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_2244;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2167;
wire n_2084;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_543;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_2310;
wire n_584;
wire n_2141;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2196;
wire n_273;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_550;
wire n_2322;
wire n_275;
wire n_652;
wire n_2154;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_2283;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_2266;
wire n_346;
wire n_1029;
wire n_1447;
wire n_2056;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_262;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_2020;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_2076;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_360;
wire n_1754;
wire n_2149;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2284;
wire n_387;
wire n_2287;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2081;
wire n_2168;
wire n_234;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_576;
wire n_1028;
wire n_2106;
wire n_472;
wire n_270;
wire n_2265;
wire n_414;
wire n_1922;
wire n_563;
wire n_2032;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_854;
wire n_1058;
wire n_2312;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_390;
wire n_1148;
wire n_2188;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_2318;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_2033;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_2071;
wire n_357;
wire n_985;
wire n_2233;
wire n_481;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_2303;
wire n_1619;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_582;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_2215;
wire n_271;
wire n_404;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_540;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_457;
wire n_2223;
wire n_2091;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_2116;
wire n_336;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_43),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_217),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_86),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_22),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_92),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_123),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_207),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_91),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_8),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_99),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_96),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_88),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_63),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_118),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_192),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_185),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_51),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_97),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_41),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_169),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_52),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_115),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_71),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_191),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_37),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_87),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_108),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_63),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_74),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_167),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_205),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_177),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_87),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_67),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_113),
.Y(n_257)
);

BUFx2_ASAP7_75t_L g258 ( 
.A(n_51),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_37),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_125),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_70),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_198),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_93),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_32),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_31),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_187),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_139),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_91),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_133),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_94),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_78),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_39),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_137),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_140),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_175),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_32),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_14),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_174),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_36),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_129),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_40),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_218),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_15),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_203),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_146),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_168),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_78),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_35),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_160),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_153),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_147),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_44),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_4),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_122),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_107),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_28),
.Y(n_300)
);

INVx2_ASAP7_75t_SL g301 ( 
.A(n_95),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_13),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g303 ( 
.A(n_55),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_194),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_159),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_190),
.Y(n_306)
);

BUFx5_ASAP7_75t_L g307 ( 
.A(n_110),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_134),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_161),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_66),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_202),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_17),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_181),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_59),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_173),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_34),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_57),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_73),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_50),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_114),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_94),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_42),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_149),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_75),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_98),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_120),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_33),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_50),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_154),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_162),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_17),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_68),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_2),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_126),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_58),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_136),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_195),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_211),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_89),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_65),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_64),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_23),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_127),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_108),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_88),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_47),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_180),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_109),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_7),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_170),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_103),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_61),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_90),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_111),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_15),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_151),
.Y(n_358)
);

BUFx10_ASAP7_75t_L g359 ( 
.A(n_40),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_206),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_182),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_155),
.Y(n_362)
);

BUFx2_ASAP7_75t_SL g363 ( 
.A(n_82),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_76),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_93),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_47),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_179),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_55),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_74),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_109),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_79),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_82),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_164),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_176),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_13),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_69),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_163),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_53),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_7),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_12),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_76),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_100),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_103),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_59),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_44),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_62),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_1),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_5),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_45),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_145),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_128),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_90),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_52),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_150),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_68),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_99),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_197),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_96),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_213),
.Y(n_400)
);

BUFx10_ASAP7_75t_L g401 ( 
.A(n_112),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_49),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_81),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_143),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_80),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_208),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_105),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_156),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_6),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_102),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_69),
.Y(n_411)
);

BUFx2_ASAP7_75t_SL g412 ( 
.A(n_61),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_30),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_107),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_135),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_105),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_34),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_84),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_178),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_102),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_142),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_165),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_81),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_157),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_60),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_98),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_209),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_4),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_95),
.Y(n_429)
);

BUFx10_ASAP7_75t_L g430 ( 
.A(n_10),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_42),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_370),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_370),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_370),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_220),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_258),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_237),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_370),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_370),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_257),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_280),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_224),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_249),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_370),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_370),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_354),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_225),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_258),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_307),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_226),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_354),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_354),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_354),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_354),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_354),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_249),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_231),
.B(n_241),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_235),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_249),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_249),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_236),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_227),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_227),
.B(n_0),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_324),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_243),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_252),
.Y(n_468)
);

NOR2xp67_ASAP7_75t_L g469 ( 
.A(n_271),
.B(n_0),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_254),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_227),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_266),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_366),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_271),
.B(n_2),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_247),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_294),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_266),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_231),
.B(n_3),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_266),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_232),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_260),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_314),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_262),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_232),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_232),
.Y(n_485)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_301),
.B(n_3),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_300),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_336),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_300),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g490 ( 
.A(n_301),
.B(n_5),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_263),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_270),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_300),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_223),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_338),
.Y(n_495)
);

INVxp67_ASAP7_75t_SL g496 ( 
.A(n_223),
.Y(n_496)
);

BUFx3_ASAP7_75t_L g497 ( 
.A(n_324),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_241),
.B(n_245),
.Y(n_498)
);

INVxp67_ASAP7_75t_L g499 ( 
.A(n_366),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_247),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_239),
.B(n_6),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_230),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_219),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_230),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_245),
.B(n_8),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_234),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_349),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_234),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_398),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_282),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_422),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_286),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_284),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_240),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_289),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_292),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_275),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_240),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_293),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_298),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_304),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_251),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_251),
.Y(n_523)
);

BUFx2_ASAP7_75t_SL g524 ( 
.A(n_324),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_273),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_305),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_275),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_312),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_273),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_281),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_267),
.B(n_9),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_316),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_327),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_246),
.B(n_268),
.Y(n_534)
);

CKINVDCx5p33_ASAP7_75t_R g535 ( 
.A(n_331),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_340),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_246),
.B(n_9),
.Y(n_537)
);

INVxp67_ASAP7_75t_SL g538 ( 
.A(n_268),
.Y(n_538)
);

INVxp33_ASAP7_75t_SL g539 ( 
.A(n_221),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_352),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_281),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_358),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_360),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_307),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_367),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_448),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_448),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_445),
.B(n_267),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_438),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_436),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_453),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_454),
.Y(n_553)
);

INVx3_ASAP7_75t_L g554 ( 
.A(n_447),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_454),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_455),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_444),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_455),
.Y(n_558)
);

CKINVDCx6p67_ASAP7_75t_R g559 ( 
.A(n_512),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_447),
.Y(n_560)
);

BUFx2_ASAP7_75t_L g561 ( 
.A(n_500),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g562 ( 
.A(n_442),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_458),
.B(n_267),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g564 ( 
.A(n_500),
.Y(n_564)
);

BUFx2_ASAP7_75t_L g565 ( 
.A(n_475),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_456),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g567 ( 
.A(n_437),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_456),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_447),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_457),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_457),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_432),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_494),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_449),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_452),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_445),
.B(n_368),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_460),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_433),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_458),
.B(n_400),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_463),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_466),
.B(n_538),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_433),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_434),
.Y(n_584)
);

BUFx6f_ASAP7_75t_L g585 ( 
.A(n_434),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_467),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_R g587 ( 
.A(n_516),
.B(n_374),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_494),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_468),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_502),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_435),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_502),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_443),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_504),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_497),
.B(n_375),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_435),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_504),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_506),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_470),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_476),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_497),
.B(n_391),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g602 ( 
.A(n_486),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_506),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_482),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_508),
.Y(n_606)
);

AND3x2_ASAP7_75t_L g607 ( 
.A(n_478),
.B(n_400),
.C(n_402),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_514),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_497),
.B(n_392),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_475),
.B(n_388),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_439),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_481),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_488),
.Y(n_613)
);

BUFx6f_ASAP7_75t_L g614 ( 
.A(n_439),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_440),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_514),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_R g617 ( 
.A(n_526),
.B(n_404),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_518),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_440),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_R g620 ( 
.A(n_532),
.B(n_406),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_483),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_518),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_441),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_461),
.B(n_400),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_503),
.B(n_277),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_491),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_495),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_492),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_480),
.B(n_274),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_L g630 ( 
.A(n_450),
.B(n_222),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_459),
.B(n_408),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_522),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_498),
.B(n_415),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_480),
.B(n_274),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_561),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_625),
.A2(n_425),
.B1(n_388),
.B2(n_501),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_548),
.B(n_484),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_595),
.B(n_510),
.Y(n_639)
);

AOI22xp33_ASAP7_75t_L g640 ( 
.A1(n_548),
.A2(n_534),
.B1(n_537),
.B2(n_505),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_629),
.B(n_461),
.Y(n_641)
);

INVx4_ASAP7_75t_L g642 ( 
.A(n_572),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_595),
.B(n_513),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_629),
.B(n_462),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_591),
.B(n_441),
.Y(n_645)
);

BUFx10_ASAP7_75t_L g646 ( 
.A(n_625),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_602),
.Y(n_647)
);

NOR2x1p5_ASAP7_75t_L g648 ( 
.A(n_550),
.B(n_465),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g649 ( 
.A(n_565),
.B(n_425),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_554),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_591),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_554),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_554),
.Y(n_653)
);

NAND3x1_ASAP7_75t_L g654 ( 
.A(n_548),
.B(n_465),
.C(n_302),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_577),
.Y(n_656)
);

AND2x6_ASAP7_75t_L g657 ( 
.A(n_591),
.B(n_253),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_554),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_577),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_631),
.B(n_539),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_557),
.B(n_515),
.Y(n_663)
);

AND2x6_ASAP7_75t_L g664 ( 
.A(n_591),
.B(n_253),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_560),
.Y(n_665)
);

INVx4_ASAP7_75t_L g666 ( 
.A(n_572),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_629),
.B(n_462),
.Y(n_667)
);

BUFx10_ASAP7_75t_L g668 ( 
.A(n_574),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_560),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_579),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_560),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_569),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_601),
.B(n_519),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_601),
.B(n_520),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_596),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_596),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_609),
.B(n_521),
.Y(n_677)
);

BUFx3_ASAP7_75t_L g678 ( 
.A(n_611),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_575),
.Y(n_679)
);

INVx4_ASAP7_75t_L g680 ( 
.A(n_572),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_596),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_578),
.B(n_528),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_569),
.Y(n_683)
);

BUFx3_ASAP7_75t_L g684 ( 
.A(n_611),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_631),
.B(n_535),
.Y(n_685)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_619),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_619),
.Y(n_688)
);

BUFx6f_ASAP7_75t_L g689 ( 
.A(n_572),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_619),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_623),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_569),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_609),
.B(n_536),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_581),
.B(n_542),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_R g695 ( 
.A(n_586),
.B(n_543),
.Y(n_695)
);

AND2x6_ASAP7_75t_L g696 ( 
.A(n_611),
.B(n_253),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_572),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_623),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_589),
.B(n_545),
.Y(n_699)
);

INVxp67_ASAP7_75t_SL g700 ( 
.A(n_611),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_602),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_623),
.Y(n_702)
);

BUFx10_ASAP7_75t_L g703 ( 
.A(n_599),
.Y(n_703)
);

BUFx6f_ASAP7_75t_L g704 ( 
.A(n_572),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_612),
.B(n_517),
.Y(n_705)
);

AND2x6_ASAP7_75t_L g706 ( 
.A(n_635),
.B(n_253),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_621),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g708 ( 
.A(n_633),
.B(n_253),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_633),
.B(n_524),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_635),
.B(n_276),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_546),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_572),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_546),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_583),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_R g715 ( 
.A(n_626),
.B(n_533),
.Y(n_715)
);

INVxp67_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_635),
.B(n_276),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_583),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_583),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_582),
.B(n_484),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_576),
.B(n_540),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_582),
.A2(n_531),
.B1(n_499),
.B2(n_473),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_583),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_583),
.B(n_446),
.Y(n_724)
);

INVx4_ASAP7_75t_L g725 ( 
.A(n_583),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_583),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_628),
.B(n_517),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_564),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_547),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_584),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_584),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_547),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_584),
.Y(n_733)
);

INVx1_ASAP7_75t_SL g734 ( 
.A(n_561),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_551),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_584),
.Y(n_736)
);

INVx2_ASAP7_75t_SL g737 ( 
.A(n_607),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_567),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_584),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_551),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_587),
.B(n_527),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_584),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_552),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_617),
.Y(n_744)
);

AND2x6_ASAP7_75t_L g745 ( 
.A(n_563),
.B(n_253),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_630),
.B(n_288),
.Y(n_746)
);

INVx4_ASAP7_75t_L g747 ( 
.A(n_584),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_576),
.B(n_527),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_585),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_585),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_552),
.Y(n_751)
);

BUFx3_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

AO21x2_ASAP7_75t_L g753 ( 
.A1(n_610),
.A2(n_306),
.B(n_288),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_553),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_553),
.Y(n_755)
);

INVx1_ASAP7_75t_SL g756 ( 
.A(n_620),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_549),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

AND2x2_ASAP7_75t_SL g759 ( 
.A(n_563),
.B(n_306),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_573),
.A2(n_499),
.B1(n_259),
.B2(n_285),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_563),
.A2(n_531),
.B1(n_501),
.B2(n_490),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_607),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_573),
.B(n_486),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_588),
.B(n_524),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_585),
.B(n_446),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_562),
.Y(n_766)
);

BUFx8_ASAP7_75t_SL g767 ( 
.A(n_593),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_588),
.B(n_485),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_600),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_590),
.B(n_485),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_585),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_585),
.Y(n_772)
);

BUFx2_ASAP7_75t_L g773 ( 
.A(n_604),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_585),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_590),
.B(n_487),
.Y(n_775)
);

BUFx6f_ASAP7_75t_L g776 ( 
.A(n_614),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_592),
.B(n_487),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_555),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_556),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_556),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_614),
.Y(n_781)
);

INVx4_ASAP7_75t_L g782 ( 
.A(n_614),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_614),
.B(n_451),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_614),
.Y(n_784)
);

INVx4_ASAP7_75t_L g785 ( 
.A(n_614),
.Y(n_785)
);

BUFx4f_ASAP7_75t_L g786 ( 
.A(n_614),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_558),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_615),
.B(n_277),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_558),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_615),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_711),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_685),
.B(n_615),
.Y(n_792)
);

OAI221xp5_ASAP7_75t_L g793 ( 
.A1(n_640),
.A2(n_469),
.B1(n_474),
.B2(n_530),
.C(n_496),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_661),
.B(n_287),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_641),
.B(n_592),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_647),
.B(n_287),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_721),
.B(n_507),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_711),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_767),
.Y(n_799)
);

AND2x6_ASAP7_75t_SL g800 ( 
.A(n_748),
.B(n_291),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_738),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_709),
.B(n_764),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_759),
.A2(n_746),
.B1(n_717),
.B2(n_710),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_647),
.B(n_701),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_759),
.A2(n_746),
.B1(n_717),
.B2(n_710),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_713),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_713),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_720),
.B(n_615),
.Y(n_808)
);

BUFx2_ASAP7_75t_L g809 ( 
.A(n_738),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_729),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_701),
.B(n_509),
.Y(n_811)
);

BUFx6f_ASAP7_75t_L g812 ( 
.A(n_651),
.Y(n_812)
);

AOI21xp5_ASAP7_75t_L g813 ( 
.A1(n_749),
.A2(n_615),
.B(n_580),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_720),
.B(n_615),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_746),
.B(n_511),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_638),
.B(n_615),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_638),
.B(n_563),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_641),
.B(n_496),
.Y(n_818)
);

NOR2xp33_ASAP7_75t_L g819 ( 
.A(n_639),
.B(n_613),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_759),
.B(n_563),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_651),
.B(n_580),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_641),
.B(n_580),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

AND2x6_ASAP7_75t_L g824 ( 
.A(n_710),
.B(n_309),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_641),
.B(n_580),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_710),
.A2(n_624),
.B1(n_580),
.B2(n_309),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_643),
.B(n_627),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_717),
.A2(n_624),
.B1(n_310),
.B2(n_332),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_737),
.A2(n_321),
.B1(n_332),
.B2(n_310),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_737),
.A2(n_421),
.B1(n_427),
.B2(n_419),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_732),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_717),
.A2(n_624),
.B1(n_321),
.B2(n_345),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_732),
.Y(n_833)
);

INVxp67_ASAP7_75t_L g834 ( 
.A(n_728),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_735),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_644),
.B(n_624),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_756),
.B(n_401),
.Y(n_837)
);

INVxp67_ASAP7_75t_L g838 ( 
.A(n_636),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_673),
.B(n_559),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_644),
.B(n_624),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_644),
.B(n_566),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_644),
.B(n_566),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_715),
.Y(n_843)
);

O2A1O1Ixp5_ASAP7_75t_L g844 ( 
.A1(n_700),
.A2(n_570),
.B(n_571),
.C(n_568),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_667),
.B(n_594),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_735),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_SL g847 ( 
.A(n_756),
.B(n_637),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_760),
.A2(n_530),
.B1(n_317),
.B2(n_342),
.C(n_278),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_667),
.B(n_568),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_740),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_740),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_637),
.B(n_401),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_667),
.B(n_489),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_646),
.B(n_401),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_667),
.B(n_570),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_646),
.B(n_401),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_753),
.A2(n_339),
.B1(n_356),
.B2(n_345),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_674),
.B(n_571),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_677),
.B(n_339),
.Y(n_859)
);

INVx5_ASAP7_75t_L g860 ( 
.A(n_657),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_753),
.A2(n_356),
.B1(n_362),
.B2(n_361),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_651),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_753),
.A2(n_361),
.B1(n_378),
.B2(n_362),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_743),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_693),
.B(n_559),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_743),
.Y(n_866)
);

BUFx3_ASAP7_75t_L g867 ( 
.A(n_744),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_753),
.B(n_761),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_751),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_744),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_751),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_679),
.B(n_559),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_754),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_646),
.B(n_250),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_754),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_646),
.B(n_250),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_762),
.B(n_278),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_768),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_755),
.B(n_378),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_695),
.B(n_490),
.Y(n_880)
);

AND2x2_ASAP7_75t_SL g881 ( 
.A(n_708),
.B(n_395),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_755),
.B(n_395),
.Y(n_882)
);

AOI22xp33_ASAP7_75t_L g883 ( 
.A1(n_758),
.A2(n_778),
.B1(n_780),
.B2(n_779),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_758),
.B(n_424),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_762),
.B(n_299),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_778),
.B(n_424),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_779),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_780),
.Y(n_888)
);

AOI22xp33_ASAP7_75t_L g889 ( 
.A1(n_787),
.A2(n_363),
.B1(n_412),
.B2(n_469),
.Y(n_889)
);

AOI22xp33_ASAP7_75t_L g890 ( 
.A1(n_787),
.A2(n_363),
.B1(n_412),
.B2(n_474),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_789),
.Y(n_891)
);

AOI22xp33_ASAP7_75t_L g892 ( 
.A1(n_789),
.A2(n_307),
.B1(n_302),
.B2(n_291),
.Y(n_892)
);

NOR2x2_ASAP7_75t_L g893 ( 
.A(n_649),
.B(n_233),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_722),
.B(n_594),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_645),
.A2(n_598),
.B(n_603),
.C(n_597),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_706),
.A2(n_788),
.B1(n_655),
.B2(n_659),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_678),
.B(n_597),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_636),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_678),
.B(n_598),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_678),
.B(n_603),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_768),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_SL g902 ( 
.A(n_649),
.B(n_668),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_716),
.B(n_299),
.Y(n_903)
);

AOI21x1_ASAP7_75t_L g904 ( 
.A1(n_645),
.A2(n_544),
.B(n_451),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_770),
.B(n_489),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_786),
.A2(n_544),
.B(n_451),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_684),
.B(n_605),
.Y(n_907)
);

INVx2_ASAP7_75t_SL g908 ( 
.A(n_770),
.Y(n_908)
);

INVx3_ASAP7_75t_L g909 ( 
.A(n_684),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_654),
.A2(n_413),
.B1(n_423),
.B2(n_303),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_648),
.A2(n_605),
.B1(n_608),
.B2(n_606),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_786),
.A2(n_544),
.B(n_606),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_665),
.Y(n_913)
);

INVx2_ASAP7_75t_SL g914 ( 
.A(n_775),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_684),
.B(n_608),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_653),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_665),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_653),
.B(n_616),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_653),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_668),
.B(n_616),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_653),
.Y(n_921)
);

NOR2xp67_ASAP7_75t_L g922 ( 
.A(n_724),
.B(n_618),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_655),
.Y(n_923)
);

AOI22xp5_ASAP7_75t_L g924 ( 
.A1(n_654),
.A2(n_634),
.B1(n_632),
.B2(n_622),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_668),
.B(n_618),
.Y(n_925)
);

OAI22xp33_ASAP7_75t_L g926 ( 
.A1(n_734),
.A2(n_342),
.B1(n_317),
.B2(n_320),
.Y(n_926)
);

NOR2xp33_ASAP7_75t_L g927 ( 
.A(n_663),
.B(n_228),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_L g928 ( 
.A(n_697),
.B(n_622),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_682),
.B(n_229),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_734),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_656),
.Y(n_931)
);

NAND2xp33_ASAP7_75t_L g932 ( 
.A(n_706),
.B(n_307),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_706),
.A2(n_307),
.B1(n_373),
.B2(n_371),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_697),
.B(n_632),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_694),
.B(n_238),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_699),
.B(n_242),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_697),
.B(n_634),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_697),
.B(n_307),
.Y(n_938)
);

NOR2xp67_ASAP7_75t_L g939 ( 
.A(n_724),
.B(n_116),
.Y(n_939)
);

INVxp67_ASAP7_75t_L g940 ( 
.A(n_686),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_741),
.B(n_244),
.Y(n_941)
);

NAND2x1_ASAP7_75t_L g942 ( 
.A(n_642),
.B(n_464),
.Y(n_942)
);

INVxp33_ASAP7_75t_L g943 ( 
.A(n_760),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_656),
.Y(n_944)
);

AOI22xp5_ASAP7_75t_L g945 ( 
.A1(n_775),
.A2(n_269),
.B1(n_248),
.B2(n_255),
.Y(n_945)
);

OAI22xp33_ASAP7_75t_L g946 ( 
.A1(n_763),
.A2(n_371),
.B1(n_315),
.B2(n_320),
.Y(n_946)
);

AOI22xp33_ASAP7_75t_L g947 ( 
.A1(n_706),
.A2(n_307),
.B1(n_397),
.B2(n_369),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_733),
.B(n_307),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_659),
.Y(n_949)
);

INVx8_ASAP7_75t_L g950 ( 
.A(n_706),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_648),
.A2(n_727),
.B1(n_705),
.B2(n_777),
.Y(n_951)
);

INVx8_ASAP7_75t_L g952 ( 
.A(n_706),
.Y(n_952)
);

NAND2x1_ASAP7_75t_L g953 ( 
.A(n_642),
.B(n_464),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_733),
.B(n_307),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_660),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_733),
.B(n_493),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_777),
.A2(n_264),
.B1(n_256),
.B2(n_261),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_668),
.B(n_265),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_703),
.B(n_272),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_660),
.Y(n_960)
);

NOR3xp33_ASAP7_75t_L g961 ( 
.A(n_773),
.B(n_493),
.C(n_283),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_773),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_799),
.B(n_757),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_909),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_803),
.B(n_703),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_916),
.Y(n_966)
);

AO221x2_ASAP7_75t_L g967 ( 
.A1(n_829),
.A2(n_926),
.B1(n_946),
.B2(n_328),
.C(n_330),
.Y(n_967)
);

BUFx6f_ASAP7_75t_L g968 ( 
.A(n_812),
.Y(n_968)
);

INVx4_ASAP7_75t_L g969 ( 
.A(n_812),
.Y(n_969)
);

NOR3xp33_ASAP7_75t_SL g970 ( 
.A(n_848),
.B(n_290),
.C(n_279),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_916),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_812),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_950),
.Y(n_973)
);

AND2x6_ASAP7_75t_L g974 ( 
.A(n_924),
.B(n_718),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_L g975 ( 
.A(n_802),
.B(n_765),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_919),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_809),
.Y(n_977)
);

BUFx4f_ASAP7_75t_L g978 ( 
.A(n_824),
.Y(n_978)
);

INVx4_ASAP7_75t_L g979 ( 
.A(n_812),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_898),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_812),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_919),
.Y(n_982)
);

BUFx3_ASAP7_75t_L g983 ( 
.A(n_809),
.Y(n_983)
);

INVx5_ASAP7_75t_L g984 ( 
.A(n_950),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_921),
.Y(n_985)
);

INVx3_ASAP7_75t_L g986 ( 
.A(n_909),
.Y(n_986)
);

AOI21x1_ASAP7_75t_L g987 ( 
.A1(n_922),
.A2(n_765),
.B(n_723),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_909),
.Y(n_988)
);

INVx3_ASAP7_75t_L g989 ( 
.A(n_862),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_801),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_862),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_858),
.B(n_662),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_878),
.B(n_662),
.Y(n_993)
);

INVx1_ASAP7_75t_SL g994 ( 
.A(n_930),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_878),
.B(n_670),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_901),
.B(n_670),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_R g997 ( 
.A(n_799),
.B(n_766),
.Y(n_997)
);

AOI22xp5_ASAP7_75t_L g998 ( 
.A1(n_805),
.A2(n_794),
.B1(n_818),
.B2(n_795),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_901),
.B(n_908),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_921),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_924),
.B(n_718),
.Y(n_1001)
);

INVx2_ASAP7_75t_SL g1002 ( 
.A(n_801),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_808),
.B(n_703),
.Y(n_1003)
);

INVx4_ASAP7_75t_L g1004 ( 
.A(n_862),
.Y(n_1004)
);

NOR2xp33_ASAP7_75t_R g1005 ( 
.A(n_843),
.B(n_769),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_908),
.B(n_675),
.Y(n_1006)
);

BUFx4f_ASAP7_75t_L g1007 ( 
.A(n_824),
.Y(n_1007)
);

AO21x2_ASAP7_75t_L g1008 ( 
.A1(n_868),
.A2(n_723),
.B(n_718),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_818),
.A2(n_707),
.B1(n_706),
.B2(n_719),
.Y(n_1009)
);

HB1xp67_ASAP7_75t_L g1010 ( 
.A(n_838),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_798),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_862),
.Y(n_1012)
);

INVx5_ASAP7_75t_L g1013 ( 
.A(n_950),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_SL g1014 ( 
.A(n_814),
.B(n_703),
.Y(n_1014)
);

AND2x4_ASAP7_75t_L g1015 ( 
.A(n_795),
.B(n_719),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_798),
.Y(n_1016)
);

NOR3xp33_ASAP7_75t_SL g1017 ( 
.A(n_847),
.B(n_296),
.C(n_295),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_806),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_806),
.Y(n_1019)
);

NOR3xp33_ASAP7_75t_SL g1020 ( 
.A(n_815),
.B(n_308),
.C(n_297),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_807),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_914),
.B(n_675),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_807),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_823),
.Y(n_1024)
);

NAND2xp33_ASAP7_75t_SL g1025 ( 
.A(n_943),
.B(n_689),
.Y(n_1025)
);

BUFx4f_ASAP7_75t_L g1026 ( 
.A(n_824),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_862),
.Y(n_1027)
);

INVx2_ASAP7_75t_L g1028 ( 
.A(n_823),
.Y(n_1028)
);

OR2x2_ASAP7_75t_L g1029 ( 
.A(n_877),
.B(n_523),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_950),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_843),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_833),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_795),
.A2(n_706),
.B1(n_742),
.B2(n_719),
.Y(n_1033)
);

NOR3xp33_ASAP7_75t_SL g1034 ( 
.A(n_885),
.B(n_313),
.C(n_311),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_962),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_833),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_792),
.B(n_723),
.Y(n_1037)
);

AOI22xp5_ASAP7_75t_L g1038 ( 
.A1(n_845),
.A2(n_742),
.B1(n_752),
.B2(n_733),
.Y(n_1038)
);

INVx5_ASAP7_75t_L g1039 ( 
.A(n_952),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_846),
.Y(n_1040)
);

BUFx4f_ASAP7_75t_L g1041 ( 
.A(n_824),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_811),
.B(n_319),
.C(n_318),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_846),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_L g1044 ( 
.A1(n_845),
.A2(n_745),
.B1(n_681),
.B2(n_687),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_850),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_914),
.B(n_676),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_850),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_791),
.B(n_676),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_866),
.Y(n_1049)
);

NAND2xp33_ASAP7_75t_R g1050 ( 
.A(n_874),
.B(n_323),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_791),
.B(n_681),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_810),
.B(n_687),
.Y(n_1052)
);

NAND3xp33_ASAP7_75t_SL g1053 ( 
.A(n_910),
.B(n_876),
.C(n_797),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_810),
.B(n_688),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_866),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_867),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_867),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_871),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_871),
.Y(n_1059)
);

BUFx6f_ASAP7_75t_L g1060 ( 
.A(n_952),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_891),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_845),
.B(n_742),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_891),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_793),
.A2(n_690),
.B(n_691),
.C(n_688),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_923),
.Y(n_1065)
);

CKINVDCx16_ASAP7_75t_R g1066 ( 
.A(n_872),
.Y(n_1066)
);

NOR3xp33_ASAP7_75t_SL g1067 ( 
.A(n_837),
.B(n_326),
.C(n_325),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_SL g1068 ( 
.A(n_852),
.B(n_333),
.C(n_329),
.Y(n_1068)
);

AOI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_912),
.A2(n_786),
.B(n_666),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_853),
.B(n_702),
.Y(n_1070)
);

OR2x2_ASAP7_75t_L g1071 ( 
.A(n_940),
.B(n_523),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

NOR2xp67_ASAP7_75t_L g1073 ( 
.A(n_834),
.B(n_690),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_831),
.B(n_691),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_931),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_931),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_952),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_870),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_944),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_944),
.Y(n_1080)
);

HAxp5_ASAP7_75t_L g1081 ( 
.A(n_800),
.B(n_343),
.CON(n_1081),
.SN(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_949),
.Y(n_1082)
);

AOI22x1_ASAP7_75t_L g1083 ( 
.A1(n_831),
.A2(n_730),
.B1(n_739),
.B2(n_784),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_870),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_SL g1085 ( 
.A(n_796),
.B(n_337),
.C(n_335),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_949),
.Y(n_1086)
);

INVxp67_ASAP7_75t_SL g1087 ( 
.A(n_821),
.Y(n_1087)
);

NOR3xp33_ASAP7_75t_SL g1088 ( 
.A(n_902),
.B(n_346),
.C(n_344),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_860),
.B(n_752),
.Y(n_1089)
);

NAND3xp33_ASAP7_75t_SL g1090 ( 
.A(n_910),
.B(n_350),
.C(n_348),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_824),
.A2(n_745),
.B1(n_698),
.B2(n_702),
.Y(n_1091)
);

CKINVDCx8_ASAP7_75t_R g1092 ( 
.A(n_819),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_955),
.Y(n_1093)
);

AND2x4_ASAP7_75t_L g1094 ( 
.A(n_853),
.B(n_752),
.Y(n_1094)
);

NAND3xp33_ASAP7_75t_SL g1095 ( 
.A(n_927),
.B(n_353),
.C(n_351),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_955),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_905),
.B(n_702),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_804),
.B(n_642),
.Y(n_1098)
);

CKINVDCx20_ASAP7_75t_R g1099 ( 
.A(n_827),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_835),
.B(n_698),
.Y(n_1100)
);

INVx4_ASAP7_75t_L g1101 ( 
.A(n_952),
.Y(n_1101)
);

BUFx3_ASAP7_75t_L g1102 ( 
.A(n_835),
.Y(n_1102)
);

BUFx4f_ASAP7_75t_L g1103 ( 
.A(n_824),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_821),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_960),
.Y(n_1105)
);

AND2x6_ASAP7_75t_SL g1106 ( 
.A(n_929),
.B(n_315),
.Y(n_1106)
);

BUFx6f_ASAP7_75t_L g1107 ( 
.A(n_821),
.Y(n_1107)
);

NOR3xp33_ASAP7_75t_SL g1108 ( 
.A(n_903),
.B(n_357),
.C(n_355),
.Y(n_1108)
);

NAND2xp33_ASAP7_75t_SL g1109 ( 
.A(n_820),
.B(n_689),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_824),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_851),
.B(n_730),
.Y(n_1111)
);

HB1xp67_ASAP7_75t_L g1112 ( 
.A(n_905),
.Y(n_1112)
);

NOR3xp33_ASAP7_75t_SL g1113 ( 
.A(n_941),
.B(n_372),
.C(n_364),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_SL g1114 ( 
.A(n_893),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_851),
.B(n_665),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_857),
.A2(n_745),
.B1(n_739),
.B2(n_774),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_893),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_864),
.B(n_730),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_960),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_913),
.Y(n_1120)
);

AOI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_817),
.A2(n_739),
.B1(n_731),
.B2(n_736),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_864),
.Y(n_1122)
);

OAI22xp5_ASAP7_75t_L g1123 ( 
.A1(n_861),
.A2(n_786),
.B1(n_731),
.B2(n_736),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_869),
.B(n_731),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_869),
.Y(n_1125)
);

INVx3_ASAP7_75t_L g1126 ( 
.A(n_913),
.Y(n_1126)
);

INVx3_ASAP7_75t_L g1127 ( 
.A(n_917),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_917),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_873),
.Y(n_1129)
);

NAND2xp33_ASAP7_75t_R g1130 ( 
.A(n_839),
.B(n_376),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_873),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_875),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_865),
.B(n_642),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_880),
.B(n_666),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_SL g1135 ( 
.A(n_816),
.B(n_736),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_945),
.B(n_525),
.Y(n_1136)
);

AND2x4_ASAP7_75t_L g1137 ( 
.A(n_875),
.B(n_750),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_887),
.Y(n_1138)
);

INVx5_ASAP7_75t_L g1139 ( 
.A(n_860),
.Y(n_1139)
);

NAND2xp33_ASAP7_75t_L g1140 ( 
.A(n_863),
.B(n_689),
.Y(n_1140)
);

INVx2_ASAP7_75t_SL g1141 ( 
.A(n_887),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_888),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_888),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_822),
.Y(n_1144)
);

BUFx2_ASAP7_75t_L g1145 ( 
.A(n_951),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_904),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_935),
.B(n_666),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_825),
.A2(n_771),
.B1(n_784),
.B2(n_750),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_859),
.B(n_750),
.Y(n_1149)
);

AND2x6_ASAP7_75t_SL g1150 ( 
.A(n_936),
.B(n_322),
.Y(n_1150)
);

AND3x2_ASAP7_75t_SL g1151 ( 
.A(n_945),
.B(n_359),
.C(n_343),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_883),
.B(n_771),
.Y(n_1152)
);

INVx4_ASAP7_75t_L g1153 ( 
.A(n_860),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_922),
.B(n_771),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_841),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_L g1156 ( 
.A(n_897),
.B(n_899),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_1144),
.A2(n_840),
.B(n_836),
.Y(n_1157)
);

AND2x4_ASAP7_75t_L g1158 ( 
.A(n_1015),
.B(n_920),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_983),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_963),
.Y(n_1160)
);

OAI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_975),
.A2(n_844),
.B(n_842),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1112),
.B(n_894),
.Y(n_1162)
);

OAI21x1_ASAP7_75t_L g1163 ( 
.A1(n_1146),
.A2(n_1083),
.B(n_987),
.Y(n_1163)
);

AO31x2_ASAP7_75t_L g1164 ( 
.A1(n_1123),
.A2(n_895),
.A3(n_882),
.B(n_884),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1132),
.A2(n_886),
.A3(n_879),
.B(n_938),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_980),
.B(n_994),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1146),
.A2(n_904),
.B(n_948),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1072),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1133),
.B(n_1155),
.Y(n_1169)
);

OAI21x1_ASAP7_75t_L g1170 ( 
.A1(n_1146),
.A2(n_954),
.B(n_813),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_1139),
.A2(n_1153),
.B(n_1069),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1139),
.A2(n_906),
.B(n_680),
.Y(n_1172)
);

INVxp67_ASAP7_75t_L g1173 ( 
.A(n_977),
.Y(n_1173)
);

HB1xp67_ASAP7_75t_L g1174 ( 
.A(n_977),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_1155),
.B(n_911),
.Y(n_1175)
);

NOR2x1_ASAP7_75t_SL g1176 ( 
.A(n_973),
.B(n_849),
.Y(n_1176)
);

BUFx12f_ASAP7_75t_L g1177 ( 
.A(n_1056),
.Y(n_1177)
);

OAI21x1_ASAP7_75t_L g1178 ( 
.A1(n_1037),
.A2(n_934),
.B(n_928),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_968),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1072),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1075),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_963),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1037),
.A2(n_1135),
.B(n_1118),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1147),
.B(n_855),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_968),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1135),
.A2(n_937),
.B(n_907),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_998),
.A2(n_1102),
.B1(n_1125),
.B2(n_1145),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_1098),
.B(n_900),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1111),
.A2(n_915),
.B(n_918),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1152),
.A2(n_1070),
.B(n_1156),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_999),
.B(n_889),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1097),
.B(n_890),
.Y(n_1192)
);

BUFx8_ASAP7_75t_SL g1193 ( 
.A(n_1031),
.Y(n_1193)
);

OA21x2_ASAP7_75t_L g1194 ( 
.A1(n_1124),
.A2(n_896),
.B(n_956),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1097),
.B(n_957),
.Y(n_1195)
);

OAI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1070),
.A2(n_1064),
.B(n_1121),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_1139),
.A2(n_680),
.B(n_666),
.Y(n_1197)
);

BUFx2_ASAP7_75t_L g1198 ( 
.A(n_983),
.Y(n_1198)
);

INVx2_ASAP7_75t_SL g1199 ( 
.A(n_990),
.Y(n_1199)
);

CKINVDCx8_ASAP7_75t_R g1200 ( 
.A(n_1031),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_997),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1075),
.Y(n_1202)
);

INVx4_ASAP7_75t_L g1203 ( 
.A(n_973),
.Y(n_1203)
);

AOI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1139),
.A2(n_712),
.B(n_680),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1131),
.A2(n_953),
.B(n_942),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_1139),
.A2(n_712),
.B(n_680),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_L g1207 ( 
.A1(n_1131),
.A2(n_953),
.B(n_942),
.Y(n_1207)
);

OAI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1148),
.A2(n_881),
.B(n_826),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_992),
.B(n_1102),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1153),
.A2(n_1140),
.B(n_984),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1131),
.A2(n_781),
.B(n_774),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1048),
.A2(n_781),
.B(n_774),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1125),
.B(n_957),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1029),
.B(n_828),
.Y(n_1214)
);

BUFx3_ASAP7_75t_L g1215 ( 
.A(n_1057),
.Y(n_1215)
);

INVxp67_ASAP7_75t_SL g1216 ( 
.A(n_968),
.Y(n_1216)
);

OR2x2_ASAP7_75t_L g1217 ( 
.A(n_1029),
.B(n_854),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1132),
.A2(n_781),
.A3(n_784),
.B(n_783),
.Y(n_1218)
);

A2O1A1Ixp33_ASAP7_75t_L g1219 ( 
.A1(n_1053),
.A2(n_1136),
.B(n_970),
.C(n_1129),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1122),
.B(n_925),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_990),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1153),
.A2(n_725),
.B(n_712),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1140),
.A2(n_725),
.B(n_712),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1138),
.B(n_832),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1092),
.B(n_1099),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1092),
.B(n_856),
.Y(n_1226)
);

NOR2xp67_ASAP7_75t_SL g1227 ( 
.A(n_973),
.B(n_860),
.Y(n_1227)
);

OAI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_965),
.A2(n_881),
.B1(n_830),
.B2(n_939),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_973),
.A2(n_726),
.B(n_725),
.Y(n_1229)
);

AOI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1003),
.A2(n_939),
.B(n_783),
.Y(n_1230)
);

OAI21x1_ASAP7_75t_L g1231 ( 
.A1(n_1051),
.A2(n_892),
.B(n_671),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1142),
.B(n_881),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_973),
.A2(n_726),
.B(n_725),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1052),
.A2(n_1074),
.B(n_1054),
.Y(n_1234)
);

O2A1O1Ixp5_ASAP7_75t_L g1235 ( 
.A1(n_1003),
.A2(n_959),
.B(n_958),
.C(n_747),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1143),
.B(n_961),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1141),
.B(n_669),
.Y(n_1237)
);

A2O1A1Ixp33_ASAP7_75t_L g1238 ( 
.A1(n_1136),
.A2(n_932),
.B(n_328),
.C(n_322),
.Y(n_1238)
);

O2A1O1Ixp5_ASAP7_75t_L g1239 ( 
.A1(n_1014),
.A2(n_726),
.B(n_747),
.C(n_782),
.Y(n_1239)
);

AO21x1_ASAP7_75t_L g1240 ( 
.A1(n_1025),
.A2(n_932),
.B(n_334),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1141),
.B(n_669),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1002),
.Y(n_1242)
);

OAI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_1149),
.A2(n_947),
.B(n_933),
.Y(n_1243)
);

AOI221xp5_ASAP7_75t_L g1244 ( 
.A1(n_1090),
.A2(n_416),
.B1(n_377),
.B2(n_379),
.C(n_380),
.Y(n_1244)
);

AOI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1014),
.A2(n_671),
.B(n_669),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1079),
.A2(n_393),
.A3(n_389),
.B(n_387),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1079),
.Y(n_1247)
);

CKINVDCx14_ASAP7_75t_R g1248 ( 
.A(n_997),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_984),
.A2(n_747),
.B(n_726),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1100),
.A2(n_672),
.B(n_671),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_984),
.A2(n_1039),
.B(n_1013),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_1005),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1080),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1035),
.Y(n_1254)
);

AOI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_984),
.A2(n_782),
.B(n_747),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_984),
.A2(n_785),
.B(n_782),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1094),
.A2(n_652),
.B(n_650),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_968),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1002),
.B(n_672),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1013),
.A2(n_785),
.B(n_782),
.Y(n_1260)
);

AOI21xp5_ASAP7_75t_L g1261 ( 
.A1(n_1013),
.A2(n_785),
.B(n_860),
.Y(n_1261)
);

OAI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1154),
.A2(n_683),
.B(n_672),
.Y(n_1262)
);

AOI21xp5_ASAP7_75t_SL g1263 ( 
.A1(n_1101),
.A2(n_785),
.B(n_704),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_1080),
.A2(n_692),
.B(n_683),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1094),
.B(n_1065),
.Y(n_1265)
);

OR2x6_ASAP7_75t_L g1266 ( 
.A(n_1107),
.B(n_689),
.Y(n_1266)
);

INVxp67_ASAP7_75t_SL g1267 ( 
.A(n_972),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1094),
.B(n_683),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1096),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1096),
.A2(n_692),
.B(n_652),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1076),
.B(n_692),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1119),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1013),
.A2(n_704),
.B(n_689),
.Y(n_1273)
);

INVx2_ASAP7_75t_SL g1274 ( 
.A(n_1010),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1082),
.B(n_650),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1119),
.A2(n_652),
.B(n_650),
.Y(n_1276)
);

INVx2_ASAP7_75t_SL g1277 ( 
.A(n_972),
.Y(n_1277)
);

OAI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_965),
.A2(n_776),
.B1(n_772),
.B2(n_714),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1086),
.Y(n_1279)
);

NOR4xp25_ASAP7_75t_L g1280 ( 
.A(n_1095),
.B(n_399),
.C(n_393),
.D(n_431),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1093),
.B(n_658),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_972),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_964),
.A2(n_658),
.B(n_472),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1105),
.Y(n_1284)
);

AO31x2_ASAP7_75t_L g1285 ( 
.A1(n_1011),
.A2(n_330),
.A3(n_334),
.B(n_341),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1011),
.B(n_658),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1016),
.A2(n_472),
.B(n_471),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_964),
.A2(n_477),
.B(n_471),
.Y(n_1288)
);

OAI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1038),
.A2(n_664),
.B(n_657),
.Y(n_1289)
);

OR2x6_ASAP7_75t_L g1290 ( 
.A(n_1107),
.B(n_689),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_964),
.A2(n_479),
.B(n_477),
.Y(n_1291)
);

A2O1A1Ixp33_ASAP7_75t_L g1292 ( 
.A1(n_1025),
.A2(n_341),
.B(n_347),
.C(n_365),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_986),
.Y(n_1293)
);

OAI21x1_ASAP7_75t_L g1294 ( 
.A1(n_986),
.A2(n_479),
.B(n_525),
.Y(n_1294)
);

OAI21xp5_ASAP7_75t_L g1295 ( 
.A1(n_1137),
.A2(n_664),
.B(n_657),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1087),
.A2(n_790),
.B1(n_776),
.B2(n_772),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_986),
.A2(n_541),
.B(n_529),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_988),
.A2(n_541),
.B(n_529),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_988),
.A2(n_428),
.B(n_365),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1023),
.Y(n_1300)
);

AOI21xp33_ASAP7_75t_L g1301 ( 
.A1(n_1050),
.A2(n_429),
.B(n_426),
.Y(n_1301)
);

AOI211x1_ASAP7_75t_L g1302 ( 
.A1(n_993),
.A2(n_396),
.B(n_428),
.C(n_409),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_SL g1303 ( 
.A(n_1107),
.B(n_704),
.Y(n_1303)
);

NOR2x1_ASAP7_75t_SL g1304 ( 
.A(n_1013),
.B(n_704),
.Y(n_1304)
);

AOI221x1_ASAP7_75t_L g1305 ( 
.A1(n_1109),
.A2(n_1134),
.B1(n_1059),
.B2(n_1058),
.C(n_1063),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1023),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_988),
.A2(n_431),
.B(n_369),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1028),
.B(n_343),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1028),
.A2(n_347),
.B(n_373),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1032),
.Y(n_1310)
);

BUFx12f_ASAP7_75t_L g1311 ( 
.A(n_1056),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1032),
.A2(n_387),
.B(n_389),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_972),
.Y(n_1313)
);

AOI211x1_ASAP7_75t_L g1314 ( 
.A1(n_995),
.A2(n_399),
.B(n_409),
.C(n_397),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1039),
.A2(n_790),
.B(n_776),
.Y(n_1315)
);

OAI22x1_ASAP7_75t_L g1316 ( 
.A1(n_1117),
.A2(n_396),
.B1(n_420),
.B2(n_418),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1049),
.A2(n_790),
.B(n_776),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1039),
.A2(n_790),
.B(n_776),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1049),
.A2(n_790),
.B(n_776),
.Y(n_1319)
);

A2O1A1Ixp33_ASAP7_75t_L g1320 ( 
.A1(n_978),
.A2(n_403),
.B(n_381),
.C(n_382),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_SL g1321 ( 
.A(n_1039),
.B(n_704),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_978),
.A2(n_407),
.B(n_383),
.C(n_384),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1055),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1039),
.A2(n_790),
.B(n_772),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_L g1325 ( 
.A(n_1099),
.B(n_1078),
.Y(n_1325)
);

INVx1_ASAP7_75t_SL g1326 ( 
.A(n_1166),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1168),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1268),
.B(n_1015),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1168),
.Y(n_1329)
);

BUFx10_ASAP7_75t_L g1330 ( 
.A(n_1325),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1163),
.A2(n_1061),
.B(n_1055),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1301),
.A2(n_1117),
.B1(n_967),
.B2(n_1114),
.Y(n_1332)
);

OAI21x1_ASAP7_75t_L g1333 ( 
.A1(n_1163),
.A2(n_1061),
.B(n_1019),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1202),
.Y(n_1334)
);

OAI221xp5_ASAP7_75t_L g1335 ( 
.A1(n_1244),
.A2(n_1050),
.B1(n_1130),
.B2(n_1034),
.C(n_1108),
.Y(n_1335)
);

OAI21x1_ASAP7_75t_L g1336 ( 
.A1(n_1317),
.A2(n_1021),
.B(n_1018),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1213),
.A2(n_967),
.B1(n_1114),
.B2(n_974),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1317),
.A2(n_1036),
.B(n_1024),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1187),
.A2(n_967),
.B1(n_1001),
.B2(n_974),
.Y(n_1339)
);

INVx3_ASAP7_75t_SL g1340 ( 
.A(n_1182),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1202),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1269),
.Y(n_1342)
);

OAI21x1_ASAP7_75t_L g1343 ( 
.A1(n_1319),
.A2(n_1043),
.B(n_1040),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1268),
.B(n_1015),
.Y(n_1344)
);

NAND3xp33_ASAP7_75t_SL g1345 ( 
.A(n_1280),
.B(n_1005),
.C(n_1113),
.Y(n_1345)
);

BUFx3_ASAP7_75t_L g1346 ( 
.A(n_1177),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1203),
.B(n_1107),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1319),
.A2(n_1047),
.B(n_1045),
.Y(n_1348)
);

AO21x2_ASAP7_75t_L g1349 ( 
.A1(n_1212),
.A2(n_1008),
.B(n_1009),
.Y(n_1349)
);

OAI21x1_ASAP7_75t_SL g1350 ( 
.A1(n_1240),
.A2(n_1006),
.B(n_996),
.Y(n_1350)
);

INVx3_ASAP7_75t_L g1351 ( 
.A(n_1203),
.Y(n_1351)
);

AND2x2_ASAP7_75t_L g1352 ( 
.A(n_1195),
.B(n_1062),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1166),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1305),
.A2(n_971),
.B(n_966),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1184),
.A2(n_1169),
.B1(n_1209),
.B2(n_1214),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1174),
.Y(n_1356)
);

OA21x2_ASAP7_75t_L g1357 ( 
.A1(n_1212),
.A2(n_982),
.B(n_976),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1217),
.B(n_1066),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1269),
.B(n_1062),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1272),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_SL g1361 ( 
.A1(n_1240),
.A2(n_1046),
.B(n_1022),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1272),
.Y(n_1362)
);

AO21x2_ASAP7_75t_L g1363 ( 
.A1(n_1196),
.A2(n_1008),
.B(n_1033),
.Y(n_1363)
);

INVx2_ASAP7_75t_L g1364 ( 
.A(n_1180),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_L g1365 ( 
.A1(n_1211),
.A2(n_1127),
.B(n_1126),
.Y(n_1365)
);

AO31x2_ASAP7_75t_L g1366 ( 
.A1(n_1292),
.A2(n_985),
.A3(n_1000),
.B(n_1120),
.Y(n_1366)
);

INVx3_ASAP7_75t_L g1367 ( 
.A(n_1203),
.Y(n_1367)
);

OAI21x1_ASAP7_75t_L g1368 ( 
.A1(n_1211),
.A2(n_1262),
.B(n_1250),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1217),
.B(n_1073),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_SL g1370 ( 
.A1(n_1210),
.A2(n_979),
.B(n_969),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1262),
.A2(n_1127),
.B(n_1126),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1158),
.A2(n_974),
.B1(n_1001),
.B2(n_1062),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_SL g1373 ( 
.A(n_1274),
.B(n_1084),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1250),
.A2(n_1127),
.B(n_1126),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1171),
.A2(n_1128),
.B(n_1120),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1181),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1227),
.B(n_969),
.Y(n_1377)
);

AO31x2_ASAP7_75t_L g1378 ( 
.A1(n_1292),
.A2(n_1008),
.A3(n_969),
.B(n_979),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1264),
.A2(n_1128),
.B(n_991),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1264),
.A2(n_1128),
.B(n_991),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1219),
.A2(n_1017),
.B(n_1020),
.C(n_1068),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_1177),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1270),
.A2(n_991),
.B(n_989),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_SL g1384 ( 
.A(n_1200),
.B(n_978),
.Y(n_1384)
);

INVx1_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1270),
.A2(n_1027),
.B(n_989),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1179),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1253),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1188),
.A2(n_1109),
.B(n_1026),
.Y(n_1389)
);

INVx4_ASAP7_75t_SL g1390 ( 
.A(n_1179),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1162),
.B(n_1071),
.Y(n_1391)
);

AND2x4_ASAP7_75t_L g1392 ( 
.A(n_1158),
.B(n_979),
.Y(n_1392)
);

OAI21x1_ASAP7_75t_L g1393 ( 
.A1(n_1297),
.A2(n_1027),
.B(n_989),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1309),
.A2(n_1115),
.B(n_1137),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1158),
.B(n_1004),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1300),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1309),
.A2(n_1312),
.B(n_1183),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1175),
.A2(n_1104),
.B1(n_1007),
.B2(n_1026),
.Y(n_1398)
);

OAI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1297),
.A2(n_1027),
.B(n_1115),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_SL g1400 ( 
.A1(n_1304),
.A2(n_1321),
.B(n_1101),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1293),
.Y(n_1401)
);

O2A1O1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1219),
.A2(n_1081),
.B(n_1042),
.C(n_1088),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1306),
.Y(n_1403)
);

OA21x2_ASAP7_75t_L g1404 ( 
.A1(n_1312),
.A2(n_1137),
.B(n_1116),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1298),
.A2(n_1276),
.B(n_1294),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_1193),
.Y(n_1406)
);

HB1xp67_ASAP7_75t_L g1407 ( 
.A(n_1254),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1310),
.Y(n_1408)
);

INVx2_ASAP7_75t_L g1409 ( 
.A(n_1323),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1271),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1279),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1311),
.Y(n_1412)
);

NAND2x1p5_ASAP7_75t_L g1413 ( 
.A(n_1293),
.B(n_1004),
.Y(n_1413)
);

AOI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1263),
.A2(n_1007),
.B(n_1026),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1226),
.B(n_1071),
.Y(n_1415)
);

OAI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1190),
.A2(n_974),
.B(n_1001),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1284),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1236),
.A2(n_974),
.B1(n_1001),
.B2(n_1110),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1265),
.A2(n_1007),
.B1(n_1041),
.B2(n_1103),
.Y(n_1419)
);

OAI21x1_ASAP7_75t_L g1420 ( 
.A1(n_1298),
.A2(n_1089),
.B(n_1091),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1232),
.A2(n_1041),
.B1(n_1103),
.B2(n_1044),
.Y(n_1421)
);

OR2x2_ASAP7_75t_L g1422 ( 
.A(n_1192),
.B(n_1191),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1276),
.A2(n_1089),
.B(n_974),
.Y(n_1423)
);

AOI221xp5_ASAP7_75t_L g1424 ( 
.A1(n_1316),
.A2(n_1085),
.B1(n_1067),
.B2(n_417),
.C(n_386),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1294),
.A2(n_1001),
.B(n_1041),
.Y(n_1425)
);

OA21x2_ASAP7_75t_L g1426 ( 
.A1(n_1183),
.A2(n_1001),
.B(n_390),
.Y(n_1426)
);

CKINVDCx11_ASAP7_75t_R g1427 ( 
.A(n_1200),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1286),
.Y(n_1428)
);

CKINVDCx5p33_ASAP7_75t_R g1429 ( 
.A(n_1193),
.Y(n_1429)
);

BUFx2_ASAP7_75t_SL g1430 ( 
.A(n_1160),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1228),
.A2(n_1130),
.B(n_1004),
.Y(n_1431)
);

NAND3xp33_ASAP7_75t_L g1432 ( 
.A(n_1302),
.B(n_1151),
.C(n_414),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1173),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1248),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1275),
.Y(n_1435)
);

INVx4_ASAP7_75t_L g1436 ( 
.A(n_1266),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1220),
.A2(n_1308),
.B1(n_1316),
.B2(n_1242),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1220),
.B(n_981),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1281),
.Y(n_1439)
);

NAND2x1p5_ASAP7_75t_L g1440 ( 
.A(n_1293),
.B(n_1101),
.Y(n_1440)
);

OAI21x1_ASAP7_75t_L g1441 ( 
.A1(n_1245),
.A2(n_1103),
.B(n_981),
.Y(n_1441)
);

OA21x2_ASAP7_75t_L g1442 ( 
.A1(n_1234),
.A2(n_385),
.B(n_394),
.Y(n_1442)
);

INVxp67_ASAP7_75t_L g1443 ( 
.A(n_1274),
.Y(n_1443)
);

AOI22x1_ASAP7_75t_L g1444 ( 
.A1(n_1161),
.A2(n_1110),
.B1(n_981),
.B2(n_1012),
.Y(n_1444)
);

AOI221xp5_ASAP7_75t_L g1445 ( 
.A1(n_1314),
.A2(n_405),
.B1(n_410),
.B2(n_1151),
.C(n_1106),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_L g1446 ( 
.A1(n_1224),
.A2(n_1208),
.B1(n_1199),
.B2(n_1238),
.Y(n_1446)
);

INVx4_ASAP7_75t_L g1447 ( 
.A(n_1266),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1266),
.B(n_981),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1237),
.Y(n_1449)
);

A2O1A1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1235),
.A2(n_1110),
.B(n_1150),
.C(n_1077),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1160),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1308),
.B(n_1081),
.Y(n_1452)
);

OAI21x1_ASAP7_75t_L g1453 ( 
.A1(n_1288),
.A2(n_1012),
.B(n_1110),
.Y(n_1453)
);

OR2x6_ASAP7_75t_L g1454 ( 
.A(n_1266),
.B(n_1012),
.Y(n_1454)
);

BUFx6f_ASAP7_75t_L g1455 ( 
.A(n_1179),
.Y(n_1455)
);

AOI21xp33_ASAP7_75t_SL g1456 ( 
.A1(n_1225),
.A2(n_10),
.B(n_11),
.Y(n_1456)
);

AO21x2_ASAP7_75t_L g1457 ( 
.A1(n_1230),
.A2(n_1012),
.B(n_745),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1241),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1288),
.A2(n_1077),
.B(n_1060),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1291),
.A2(n_1077),
.B(n_1060),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1238),
.B(n_1030),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1199),
.A2(n_1077),
.B1(n_1060),
.B2(n_1030),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1291),
.A2(n_1060),
.B(n_1030),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1170),
.A2(n_1030),
.B(n_772),
.Y(n_1464)
);

OAI211xp5_ASAP7_75t_SL g1465 ( 
.A1(n_1320),
.A2(n_430),
.B(n_411),
.C(n_359),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1285),
.Y(n_1466)
);

BUFx12f_ASAP7_75t_L g1467 ( 
.A(n_1311),
.Y(n_1467)
);

HB1xp67_ASAP7_75t_L g1468 ( 
.A(n_1198),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1170),
.A2(n_772),
.B(n_714),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1167),
.A2(n_772),
.B(n_714),
.Y(n_1470)
);

INVx2_ASAP7_75t_SL g1471 ( 
.A(n_1215),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1167),
.A2(n_714),
.B(n_704),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1221),
.B(n_745),
.Y(n_1473)
);

OAI21xp5_ASAP7_75t_L g1474 ( 
.A1(n_1157),
.A2(n_745),
.B(n_657),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1159),
.A2(n_343),
.B1(n_359),
.B2(n_411),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1164),
.B(n_1259),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1164),
.B(n_359),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1215),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1285),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1164),
.B(n_411),
.Y(n_1480)
);

OAI21x1_ASAP7_75t_L g1481 ( 
.A1(n_1283),
.A2(n_1178),
.B(n_1186),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1218),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1159),
.Y(n_1483)
);

OAI21x1_ASAP7_75t_L g1484 ( 
.A1(n_1283),
.A2(n_714),
.B(n_745),
.Y(n_1484)
);

OR2x2_ASAP7_75t_L g1485 ( 
.A(n_1165),
.B(n_11),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1285),
.Y(n_1486)
);

OAI21x1_ASAP7_75t_L g1487 ( 
.A1(n_1178),
.A2(n_714),
.B(n_745),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1165),
.B(n_12),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1182),
.Y(n_1489)
);

BUFx16f_ASAP7_75t_R g1490 ( 
.A(n_1248),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1285),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1186),
.A2(n_696),
.B(n_664),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1285),
.Y(n_1493)
);

A2O1A1Ixp33_ASAP7_75t_L g1494 ( 
.A1(n_1320),
.A2(n_430),
.B(n_411),
.C(n_19),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1218),
.Y(n_1495)
);

AND2x6_ASAP7_75t_L g1496 ( 
.A(n_1179),
.B(n_117),
.Y(n_1496)
);

AOI22xp33_ASAP7_75t_L g1497 ( 
.A1(n_1252),
.A2(n_430),
.B1(n_664),
.B2(n_657),
.Y(n_1497)
);

OAI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1231),
.A2(n_696),
.B(n_664),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1234),
.A2(n_696),
.B(n_664),
.Y(n_1499)
);

O2A1O1Ixp33_ASAP7_75t_SL g1500 ( 
.A1(n_1322),
.A2(n_172),
.B(n_121),
.C(n_124),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1231),
.A2(n_696),
.B(n_664),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1223),
.A2(n_696),
.B(n_664),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1246),
.Y(n_1503)
);

AOI21xp5_ASAP7_75t_L g1504 ( 
.A1(n_1263),
.A2(n_696),
.B(n_657),
.Y(n_1504)
);

NAND2x1_ASAP7_75t_L g1505 ( 
.A(n_1400),
.B(n_1290),
.Y(n_1505)
);

BUFx2_ASAP7_75t_SL g1506 ( 
.A(n_1451),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1411),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1391),
.A2(n_1201),
.B1(n_1252),
.B2(n_1290),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1414),
.A2(n_1251),
.B(n_1176),
.Y(n_1509)
);

INVx1_ASAP7_75t_SL g1510 ( 
.A(n_1326),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1415),
.A2(n_1201),
.B1(n_1322),
.B2(n_1290),
.Y(n_1511)
);

OAI22xp5_ASAP7_75t_L g1512 ( 
.A1(n_1339),
.A2(n_1290),
.B1(n_1216),
.B2(n_1258),
.Y(n_1512)
);

INVx8_ASAP7_75t_L g1513 ( 
.A(n_1448),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1452),
.B(n_1246),
.Y(n_1514)
);

AOI22xp33_ASAP7_75t_L g1515 ( 
.A1(n_1335),
.A2(n_430),
.B1(n_1243),
.B2(n_1194),
.Y(n_1515)
);

BUFx2_ASAP7_75t_L g1516 ( 
.A(n_1478),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1452),
.B(n_1246),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1353),
.Y(n_1518)
);

BUFx2_ASAP7_75t_L g1519 ( 
.A(n_1478),
.Y(n_1519)
);

O2A1O1Ixp33_ASAP7_75t_L g1520 ( 
.A1(n_1456),
.A2(n_1303),
.B(n_1278),
.C(n_1289),
.Y(n_1520)
);

NAND2xp33_ASAP7_75t_SL g1521 ( 
.A(n_1416),
.B(n_1185),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_L g1522 ( 
.A(n_1358),
.B(n_1303),
.Y(n_1522)
);

INVx4_ASAP7_75t_L g1523 ( 
.A(n_1448),
.Y(n_1523)
);

AOI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1389),
.A2(n_1324),
.B(n_1318),
.Y(n_1524)
);

OR2x6_ASAP7_75t_L g1525 ( 
.A(n_1448),
.B(n_1299),
.Y(n_1525)
);

AOI22xp5_ASAP7_75t_L g1526 ( 
.A1(n_1345),
.A2(n_1267),
.B1(n_1313),
.B2(n_1282),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1445),
.A2(n_1194),
.B1(n_1189),
.B2(n_1257),
.Y(n_1527)
);

BUFx8_ASAP7_75t_SL g1528 ( 
.A(n_1406),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_SL g1529 ( 
.A1(n_1496),
.A2(n_1307),
.B1(n_1299),
.B2(n_1194),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1436),
.Y(n_1530)
);

AOI22xp33_ASAP7_75t_L g1531 ( 
.A1(n_1465),
.A2(n_1189),
.B1(n_1307),
.B2(n_1313),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1432),
.A2(n_1277),
.B1(n_1282),
.B2(n_1185),
.Y(n_1532)
);

AOI22xp33_ASAP7_75t_L g1533 ( 
.A1(n_1432),
.A2(n_1337),
.B1(n_1332),
.B2(n_1355),
.Y(n_1533)
);

OAI21xp33_ASAP7_75t_SL g1534 ( 
.A1(n_1418),
.A2(n_1207),
.B(n_1205),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1411),
.Y(n_1535)
);

AND2x4_ASAP7_75t_L g1536 ( 
.A(n_1328),
.B(n_1277),
.Y(n_1536)
);

AOI221xp5_ASAP7_75t_L g1537 ( 
.A1(n_1402),
.A2(n_1296),
.B1(n_1295),
.B2(n_1239),
.C(n_1172),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1328),
.B(n_1185),
.Y(n_1538)
);

INVxp67_ASAP7_75t_L g1539 ( 
.A(n_1407),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1422),
.B(n_1165),
.Y(n_1540)
);

BUFx2_ASAP7_75t_L g1541 ( 
.A(n_1468),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1417),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1422),
.B(n_1165),
.Y(n_1543)
);

CKINVDCx6p67_ASAP7_75t_R g1544 ( 
.A(n_1427),
.Y(n_1544)
);

AOI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1477),
.A2(n_1480),
.B1(n_1431),
.B2(n_1424),
.Y(n_1545)
);

BUFx3_ASAP7_75t_L g1546 ( 
.A(n_1471),
.Y(n_1546)
);

AO21x2_ASAP7_75t_L g1547 ( 
.A1(n_1431),
.A2(n_1287),
.B(n_1315),
.Y(n_1547)
);

AO32x2_ASAP7_75t_L g1548 ( 
.A1(n_1446),
.A2(n_1246),
.A3(n_1165),
.B1(n_1218),
.B2(n_1164),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1342),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1417),
.Y(n_1550)
);

BUFx2_ASAP7_75t_L g1551 ( 
.A(n_1356),
.Y(n_1551)
);

BUFx2_ASAP7_75t_R g1552 ( 
.A(n_1406),
.Y(n_1552)
);

OAI21x1_ASAP7_75t_L g1553 ( 
.A1(n_1368),
.A2(n_1207),
.B(n_1205),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1376),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1471),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1437),
.A2(n_1273),
.B1(n_1222),
.B2(n_1197),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1496),
.A2(n_16),
.B1(n_18),
.B2(n_19),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1344),
.B(n_1359),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1352),
.B(n_1359),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1369),
.B(n_1218),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1352),
.B(n_1449),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1366),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1433),
.Y(n_1563)
);

AND2x4_ASAP7_75t_L g1564 ( 
.A(n_1392),
.B(n_1261),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1433),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1381),
.A2(n_657),
.B1(n_696),
.B2(n_1255),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1438),
.B(n_16),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_L g1568 ( 
.A1(n_1477),
.A2(n_1260),
.B1(n_1256),
.B2(n_1249),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1436),
.Y(n_1569)
);

CKINVDCx11_ASAP7_75t_R g1570 ( 
.A(n_1490),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1436),
.Y(n_1571)
);

OAI22xp33_ASAP7_75t_SL g1572 ( 
.A1(n_1384),
.A2(n_18),
.B1(n_20),
.B2(n_21),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_1342),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1372),
.A2(n_1206),
.B1(n_1204),
.B2(n_1233),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1376),
.Y(n_1575)
);

OAI21x1_ASAP7_75t_L g1576 ( 
.A1(n_1368),
.A2(n_1229),
.B(n_696),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1400),
.A2(n_183),
.B(n_216),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1385),
.Y(n_1578)
);

NAND3xp33_ASAP7_75t_L g1579 ( 
.A(n_1456),
.B(n_20),
.C(n_21),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1430),
.B(n_22),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1385),
.Y(n_1581)
);

CKINVDCx5p33_ASAP7_75t_R g1582 ( 
.A(n_1429),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1480),
.A2(n_657),
.B1(n_24),
.B2(n_25),
.Y(n_1583)
);

OAI22xp5_ASAP7_75t_L g1584 ( 
.A1(n_1443),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_1584)
);

AOI221xp5_ASAP7_75t_L g1585 ( 
.A1(n_1494),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.C(n_29),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1449),
.B(n_26),
.Y(n_1586)
);

NAND2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1436),
.B(n_214),
.Y(n_1587)
);

BUFx6f_ASAP7_75t_L g1588 ( 
.A(n_1387),
.Y(n_1588)
);

OAI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1333),
.A2(n_212),
.B(n_210),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1496),
.A2(n_1384),
.B1(n_1430),
.B2(n_1330),
.Y(n_1590)
);

OAI22x1_ASAP7_75t_L g1591 ( 
.A1(n_1444),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1388),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1373),
.A2(n_1340),
.B1(n_1450),
.B2(n_1489),
.Y(n_1593)
);

OAI22xp5_ASAP7_75t_L g1594 ( 
.A1(n_1340),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_1594)
);

CKINVDCx6p67_ASAP7_75t_R g1595 ( 
.A(n_1340),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1360),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1350),
.A2(n_204),
.B(n_201),
.Y(n_1597)
);

AOI22xp33_ASAP7_75t_L g1598 ( 
.A1(n_1485),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_1598)
);

HB1xp67_ASAP7_75t_L g1599 ( 
.A(n_1366),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1483),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1396),
.Y(n_1601)
);

BUFx12f_ASAP7_75t_L g1602 ( 
.A(n_1467),
.Y(n_1602)
);

NAND2xp33_ASAP7_75t_R g1603 ( 
.A(n_1404),
.B(n_200),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1396),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1403),
.Y(n_1605)
);

AOI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1350),
.A2(n_38),
.B(n_43),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1421),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_1607)
);

INVx4_ASAP7_75t_SL g1608 ( 
.A(n_1496),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1475),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1609)
);

AOI22xp33_ASAP7_75t_L g1610 ( 
.A1(n_1485),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1447),
.Y(n_1611)
);

OAI21xp33_ASAP7_75t_L g1612 ( 
.A1(n_1488),
.A2(n_54),
.B(n_57),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1330),
.B(n_1392),
.Y(n_1613)
);

CKINVDCx5p33_ASAP7_75t_R g1614 ( 
.A(n_1429),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1448),
.A2(n_58),
.B1(n_60),
.B2(n_62),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1458),
.B(n_64),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1330),
.B(n_65),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1458),
.B(n_66),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1392),
.B(n_193),
.Y(n_1619)
);

AOI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1361),
.A2(n_67),
.B(n_70),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1403),
.Y(n_1621)
);

AOI222xp33_ASAP7_75t_L g1622 ( 
.A1(n_1467),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.C1(n_77),
.C2(n_79),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_L g1623 ( 
.A1(n_1488),
.A2(n_72),
.B1(n_77),
.B2(n_80),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1364),
.B(n_83),
.Y(n_1624)
);

NAND2xp33_ASAP7_75t_SL g1625 ( 
.A(n_1447),
.B(n_83),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1435),
.B(n_84),
.Y(n_1626)
);

AO31x2_ASAP7_75t_L g1627 ( 
.A1(n_1503),
.A2(n_85),
.A3(n_86),
.B(n_89),
.Y(n_1627)
);

OAI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1435),
.A2(n_85),
.B1(n_92),
.B2(n_97),
.C1(n_100),
.C2(n_101),
.Y(n_1628)
);

AOI22xp33_ASAP7_75t_L g1629 ( 
.A1(n_1476),
.A2(n_101),
.B1(n_104),
.B2(n_106),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1360),
.Y(n_1630)
);

BUFx2_ASAP7_75t_L g1631 ( 
.A(n_1434),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1448),
.A2(n_104),
.B1(n_106),
.B2(n_119),
.Y(n_1632)
);

AO31x2_ASAP7_75t_L g1633 ( 
.A1(n_1503),
.A2(n_130),
.A3(n_131),
.B(n_132),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1439),
.B(n_189),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1447),
.Y(n_1635)
);

INVx8_ASAP7_75t_L g1636 ( 
.A(n_1454),
.Y(n_1636)
);

AO21x2_ASAP7_75t_L g1637 ( 
.A1(n_1361),
.A2(n_1481),
.B(n_1333),
.Y(n_1637)
);

OA21x2_ASAP7_75t_L g1638 ( 
.A1(n_1331),
.A2(n_138),
.B(n_141),
.Y(n_1638)
);

OAI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1331),
.A2(n_144),
.B(n_148),
.Y(n_1639)
);

OAI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1497),
.A2(n_1398),
.B1(n_1346),
.B2(n_1382),
.C(n_1412),
.Y(n_1640)
);

BUFx3_ASAP7_75t_L g1641 ( 
.A(n_1346),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1434),
.Y(n_1642)
);

AO31x2_ASAP7_75t_L g1643 ( 
.A1(n_1466),
.A2(n_152),
.A3(n_158),
.B(n_166),
.Y(n_1643)
);

AOI222xp33_ASAP7_75t_L g1644 ( 
.A1(n_1330),
.A2(n_186),
.B1(n_1382),
.B2(n_1412),
.C1(n_1346),
.C2(n_1496),
.Y(n_1644)
);

AOI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1392),
.A2(n_1395),
.B1(n_1461),
.B2(n_1412),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1408),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_SL g1647 ( 
.A1(n_1496),
.A2(n_1444),
.B1(n_1382),
.B2(n_1363),
.Y(n_1647)
);

AND2x6_ASAP7_75t_SL g1648 ( 
.A(n_1473),
.B(n_1395),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1408),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1395),
.B(n_1447),
.Y(n_1650)
);

AND2x4_ASAP7_75t_SL g1651 ( 
.A(n_1395),
.B(n_1454),
.Y(n_1651)
);

INVx6_ASAP7_75t_L g1652 ( 
.A(n_1390),
.Y(n_1652)
);

HB1xp67_ASAP7_75t_L g1653 ( 
.A(n_1366),
.Y(n_1653)
);

AND2x4_ASAP7_75t_L g1654 ( 
.A(n_1390),
.B(n_1454),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1476),
.A2(n_1496),
.B1(n_1363),
.B2(n_1439),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1409),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1410),
.B(n_1461),
.Y(n_1657)
);

AND2x4_ASAP7_75t_L g1658 ( 
.A(n_1390),
.B(n_1454),
.Y(n_1658)
);

INVx2_ASAP7_75t_SL g1659 ( 
.A(n_1387),
.Y(n_1659)
);

AO31x2_ASAP7_75t_L g1660 ( 
.A1(n_1466),
.A2(n_1493),
.A3(n_1491),
.B(n_1486),
.Y(n_1660)
);

OR2x6_ASAP7_75t_L g1661 ( 
.A(n_1454),
.B(n_1347),
.Y(n_1661)
);

CKINVDCx6p67_ASAP7_75t_R g1662 ( 
.A(n_1387),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1327),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1419),
.A2(n_1363),
.B(n_1474),
.Y(n_1664)
);

OR2x2_ASAP7_75t_L g1665 ( 
.A(n_1327),
.B(n_1329),
.Y(n_1665)
);

CKINVDCx6p67_ASAP7_75t_R g1666 ( 
.A(n_1387),
.Y(n_1666)
);

AOI22xp33_ASAP7_75t_SL g1667 ( 
.A1(n_1404),
.A2(n_1410),
.B1(n_1425),
.B2(n_1428),
.Y(n_1667)
);

AOI22xp5_ASAP7_75t_L g1668 ( 
.A1(n_1428),
.A2(n_1462),
.B1(n_1500),
.B2(n_1401),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1329),
.A2(n_1334),
.B1(n_1362),
.B2(n_1341),
.Y(n_1669)
);

OAI22xp5_ASAP7_75t_L g1670 ( 
.A1(n_1377),
.A2(n_1347),
.B1(n_1362),
.B2(n_1334),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_L g1671 ( 
.A1(n_1479),
.A2(n_1491),
.B1(n_1486),
.B2(n_1493),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1347),
.B(n_1425),
.Y(n_1672)
);

AND2x4_ASAP7_75t_L g1673 ( 
.A(n_1390),
.B(n_1401),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1341),
.B(n_1401),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1387),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1479),
.A2(n_1354),
.B1(n_1495),
.B2(n_1482),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1366),
.Y(n_1677)
);

AND2x4_ASAP7_75t_L g1678 ( 
.A(n_1401),
.B(n_1455),
.Y(n_1678)
);

OAI21x1_ASAP7_75t_L g1679 ( 
.A1(n_1464),
.A2(n_1481),
.B(n_1469),
.Y(n_1679)
);

AOI22xp33_ASAP7_75t_L g1680 ( 
.A1(n_1354),
.A2(n_1426),
.B1(n_1404),
.B2(n_1394),
.Y(n_1680)
);

OAI21x1_ASAP7_75t_L g1681 ( 
.A1(n_1464),
.A2(n_1469),
.B(n_1405),
.Y(n_1681)
);

AOI21xp33_ASAP7_75t_L g1682 ( 
.A1(n_1426),
.A2(n_1349),
.B(n_1354),
.Y(n_1682)
);

BUFx2_ASAP7_75t_SL g1683 ( 
.A(n_1455),
.Y(n_1683)
);

INVx2_ASAP7_75t_SL g1684 ( 
.A(n_1455),
.Y(n_1684)
);

NOR2xp33_ASAP7_75t_L g1685 ( 
.A(n_1413),
.B(n_1455),
.Y(n_1685)
);

AO21x2_ASAP7_75t_L g1686 ( 
.A1(n_1470),
.A2(n_1472),
.B(n_1349),
.Y(n_1686)
);

AND2x4_ASAP7_75t_L g1687 ( 
.A(n_1455),
.B(n_1351),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1366),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1354),
.B(n_1413),
.Y(n_1689)
);

AND2x4_ASAP7_75t_L g1690 ( 
.A(n_1351),
.B(n_1367),
.Y(n_1690)
);

AOI22xp5_ASAP7_75t_L g1691 ( 
.A1(n_1622),
.A2(n_1367),
.B1(n_1351),
.B2(n_1426),
.Y(n_1691)
);

AOI221xp5_ASAP7_75t_SL g1692 ( 
.A1(n_1629),
.A2(n_1504),
.B1(n_1367),
.B2(n_1351),
.C(n_1442),
.Y(n_1692)
);

NOR2x1_ASAP7_75t_R g1693 ( 
.A(n_1570),
.B(n_1602),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1585),
.A2(n_1426),
.B1(n_1394),
.B2(n_1404),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1561),
.B(n_1413),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_L g1696 ( 
.A(n_1522),
.B(n_1442),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1557),
.A2(n_1442),
.B1(n_1377),
.B2(n_1440),
.Y(n_1697)
);

OAI221xp5_ASAP7_75t_L g1698 ( 
.A1(n_1557),
.A2(n_1442),
.B1(n_1377),
.B2(n_1440),
.C(n_1367),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1559),
.B(n_1378),
.Y(n_1699)
);

INVx2_ASAP7_75t_SL g1700 ( 
.A(n_1641),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1612),
.A2(n_1394),
.B1(n_1349),
.B2(n_1357),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1598),
.A2(n_1394),
.B1(n_1357),
.B2(n_1397),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1598),
.A2(n_1357),
.B1(n_1397),
.B2(n_1370),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1518),
.B(n_1514),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1518),
.B(n_1378),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1533),
.A2(n_1440),
.B1(n_1357),
.B2(n_1397),
.Y(n_1706)
);

CKINVDCx6p67_ASAP7_75t_R g1707 ( 
.A(n_1544),
.Y(n_1707)
);

INVx2_ASAP7_75t_L g1708 ( 
.A(n_1554),
.Y(n_1708)
);

AO31x2_ASAP7_75t_L g1709 ( 
.A1(n_1664),
.A2(n_1397),
.A3(n_1470),
.B(n_1472),
.Y(n_1709)
);

HB1xp67_ASAP7_75t_L g1710 ( 
.A(n_1551),
.Y(n_1710)
);

BUFx6f_ASAP7_75t_L g1711 ( 
.A(n_1652),
.Y(n_1711)
);

OAI22xp5_ASAP7_75t_L g1712 ( 
.A1(n_1533),
.A2(n_1499),
.B1(n_1370),
.B2(n_1378),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1629),
.A2(n_1499),
.B(n_1338),
.C(n_1343),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1528),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_L g1715 ( 
.A1(n_1610),
.A2(n_1623),
.B1(n_1579),
.B2(n_1609),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_L g1716 ( 
.A(n_1545),
.B(n_1499),
.C(n_1378),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1535),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1650),
.B(n_1378),
.Y(n_1718)
);

A2O1A1Ixp33_ASAP7_75t_L g1719 ( 
.A1(n_1545),
.A2(n_1423),
.B(n_1441),
.C(n_1420),
.Y(n_1719)
);

AOI221xp5_ASAP7_75t_L g1720 ( 
.A1(n_1607),
.A2(n_1457),
.B1(n_1338),
.B2(n_1343),
.C(n_1348),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1522),
.A2(n_1499),
.B1(n_1423),
.B2(n_1441),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1558),
.B(n_1399),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1610),
.A2(n_1336),
.B(n_1348),
.C(n_1375),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1542),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1623),
.A2(n_1457),
.B1(n_1399),
.B2(n_1375),
.Y(n_1725)
);

AOI221xp5_ASAP7_75t_L g1726 ( 
.A1(n_1584),
.A2(n_1457),
.B1(n_1336),
.B2(n_1374),
.C(n_1487),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1628),
.A2(n_1374),
.B1(n_1487),
.B2(n_1371),
.C(n_1498),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1550),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1628),
.A2(n_1371),
.B1(n_1501),
.B2(n_1498),
.C(n_1393),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1640),
.A2(n_1420),
.B1(n_1453),
.B2(n_1463),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1510),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1625),
.A2(n_1463),
.B(n_1460),
.C(n_1459),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1575),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1517),
.B(n_1501),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_SL g1735 ( 
.A1(n_1590),
.A2(n_1460),
.B1(n_1459),
.B2(n_1453),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1578),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1606),
.A2(n_1393),
.B1(n_1379),
.B2(n_1380),
.C(n_1383),
.Y(n_1737)
);

AOI21xp5_ASAP7_75t_L g1738 ( 
.A1(n_1509),
.A2(n_1484),
.B(n_1365),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1644),
.A2(n_1379),
.B1(n_1380),
.B2(n_1365),
.Y(n_1739)
);

A2O1A1Ixp33_ASAP7_75t_L g1740 ( 
.A1(n_1625),
.A2(n_1502),
.B(n_1405),
.C(n_1492),
.Y(n_1740)
);

HB1xp67_ASAP7_75t_L g1741 ( 
.A(n_1516),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1594),
.A2(n_1383),
.B1(n_1386),
.B2(n_1502),
.Y(n_1742)
);

OAI22xp5_ASAP7_75t_SL g1743 ( 
.A1(n_1590),
.A2(n_1386),
.B1(n_1492),
.B2(n_1484),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1620),
.A2(n_1615),
.B1(n_1572),
.B2(n_1583),
.C(n_1567),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1652),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1583),
.A2(n_1567),
.B1(n_1515),
.B2(n_1632),
.Y(n_1746)
);

OR2x6_ASAP7_75t_L g1747 ( 
.A(n_1513),
.B(n_1636),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1515),
.A2(n_1591),
.B1(n_1626),
.B2(n_1586),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1617),
.B(n_1538),
.Y(n_1749)
);

BUFx2_ASAP7_75t_L g1750 ( 
.A(n_1519),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1508),
.B(n_1657),
.Y(n_1751)
);

OAI211xp5_ASAP7_75t_SL g1752 ( 
.A1(n_1539),
.A2(n_1563),
.B(n_1580),
.C(n_1565),
.Y(n_1752)
);

INVx8_ASAP7_75t_L g1753 ( 
.A(n_1513),
.Y(n_1753)
);

AOI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1593),
.A2(n_1511),
.B1(n_1508),
.B2(n_1506),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1581),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1539),
.A2(n_1616),
.B(n_1618),
.C(n_1532),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1532),
.A2(n_1526),
.B1(n_1563),
.B2(n_1577),
.C(n_1531),
.Y(n_1757)
);

CKINVDCx5p33_ASAP7_75t_R g1758 ( 
.A(n_1528),
.Y(n_1758)
);

AOI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1520),
.A2(n_1657),
.B1(n_1600),
.B2(n_1541),
.C(n_1655),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1624),
.A2(n_1570),
.B1(n_1631),
.B2(n_1595),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1619),
.A2(n_1521),
.B1(n_1537),
.B2(n_1536),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1592),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1619),
.A2(n_1521),
.B1(n_1560),
.B2(n_1527),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_SL g1764 ( 
.A1(n_1513),
.A2(n_1636),
.B1(n_1587),
.B2(n_1641),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1527),
.A2(n_1634),
.B1(n_1540),
.B2(n_1543),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1655),
.A2(n_1597),
.B1(n_1613),
.B2(n_1647),
.Y(n_1766)
);

AND2x2_ASAP7_75t_L g1767 ( 
.A(n_1650),
.B(n_1645),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1647),
.A2(n_1555),
.B1(n_1546),
.B2(n_1668),
.Y(n_1768)
);

AOI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1613),
.A2(n_1642),
.B1(n_1564),
.B2(n_1587),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1601),
.Y(n_1770)
);

AOI222xp33_ASAP7_75t_L g1771 ( 
.A1(n_1608),
.A2(n_1646),
.B1(n_1656),
.B2(n_1621),
.C1(n_1605),
.C2(n_1604),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1649),
.B(n_1549),
.Y(n_1772)
);

AOI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1597),
.A2(n_1546),
.B1(n_1555),
.B2(n_1608),
.Y(n_1773)
);

AOI22xp33_ASAP7_75t_L g1774 ( 
.A1(n_1608),
.A2(n_1564),
.B1(n_1663),
.B2(n_1636),
.Y(n_1774)
);

OAI211xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1531),
.A2(n_1667),
.B(n_1682),
.C(n_1534),
.Y(n_1775)
);

OAI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1556),
.A2(n_1603),
.B1(n_1566),
.B2(n_1568),
.C(n_1524),
.Y(n_1776)
);

AOI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1669),
.A2(n_1653),
.B1(n_1562),
.B2(n_1599),
.C(n_1677),
.Y(n_1777)
);

AOI221xp5_ASAP7_75t_L g1778 ( 
.A1(n_1669),
.A2(n_1653),
.B1(n_1562),
.B2(n_1599),
.C(n_1512),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1673),
.Y(n_1779)
);

OAI211xp5_ASAP7_75t_L g1780 ( 
.A1(n_1667),
.A2(n_1529),
.B(n_1680),
.C(n_1671),
.Y(n_1780)
);

OA21x2_ASAP7_75t_L g1781 ( 
.A1(n_1680),
.A2(n_1681),
.B(n_1679),
.Y(n_1781)
);

INVx3_ASAP7_75t_L g1782 ( 
.A(n_1652),
.Y(n_1782)
);

AOI21xp5_ASAP7_75t_L g1783 ( 
.A1(n_1505),
.A2(n_1574),
.B(n_1568),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1651),
.B(n_1674),
.Y(n_1784)
);

CKINVDCx5p33_ASAP7_75t_R g1785 ( 
.A(n_1582),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_L g1786 ( 
.A1(n_1523),
.A2(n_1630),
.B1(n_1596),
.B2(n_1573),
.Y(n_1786)
);

NOR2x1_ASAP7_75t_R g1787 ( 
.A(n_1614),
.B(n_1552),
.Y(n_1787)
);

OAI211xp5_ASAP7_75t_SL g1788 ( 
.A1(n_1671),
.A2(n_1529),
.B(n_1689),
.C(n_1676),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1660),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1523),
.A2(n_1654),
.B1(n_1658),
.B2(n_1603),
.Y(n_1790)
);

AOI221xp5_ASAP7_75t_L g1791 ( 
.A1(n_1670),
.A2(n_1688),
.B1(n_1676),
.B2(n_1685),
.C(n_1569),
.Y(n_1791)
);

AOI221x1_ASAP7_75t_SL g1792 ( 
.A1(n_1627),
.A2(n_1658),
.B1(n_1685),
.B2(n_1673),
.C(n_1678),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1665),
.Y(n_1793)
);

OR2x2_ASAP7_75t_L g1794 ( 
.A(n_1661),
.B(n_1569),
.Y(n_1794)
);

AND2x4_ASAP7_75t_L g1795 ( 
.A(n_1661),
.B(n_1571),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1661),
.A2(n_1525),
.B1(n_1530),
.B2(n_1635),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1525),
.A2(n_1530),
.B1(n_1611),
.B2(n_1635),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1690),
.B(n_1687),
.Y(n_1798)
);

AND2x4_ASAP7_75t_L g1799 ( 
.A(n_1571),
.B(n_1611),
.Y(n_1799)
);

OAI211xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1675),
.A2(n_1684),
.B(n_1659),
.C(n_1648),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1525),
.A2(n_1547),
.B1(n_1638),
.B2(n_1690),
.Y(n_1801)
);

HB1xp67_ASAP7_75t_L g1802 ( 
.A(n_1687),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1675),
.B(n_1627),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1588),
.Y(n_1804)
);

OAI21xp33_ASAP7_75t_SL g1805 ( 
.A1(n_1589),
.A2(n_1639),
.B(n_1672),
.Y(n_1805)
);

OAI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1576),
.A2(n_1553),
.B(n_1638),
.Y(n_1806)
);

OAI211xp5_ASAP7_75t_L g1807 ( 
.A1(n_1638),
.A2(n_1627),
.B(n_1643),
.C(n_1633),
.Y(n_1807)
);

AOI21xp33_ASAP7_75t_L g1808 ( 
.A1(n_1547),
.A2(n_1637),
.B(n_1672),
.Y(n_1808)
);

AOI221xp5_ASAP7_75t_L g1809 ( 
.A1(n_1637),
.A2(n_1588),
.B1(n_1683),
.B2(n_1627),
.C(n_1686),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1643),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1588),
.A2(n_1672),
.B1(n_1643),
.B2(n_1633),
.Y(n_1811)
);

AOI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1588),
.A2(n_1686),
.B1(n_1643),
.B2(n_1633),
.C(n_1548),
.Y(n_1812)
);

AND2x4_ASAP7_75t_L g1813 ( 
.A(n_1633),
.B(n_1666),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_SL g1814 ( 
.A1(n_1548),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1548),
.A2(n_1053),
.B1(n_794),
.B2(n_1301),
.C(n_848),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1548),
.Y(n_1816)
);

AOI222xp33_ASAP7_75t_L g1817 ( 
.A1(n_1662),
.A2(n_1053),
.B1(n_1090),
.B2(n_852),
.C1(n_848),
.C2(n_794),
.Y(n_1817)
);

OA21x2_ASAP7_75t_L g1818 ( 
.A1(n_1682),
.A2(n_1664),
.B(n_1368),
.Y(n_1818)
);

OAI221xp5_ASAP7_75t_L g1819 ( 
.A1(n_1622),
.A2(n_797),
.B1(n_1092),
.B2(n_661),
.C(n_721),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_SL g1820 ( 
.A1(n_1579),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1518),
.Y(n_1821)
);

AOI222xp33_ASAP7_75t_L g1822 ( 
.A1(n_1585),
.A2(n_1053),
.B1(n_1090),
.B2(n_852),
.C1(n_848),
.C2(n_794),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1561),
.B(n_1353),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1507),
.Y(n_1824)
);

INVxp33_ASAP7_75t_L g1825 ( 
.A(n_1541),
.Y(n_1825)
);

HB1xp67_ASAP7_75t_L g1826 ( 
.A(n_1518),
.Y(n_1826)
);

OR2x2_ASAP7_75t_L g1827 ( 
.A(n_1518),
.B(n_1514),
.Y(n_1827)
);

OAI221xp5_ASAP7_75t_L g1828 ( 
.A1(n_1622),
.A2(n_797),
.B1(n_1092),
.B2(n_661),
.C(n_721),
.Y(n_1828)
);

AOI221xp5_ASAP7_75t_L g1829 ( 
.A1(n_1585),
.A2(n_1053),
.B1(n_794),
.B2(n_1301),
.C(n_848),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_SL g1830 ( 
.A1(n_1579),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1830)
);

INVx1_ASAP7_75t_SL g1831 ( 
.A(n_1510),
.Y(n_1831)
);

OAI21x1_ASAP7_75t_L g1832 ( 
.A1(n_1509),
.A2(n_1524),
.B(n_1553),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1561),
.B(n_1353),
.Y(n_1833)
);

AOI22xp33_ASAP7_75t_SL g1834 ( 
.A1(n_1579),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1834)
);

AOI22xp33_ASAP7_75t_L g1835 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1835)
);

AOI222xp33_ASAP7_75t_L g1836 ( 
.A1(n_1585),
.A2(n_1053),
.B1(n_1090),
.B2(n_852),
.C1(n_848),
.C2(n_794),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1837)
);

OAI22xp33_ASAP7_75t_L g1838 ( 
.A1(n_1579),
.A2(n_1130),
.B1(n_1050),
.B2(n_1092),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1559),
.B(n_1558),
.Y(n_1839)
);

AOI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1533),
.A2(n_1092),
.B1(n_1099),
.B2(n_1332),
.Y(n_1841)
);

AOI22xp33_ASAP7_75t_L g1842 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1843)
);

AOI22xp33_ASAP7_75t_L g1844 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1844)
);

AOI22xp33_ASAP7_75t_SL g1845 ( 
.A1(n_1579),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_SL g1846 ( 
.A1(n_1579),
.A2(n_797),
.B1(n_1335),
.B2(n_1099),
.Y(n_1846)
);

BUFx6f_ASAP7_75t_L g1847 ( 
.A(n_1652),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1533),
.A2(n_1092),
.B1(n_1099),
.B2(n_1332),
.Y(n_1848)
);

OAI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1545),
.A2(n_797),
.B(n_661),
.Y(n_1849)
);

OAI22xp33_ASAP7_75t_L g1850 ( 
.A1(n_1579),
.A2(n_1130),
.B1(n_1050),
.B2(n_1092),
.Y(n_1850)
);

AOI22xp33_ASAP7_75t_L g1851 ( 
.A1(n_1622),
.A2(n_1053),
.B1(n_1585),
.B2(n_1612),
.Y(n_1851)
);

BUFx6f_ASAP7_75t_L g1852 ( 
.A(n_1652),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1541),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1533),
.A2(n_1053),
.B(n_1402),
.C(n_797),
.Y(n_1854)
);

NOR2xp33_ASAP7_75t_L g1855 ( 
.A(n_1731),
.B(n_1831),
.Y(n_1855)
);

AO31x2_ASAP7_75t_L g1856 ( 
.A1(n_1706),
.A2(n_1810),
.A3(n_1696),
.B(n_1712),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1699),
.B(n_1718),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1783),
.B(n_1738),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1718),
.B(n_1734),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1718),
.B(n_1803),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1789),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1705),
.B(n_1704),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1708),
.Y(n_1863)
);

BUFx3_ASAP7_75t_L g1864 ( 
.A(n_1795),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1827),
.B(n_1821),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1696),
.B(n_1826),
.Y(n_1866)
);

BUFx6f_ASAP7_75t_L g1867 ( 
.A(n_1781),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1733),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1733),
.Y(n_1869)
);

OAI33xp33_ASAP7_75t_L g1870 ( 
.A1(n_1838),
.A2(n_1850),
.A3(n_1848),
.B1(n_1841),
.B2(n_1752),
.B3(n_1823),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1819),
.A2(n_1828),
.B1(n_1851),
.B2(n_1837),
.Y(n_1871)
);

OAI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1849),
.A2(n_1835),
.B1(n_1851),
.B2(n_1837),
.C(n_1840),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1710),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1755),
.Y(n_1874)
);

NOR4xp25_ASAP7_75t_SL g1875 ( 
.A(n_1815),
.B(n_1854),
.C(n_1800),
.D(n_1744),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1762),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1781),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1717),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1724),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1793),
.B(n_1728),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1736),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1816),
.B(n_1812),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1770),
.Y(n_1883)
);

AND2x2_ASAP7_75t_L g1884 ( 
.A(n_1722),
.B(n_1781),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1818),
.B(n_1709),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1716),
.B(n_1741),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1835),
.A2(n_1840),
.B1(n_1844),
.B2(n_1843),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1824),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1765),
.B(n_1751),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1807),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1765),
.B(n_1792),
.Y(n_1891)
);

BUFx2_ASAP7_75t_L g1892 ( 
.A(n_1813),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1751),
.B(n_1811),
.Y(n_1893)
);

INVx3_ASAP7_75t_L g1894 ( 
.A(n_1795),
.Y(n_1894)
);

INVx2_ASAP7_75t_L g1895 ( 
.A(n_1709),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1776),
.A2(n_1723),
.B(n_1732),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1713),
.A2(n_1697),
.B(n_1698),
.Y(n_1897)
);

INVx1_ASAP7_75t_SL g1898 ( 
.A(n_1750),
.Y(n_1898)
);

INVx2_ASAP7_75t_SL g1899 ( 
.A(n_1794),
.Y(n_1899)
);

INVxp67_ASAP7_75t_SL g1900 ( 
.A(n_1809),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1766),
.B(n_1767),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1766),
.B(n_1796),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1796),
.B(n_1839),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1709),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1709),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1772),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1778),
.B(n_1763),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1842),
.A2(n_1844),
.B1(n_1843),
.B2(n_1746),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1763),
.B(n_1814),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1777),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1813),
.Y(n_1911)
);

INVxp67_ASAP7_75t_SL g1912 ( 
.A(n_1797),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1813),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1788),
.Y(n_1914)
);

OA21x2_ASAP7_75t_L g1915 ( 
.A1(n_1692),
.A2(n_1808),
.B(n_1832),
.Y(n_1915)
);

OAI222xp33_ASAP7_75t_L g1916 ( 
.A1(n_1842),
.A2(n_1746),
.B1(n_1715),
.B2(n_1754),
.C1(n_1691),
.C2(n_1830),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1818),
.B(n_1801),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1833),
.B(n_1759),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1695),
.B(n_1791),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1748),
.B(n_1771),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1818),
.Y(n_1921)
);

INVx3_ASAP7_75t_L g1922 ( 
.A(n_1799),
.Y(n_1922)
);

INVx1_ASAP7_75t_SL g1923 ( 
.A(n_1804),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1780),
.B(n_1802),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1749),
.B(n_1702),
.Y(n_1925)
);

INVx2_ASAP7_75t_L g1926 ( 
.A(n_1735),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1721),
.Y(n_1927)
);

BUFx2_ASAP7_75t_L g1928 ( 
.A(n_1805),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1753),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1730),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1719),
.B(n_1747),
.Y(n_1931)
);

AND2x2_ASAP7_75t_L g1932 ( 
.A(n_1702),
.B(n_1784),
.Y(n_1932)
);

INVxp67_ASAP7_75t_L g1933 ( 
.A(n_1768),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1748),
.B(n_1701),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1806),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1701),
.B(n_1756),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1801),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1775),
.Y(n_1938)
);

NAND2x1p5_ASAP7_75t_L g1939 ( 
.A(n_1769),
.B(n_1700),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1786),
.B(n_1773),
.Y(n_1940)
);

AO31x2_ASAP7_75t_L g1941 ( 
.A1(n_1740),
.A2(n_1703),
.A3(n_1720),
.B(n_1694),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1703),
.Y(n_1942)
);

AOI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1829),
.A2(n_1715),
.B1(n_1836),
.B2(n_1822),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1743),
.Y(n_1944)
);

BUFx2_ASAP7_75t_L g1945 ( 
.A(n_1779),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1798),
.Y(n_1946)
);

INVx2_ASAP7_75t_L g1947 ( 
.A(n_1747),
.Y(n_1947)
);

INVx2_ASAP7_75t_L g1948 ( 
.A(n_1757),
.Y(n_1948)
);

OAI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1820),
.A2(n_1834),
.B1(n_1846),
.B2(n_1845),
.C(n_1817),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1873),
.Y(n_1950)
);

OAI22xp5_ASAP7_75t_L g1951 ( 
.A1(n_1943),
.A2(n_1761),
.B1(n_1790),
.B2(n_1760),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1914),
.B(n_1825),
.Y(n_1952)
);

INVx1_ASAP7_75t_SL g1953 ( 
.A(n_1898),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1872),
.A2(n_1761),
.B1(n_1764),
.B2(n_1774),
.Y(n_1954)
);

NAND2xp5_ASAP7_75t_L g1955 ( 
.A(n_1866),
.B(n_1853),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1866),
.B(n_1786),
.Y(n_1956)
);

AND2x2_ASAP7_75t_L g1957 ( 
.A(n_1857),
.B(n_1773),
.Y(n_1957)
);

OAI22xp5_ASAP7_75t_L g1958 ( 
.A1(n_1887),
.A2(n_1760),
.B1(n_1774),
.B2(n_1694),
.Y(n_1958)
);

AOI22xp33_ASAP7_75t_L g1959 ( 
.A1(n_1872),
.A2(n_1725),
.B1(n_1707),
.B2(n_1753),
.Y(n_1959)
);

NOR2x1_ASAP7_75t_L g1960 ( 
.A(n_1886),
.B(n_1782),
.Y(n_1960)
);

AOI22xp5_ASAP7_75t_L g1961 ( 
.A1(n_1908),
.A2(n_1782),
.B1(n_1711),
.B2(n_1847),
.Y(n_1961)
);

OAI211xp5_ASAP7_75t_L g1962 ( 
.A1(n_1871),
.A2(n_1725),
.B(n_1739),
.C(n_1742),
.Y(n_1962)
);

AOI33xp33_ASAP7_75t_L g1963 ( 
.A1(n_1914),
.A2(n_1742),
.A3(n_1739),
.B1(n_1729),
.B2(n_1727),
.B3(n_1726),
.Y(n_1963)
);

OAI33xp33_ASAP7_75t_L g1964 ( 
.A1(n_1891),
.A2(n_1758),
.A3(n_1714),
.B1(n_1785),
.B2(n_1693),
.B3(n_1787),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1878),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1879),
.Y(n_1966)
);

OAI22xp5_ASAP7_75t_L g1967 ( 
.A1(n_1908),
.A2(n_1711),
.B1(n_1745),
.B2(n_1847),
.Y(n_1967)
);

OAI21xp5_ASAP7_75t_L g1968 ( 
.A1(n_1949),
.A2(n_1737),
.B(n_1745),
.Y(n_1968)
);

HB1xp67_ASAP7_75t_L g1969 ( 
.A(n_1873),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1879),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1949),
.A2(n_1847),
.B1(n_1852),
.B2(n_1948),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1948),
.B(n_1847),
.Y(n_1972)
);

AOI22xp5_ASAP7_75t_L g1973 ( 
.A1(n_1948),
.A2(n_1852),
.B1(n_1870),
.B2(n_1889),
.Y(n_1973)
);

AOI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1870),
.A2(n_1916),
.B1(n_1938),
.B2(n_1900),
.C(n_1889),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1938),
.B(n_1852),
.Y(n_1975)
);

BUFx2_ASAP7_75t_L g1976 ( 
.A(n_1864),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1881),
.Y(n_1977)
);

OR2x2_ASAP7_75t_L g1978 ( 
.A(n_1862),
.B(n_1852),
.Y(n_1978)
);

OAI22xp5_ASAP7_75t_L g1979 ( 
.A1(n_1933),
.A2(n_1920),
.B1(n_1875),
.B2(n_1909),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1863),
.Y(n_1980)
);

OR2x6_ASAP7_75t_SL g1981 ( 
.A(n_1891),
.B(n_1920),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1933),
.A2(n_1875),
.B1(n_1909),
.B2(n_1918),
.Y(n_1982)
);

BUFx3_ASAP7_75t_L g1983 ( 
.A(n_1945),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1900),
.A2(n_1896),
.B1(n_1934),
.B2(n_1897),
.C(n_1936),
.Y(n_1984)
);

AND4x1_ASAP7_75t_L g1985 ( 
.A(n_1896),
.B(n_1897),
.C(n_1944),
.D(n_1907),
.Y(n_1985)
);

NAND3xp33_ASAP7_75t_SL g1986 ( 
.A(n_1936),
.B(n_1918),
.C(n_1934),
.Y(n_1986)
);

OAI33xp33_ASAP7_75t_L g1987 ( 
.A1(n_1910),
.A2(n_1890),
.A3(n_1944),
.B1(n_1919),
.B2(n_1886),
.B3(n_1880),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1862),
.B(n_1865),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1863),
.Y(n_1989)
);

AOI222xp33_ASAP7_75t_L g1990 ( 
.A1(n_1916),
.A2(n_1907),
.B1(n_1910),
.B2(n_1893),
.C1(n_1919),
.C2(n_1902),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1883),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1893),
.A2(n_1898),
.B1(n_1939),
.B2(n_1912),
.Y(n_1992)
);

AO21x2_ASAP7_75t_L g1993 ( 
.A1(n_1921),
.A2(n_1905),
.B(n_1895),
.Y(n_1993)
);

NAND2x1_ASAP7_75t_L g1994 ( 
.A(n_1922),
.B(n_1894),
.Y(n_1994)
);

AOI22xp33_ASAP7_75t_L g1995 ( 
.A1(n_1902),
.A2(n_1942),
.B1(n_1890),
.B2(n_1901),
.Y(n_1995)
);

INVxp67_ASAP7_75t_L g1996 ( 
.A(n_1855),
.Y(n_1996)
);

OAI211xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1926),
.A2(n_1937),
.B(n_1940),
.C(n_1942),
.Y(n_1997)
);

OAI33xp33_ASAP7_75t_L g1998 ( 
.A1(n_1880),
.A2(n_1861),
.A3(n_1883),
.B1(n_1888),
.B2(n_1937),
.B3(n_1906),
.Y(n_1998)
);

INVx2_ASAP7_75t_SL g1999 ( 
.A(n_1864),
.Y(n_1999)
);

INVx3_ASAP7_75t_L g2000 ( 
.A(n_1894),
.Y(n_2000)
);

AOI322xp5_ASAP7_75t_L g2001 ( 
.A1(n_1901),
.A2(n_1882),
.A3(n_1926),
.B1(n_1912),
.B2(n_1924),
.C1(n_1940),
.C2(n_1925),
.Y(n_2001)
);

OAI22xp33_ASAP7_75t_L g2002 ( 
.A1(n_1926),
.A2(n_1939),
.B1(n_1858),
.B2(n_1947),
.Y(n_2002)
);

AO21x2_ASAP7_75t_L g2003 ( 
.A1(n_1895),
.A2(n_1905),
.B(n_1885),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1857),
.B(n_1860),
.Y(n_2004)
);

OAI21xp5_ASAP7_75t_L g2005 ( 
.A1(n_1935),
.A2(n_1939),
.B(n_1858),
.Y(n_2005)
);

AOI211xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1931),
.A2(n_1924),
.B(n_1913),
.C(n_1927),
.Y(n_2006)
);

AOI221xp5_ASAP7_75t_L g2007 ( 
.A1(n_1935),
.A2(n_1882),
.B1(n_1946),
.B2(n_1917),
.C(n_1930),
.Y(n_2007)
);

OAI21xp33_ASAP7_75t_L g2008 ( 
.A1(n_1858),
.A2(n_1917),
.B(n_1925),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1868),
.Y(n_2009)
);

AOI221xp5_ASAP7_75t_L g2010 ( 
.A1(n_1882),
.A2(n_1946),
.B1(n_1917),
.B2(n_1930),
.C(n_1906),
.Y(n_2010)
);

AOI22xp33_ASAP7_75t_L g2011 ( 
.A1(n_1930),
.A2(n_1858),
.B1(n_1927),
.B2(n_1903),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_1858),
.A2(n_1927),
.B1(n_1903),
.B2(n_1932),
.Y(n_2012)
);

INVx4_ASAP7_75t_L g2013 ( 
.A(n_1929),
.Y(n_2013)
);

AO21x2_ASAP7_75t_L g2014 ( 
.A1(n_1895),
.A2(n_1905),
.B(n_1885),
.Y(n_2014)
);

OAI222xp33_ASAP7_75t_L g2015 ( 
.A1(n_1939),
.A2(n_1932),
.B1(n_1858),
.B2(n_1911),
.C1(n_1892),
.C2(n_1899),
.Y(n_2015)
);

OR2x2_ASAP7_75t_L g2016 ( 
.A(n_1988),
.B(n_1904),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_2010),
.B(n_2007),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_2004),
.B(n_1884),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1980),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1957),
.B(n_1884),
.Y(n_2020)
);

AOI222xp33_ASAP7_75t_L g2021 ( 
.A1(n_1974),
.A2(n_1931),
.B1(n_1874),
.B2(n_1876),
.C1(n_1869),
.C2(n_1945),
.Y(n_2021)
);

INVx3_ASAP7_75t_L g2022 ( 
.A(n_1993),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_1957),
.B(n_1928),
.Y(n_2023)
);

INVx1_ASAP7_75t_L g2024 ( 
.A(n_1980),
.Y(n_2024)
);

INVx2_ASAP7_75t_L g2025 ( 
.A(n_1993),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2003),
.B(n_1928),
.Y(n_2026)
);

AND2x2_ASAP7_75t_L g2027 ( 
.A(n_2014),
.B(n_1885),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1989),
.Y(n_2028)
);

OR2x2_ASAP7_75t_L g2029 ( 
.A(n_2014),
.B(n_1856),
.Y(n_2029)
);

AND2x2_ASAP7_75t_L g2030 ( 
.A(n_2008),
.B(n_1860),
.Y(n_2030)
);

AND2x4_ASAP7_75t_L g2031 ( 
.A(n_2000),
.B(n_1994),
.Y(n_2031)
);

INVx2_ASAP7_75t_L g2032 ( 
.A(n_1993),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2000),
.B(n_1856),
.Y(n_2033)
);

AND2x2_ASAP7_75t_L g2034 ( 
.A(n_2000),
.B(n_1856),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_2012),
.B(n_1856),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_2009),
.B(n_1956),
.Y(n_2036)
);

OR2x2_ASAP7_75t_L g2037 ( 
.A(n_1950),
.B(n_1856),
.Y(n_2037)
);

INVx3_ASAP7_75t_SL g2038 ( 
.A(n_2013),
.Y(n_2038)
);

AND2x2_ASAP7_75t_SL g2039 ( 
.A(n_1963),
.B(n_1931),
.Y(n_2039)
);

INVxp67_ASAP7_75t_L g2040 ( 
.A(n_1981),
.Y(n_2040)
);

NOR2xp67_ASAP7_75t_L g2041 ( 
.A(n_1984),
.B(n_1877),
.Y(n_2041)
);

INVx2_ASAP7_75t_L g2042 ( 
.A(n_1965),
.Y(n_2042)
);

AND2x2_ASAP7_75t_L g2043 ( 
.A(n_2012),
.B(n_1856),
.Y(n_2043)
);

BUFx2_ASAP7_75t_L g2044 ( 
.A(n_1960),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1966),
.B(n_1923),
.Y(n_2045)
);

AND2x2_ASAP7_75t_L g2046 ( 
.A(n_2005),
.B(n_1856),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1970),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_L g2048 ( 
.A(n_1990),
.B(n_1915),
.C(n_1947),
.Y(n_2048)
);

AND2x2_ASAP7_75t_L g2049 ( 
.A(n_2011),
.B(n_1867),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1977),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1991),
.B(n_1923),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_2011),
.B(n_1867),
.Y(n_2052)
);

HB1xp67_ASAP7_75t_L g2053 ( 
.A(n_1969),
.Y(n_2053)
);

BUFx3_ASAP7_75t_L g2054 ( 
.A(n_1983),
.Y(n_2054)
);

NOR2xp67_ASAP7_75t_L g2055 ( 
.A(n_1986),
.B(n_1877),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1983),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1955),
.B(n_1899),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1995),
.B(n_1953),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_2025),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_2036),
.B(n_2001),
.Y(n_2060)
);

AND2x2_ASAP7_75t_L g2061 ( 
.A(n_2033),
.B(n_2006),
.Y(n_2061)
);

AND2x2_ASAP7_75t_L g2062 ( 
.A(n_2033),
.B(n_1976),
.Y(n_2062)
);

NAND2x1p5_ASAP7_75t_L g2063 ( 
.A(n_2044),
.B(n_1931),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2033),
.B(n_1999),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2042),
.Y(n_2065)
);

INVxp33_ASAP7_75t_L g2066 ( 
.A(n_2041),
.Y(n_2066)
);

AOI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_2039),
.A2(n_1971),
.B1(n_1951),
.B2(n_1979),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_2034),
.B(n_1999),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2036),
.B(n_1995),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2042),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_2023),
.B(n_1981),
.Y(n_2071)
);

BUFx2_ASAP7_75t_L g2072 ( 
.A(n_2044),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2042),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_2019),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2023),
.B(n_1992),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2025),
.Y(n_2076)
);

INVxp67_ASAP7_75t_L g2077 ( 
.A(n_2040),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_2034),
.B(n_1877),
.Y(n_2078)
);

OAI21xp33_ASAP7_75t_L g2079 ( 
.A1(n_2017),
.A2(n_1985),
.B(n_1982),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_2025),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_2037),
.B(n_1978),
.Y(n_2081)
);

INVxp67_ASAP7_75t_SL g2082 ( 
.A(n_2029),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2034),
.B(n_1877),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_L g2084 ( 
.A(n_2023),
.B(n_1963),
.Y(n_2084)
);

INVx2_ASAP7_75t_L g2085 ( 
.A(n_2032),
.Y(n_2085)
);

INVxp67_ASAP7_75t_SL g2086 ( 
.A(n_2029),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_2019),
.Y(n_2087)
);

AND2x2_ASAP7_75t_L g2088 ( 
.A(n_2026),
.B(n_1859),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2032),
.Y(n_2089)
);

BUFx2_ASAP7_75t_L g2090 ( 
.A(n_2038),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2026),
.B(n_1859),
.Y(n_2091)
);

AND2x2_ASAP7_75t_L g2092 ( 
.A(n_2026),
.B(n_1941),
.Y(n_2092)
);

AND2x4_ASAP7_75t_L g2093 ( 
.A(n_2031),
.B(n_2013),
.Y(n_2093)
);

OR3x2_ASAP7_75t_L g2094 ( 
.A(n_2040),
.B(n_1964),
.C(n_1987),
.Y(n_2094)
);

NOR2xp33_ASAP7_75t_L g2095 ( 
.A(n_2017),
.B(n_1952),
.Y(n_2095)
);

AOI33xp33_ASAP7_75t_L g2096 ( 
.A1(n_2035),
.A2(n_1973),
.A3(n_2002),
.B1(n_1959),
.B2(n_1954),
.B3(n_1997),
.Y(n_2096)
);

INVx3_ASAP7_75t_SL g2097 ( 
.A(n_2038),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2041),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2047),
.B(n_1952),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2024),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2047),
.B(n_2050),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2027),
.B(n_1941),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2024),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2031),
.B(n_2013),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2050),
.B(n_1962),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2037),
.B(n_1941),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2028),
.Y(n_2107)
);

OR2x2_ASAP7_75t_L g2108 ( 
.A(n_2037),
.B(n_1941),
.Y(n_2108)
);

INVx2_ASAP7_75t_L g2109 ( 
.A(n_2032),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_2038),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2028),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2095),
.B(n_2039),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2101),
.Y(n_2113)
);

AOI22xp5_ASAP7_75t_L g2114 ( 
.A1(n_2079),
.A2(n_2039),
.B1(n_2035),
.B2(n_2043),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2077),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2077),
.B(n_2016),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_L g2117 ( 
.A(n_2095),
.B(n_2039),
.Y(n_2117)
);

NAND4xp25_ASAP7_75t_L g2118 ( 
.A(n_2079),
.B(n_2048),
.C(n_2021),
.D(n_1968),
.Y(n_2118)
);

AND3x1_ASAP7_75t_L g2119 ( 
.A(n_2096),
.B(n_2084),
.C(n_2071),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2061),
.B(n_2020),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2061),
.B(n_2020),
.Y(n_2121)
);

INVx1_ASAP7_75t_SL g2122 ( 
.A(n_2071),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_L g2123 ( 
.A(n_2084),
.B(n_2058),
.Y(n_2123)
);

HB1xp67_ASAP7_75t_L g2124 ( 
.A(n_2072),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2061),
.B(n_2020),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_2105),
.B(n_2058),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_R g2127 ( 
.A(n_2067),
.B(n_1929),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2101),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2074),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_2074),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2088),
.B(n_2018),
.Y(n_2131)
);

INVx5_ASAP7_75t_L g2132 ( 
.A(n_2090),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2105),
.B(n_2055),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2087),
.Y(n_2134)
);

AND2x2_ASAP7_75t_L g2135 ( 
.A(n_2088),
.B(n_2091),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2088),
.B(n_2018),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_2081),
.B(n_2016),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2081),
.B(n_2106),
.Y(n_2138)
);

OR2x2_ASAP7_75t_L g2139 ( 
.A(n_2081),
.B(n_2016),
.Y(n_2139)
);

OR2x6_ASAP7_75t_L g2140 ( 
.A(n_2090),
.B(n_2055),
.Y(n_2140)
);

INVx2_ASAP7_75t_L g2141 ( 
.A(n_2059),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2069),
.B(n_2030),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2111),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_SL g2144 ( 
.A(n_2096),
.B(n_2021),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2069),
.B(n_2030),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2111),
.Y(n_2146)
);

AND2x4_ASAP7_75t_L g2147 ( 
.A(n_2093),
.B(n_2031),
.Y(n_2147)
);

OAI211xp5_ASAP7_75t_SL g2148 ( 
.A1(n_2067),
.A2(n_2098),
.B(n_2060),
.C(n_2099),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2099),
.B(n_2030),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2060),
.B(n_2075),
.Y(n_2150)
);

INVx1_ASAP7_75t_L g2151 ( 
.A(n_2087),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2075),
.B(n_2057),
.Y(n_2152)
);

BUFx2_ASAP7_75t_L g2153 ( 
.A(n_2097),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2100),
.Y(n_2154)
);

OR2x2_ASAP7_75t_L g2155 ( 
.A(n_2106),
.B(n_2048),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2100),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2103),
.Y(n_2157)
);

INVx3_ASAP7_75t_L g2158 ( 
.A(n_2093),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_2103),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_2092),
.B(n_2057),
.Y(n_2160)
);

INVx3_ASAP7_75t_L g2161 ( 
.A(n_2132),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2115),
.Y(n_2162)
);

AOI221xp5_ASAP7_75t_L g2163 ( 
.A1(n_2119),
.A2(n_2094),
.B1(n_2046),
.B2(n_2066),
.C(n_2092),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2120),
.B(n_2121),
.Y(n_2164)
);

OAI21xp33_ASAP7_75t_L g2165 ( 
.A1(n_2144),
.A2(n_2046),
.B(n_2066),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_2123),
.B(n_2098),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2129),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2129),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_L g2169 ( 
.A(n_2112),
.B(n_2091),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2130),
.Y(n_2170)
);

OAI221xp5_ASAP7_75t_L g2171 ( 
.A1(n_2144),
.A2(n_2097),
.B1(n_2063),
.B2(n_2106),
.C(n_2108),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_L g2172 ( 
.A(n_2117),
.B(n_2126),
.Y(n_2172)
);

AOI222xp33_ASAP7_75t_L g2173 ( 
.A1(n_2148),
.A2(n_2035),
.B1(n_2043),
.B2(n_2046),
.C1(n_2092),
.C2(n_2102),
.Y(n_2173)
);

OAI22xp33_ASAP7_75t_SL g2174 ( 
.A1(n_2114),
.A2(n_2097),
.B1(n_2110),
.B2(n_2072),
.Y(n_2174)
);

NAND3xp33_ASAP7_75t_L g2175 ( 
.A(n_2118),
.B(n_2043),
.C(n_2110),
.Y(n_2175)
);

AND2x2_ASAP7_75t_L g2176 ( 
.A(n_2120),
.B(n_2093),
.Y(n_2176)
);

OAI22xp33_ASAP7_75t_SL g2177 ( 
.A1(n_2153),
.A2(n_2155),
.B1(n_2140),
.B2(n_2150),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_2130),
.Y(n_2178)
);

BUFx3_ASAP7_75t_L g2179 ( 
.A(n_2153),
.Y(n_2179)
);

NOR2xp67_ASAP7_75t_L g2180 ( 
.A(n_2132),
.B(n_2093),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_2134),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2143),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2122),
.B(n_2091),
.Y(n_2183)
);

NAND2xp5_ASAP7_75t_L g2184 ( 
.A(n_2133),
.B(n_2102),
.Y(n_2184)
);

AOI21xp5_ASAP7_75t_L g2185 ( 
.A1(n_2142),
.A2(n_1958),
.B(n_2102),
.Y(n_2185)
);

OAI22xp5_ASAP7_75t_L g2186 ( 
.A1(n_2152),
.A2(n_2094),
.B1(n_2063),
.B2(n_1959),
.Y(n_2186)
);

INVx1_ASAP7_75t_SL g2187 ( 
.A(n_2127),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2145),
.B(n_2149),
.Y(n_2188)
);

OR2x2_ASAP7_75t_L g2189 ( 
.A(n_2116),
.B(n_2108),
.Y(n_2189)
);

INVxp67_ASAP7_75t_L g2190 ( 
.A(n_2124),
.Y(n_2190)
);

NOR2xp33_ASAP7_75t_L g2191 ( 
.A(n_2132),
.B(n_1996),
.Y(n_2191)
);

AOI222xp33_ASAP7_75t_L g2192 ( 
.A1(n_2121),
.A2(n_2052),
.B1(n_2049),
.B2(n_2094),
.C1(n_2015),
.C2(n_2082),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2146),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_2132),
.B(n_2097),
.Y(n_2194)
);

OA21x2_ASAP7_75t_L g2195 ( 
.A1(n_2141),
.A2(n_2109),
.B(n_2059),
.Y(n_2195)
);

OAI221xp5_ASAP7_75t_L g2196 ( 
.A1(n_2155),
.A2(n_2063),
.B1(n_2108),
.B2(n_2029),
.C(n_2086),
.Y(n_2196)
);

INVx2_ASAP7_75t_SL g2197 ( 
.A(n_2132),
.Y(n_2197)
);

INVxp67_ASAP7_75t_L g2198 ( 
.A(n_2116),
.Y(n_2198)
);

AOI22xp33_ASAP7_75t_L g2199 ( 
.A1(n_2125),
.A2(n_2049),
.B1(n_2052),
.B2(n_1998),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2167),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2168),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2170),
.Y(n_2202)
);

OAI21xp5_ASAP7_75t_L g2203 ( 
.A1(n_2175),
.A2(n_2140),
.B(n_2113),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2178),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2181),
.Y(n_2205)
);

AND2x4_ASAP7_75t_L g2206 ( 
.A(n_2180),
.B(n_2125),
.Y(n_2206)
);

AOI221xp5_ASAP7_75t_SL g2207 ( 
.A1(n_2163),
.A2(n_2174),
.B1(n_2165),
.B2(n_2177),
.C(n_2186),
.Y(n_2207)
);

NAND2xp33_ASAP7_75t_SL g2208 ( 
.A(n_2166),
.B(n_2038),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2192),
.A2(n_2140),
.B1(n_2147),
.B2(n_2104),
.Y(n_2209)
);

NOR2xp33_ASAP7_75t_L g2210 ( 
.A(n_2187),
.B(n_2158),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2182),
.Y(n_2211)
);

AND2x2_ASAP7_75t_L g2212 ( 
.A(n_2164),
.B(n_2158),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2161),
.Y(n_2213)
);

INVx2_ASAP7_75t_SL g2214 ( 
.A(n_2161),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2193),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2179),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2162),
.Y(n_2217)
);

O2A1O1Ixp33_ASAP7_75t_SL g2218 ( 
.A1(n_2197),
.A2(n_2082),
.B(n_2086),
.C(n_2056),
.Y(n_2218)
);

AOI21xp33_ASAP7_75t_SL g2219 ( 
.A1(n_2191),
.A2(n_2140),
.B(n_2063),
.Y(n_2219)
);

NAND2xp5_ASAP7_75t_L g2220 ( 
.A(n_2179),
.B(n_2128),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2183),
.B(n_2160),
.Y(n_2221)
);

INVxp67_ASAP7_75t_L g2222 ( 
.A(n_2191),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_2172),
.B(n_2158),
.Y(n_2223)
);

AND2x2_ASAP7_75t_L g2224 ( 
.A(n_2176),
.B(n_2147),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_2190),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2198),
.Y(n_2226)
);

OAI221xp5_ASAP7_75t_L g2227 ( 
.A1(n_2171),
.A2(n_2128),
.B1(n_2138),
.B2(n_2137),
.C(n_2139),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2176),
.B(n_2147),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2200),
.Y(n_2229)
);

OR2x2_ASAP7_75t_L g2230 ( 
.A(n_2225),
.B(n_2169),
.Y(n_2230)
);

OAI221xp5_ASAP7_75t_L g2231 ( 
.A1(n_2207),
.A2(n_2173),
.B1(n_2199),
.B2(n_2196),
.C(n_2185),
.Y(n_2231)
);

AND2x4_ASAP7_75t_SL g2232 ( 
.A(n_2206),
.B(n_2161),
.Y(n_2232)
);

NOR3xp33_ASAP7_75t_SL g2233 ( 
.A(n_2208),
.B(n_2194),
.C(n_2188),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2200),
.Y(n_2234)
);

AND2x2_ASAP7_75t_L g2235 ( 
.A(n_2224),
.B(n_2194),
.Y(n_2235)
);

AND2x2_ASAP7_75t_L g2236 ( 
.A(n_2224),
.B(n_2197),
.Y(n_2236)
);

INVxp67_ASAP7_75t_L g2237 ( 
.A(n_2210),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2202),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2222),
.B(n_2188),
.Y(n_2239)
);

INVx2_ASAP7_75t_SL g2240 ( 
.A(n_2206),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_2219),
.B(n_2206),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2202),
.Y(n_2242)
);

NOR3xp33_ASAP7_75t_SL g2243 ( 
.A(n_2208),
.B(n_2184),
.C(n_1975),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2201),
.Y(n_2244)
);

OAI21xp5_ASAP7_75t_L g2245 ( 
.A1(n_2209),
.A2(n_2199),
.B(n_2189),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2204),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_2213),
.Y(n_2247)
);

INVx2_ASAP7_75t_L g2248 ( 
.A(n_2214),
.Y(n_2248)
);

NAND2x1p5_ASAP7_75t_L g2249 ( 
.A(n_2216),
.B(n_2195),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2228),
.B(n_2135),
.Y(n_2250)
);

NOR3xp33_ASAP7_75t_SL g2251 ( 
.A(n_2203),
.B(n_1975),
.C(n_1967),
.Y(n_2251)
);

NOR3xp33_ASAP7_75t_L g2252 ( 
.A(n_2237),
.B(n_2216),
.C(n_2226),
.Y(n_2252)
);

NAND2x1_ASAP7_75t_L g2253 ( 
.A(n_2240),
.B(n_2214),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_SL g2254 ( 
.A(n_2233),
.B(n_2223),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_2247),
.Y(n_2255)
);

AOI21xp5_ASAP7_75t_L g2256 ( 
.A1(n_2231),
.A2(n_2218),
.B(n_2227),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2248),
.Y(n_2257)
);

OAI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_2243),
.A2(n_2217),
.B1(n_2220),
.B2(n_2211),
.Y(n_2258)
);

NAND3xp33_ASAP7_75t_SL g2259 ( 
.A(n_2245),
.B(n_2239),
.C(n_2241),
.Y(n_2259)
);

NOR2xp67_ASAP7_75t_L g2260 ( 
.A(n_2240),
.B(n_2248),
.Y(n_2260)
);

NOR3xp33_ASAP7_75t_SL g2261 ( 
.A(n_2244),
.B(n_2205),
.C(n_2215),
.Y(n_2261)
);

OAI21xp33_ASAP7_75t_L g2262 ( 
.A1(n_2235),
.A2(n_2236),
.B(n_2251),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2232),
.Y(n_2263)
);

NOR3xp33_ASAP7_75t_L g2264 ( 
.A(n_2235),
.B(n_2213),
.C(n_2218),
.Y(n_2264)
);

AND2x2_ASAP7_75t_L g2265 ( 
.A(n_2236),
.B(n_2228),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2250),
.B(n_2212),
.Y(n_2266)
);

AOI211xp5_ASAP7_75t_L g2267 ( 
.A1(n_2256),
.A2(n_2259),
.B(n_2264),
.C(n_2258),
.Y(n_2267)
);

NOR2x1p5_ASAP7_75t_L g2268 ( 
.A(n_2253),
.B(n_2230),
.Y(n_2268)
);

AOI211xp5_ASAP7_75t_L g2269 ( 
.A1(n_2258),
.A2(n_2230),
.B(n_2246),
.C(n_2244),
.Y(n_2269)
);

NAND5xp2_ASAP7_75t_L g2270 ( 
.A(n_2262),
.B(n_2246),
.C(n_2229),
.D(n_2249),
.E(n_2242),
.Y(n_2270)
);

NAND4xp25_ASAP7_75t_SL g2271 ( 
.A(n_2266),
.B(n_2250),
.C(n_2212),
.D(n_2221),
.Y(n_2271)
);

AND2x2_ASAP7_75t_L g2272 ( 
.A(n_2265),
.B(n_2232),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_SL g2273 ( 
.A(n_2263),
.B(n_2249),
.Y(n_2273)
);

OAI211xp5_ASAP7_75t_L g2274 ( 
.A1(n_2254),
.A2(n_2242),
.B(n_2238),
.C(n_2234),
.Y(n_2274)
);

AOI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2252),
.A2(n_2238),
.B1(n_2234),
.B2(n_2221),
.Y(n_2275)
);

AOI331xp33_ASAP7_75t_L g2276 ( 
.A1(n_2257),
.A2(n_2249),
.A3(n_2159),
.B1(n_2151),
.B2(n_2157),
.B3(n_2154),
.C1(n_2156),
.Y(n_2276)
);

OAI22xp5_ASAP7_75t_L g2277 ( 
.A1(n_2261),
.A2(n_2260),
.B1(n_2255),
.B2(n_2104),
.Y(n_2277)
);

OAI21xp33_ASAP7_75t_SL g2278 ( 
.A1(n_2256),
.A2(n_2135),
.B(n_2138),
.Y(n_2278)
);

OAI21xp33_ASAP7_75t_L g2279 ( 
.A1(n_2262),
.A2(n_2139),
.B(n_2137),
.Y(n_2279)
);

NAND4xp25_ASAP7_75t_L g2280 ( 
.A(n_2256),
.B(n_1961),
.C(n_2052),
.D(n_2049),
.Y(n_2280)
);

OAI21xp5_ASAP7_75t_L g2281 ( 
.A1(n_2256),
.A2(n_2093),
.B(n_2104),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_R g2282 ( 
.A(n_2272),
.B(n_2054),
.Y(n_2282)
);

AOI211xp5_ASAP7_75t_L g2283 ( 
.A1(n_2267),
.A2(n_2104),
.B(n_2141),
.C(n_2056),
.Y(n_2283)
);

OR2x2_ASAP7_75t_L g2284 ( 
.A(n_2271),
.B(n_2131),
.Y(n_2284)
);

AOI21xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2268),
.A2(n_2273),
.B(n_2277),
.Y(n_2285)
);

NAND4xp75_ASAP7_75t_L g2286 ( 
.A(n_2278),
.B(n_2195),
.C(n_1972),
.D(n_2131),
.Y(n_2286)
);

NOR3x1_ASAP7_75t_L g2287 ( 
.A(n_2281),
.B(n_1972),
.C(n_2045),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2275),
.Y(n_2288)
);

AOI22xp5_ASAP7_75t_L g2289 ( 
.A1(n_2279),
.A2(n_2104),
.B1(n_2136),
.B2(n_2054),
.Y(n_2289)
);

AO22x2_ASAP7_75t_L g2290 ( 
.A1(n_2274),
.A2(n_2270),
.B1(n_2269),
.B2(n_2276),
.Y(n_2290)
);

INVx2_ASAP7_75t_L g2291 ( 
.A(n_2274),
.Y(n_2291)
);

NOR2xp33_ASAP7_75t_R g2292 ( 
.A(n_2280),
.B(n_2054),
.Y(n_2292)
);

AND2x4_ASAP7_75t_L g2293 ( 
.A(n_2288),
.B(n_2136),
.Y(n_2293)
);

OAI22xp5_ASAP7_75t_L g2294 ( 
.A1(n_2290),
.A2(n_2053),
.B1(n_2068),
.B2(n_2064),
.Y(n_2294)
);

OR2x2_ASAP7_75t_L g2295 ( 
.A(n_2284),
.B(n_2053),
.Y(n_2295)
);

OR2x2_ASAP7_75t_L g2296 ( 
.A(n_2291),
.B(n_2195),
.Y(n_2296)
);

NOR2xp33_ASAP7_75t_L g2297 ( 
.A(n_2285),
.B(n_2107),
.Y(n_2297)
);

CKINVDCx16_ASAP7_75t_R g2298 ( 
.A(n_2282),
.Y(n_2298)
);

NOR3xp33_ASAP7_75t_SL g2299 ( 
.A(n_2286),
.B(n_2045),
.C(n_2051),
.Y(n_2299)
);

INVxp67_ASAP7_75t_L g2300 ( 
.A(n_2290),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2292),
.Y(n_2301)
);

AOI21xp5_ASAP7_75t_L g2302 ( 
.A1(n_2283),
.A2(n_2109),
.B(n_2059),
.Y(n_2302)
);

NAND2xp5_ASAP7_75t_L g2303 ( 
.A(n_2298),
.B(n_2287),
.Y(n_2303)
);

NAND5xp2_ASAP7_75t_L g2304 ( 
.A(n_2301),
.B(n_2289),
.C(n_2062),
.D(n_2064),
.E(n_2068),
.Y(n_2304)
);

HB1xp67_ASAP7_75t_L g2305 ( 
.A(n_2296),
.Y(n_2305)
);

INVx4_ASAP7_75t_L g2306 ( 
.A(n_2293),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_2295),
.Y(n_2307)
);

AOI22xp5_ASAP7_75t_SL g2308 ( 
.A1(n_2300),
.A2(n_2031),
.B1(n_2062),
.B2(n_2068),
.Y(n_2308)
);

NAND3xp33_ASAP7_75t_SL g2309 ( 
.A(n_2297),
.B(n_2062),
.C(n_2109),
.Y(n_2309)
);

AND2x4_ASAP7_75t_L g2310 ( 
.A(n_2299),
.B(n_2064),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2306),
.Y(n_2311)
);

AOI311xp33_ASAP7_75t_L g2312 ( 
.A1(n_2307),
.A2(n_2294),
.A3(n_2302),
.B(n_2065),
.C(n_2070),
.Y(n_2312)
);

CKINVDCx5p33_ASAP7_75t_R g2313 ( 
.A(n_2305),
.Y(n_2313)
);

CKINVDCx5p33_ASAP7_75t_R g2314 ( 
.A(n_2303),
.Y(n_2314)
);

AOI22x1_ASAP7_75t_L g2315 ( 
.A1(n_2313),
.A2(n_2308),
.B1(n_2310),
.B2(n_2309),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2311),
.Y(n_2316)
);

INVx4_ASAP7_75t_L g2317 ( 
.A(n_2316),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2315),
.A2(n_2311),
.B(n_2314),
.Y(n_2318)
);

HB1xp67_ASAP7_75t_L g2319 ( 
.A(n_2317),
.Y(n_2319)
);

AND3x1_ASAP7_75t_L g2320 ( 
.A(n_2318),
.B(n_2304),
.C(n_2312),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2317),
.Y(n_2321)
);

AOI222xp33_ASAP7_75t_L g2322 ( 
.A1(n_2321),
.A2(n_2310),
.B1(n_2076),
.B2(n_2089),
.C1(n_2085),
.C2(n_2080),
.Y(n_2322)
);

AOI222xp33_ASAP7_75t_L g2323 ( 
.A1(n_2319),
.A2(n_2080),
.B1(n_2089),
.B2(n_2085),
.C1(n_2076),
.C2(n_2073),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2322),
.A2(n_2320),
.B1(n_2089),
.B2(n_2085),
.Y(n_2324)
);

AOI22xp33_ASAP7_75t_L g2325 ( 
.A1(n_2323),
.A2(n_2080),
.B1(n_2076),
.B2(n_2031),
.Y(n_2325)
);

AOI22xp33_ASAP7_75t_SL g2326 ( 
.A1(n_2324),
.A2(n_2083),
.B1(n_2078),
.B2(n_2022),
.Y(n_2326)
);

AOI221xp5_ASAP7_75t_L g2327 ( 
.A1(n_2326),
.A2(n_2325),
.B1(n_2065),
.B2(n_2073),
.C(n_2070),
.Y(n_2327)
);

AOI211xp5_ASAP7_75t_L g2328 ( 
.A1(n_2327),
.A2(n_2107),
.B(n_2051),
.C(n_1929),
.Y(n_2328)
);


endmodule