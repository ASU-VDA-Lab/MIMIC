module fake_jpeg_7315_n_138 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_138);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_138;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx3_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_28),
.Y(n_37)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_30),
.Y(n_47)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_34),
.C(n_25),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_13),
.B(n_0),
.C(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_18),
.B1(n_22),
.B2(n_13),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_35),
.A2(n_38),
.B1(n_39),
.B2(n_43),
.Y(n_54)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_31),
.A2(n_22),
.B1(n_18),
.B2(n_25),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_22),
.B1(n_18),
.B2(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_34),
.Y(n_55)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_27),
.A2(n_24),
.B1(n_30),
.B2(n_28),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_24),
.B1(n_21),
.B2(n_14),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_46),
.A2(n_34),
.B1(n_15),
.B2(n_21),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_57),
.B1(n_35),
.B2(n_38),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_46),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_59),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_55),
.B(n_41),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_60),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_33),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_47),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_62),
.B(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_73),
.Y(n_78)
);

OR2x2_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_37),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_72),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_68),
.A2(n_70),
.B1(n_77),
.B2(n_67),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_77),
.C(n_29),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_54),
.A2(n_40),
.B1(n_42),
.B2(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_62),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_12),
.Y(n_75)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_52),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_83),
.B(n_85),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_73),
.A2(n_12),
.B1(n_43),
.B2(n_15),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_71),
.A2(n_29),
.B(n_61),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_90),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_88),
.C(n_68),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_52),
.C(n_30),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_89),
.A2(n_45),
.B1(n_36),
.B2(n_32),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_71),
.A2(n_17),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_81),
.B(n_65),
.Y(n_91)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_87),
.C(n_85),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_SL g93 ( 
.A1(n_83),
.A2(n_65),
.A3(n_11),
.B1(n_10),
.B2(n_70),
.C1(n_7),
.C2(n_8),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_93),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_78),
.Y(n_95)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_80),
.B(n_17),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_79),
.B(n_76),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_98),
.A2(n_20),
.B(n_16),
.Y(n_111)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_100),
.B1(n_45),
.B2(n_63),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_106),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_92),
.C(n_97),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_82),
.C(n_26),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_109),
.Y(n_119)
);

HB1xp67_ASAP7_75t_L g110 ( 
.A(n_100),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_110),
.A2(n_101),
.B1(n_94),
.B2(n_63),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_3),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_113),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_101),
.B1(n_82),
.B2(n_64),
.Y(n_114)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g115 ( 
.A1(n_106),
.A2(n_36),
.A3(n_16),
.B1(n_20),
.B2(n_32),
.C1(n_45),
.C2(n_44),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_116),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_102),
.A2(n_44),
.B1(n_58),
.B2(n_48),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_44),
.B1(n_20),
.B2(n_48),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_117),
.A2(n_118),
.B(n_111),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_121),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_112),
.B(n_119),
.C(n_116),
.Y(n_124)
);

NOR2xp67_ASAP7_75t_L g125 ( 
.A(n_114),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_125),
.B(n_105),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_123),
.A2(n_107),
.B1(n_119),
.B2(n_118),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_128),
.B1(n_130),
.B2(n_122),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_120),
.B(n_112),
.Y(n_129)
);

OAI221xp5_ASAP7_75t_L g133 ( 
.A1(n_129),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.C(n_8),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_122),
.A2(n_48),
.B1(n_11),
.B2(n_5),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_8),
.C(n_9),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_L g132 ( 
.A1(n_127),
.A2(n_124),
.B1(n_126),
.B2(n_5),
.C(n_6),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g135 ( 
.A1(n_132),
.A2(n_133),
.B(n_9),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g136 ( 
.A(n_134),
.B(n_135),
.CI(n_9),
.CON(n_136),
.SN(n_136)
);

NAND2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_135),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_136),
.Y(n_138)
);


endmodule