module fake_jpeg_12984_n_242 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_16),
.B(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_14),
.B(n_10),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx11_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_40),
.B(n_56),
.Y(n_95)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_46),
.B(n_61),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_52),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_28),
.Y(n_57)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

AOI21xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_1),
.B(n_2),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_58),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_18),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

BUFx24_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_35),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_63),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_61),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_65),
.B(n_71),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_45),
.A2(n_17),
.B1(n_33),
.B2(n_18),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_73),
.B1(n_76),
.B2(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_29),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_L g125 ( 
.A1(n_72),
.A2(n_85),
.B(n_86),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_42),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_53),
.A2(n_20),
.B1(n_31),
.B2(n_30),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_75),
.A2(n_87),
.B1(n_88),
.B2(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_52),
.A2(n_34),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_55),
.A2(n_25),
.B1(n_22),
.B2(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_22),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_15),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_14),
.Y(n_89)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_11),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_93),
.B(n_6),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_98),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_51),
.B1(n_47),
.B2(n_39),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_99),
.A2(n_111),
.B1(n_116),
.B2(n_118),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_100),
.B(n_95),
.Y(n_127)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_67),
.Y(n_101)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_101),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_108),
.Y(n_128)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_103),
.Y(n_149)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g129 ( 
.A(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_97),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_109),
.Y(n_147)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_47),
.B(n_49),
.C(n_48),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_112),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_60),
.B1(n_57),
.B2(n_8),
.Y(n_111)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_113),
.B(n_114),
.Y(n_140)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_117),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_81),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_74),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_10),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_124),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_91),
.A2(n_75),
.B1(n_64),
.B2(n_90),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_121),
.A2(n_103),
.B1(n_108),
.B2(n_115),
.Y(n_146)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_122),
.B(n_126),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_13),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_127),
.B(n_148),
.Y(n_160)
);

NAND2x1_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_90),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_130),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_88),
.B1(n_66),
.B2(n_84),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_131),
.B(n_138),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_134),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_125),
.A2(n_91),
.B(n_69),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_137),
.A2(n_143),
.B(n_139),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_104),
.A2(n_66),
.B1(n_84),
.B2(n_94),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_123),
.B(n_64),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_141),
.B(n_150),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_120),
.A2(n_69),
.B(n_83),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_110),
.B1(n_101),
.B2(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_144),
.A2(n_146),
.B1(n_105),
.B2(n_139),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_119),
.B(n_124),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_112),
.A2(n_114),
.B1(n_122),
.B2(n_117),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_130),
.Y(n_161)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_147),
.Y(n_153)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_141),
.B(n_107),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_154),
.A2(n_169),
.B(n_170),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_156),
.A2(n_173),
.B1(n_133),
.B2(n_142),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_132),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_147),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_158),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx13_ASAP7_75t_L g162 ( 
.A(n_149),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_162),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_145),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_132),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_164),
.B(n_165),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_150),
.B(n_128),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_168),
.Y(n_179)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_128),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_140),
.B(n_138),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_172),
.A2(n_161),
.B(n_169),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_131),
.B1(n_130),
.B2(n_146),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_182),
.B1(n_167),
.B2(n_155),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_140),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_183),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_153),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_171),
.A2(n_151),
.B1(n_135),
.B2(n_149),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_165),
.B(n_148),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_164),
.A2(n_127),
.B1(n_129),
.B2(n_134),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_185),
.B(n_190),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_129),
.B1(n_134),
.B2(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_199),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_157),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_192),
.B(n_175),
.C(n_186),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_189),
.A2(n_167),
.B(n_154),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_193),
.B(n_175),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_194),
.A2(n_198),
.B1(n_185),
.B2(n_187),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_181),
.A2(n_173),
.B(n_166),
.Y(n_196)
);

O2A1O1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_197),
.B(n_187),
.C(n_184),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_189),
.A2(n_159),
.B1(n_158),
.B2(n_172),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_179),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_174),
.Y(n_203)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_204),
.C(n_160),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_205),
.B(n_196),
.C(n_193),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_206),
.A2(n_213),
.B(n_203),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_210),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_209),
.B(n_211),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_192),
.B(n_176),
.Y(n_210)
);

XOR2x2_ASAP7_75t_L g211 ( 
.A(n_197),
.B(n_176),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_212),
.A2(n_177),
.B1(n_201),
.B2(n_214),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_172),
.B(n_178),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_221),
.C(n_188),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_208),
.B(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_219),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_206),
.B(n_195),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_198),
.C(n_201),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_222),
.A2(n_211),
.B1(n_190),
.B2(n_213),
.Y(n_223)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_217),
.A2(n_182),
.B1(n_210),
.B2(n_191),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_225),
.Y(n_229)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_226),
.B(n_218),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_228),
.B(n_216),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NOR2xp67_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_218),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_232),
.A2(n_224),
.B1(n_225),
.B2(n_231),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_229),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_237),
.B(n_238),
.C(n_234),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_235),
.B(n_229),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_239),
.A2(n_228),
.B(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_240),
.B(n_152),
.C(n_129),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_162),
.Y(n_242)
);


endmodule