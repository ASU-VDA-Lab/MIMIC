module fake_aes_11788_n_663 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_663);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_663;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_581;
wire n_458;
wire n_504;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_13), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_68), .Y(n_81) );
BUFx5_ASAP7_75t_L g82 ( .A(n_38), .Y(n_82) );
INVxp67_ASAP7_75t_L g83 ( .A(n_35), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_65), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_75), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_17), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_8), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_25), .Y(n_88) );
INVx1_ASAP7_75t_SL g89 ( .A(n_30), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_28), .Y(n_90) );
BUFx6f_ASAP7_75t_L g91 ( .A(n_42), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_18), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
BUFx3_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_77), .Y(n_95) );
INVx3_ASAP7_75t_L g96 ( .A(n_44), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_29), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_48), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_62), .Y(n_99) );
INVxp33_ASAP7_75t_SL g100 ( .A(n_55), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_8), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_2), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_57), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_0), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_72), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_53), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_22), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_59), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_14), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_51), .Y(n_110) );
INVx3_ASAP7_75t_L g111 ( .A(n_46), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_40), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_37), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_50), .Y(n_114) );
CKINVDCx14_ASAP7_75t_R g115 ( .A(n_58), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_61), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_13), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_64), .Y(n_118) );
NOR2xp33_ASAP7_75t_L g119 ( .A(n_36), .B(n_33), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_90), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_94), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_94), .Y(n_123) );
HB1xp67_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_96), .B(n_0), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_96), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_96), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_81), .Y(n_128) );
BUFx8_ASAP7_75t_L g129 ( .A(n_82), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_98), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_88), .Y(n_131) );
INVxp67_ASAP7_75t_L g132 ( .A(n_80), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_111), .B(n_1), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_98), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_111), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_86), .Y(n_136) );
INVx3_ASAP7_75t_L g137 ( .A(n_111), .Y(n_137) );
NAND2xp33_ASAP7_75t_L g138 ( .A(n_82), .B(n_79), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_115), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_85), .Y(n_140) );
AOI22xp5_ASAP7_75t_L g141 ( .A1(n_102), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_141) );
INVx2_ASAP7_75t_SL g142 ( .A(n_95), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_103), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_99), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_84), .Y(n_145) );
NOR2xp33_ASAP7_75t_R g146 ( .A(n_84), .B(n_34), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_82), .Y(n_147) );
CKINVDCx5p33_ASAP7_75t_R g148 ( .A(n_92), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_82), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_112), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_95), .B(n_3), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
NOR2xp33_ASAP7_75t_R g153 ( .A(n_92), .B(n_39), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_130), .Y(n_154) );
BUFx10_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
INVx2_ASAP7_75t_L g156 ( .A(n_131), .Y(n_156) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_123), .B(n_137), .Y(n_157) );
BUFx3_ASAP7_75t_L g158 ( .A(n_129), .Y(n_158) );
BUFx2_ASAP7_75t_L g159 ( .A(n_148), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_147), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_151), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_151), .B(n_110), .Y(n_162) );
BUFx4f_ASAP7_75t_L g163 ( .A(n_151), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_137), .B(n_105), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_128), .B(n_82), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_131), .Y(n_167) );
AND2x6_ASAP7_75t_L g168 ( .A(n_151), .B(n_110), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_149), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_128), .B(n_83), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_129), .B(n_106), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_129), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_131), .Y(n_174) );
OR2x2_ASAP7_75t_L g175 ( .A(n_124), .B(n_104), .Y(n_175) );
INVx2_ASAP7_75t_SL g176 ( .A(n_129), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_137), .B(n_118), .Y(n_177) );
CKINVDCx11_ASAP7_75t_R g178 ( .A(n_139), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
INVx4_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
INVx5_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_126), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
AO21x2_ASAP7_75t_L g184 ( .A1(n_138), .A2(n_114), .B(n_99), .Y(n_184) );
AND2x2_ASAP7_75t_L g185 ( .A(n_136), .B(n_105), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_126), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_140), .B(n_97), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_141), .A2(n_102), .B1(n_100), .B2(n_93), .Y(n_188) );
INVxp67_ASAP7_75t_SL g189 ( .A(n_132), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_127), .Y(n_190) );
BUFx8_ASAP7_75t_SL g191 ( .A(n_134), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_127), .Y(n_192) );
INVx3_ASAP7_75t_L g193 ( .A(n_135), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_120), .A2(n_121), .B1(n_152), .B2(n_150), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_189), .B(n_161), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_180), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_180), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_180), .Y(n_198) );
BUFx8_ASAP7_75t_L g199 ( .A(n_159), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_163), .B(n_172), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_185), .B(n_140), .Y(n_201) );
NOR2x1p5_ASAP7_75t_L g202 ( .A(n_154), .B(n_106), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_185), .A2(n_142), .B1(n_141), .B2(n_133), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_157), .B(n_120), .Y(n_204) );
AND2x6_ASAP7_75t_L g205 ( .A(n_158), .B(n_135), .Y(n_205) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_158), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_165), .B(n_121), .Y(n_207) );
NAND3xp33_ASAP7_75t_SL g208 ( .A(n_188), .B(n_116), .C(n_146), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_180), .B(n_143), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_182), .Y(n_210) );
NOR3xp33_ASAP7_75t_L g211 ( .A(n_188), .B(n_117), .C(n_101), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_194), .B(n_143), .Y(n_212) );
INVx2_ASAP7_75t_L g213 ( .A(n_186), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g214 ( .A(n_155), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_186), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_163), .B(n_152), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_170), .B(n_150), .Y(n_217) );
CKINVDCx11_ASAP7_75t_R g218 ( .A(n_178), .Y(n_218) );
BUFx12f_ASAP7_75t_L g219 ( .A(n_155), .Y(n_219) );
HB1xp67_ASAP7_75t_L g220 ( .A(n_159), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_163), .B(n_100), .Y(n_221) );
NAND2x2_ASAP7_75t_L g222 ( .A(n_175), .B(n_142), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_182), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_191), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_158), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_190), .Y(n_226) );
INVxp67_ASAP7_75t_L g227 ( .A(n_155), .Y(n_227) );
INVx2_ASAP7_75t_SL g228 ( .A(n_175), .Y(n_228) );
INVx5_ASAP7_75t_L g229 ( .A(n_162), .Y(n_229) );
NOR3xp33_ASAP7_75t_SL g230 ( .A(n_187), .B(n_116), .C(n_109), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_190), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_186), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_161), .B(n_122), .Y(n_233) );
BUFx3_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_163), .A2(n_125), .B1(n_122), .B2(n_144), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_186), .Y(n_236) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_176), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_161), .B(n_153), .Y(n_238) );
AND2x6_ASAP7_75t_SL g239 ( .A(n_155), .B(n_87), .Y(n_239) );
AO22x1_ASAP7_75t_L g240 ( .A1(n_162), .A2(n_108), .B1(n_89), .B2(n_107), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
CKINVDCx5p33_ASAP7_75t_R g242 ( .A(n_177), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_161), .B(n_144), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_162), .B(n_144), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_193), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_192), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_201), .B(n_162), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_228), .B(n_220), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_217), .B(n_176), .Y(n_249) );
OAI22xp5_ASAP7_75t_L g250 ( .A1(n_242), .A2(n_171), .B1(n_192), .B2(n_193), .Y(n_250) );
NAND2xp33_ASAP7_75t_L g251 ( .A(n_225), .B(n_168), .Y(n_251) );
BUFx12f_ASAP7_75t_L g252 ( .A(n_218), .Y(n_252) );
AND2x2_ASAP7_75t_L g253 ( .A(n_217), .B(n_193), .Y(n_253) );
AND2x4_ASAP7_75t_L g254 ( .A(n_229), .B(n_168), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_196), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_196), .Y(n_256) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_214), .B(n_162), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_218), .Y(n_258) );
INVx5_ASAP7_75t_L g259 ( .A(n_206), .Y(n_259) );
INVx3_ASAP7_75t_L g260 ( .A(n_198), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_204), .B(n_168), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_210), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_198), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_199), .Y(n_264) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_206), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_199), .Y(n_266) );
AOI21x1_ASAP7_75t_L g267 ( .A1(n_240), .A2(n_173), .B(n_160), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_195), .B(n_168), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_223), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_195), .B(n_168), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_234), .B(n_160), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_229), .B(n_168), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_195), .B(n_168), .Y(n_273) );
O2A1O1Ixp33_ASAP7_75t_L g274 ( .A1(n_211), .A2(n_166), .B(n_169), .C(n_173), .Y(n_274) );
INVx2_ASAP7_75t_L g275 ( .A(n_226), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_199), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_208), .A2(n_162), .B1(n_177), .B2(n_184), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_229), .B(n_227), .Y(n_278) );
INVx5_ASAP7_75t_L g279 ( .A(n_206), .Y(n_279) );
INVx5_ASAP7_75t_SL g280 ( .A(n_206), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
O2A1O1Ixp5_ASAP7_75t_L g282 ( .A1(n_200), .A2(n_164), .B(n_169), .C(n_107), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_203), .B(n_184), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_207), .B(n_162), .Y(n_284) );
INVx4_ASAP7_75t_L g285 ( .A(n_229), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g286 ( .A(n_219), .Y(n_286) );
INVx3_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_200), .A2(n_184), .B(n_164), .Y(n_288) );
AND2x4_ASAP7_75t_L g289 ( .A(n_234), .B(n_177), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_237), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_246), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_225), .Y(n_292) );
OR2x2_ASAP7_75t_L g293 ( .A(n_202), .B(n_144), .Y(n_293) );
HB1xp67_ASAP7_75t_L g294 ( .A(n_222), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_213), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_268), .Y(n_296) );
OAI22xp33_ASAP7_75t_L g297 ( .A1(n_264), .A2(n_219), .B1(n_222), .B2(n_242), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_267), .A2(n_244), .B(n_216), .Y(n_298) );
OAI21x1_ASAP7_75t_L g299 ( .A1(n_288), .A2(n_235), .B(n_216), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_267), .A2(n_245), .B(n_215), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_255), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_281), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_283), .B(n_212), .Y(n_303) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_284), .A2(n_209), .B(n_233), .Y(n_304) );
OA21x2_ASAP7_75t_L g305 ( .A1(n_282), .A2(n_243), .B(n_245), .Y(n_305) );
OAI21x1_ASAP7_75t_L g306 ( .A1(n_287), .A2(n_241), .B(n_213), .Y(n_306) );
INVx4_ASAP7_75t_L g307 ( .A(n_259), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_268), .B(n_197), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_281), .Y(n_309) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_248), .A2(n_221), .B1(n_177), .B2(n_205), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_255), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_281), .Y(n_312) );
OAI21x1_ASAP7_75t_L g313 ( .A1(n_287), .A2(n_241), .B(n_215), .Y(n_313) );
OAI21x1_ASAP7_75t_L g314 ( .A1(n_287), .A2(n_232), .B(n_236), .Y(n_314) );
AO21x1_ASAP7_75t_L g315 ( .A1(n_283), .A2(n_221), .B(n_236), .Y(n_315) );
HB1xp67_ASAP7_75t_L g316 ( .A(n_264), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_270), .Y(n_317) );
BUFx2_ASAP7_75t_L g318 ( .A(n_270), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_265), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_287), .A2(n_232), .B(n_238), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_249), .A2(n_177), .B1(n_205), .B2(n_237), .Y(n_321) );
OAI21x1_ASAP7_75t_L g322 ( .A1(n_290), .A2(n_156), .B(n_167), .Y(n_322) );
AO32x2_ASAP7_75t_L g323 ( .A1(n_250), .A2(n_285), .A3(n_277), .B1(n_230), .B2(n_279), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_262), .Y(n_324) );
BUFx6f_ASAP7_75t_L g325 ( .A(n_265), .Y(n_325) );
AO21x2_ASAP7_75t_L g326 ( .A1(n_262), .A2(n_174), .B(n_156), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_290), .A2(n_275), .B(n_295), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_289), .B(n_237), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_SL g330 ( .A1(n_271), .A2(n_119), .B(n_156), .C(n_183), .Y(n_330) );
AOI21xp5_ASAP7_75t_L g331 ( .A1(n_330), .A2(n_251), .B(n_249), .Y(n_331) );
NAND3xp33_ASAP7_75t_L g332 ( .A(n_310), .B(n_294), .C(n_293), .Y(n_332) );
BUFx4f_ASAP7_75t_SL g333 ( .A(n_327), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g334 ( .A1(n_303), .A2(n_266), .B1(n_276), .B2(n_257), .Y(n_334) );
AOI21xp5_ASAP7_75t_L g335 ( .A1(n_301), .A2(n_269), .B(n_291), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_324), .B(n_253), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_301), .A2(n_269), .B(n_291), .Y(n_337) );
OR2x6_ASAP7_75t_L g338 ( .A(n_327), .B(n_252), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g339 ( .A1(n_297), .A2(n_253), .B1(n_293), .B2(n_274), .C(n_286), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_301), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g341 ( .A1(n_302), .A2(n_275), .B1(n_247), .B2(n_261), .Y(n_341) );
AO21x2_ASAP7_75t_L g342 ( .A1(n_300), .A2(n_315), .B(n_328), .Y(n_342) );
O2A1O1Ixp33_ASAP7_75t_L g343 ( .A1(n_303), .A2(n_273), .B(n_261), .C(n_260), .Y(n_343) );
OAI22xp5_ASAP7_75t_L g344 ( .A1(n_302), .A2(n_280), .B1(n_289), .B2(n_292), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g345 ( .A1(n_316), .A2(n_224), .B1(n_258), .B2(n_252), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_296), .B(n_255), .Y(n_346) );
A2O1A1Ixp33_ASAP7_75t_L g347 ( .A1(n_309), .A2(n_263), .B(n_256), .C(n_295), .Y(n_347) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_309), .A2(n_224), .B1(n_289), .B2(n_177), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_296), .B(n_263), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_324), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_318), .B(n_263), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_312), .B(n_260), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_312), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_300), .A2(n_290), .B(n_295), .Y(n_354) );
NOR2x1_ASAP7_75t_L g355 ( .A(n_307), .B(n_278), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_317), .B(n_260), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_318), .B(n_239), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_307), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_353), .B(n_311), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_340), .B(n_311), .Y(n_360) );
OR2x2_ASAP7_75t_L g361 ( .A(n_340), .B(n_311), .Y(n_361) );
NAND4xp25_ASAP7_75t_L g362 ( .A(n_357), .B(n_317), .C(n_308), .D(n_321), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_354), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_342), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_350), .Y(n_365) );
INVx4_ASAP7_75t_L g366 ( .A(n_358), .Y(n_366) );
AND2x2_ASAP7_75t_L g367 ( .A(n_346), .B(n_315), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_349), .B(n_307), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_342), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_352), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_351), .B(n_307), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_335), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_333), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_347), .B(n_328), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_357), .A2(n_308), .B1(n_304), .B2(n_278), .Y(n_376) );
NOR4xp25_ASAP7_75t_SL g377 ( .A(n_339), .B(n_323), .C(n_320), .D(n_82), .Y(n_377) );
AND2x4_ASAP7_75t_L g378 ( .A(n_355), .B(n_319), .Y(n_378) );
NOR2xp33_ASAP7_75t_L g379 ( .A(n_333), .B(n_308), .Y(n_379) );
BUFx2_ASAP7_75t_L g380 ( .A(n_338), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_331), .A2(n_320), .B(n_306), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_336), .Y(n_382) );
INVxp67_ASAP7_75t_SL g383 ( .A(n_337), .Y(n_383) );
NOR2x1_ASAP7_75t_L g384 ( .A(n_332), .B(n_298), .Y(n_384) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_347), .Y(n_385) );
OAI22xp33_ASAP7_75t_L g386 ( .A1(n_334), .A2(n_329), .B1(n_304), .B2(n_319), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_338), .B(n_308), .Y(n_387) );
AND2x4_ASAP7_75t_L g388 ( .A(n_356), .B(n_319), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_344), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
NAND3xp33_ASAP7_75t_SL g392 ( .A(n_380), .B(n_345), .C(n_348), .Y(n_392) );
AND2x4_ASAP7_75t_L g393 ( .A(n_367), .B(n_326), .Y(n_393) );
OAI21xp5_ASAP7_75t_L g394 ( .A1(n_376), .A2(n_343), .B(n_299), .Y(n_394) );
INVxp67_ASAP7_75t_SL g395 ( .A(n_361), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_367), .B(n_323), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
INVx5_ASAP7_75t_SL g398 ( .A(n_378), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_367), .B(n_323), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_362), .A2(n_338), .B1(n_341), .B2(n_88), .C(n_91), .Y(n_400) );
NAND3xp33_ASAP7_75t_L g401 ( .A(n_362), .B(n_88), .C(n_91), .Y(n_401) );
INVx3_ASAP7_75t_L g402 ( .A(n_378), .Y(n_402) );
OR2x2_ASAP7_75t_L g403 ( .A(n_359), .B(n_298), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_364), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_360), .B(n_323), .Y(n_405) );
AOI221xp5_ASAP7_75t_L g406 ( .A1(n_386), .A2(n_88), .B1(n_91), .B2(n_260), .C(n_278), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_370), .Y(n_408) );
INVxp67_ASAP7_75t_SL g409 ( .A(n_359), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_365), .B(n_298), .Y(n_411) );
NAND4xp25_ASAP7_75t_L g412 ( .A(n_380), .B(n_4), .C(n_5), .D(n_6), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_369), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_360), .Y(n_414) );
XNOR2xp5_ASAP7_75t_L g415 ( .A(n_374), .B(n_278), .Y(n_415) );
NAND4xp25_ASAP7_75t_L g416 ( .A(n_374), .B(n_4), .C(n_5), .D(n_6), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_373), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_382), .B(n_298), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_369), .Y(n_419) );
OAI22xp5_ASAP7_75t_SL g420 ( .A1(n_374), .A2(n_329), .B1(n_323), .B2(n_325), .Y(n_420) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_387), .B(n_7), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_382), .B(n_299), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_368), .B(n_323), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_373), .Y(n_424) );
INVx3_ASAP7_75t_L g425 ( .A(n_378), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_368), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_372), .B(n_82), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_375), .B(n_326), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_382), .B(n_326), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_369), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_363), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_372), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_401), .A2(n_379), .B(n_387), .C(n_383), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_426), .B(n_371), .Y(n_435) );
AOI221xp5_ASAP7_75t_L g436 ( .A1(n_412), .A2(n_386), .B1(n_385), .B2(n_88), .C(n_91), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_390), .Y(n_437) );
NAND2xp5_ASAP7_75t_SL g438 ( .A(n_401), .B(n_366), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_432), .B(n_371), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_409), .B(n_371), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_407), .Y(n_441) );
INVx3_ASAP7_75t_L g442 ( .A(n_398), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_408), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_391), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_423), .B(n_375), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_414), .B(n_366), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_423), .B(n_375), .Y(n_448) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_416), .A2(n_366), .B1(n_389), .B2(n_378), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_427), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_395), .B(n_366), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_396), .B(n_385), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_427), .B(n_388), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_397), .B(n_388), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_397), .B(n_388), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_396), .B(n_388), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_412), .B(n_389), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_393), .B(n_383), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_399), .B(n_389), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_399), .B(n_384), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_393), .B(n_384), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_403), .B(n_363), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_402), .B(n_363), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_416), .B(n_7), .C(n_9), .D(n_10), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_393), .B(n_377), .Y(n_465) );
HB1xp67_ASAP7_75t_L g466 ( .A(n_429), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_391), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_417), .Y(n_468) );
INVx3_ASAP7_75t_L g469 ( .A(n_398), .Y(n_469) );
OR2x2_ASAP7_75t_L g470 ( .A(n_403), .B(n_10), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_415), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_417), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_393), .B(n_377), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_424), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_402), .B(n_381), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_405), .B(n_381), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_405), .B(n_381), .Y(n_477) );
OAI21x1_ASAP7_75t_L g478 ( .A1(n_394), .A2(n_306), .B(n_313), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_404), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_421), .B(n_11), .Y(n_480) );
OAI221xp5_ASAP7_75t_L g481 ( .A1(n_400), .A2(n_91), .B1(n_329), .B2(n_290), .C(n_256), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_428), .B(n_82), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_424), .Y(n_483) );
INVxp67_ASAP7_75t_L g484 ( .A(n_392), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_420), .B(n_319), .Y(n_485) );
OR2x2_ASAP7_75t_L g486 ( .A(n_398), .B(n_11), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_411), .B(n_12), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_404), .Y(n_488) );
AND2x2_ASAP7_75t_L g489 ( .A(n_428), .B(n_326), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_441), .B(n_411), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_444), .Y(n_491) );
INVx4_ASAP7_75t_L g492 ( .A(n_442), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_443), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_435), .B(n_418), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_482), .B(n_402), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_438), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_434), .Y(n_497) );
OAI31xp33_ASAP7_75t_L g498 ( .A1(n_464), .A2(n_420), .A3(n_415), .B(n_425), .Y(n_498) );
NOR2x1_ASAP7_75t_SL g499 ( .A(n_486), .B(n_404), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_471), .Y(n_500) );
NAND4xp25_ASAP7_75t_SL g501 ( .A(n_436), .B(n_406), .C(n_398), .D(n_422), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_484), .B(n_402), .C(n_425), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_482), .B(n_425), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_452), .B(n_428), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_437), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_468), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_472), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_474), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_439), .B(n_425), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_483), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_440), .B(n_398), .Y(n_512) );
INVx1_ASAP7_75t_SL g513 ( .A(n_447), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_466), .Y(n_514) );
NOR2x1_ASAP7_75t_L g515 ( .A(n_438), .B(n_428), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_445), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_470), .Y(n_517) );
OAI31xp33_ASAP7_75t_L g518 ( .A1(n_433), .A2(n_419), .A3(n_430), .B(n_410), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_446), .B(n_430), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_446), .B(n_413), .Y(n_520) );
INVxp67_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_451), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_448), .B(n_413), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_452), .B(n_410), .Y(n_524) );
AOI221xp5_ASAP7_75t_L g525 ( .A1(n_457), .A2(n_419), .B1(n_431), .B2(n_16), .C(n_17), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_454), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_455), .Y(n_527) );
INVxp67_ASAP7_75t_L g528 ( .A(n_485), .Y(n_528) );
O2A1O1Ixp33_ASAP7_75t_L g529 ( .A1(n_433), .A2(n_419), .B(n_431), .C(n_329), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_448), .B(n_431), .Y(n_530) );
NAND2x1p5_ASAP7_75t_L g531 ( .A(n_442), .B(n_325), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_456), .B(n_12), .Y(n_532) );
OR2x2_ASAP7_75t_L g533 ( .A(n_453), .B(n_15), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_487), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_459), .B(n_15), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_450), .B(n_16), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_462), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_457), .B(n_305), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_445), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_467), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_460), .B(n_305), .Y(n_541) );
OR2x2_ASAP7_75t_L g542 ( .A(n_458), .B(n_314), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_489), .B(n_314), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_449), .B(n_19), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_467), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_479), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_489), .B(n_476), .Y(n_547) );
INVxp67_ASAP7_75t_L g548 ( .A(n_458), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_493), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_514), .Y(n_550) );
OAI321xp33_ASAP7_75t_L g551 ( .A1(n_521), .A2(n_480), .A3(n_461), .B1(n_481), .B2(n_465), .C(n_460), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_500), .B(n_442), .Y(n_552) );
AOI221xp5_ASAP7_75t_SL g553 ( .A1(n_521), .A2(n_461), .B1(n_477), .B2(n_476), .C(n_473), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_547), .B(n_477), .Y(n_554) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_498), .A2(n_473), .B(n_475), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g556 ( .A1(n_525), .A2(n_469), .B(n_475), .Y(n_556) );
NOR2xp33_ASAP7_75t_L g557 ( .A(n_500), .B(n_469), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_522), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_525), .A2(n_475), .B1(n_469), .B2(n_463), .Y(n_559) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_502), .A2(n_479), .B1(n_488), .B2(n_329), .C(n_279), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_517), .B(n_488), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_497), .Y(n_562) );
CKINVDCx14_ASAP7_75t_R g563 ( .A(n_519), .Y(n_563) );
AOI32xp33_ASAP7_75t_L g564 ( .A1(n_502), .A2(n_463), .A3(n_478), .B1(n_289), .B2(n_254), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_526), .B(n_463), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_505), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_534), .A2(n_167), .B1(n_174), .B2(n_183), .C(n_179), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_527), .B(n_478), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_548), .B(n_305), .Y(n_569) );
O2A1O1Ixp33_ASAP7_75t_L g570 ( .A1(n_529), .A2(n_183), .B(n_174), .C(n_167), .Y(n_570) );
INVxp67_ASAP7_75t_L g571 ( .A(n_499), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_506), .Y(n_572) );
OAI211xp5_ASAP7_75t_L g573 ( .A1(n_496), .A2(n_259), .B(n_279), .C(n_285), .Y(n_573) );
OAI32xp33_ASAP7_75t_L g574 ( .A1(n_528), .A2(n_285), .A3(n_21), .B1(n_23), .B2(n_24), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g575 ( .A1(n_528), .A2(n_325), .B1(n_319), .B2(n_280), .Y(n_575) );
NOR2xp33_ASAP7_75t_R g576 ( .A(n_492), .B(n_20), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_491), .B(n_513), .Y(n_577) );
OAI322xp33_ASAP7_75t_L g578 ( .A1(n_548), .A2(n_179), .A3(n_325), .B1(n_319), .B2(n_285), .C1(n_265), .C2(n_43), .Y(n_578) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_515), .A2(n_272), .A3(n_254), .B1(n_313), .B2(n_322), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_537), .B(n_305), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g581 ( .A1(n_529), .A2(n_325), .B(n_259), .Y(n_581) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_492), .A2(n_496), .B1(n_512), .B2(n_533), .Y(n_582) );
OAI322xp33_ASAP7_75t_L g583 ( .A1(n_535), .A2(n_325), .A3(n_265), .B1(n_31), .B2(n_32), .C1(n_41), .C2(n_45), .Y(n_583) );
INVxp67_ASAP7_75t_L g584 ( .A(n_490), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_493), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_507), .Y(n_586) );
NAND3x2_ASAP7_75t_L g587 ( .A(n_532), .B(n_272), .C(n_254), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_510), .Y(n_588) );
OAI21xp5_ASAP7_75t_L g589 ( .A1(n_544), .A2(n_205), .B(n_254), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_509), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_520), .B(n_26), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_511), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_536), .A2(n_177), .B1(n_205), .B2(n_272), .C1(n_280), .C2(n_279), .Y(n_593) );
AOI21xp5_ASAP7_75t_L g594 ( .A1(n_581), .A2(n_518), .B(n_492), .Y(n_594) );
OAI21xp33_ASAP7_75t_L g595 ( .A1(n_555), .A2(n_504), .B(n_524), .Y(n_595) );
INVxp67_ASAP7_75t_SL g596 ( .A(n_571), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
OAI22xp5_ASAP7_75t_L g598 ( .A1(n_563), .A2(n_494), .B1(n_523), .B2(n_544), .Y(n_598) );
O2A1O1Ixp33_ASAP7_75t_L g599 ( .A1(n_551), .A2(n_538), .B(n_542), .C(n_531), .Y(n_599) );
INVx2_ASAP7_75t_SL g600 ( .A(n_576), .Y(n_600) );
A2O1A1Ixp33_ASAP7_75t_L g601 ( .A1(n_553), .A2(n_495), .B(n_503), .C(n_530), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_582), .A2(n_501), .B1(n_543), .B2(n_541), .Y(n_602) );
OAI31xp33_ASAP7_75t_L g603 ( .A1(n_560), .A2(n_531), .A3(n_546), .B(n_540), .Y(n_603) );
INVx1_ASAP7_75t_SL g604 ( .A(n_577), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_558), .Y(n_605) );
XNOR2x1_ASAP7_75t_L g606 ( .A(n_587), .B(n_550), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_549), .Y(n_607) );
INVxp67_ASAP7_75t_L g608 ( .A(n_568), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_584), .B(n_539), .Y(n_609) );
NOR2xp67_ASAP7_75t_L g610 ( .A(n_581), .B(n_545), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_562), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_588), .B(n_545), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_554), .B(n_516), .Y(n_613) );
INVxp33_ASAP7_75t_SL g614 ( .A(n_552), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_565), .B(n_516), .Y(n_615) );
OAI21xp33_ASAP7_75t_L g616 ( .A1(n_559), .A2(n_508), .B(n_272), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_570), .B(n_508), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_566), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_572), .B(n_27), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_586), .B(n_47), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_590), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_597), .B(n_595), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_596), .A2(n_570), .B(n_573), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g624 ( .A1(n_596), .A2(n_556), .B(n_573), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_609), .Y(n_625) );
INVx3_ASAP7_75t_L g626 ( .A(n_600), .Y(n_626) );
INVxp67_ASAP7_75t_L g627 ( .A(n_606), .Y(n_627) );
CKINVDCx20_ASAP7_75t_L g628 ( .A(n_614), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_602), .A2(n_557), .B1(n_592), .B2(n_591), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_601), .A2(n_564), .B(n_589), .C(n_579), .Y(n_630) );
AOI21xp33_ASAP7_75t_L g631 ( .A1(n_599), .A2(n_574), .B(n_575), .Y(n_631) );
A2O1A1Ixp33_ASAP7_75t_L g632 ( .A1(n_601), .A2(n_585), .B(n_569), .C(n_567), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_604), .Y(n_633) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_608), .A2(n_583), .B1(n_578), .B2(n_567), .C(n_580), .Y(n_634) );
AOI322xp5_ASAP7_75t_L g635 ( .A1(n_616), .A2(n_593), .A3(n_279), .B1(n_259), .B2(n_265), .C1(n_60), .C2(n_63), .Y(n_635) );
NOR3xp33_ASAP7_75t_L g636 ( .A(n_598), .B(n_322), .C(n_52), .Y(n_636) );
A2O1A1Ixp33_ASAP7_75t_L g637 ( .A1(n_594), .A2(n_279), .B(n_259), .C(n_292), .Y(n_637) );
OAI221xp5_ASAP7_75t_SL g638 ( .A1(n_627), .A2(n_603), .B1(n_608), .B2(n_612), .C(n_605), .Y(n_638) );
NAND3xp33_ASAP7_75t_L g639 ( .A(n_632), .B(n_617), .C(n_620), .Y(n_639) );
AOI211xp5_ASAP7_75t_L g640 ( .A1(n_631), .A2(n_610), .B(n_617), .C(n_612), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_633), .A2(n_621), .B1(n_618), .B2(n_611), .C(n_615), .Y(n_641) );
AOI222xp33_ASAP7_75t_L g642 ( .A1(n_624), .A2(n_607), .B1(n_613), .B2(n_619), .C1(n_205), .C2(n_280), .Y(n_642) );
NOR3xp33_ASAP7_75t_L g643 ( .A(n_630), .B(n_49), .C(n_54), .Y(n_643) );
OAI211xp5_ASAP7_75t_L g644 ( .A1(n_626), .A2(n_259), .B(n_292), .C(n_181), .Y(n_644) );
OAI221xp5_ASAP7_75t_SL g645 ( .A1(n_629), .A2(n_626), .B1(n_637), .B2(n_623), .C(n_622), .Y(n_645) );
OAI21xp5_ASAP7_75t_L g646 ( .A1(n_636), .A2(n_280), .B(n_181), .Y(n_646) );
NOR3xp33_ASAP7_75t_L g647 ( .A(n_634), .B(n_56), .C(n_66), .Y(n_647) );
NOR2x1_ASAP7_75t_R g648 ( .A(n_643), .B(n_628), .Y(n_648) );
BUFx12f_ASAP7_75t_L g649 ( .A(n_645), .Y(n_649) );
OAI211xp5_ASAP7_75t_SL g650 ( .A1(n_640), .A2(n_635), .B(n_625), .C(n_70), .Y(n_650) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_638), .A2(n_292), .B(n_181), .Y(n_651) );
NAND4xp25_ASAP7_75t_L g652 ( .A(n_647), .B(n_67), .C(n_69), .D(n_71), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_648), .Y(n_653) );
XNOR2x1_ASAP7_75t_L g654 ( .A(n_649), .B(n_639), .Y(n_654) );
NOR4xp25_ASAP7_75t_L g655 ( .A(n_650), .B(n_641), .C(n_644), .D(n_646), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_653), .B(n_642), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_654), .B(n_651), .Y(n_657) );
INVx3_ASAP7_75t_L g658 ( .A(n_656), .Y(n_658) );
OAI22xp5_ASAP7_75t_SL g659 ( .A1(n_657), .A2(n_655), .B1(n_652), .B2(n_292), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_659), .A2(n_181), .B1(n_74), .B2(n_76), .Y(n_660) );
AOI31xp33_ASAP7_75t_L g661 ( .A1(n_660), .A2(n_658), .A3(n_78), .B(n_73), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_661), .Y(n_662) );
AOI21xp5_ASAP7_75t_L g663 ( .A1(n_662), .A2(n_181), .B(n_657), .Y(n_663) );
endmodule