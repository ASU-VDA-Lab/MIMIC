module fake_jpeg_5423_n_279 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx8_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_9),
.B(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_17),
.B(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_34),
.B(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_26),
.Y(n_38)
);

BUFx2_ASAP7_75t_SL g55 ( 
.A(n_38),
.Y(n_55)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_23),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_35),
.A2(n_16),
.B(n_30),
.C(n_24),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_42),
.B(n_45),
.Y(n_77)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_44),
.B(n_49),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_35),
.Y(n_45)
);

INVx4_ASAP7_75t_SL g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_32),
.A2(n_24),
.B1(n_30),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_50),
.A2(n_18),
.B1(n_19),
.B2(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_28),
.Y(n_54)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_28),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_56),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_34),
.B(n_22),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_62),
.Y(n_82)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_34),
.B(n_30),
.Y(n_63)
);

NAND3xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_41),
.C(n_34),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_66),
.A2(n_75),
.B1(n_87),
.B2(n_63),
.Y(n_90)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_70),
.Y(n_89)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_83),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_42),
.A2(n_39),
.B1(n_32),
.B2(n_34),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_45),
.A2(n_32),
.B1(n_44),
.B2(n_39),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_61),
.B1(n_53),
.B2(n_51),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_36),
.B(n_16),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_25),
.B1(n_36),
.B2(n_32),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_85),
.A2(n_60),
.B1(n_25),
.B2(n_53),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_47),
.A2(n_41),
.B1(n_17),
.B2(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_88),
.B(n_90),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_47),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_91),
.B(n_95),
.Y(n_119)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_76),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_94),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_81),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_96),
.A2(n_101),
.B1(n_69),
.B2(n_80),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_71),
.A2(n_51),
.B1(n_61),
.B2(n_60),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_98),
.Y(n_113)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_103),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_77),
.A2(n_74),
.B1(n_68),
.B2(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_62),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_102),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_67),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_84),
.B(n_65),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_68),
.B(n_49),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_106),
.A2(n_27),
.B(n_19),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_64),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_107),
.B(n_110),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_23),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_41),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_109),
.A2(n_111),
.B1(n_97),
.B2(n_78),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_64),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_25),
.B1(n_59),
.B2(n_22),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_111),
.A2(n_80),
.B1(n_19),
.B2(n_18),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_96),
.A2(n_40),
.B(n_46),
.C(n_64),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_112),
.A2(n_123),
.B1(n_126),
.B2(n_106),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_118),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_116),
.A2(n_124),
.B1(n_129),
.B2(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_108),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_99),
.A2(n_103),
.B1(n_95),
.B2(n_101),
.Y(n_124)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_128),
.B(n_131),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_100),
.A2(n_46),
.B1(n_40),
.B2(n_33),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_91),
.B(n_29),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_130),
.B(n_134),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_52),
.C(n_46),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_52),
.C(n_72),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_72),
.C(n_40),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_127),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_142),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_124),
.A2(n_90),
.B1(n_109),
.B2(n_102),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_139),
.A2(n_150),
.B1(n_126),
.B2(n_112),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_153),
.B1(n_157),
.B2(n_116),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_117),
.A2(n_94),
.B(n_105),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_135),
.Y(n_170)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_145),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_104),
.Y(n_146)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_146),
.Y(n_165)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_113),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_109),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_149),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_108),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_98),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_156),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_121),
.A2(n_29),
.B(n_20),
.Y(n_153)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_113),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_154),
.B(n_155),
.Y(n_182)
);

INVx13_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_117),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_125),
.A2(n_29),
.B(n_20),
.Y(n_157)
);

XOR2x2_ASAP7_75t_SL g158 ( 
.A(n_120),
.B(n_41),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_158),
.B(n_135),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g159 ( 
.A(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_137),
.B(n_133),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_162),
.B(n_170),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_137),
.B(n_155),
.C(n_138),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_164),
.B(n_176),
.C(n_177),
.Y(n_186)
);

NOR2xp67_ASAP7_75t_R g169 ( 
.A(n_158),
.B(n_120),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_169),
.A2(n_184),
.B1(n_178),
.B2(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_173),
.A2(n_184),
.B1(n_157),
.B2(n_147),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_174),
.A2(n_175),
.B1(n_179),
.B2(n_180),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_140),
.A2(n_129),
.B1(n_130),
.B2(n_112),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_138),
.C(n_156),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_123),
.C(n_128),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_159),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_150),
.A2(n_131),
.B1(n_40),
.B2(n_20),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_139),
.A2(n_131),
.B1(n_40),
.B2(n_22),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_149),
.B(n_92),
.Y(n_181)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_181),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_15),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_183),
.B(n_142),
.C(n_136),
.Y(n_196)
);

OAI22x1_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_160),
.B1(n_159),
.B2(n_145),
.Y(n_184)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_160),
.Y(n_191)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_191),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_192),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_201),
.C(n_15),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_163),
.B(n_152),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NOR3xp33_ASAP7_75t_L g206 ( 
.A(n_198),
.B(n_199),
.C(n_205),
.Y(n_206)
);

CKINVDCx14_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_159),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_200),
.A2(n_202),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_141),
.C(n_152),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_203),
.A2(n_18),
.B1(n_154),
.B2(n_31),
.Y(n_216)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_195),
.B(n_173),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_209),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_189),
.A2(n_167),
.B1(n_182),
.B2(n_176),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_208),
.A2(n_211),
.B1(n_215),
.B2(n_213),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_162),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_165),
.B1(n_88),
.B2(n_27),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_154),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_214),
.B(n_217),
.C(n_196),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_216),
.A2(n_222),
.B1(n_193),
.B2(n_188),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_15),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_219),
.B(n_200),
.Y(n_232)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_15),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_15),
.B1(n_2),
.B2(n_3),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_185),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_98),
.B1(n_40),
.B2(n_31),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_236),
.B1(n_237),
.B2(n_10),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_235),
.C(n_237),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_228),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_212),
.A2(n_198),
.B(n_191),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_229),
.B(n_233),
.Y(n_249)
);

BUFx24_ASAP7_75t_SL g230 ( 
.A(n_214),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_230),
.B(n_234),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_211),
.A2(n_200),
.B1(n_187),
.B2(n_31),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_231),
.A2(n_216),
.B1(n_222),
.B2(n_210),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_238),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_218),
.A2(n_9),
.B(n_14),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_223),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_37),
.C(n_15),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_217),
.B(n_37),
.C(n_2),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_37),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_235),
.C(n_238),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_241),
.B(n_245),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_232),
.A2(n_206),
.B1(n_219),
.B2(n_220),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_243),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_247),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_226),
.B(n_37),
.C(n_4),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_226),
.B(n_9),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_7),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_246),
.B(n_8),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_255),
.C(n_257),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_256),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_10),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_6),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_7),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_250),
.B(n_5),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_11),
.A3(n_12),
.B1(n_13),
.B2(n_14),
.C1(n_246),
.C2(n_254),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_253),
.A2(n_241),
.B(n_239),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_264),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_251),
.A2(n_239),
.B1(n_245),
.B2(n_243),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_11),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_248),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_12),
.B(n_13),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_258),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_268),
.A2(n_269),
.B(n_270),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_11),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_SL g273 ( 
.A(n_267),
.B(n_261),
.C(n_262),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_272),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_276),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_277),
.B(n_275),
.Y(n_278)
);

XNOR2x2_ASAP7_75t_SL g279 ( 
.A(n_278),
.B(n_274),
.Y(n_279)
);


endmodule