module fake_jpeg_619_n_445 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_445);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_445;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx3_ASAP7_75t_SL g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx4f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_45),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_8),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_46),
.B(n_70),
.Y(n_128)
);

BUFx24_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_56),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_49),
.Y(n_127)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_51),
.Y(n_134)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_23),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_53),
.A2(n_35),
.B1(n_33),
.B2(n_18),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_54),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_23),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_21),
.B(n_8),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_62),
.Y(n_100)
);

HB1xp67_ASAP7_75t_L g59 ( 
.A(n_17),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_59),
.Y(n_108)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_61),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_26),
.B(n_8),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_65),
.Y(n_94)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_66),
.Y(n_135)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_15),
.B(n_9),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_72),
.B(n_75),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_22),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_77),
.Y(n_117)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_78),
.B(n_85),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_9),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_84),
.Y(n_103)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_17),
.Y(n_80)
);

NAND2xp33_ASAP7_75t_SL g110 ( 
.A(n_80),
.B(n_82),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_81),
.B(n_83),
.Y(n_133)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_18),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_17),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_31),
.Y(n_84)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_27),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_86),
.B(n_43),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_88),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_44),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_93),
.B(n_105),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_66),
.A2(n_20),
.B1(n_43),
.B2(n_40),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_104),
.A2(n_109),
.B1(n_119),
.B2(n_126),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_53),
.B(n_35),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_122),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_20),
.B1(n_43),
.B2(n_40),
.Y(n_109)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_44),
.B(n_39),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g158 ( 
.A1(n_112),
.A2(n_47),
.B(n_15),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_52),
.B(n_19),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_86),
.B(n_19),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_114),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_55),
.A2(n_39),
.B1(n_37),
.B2(n_18),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_115),
.A2(n_41),
.B1(n_28),
.B2(n_29),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_43),
.B1(n_40),
.B2(n_18),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_57),
.B1(n_54),
.B2(n_61),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_40),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_63),
.B(n_41),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_123),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_64),
.B(n_33),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_18),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_73),
.B(n_18),
.C(n_37),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_81),
.C(n_77),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_74),
.A2(n_18),
.B1(n_36),
.B2(n_34),
.Y(n_126)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_111),
.Y(n_138)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_138),
.Y(n_183)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_139),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_140),
.B(n_161),
.Y(n_218)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_141),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_142),
.B(n_170),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_36),
.B1(n_28),
.B2(n_34),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_143),
.A2(n_144),
.B1(n_178),
.B2(n_179),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_51),
.B1(n_45),
.B2(n_49),
.Y(n_144)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_146),
.Y(n_198)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_95),
.Y(n_147)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_147),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_156),
.B1(n_117),
.B2(n_97),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_93),
.B(n_87),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_149),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g151 ( 
.A(n_97),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_151),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_152),
.B(n_122),
.C(n_118),
.Y(n_190)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_153),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_154),
.Y(n_199)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_158),
.B(n_177),
.Y(n_212)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_99),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_100),
.A2(n_29),
.B1(n_83),
.B2(n_69),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_110),
.A2(n_47),
.B(n_65),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_168),
.B(n_118),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_105),
.A2(n_71),
.B1(n_24),
.B2(n_10),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_164),
.A2(n_127),
.B1(n_107),
.B2(n_131),
.Y(n_210)
);

A2O1A1Ixp33_ASAP7_75t_L g165 ( 
.A1(n_103),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_165)
);

A2O1A1Ixp33_ASAP7_75t_L g222 ( 
.A1(n_165),
.A2(n_180),
.B(n_101),
.C(n_13),
.Y(n_222)
);

INVx6_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_167),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_110),
.A2(n_24),
.B(n_10),
.Y(n_168)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_99),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_91),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_91),
.Y(n_172)
);

AO22x1_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_24),
.B1(n_2),
.B2(n_1),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_98),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_125),
.B(n_3),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_175),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_98),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_118),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_102),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_128),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_117),
.A2(n_3),
.B1(n_6),
.B2(n_10),
.Y(n_179)
);

AOI21xp33_ASAP7_75t_L g180 ( 
.A1(n_128),
.A2(n_3),
.B(n_10),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_108),
.B(n_122),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_181),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_90),
.B(n_11),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_186),
.A2(n_210),
.B1(n_211),
.B2(n_147),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_196),
.C(n_138),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_139),
.A2(n_115),
.B1(n_137),
.B2(n_136),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_192),
.A2(n_193),
.B1(n_200),
.B2(n_221),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_148),
.A2(n_90),
.B1(n_137),
.B2(n_134),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_108),
.C(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_142),
.A2(n_134),
.B1(n_120),
.B2(n_127),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_154),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_214),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_166),
.A2(n_133),
.B(n_130),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g238 ( 
.A1(n_204),
.A2(n_207),
.B(n_162),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_144),
.A2(n_134),
.B1(n_120),
.B2(n_127),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_209),
.A2(n_215),
.B1(n_171),
.B2(n_172),
.Y(n_245)
);

AOI22x1_ASAP7_75t_SL g211 ( 
.A1(n_153),
.A2(n_107),
.B1(n_101),
.B2(n_135),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_152),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_169),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_181),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_166),
.A2(n_159),
.B1(n_170),
.B2(n_169),
.Y(n_215)
);

OA22x2_ASAP7_75t_L g216 ( 
.A1(n_145),
.A2(n_135),
.B1(n_132),
.B2(n_116),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_216),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_154),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_220),
.B(n_151),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_168),
.A2(n_92),
.B1(n_116),
.B2(n_132),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_222),
.B(n_95),
.Y(n_250)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

HB1xp67_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_228),
.B(n_249),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_173),
.B1(n_163),
.B2(n_150),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_229),
.A2(n_238),
.B(n_241),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_165),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_244),
.Y(n_271)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_195),
.Y(n_231)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_231),
.Y(n_286)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_195),
.Y(n_232)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_198),
.Y(n_233)
);

INVx13_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_207),
.A2(n_162),
.B(n_181),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_211),
.B(n_218),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_206),
.B(n_149),
.Y(n_236)
);

NOR3xp33_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_239),
.C(n_246),
.Y(n_276)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_189),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_237),
.B(n_219),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_206),
.B(n_149),
.Y(n_239)
);

MAJx2_ASAP7_75t_L g240 ( 
.A(n_205),
.B(n_213),
.C(n_187),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_146),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_204),
.A2(n_157),
.B(n_178),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_183),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_242),
.B(n_258),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_177),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_243),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_187),
.B(n_165),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_245),
.A2(n_248),
.B1(n_193),
.B2(n_184),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_180),
.Y(n_246)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_203),
.B(n_173),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_247),
.Y(n_266)
);

AND2x2_ASAP7_75t_SL g249 ( 
.A(n_196),
.B(n_194),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_250),
.A2(n_251),
.B(n_255),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_194),
.A2(n_176),
.B(n_174),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_203),
.B(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_253),
.Y(n_273)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_212),
.B(n_201),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_259),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_201),
.A2(n_96),
.B1(n_131),
.B2(n_151),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_256),
.B(n_161),
.C(n_223),
.Y(n_284)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_190),
.B(n_141),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_199),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_260),
.B(n_188),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_249),
.A2(n_186),
.B1(n_209),
.B2(n_215),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_261),
.A2(n_268),
.B1(n_277),
.B2(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_226),
.A2(n_184),
.B1(n_192),
.B2(n_200),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_270),
.B1(n_278),
.B2(n_283),
.Y(n_300)
);

OA21x2_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_221),
.B(n_216),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_263),
.B(n_290),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_238),
.A2(n_222),
.B(n_197),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_264),
.A2(n_267),
.B(n_250),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_257),
.A2(n_217),
.B1(n_185),
.B2(n_191),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_234),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_275),
.B(n_243),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_249),
.A2(n_217),
.B1(n_216),
.B2(n_191),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_257),
.A2(n_216),
.B1(n_211),
.B2(n_220),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_279),
.Y(n_308)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_254),
.B(n_216),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_241),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_226),
.A2(n_202),
.B1(n_199),
.B2(n_223),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_249),
.C(n_240),
.Y(n_322)
);

INVx13_ASAP7_75t_L g285 ( 
.A(n_233),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g318 ( 
.A(n_285),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_247),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_245),
.A2(n_92),
.B1(n_188),
.B2(n_96),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_231),
.B(n_219),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_293),
.B(n_295),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_228),
.B(n_155),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_265),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_302),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_313),
.B(n_319),
.Y(n_347)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_265),
.Y(n_298)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_298),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_299),
.B(n_270),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_294),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_269),
.B(n_232),
.Y(n_303)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_303),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_314),
.B1(n_317),
.B2(n_266),
.Y(n_336)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_274),
.B(n_240),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_322),
.C(n_323),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_286),
.B(n_251),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_310),
.B(n_311),
.Y(n_349)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_267),
.A2(n_288),
.B(n_282),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_227),
.B1(n_259),
.B2(n_256),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_286),
.B(n_227),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_315),
.B(n_320),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_316),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_277),
.A2(n_252),
.B1(n_247),
.B2(n_246),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_288),
.A2(n_225),
.B(n_224),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_282),
.A2(n_229),
.B(n_225),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_324),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_274),
.B(n_230),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_280),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_284),
.B(n_244),
.C(n_236),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_325),
.B(n_273),
.C(n_271),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_300),
.A2(n_266),
.B1(n_275),
.B2(n_281),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_326),
.A2(n_336),
.B1(n_340),
.B2(n_344),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_291),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_330),
.B(n_346),
.Y(n_353)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_307),
.A2(n_263),
.B(n_278),
.C(n_273),
.Y(n_332)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_332),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_301),
.A2(n_268),
.B1(n_280),
.B2(n_287),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_333),
.A2(n_345),
.B1(n_312),
.B2(n_302),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_338),
.B(n_325),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_276),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_339),
.B(n_342),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_300),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_340)
);

XNOR2x1_ASAP7_75t_L g341 ( 
.A(n_314),
.B(n_299),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_341),
.B(n_343),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_271),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_301),
.A2(n_263),
.B1(n_283),
.B2(n_292),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_303),
.A2(n_239),
.B1(n_290),
.B2(n_255),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_258),
.Y(n_346)
);

AND2x4_ASAP7_75t_SL g350 ( 
.A(n_310),
.B(n_285),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_350),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_296),
.A2(n_237),
.B1(n_272),
.B2(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_318),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_357),
.B(n_372),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_341),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_362),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_307),
.B1(n_298),
.B2(n_313),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_349),
.B1(n_350),
.B2(n_344),
.Y(n_376)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_360),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_327),
.B(n_323),
.C(n_317),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_361),
.B(n_364),
.C(n_370),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_321),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_319),
.B(n_297),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_363),
.A2(n_374),
.B(n_347),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_305),
.C(n_306),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_337),
.Y(n_365)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_365),
.Y(n_386)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_366),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_315),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_368),
.B(n_353),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_343),
.B(n_311),
.C(n_320),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_337),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_328),
.B1(n_340),
.B2(n_349),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_332),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_376),
.A2(n_382),
.B1(n_388),
.B2(n_355),
.Y(n_394)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_380),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_354),
.B(n_312),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_381),
.B(n_383),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_367),
.A2(n_355),
.B1(n_359),
.B2(n_350),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_347),
.C(n_326),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_364),
.B(n_348),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_384),
.B(n_389),
.Y(n_399)
);

MAJx2_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_391),
.C(n_272),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_362),
.B(n_351),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_353),
.B(n_329),
.C(n_318),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_361),
.C(n_368),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_358),
.B(n_332),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_394),
.A2(n_403),
.B1(n_147),
.B2(n_146),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_401),
.Y(n_409)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_356),
.Y(n_396)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_396),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_387),
.A2(n_332),
.B1(n_369),
.B2(n_370),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_397),
.A2(n_389),
.B1(n_383),
.B2(n_386),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_369),
.C(n_366),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_400),
.B(n_375),
.C(n_377),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_329),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_242),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_405),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_387),
.A2(n_260),
.B1(n_253),
.B2(n_272),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_378),
.Y(n_404)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_404),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_376),
.A2(n_233),
.B(n_155),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_406),
.A2(n_382),
.B(n_403),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_398),
.B(n_379),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_407),
.B(n_410),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_411),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_377),
.C(n_392),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_412),
.B(n_416),
.Y(n_425)
);

OAI22x1_ASAP7_75t_L g414 ( 
.A1(n_393),
.A2(n_167),
.B1(n_95),
.B2(n_129),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_414),
.B(n_415),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_401),
.B(n_167),
.C(n_129),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_399),
.Y(n_418)
);

AOI322xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_396),
.A3(n_406),
.B1(n_397),
.B2(n_405),
.C1(n_129),
.C2(n_12),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_412),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_421),
.B(n_422),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_400),
.C(n_402),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_427),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_409),
.B(n_396),
.C(n_129),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_417),
.A2(n_12),
.B(n_14),
.Y(n_428)
);

OAI21x1_ASAP7_75t_L g436 ( 
.A1(n_428),
.A2(n_415),
.B(n_14),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_413),
.A2(n_12),
.B(n_14),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_429),
.B(n_419),
.Y(n_434)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_423),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_430),
.B(n_431),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_425),
.Y(n_431)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_434),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_416),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_435),
.A2(n_436),
.B(n_428),
.Y(n_438)
);

AO21x1_ASAP7_75t_L g441 ( 
.A1(n_438),
.A2(n_434),
.B(n_414),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g439 ( 
.A1(n_433),
.A2(n_432),
.B(n_420),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_439),
.A2(n_422),
.B(n_427),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_441),
.B(n_442),
.C(n_437),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_443),
.A2(n_440),
.B(n_424),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_424),
.Y(n_445)
);


endmodule