module real_jpeg_18258_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_412;
wire n_120;
wire n_155;
wire n_405;
wire n_319;
wire n_493;
wire n_93;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_524),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_0),
.B(n_525),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_1),
.A2(n_113),
.B1(n_298),
.B2(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_1),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_1),
.A2(n_300),
.B1(n_413),
.B2(n_416),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_SL g470 ( 
.A1(n_1),
.A2(n_300),
.B1(n_471),
.B2(n_476),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_2),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_2),
.Y(n_132)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_2),
.Y(n_209)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_3),
.Y(n_70)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_3),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_3),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_118),
.B1(n_121),
.B2(n_122),
.Y(n_117)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_4),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_4),
.A2(n_121),
.B1(n_138),
.B2(n_142),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_4),
.A2(n_121),
.B1(n_213),
.B2(n_304),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_4),
.A2(n_121),
.B1(n_392),
.B2(n_395),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_5),
.A2(n_322),
.B1(n_324),
.B2(n_325),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_5),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_L g426 ( 
.A1(n_5),
.A2(n_325),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_5),
.A2(n_228),
.B1(n_325),
.B2(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_6),
.A2(n_81),
.B1(n_83),
.B2(n_84),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_6),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_83),
.B1(n_162),
.B2(n_165),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_83),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g363 ( 
.A1(n_6),
.A2(n_83),
.B1(n_364),
.B2(n_366),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g100 ( 
.A(n_7),
.Y(n_100)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g152 ( 
.A(n_7),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_7),
.Y(n_256)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_8),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_8),
.Y(n_244)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_8),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_8),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_9),
.A2(n_258),
.B1(n_262),
.B2(n_263),
.Y(n_257)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_9),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_9),
.A2(n_193),
.B1(n_262),
.B2(n_379),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_9),
.A2(n_262),
.B1(n_445),
.B2(n_446),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_9),
.A2(n_262),
.B1(n_516),
.B2(n_517),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_10),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_10),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_10),
.A2(n_91),
.B1(n_188),
.B2(n_192),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g370 ( 
.A1(n_10),
.A2(n_91),
.B1(n_371),
.B2(n_374),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_10),
.A2(n_91),
.B1(n_362),
.B2(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_11),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_11),
.Y(n_360)
);

BUFx8_ASAP7_75t_L g394 ( 
.A(n_11),
.Y(n_394)
);

BUFx5_ASAP7_75t_L g518 ( 
.A(n_11),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_12),
.A2(n_109),
.B1(n_111),
.B2(n_112),
.Y(n_108)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_12),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_12),
.A2(n_111),
.B1(n_122),
.B2(n_279),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_12),
.A2(n_111),
.B1(n_220),
.B2(n_402),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g482 ( 
.A1(n_12),
.A2(n_111),
.B1(n_483),
.B2(n_485),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_13),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_13),
.Y(n_345)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_13),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_14),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_15),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_16),
.Y(n_95)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_17),
.B(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_17),
.B(n_151),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_17),
.B(n_79),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_17),
.A2(n_44),
.B1(n_213),
.B2(n_217),
.Y(n_212)
);

OAI32xp33_ASAP7_75t_L g231 ( 
.A1(n_17),
.A2(n_232),
.A3(n_236),
.B1(n_240),
.B2(n_245),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_17),
.B(n_288),
.Y(n_287)
);

OAI32xp33_ASAP7_75t_L g326 ( 
.A1(n_17),
.A2(n_327),
.A3(n_331),
.B1(n_336),
.B2(n_339),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_L g357 ( 
.A1(n_17),
.A2(n_44),
.B1(n_358),
.B2(n_361),
.Y(n_357)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_493),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_456),
.B(n_490),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_381),
.B(n_453),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

OAI21x1_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_309),
.B(n_380),
.Y(n_24)
);

AOI21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_268),
.B(n_308),
.Y(n_25)
);

OAI21x1_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_180),
.B(n_267),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_133),
.B(n_179),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_87),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_29),
.B(n_87),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_53),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_30),
.A2(n_53),
.B1(n_54),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_30),
.Y(n_154)
);

OAI32xp33_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.A3(n_39),
.B1(n_43),
.B2(n_47),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AO22x2_ASAP7_75t_L g128 ( 
.A1(n_33),
.A2(n_82),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_37),
.Y(n_145)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI21xp33_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_44),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_44),
.A2(n_96),
.B1(n_158),
.B2(n_161),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_44),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_44),
.B(n_337),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_46),
.Y(n_71)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_46),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_46),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_50),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_79),
.B2(n_80),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_60),
.A2(n_79),
.B1(n_80),
.B2(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_60),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_60),
.A2(n_276),
.B(n_277),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_60),
.B(n_378),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_72),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_67),
.B2(n_71),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g184 ( 
.A1(n_72),
.A2(n_185),
.B1(n_186),
.B2(n_187),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_72),
.B(n_278),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_72),
.A2(n_185),
.B1(n_425),
.B2(n_426),
.Y(n_424)
);

OA22x2_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_78),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_73),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_76),
.Y(n_171)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_77),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_79),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_79),
.B(n_412),
.Y(n_411)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_86),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g428 ( 
.A(n_86),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_115),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_88),
.B(n_116),
.C(n_127),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_96),
.B(n_101),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_94),
.Y(n_299)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_94),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_95),
.Y(n_266)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_96),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_96),
.A2(n_137),
.B1(n_161),
.B2(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_96),
.B(n_257),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_96),
.A2(n_108),
.B(n_149),
.Y(n_462)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_99),
.Y(n_96)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_99),
.A2(n_297),
.B(n_301),
.Y(n_296)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_102),
.B(n_301),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_105),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_105),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_107),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_108),
.Y(n_252)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_127),
.Y(n_115)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_117),
.Y(n_186)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_126),
.Y(n_191)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_126),
.Y(n_239)
);

OR2x2_ASAP7_75t_L g196 ( 
.A(n_128),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_128),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_128),
.B(n_444),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_128),
.A2(n_398),
.B1(n_503),
.B2(n_504),
.Y(n_502)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_132),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_155),
.B(n_178),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_153),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g178 ( 
.A(n_135),
.B(n_153),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_146),
.A2(n_252),
.B(n_253),
.Y(n_251)
);

OAI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_146),
.A2(n_297),
.B1(n_319),
.B2(n_321),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_146),
.A2(n_253),
.B(n_321),
.Y(n_409)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_172),
.B(n_177),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_168),
.Y(n_156)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_181),
.B(n_182),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_230),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_195),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_184),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_185),
.A2(n_278),
.B(n_377),
.Y(n_376)
);

OA21x2_ASAP7_75t_L g464 ( 
.A1(n_185),
.A2(n_377),
.B(n_426),
.Y(n_464)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_187),
.Y(n_276)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g379 ( 
.A(n_190),
.Y(n_379)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_195),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_196),
.A2(n_212),
.B1(n_222),
.B2(n_229),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_196),
.A2(n_222),
.B1(n_229),
.B2(n_303),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_196),
.A2(n_229),
.B1(n_303),
.B2(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_196),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_SL g442 ( 
.A1(n_196),
.A2(n_401),
.B(n_443),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_196),
.A2(n_229),
.B1(n_469),
.B2(n_470),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_201),
.B1(n_205),
.B2(n_210),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_202),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_204),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_204),
.Y(n_475)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_210),
.Y(n_228)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_211),
.Y(n_445)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_216),
.Y(n_338)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

AO22x2_ASAP7_75t_L g288 ( 
.A1(n_225),
.A2(n_289),
.B1(n_291),
.B2(n_294),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g405 ( 
.A(n_226),
.Y(n_405)
);

INVx3_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

NOR2xp67_ASAP7_75t_SL g400 ( 
.A(n_229),
.B(n_401),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_230),
.B(n_270),
.C(n_271),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_251),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_235),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g447 ( 
.A(n_235),
.Y(n_447)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_235),
.Y(n_506)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVx6_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_264),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_269),
.B(n_272),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_283),
.B1(n_284),
.B2(n_307),
.Y(n_272)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

XOR2x1_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_274),
.B(n_275),
.C(n_283),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_277),
.B(n_508),
.Y(n_507)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_302),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_295),
.B2(n_296),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_302),
.C(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

OR2x6_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_349),
.Y(n_348)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_288),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_288),
.A2(n_388),
.B1(n_389),
.B2(n_390),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_288),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_288),
.B(n_515),
.Y(n_514)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_290),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_290),
.Y(n_375)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_293),
.Y(n_294)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_293),
.Y(n_350)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_296),
.Y(n_315)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_311),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_310),
.B(n_311),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_346),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_313),
.A2(n_314),
.B1(n_316),
.B2(n_317),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_314),
.B(n_316),
.C(n_346),
.Y(n_450)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_326),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_326),
.Y(n_406)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx3_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx5_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_334),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_368),
.Y(n_346)
);

MAJx2_ASAP7_75t_L g407 ( 
.A(n_347),
.B(n_369),
.C(n_376),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_348),
.A2(n_357),
.B1(n_363),
.B2(n_367),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_348),
.Y(n_389)
);

OAI22x1_ASAP7_75t_SL g437 ( 
.A1(n_348),
.A2(n_367),
.B1(n_391),
.B2(n_438),
.Y(n_437)
);

OAI21x1_ASAP7_75t_SL g480 ( 
.A1(n_348),
.A2(n_438),
.B(n_481),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_348),
.A2(n_513),
.B(n_514),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_350),
.A2(n_351),
.B1(n_353),
.B2(n_354),
.Y(n_349)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_351),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_351),
.Y(n_365)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_352),
.Y(n_366)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_360),
.Y(n_441)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_363),
.Y(n_388)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_376),
.Y(n_368)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_370),
.Y(n_399)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_449),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_419),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_384),
.B(n_419),
.C(n_455),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_407),
.C(n_408),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_385),
.B(n_452),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_406),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_397),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_387),
.B(n_397),
.C(n_406),
.Y(n_420)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

BUFx12f_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_394),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_394),
.Y(n_485)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_398),
.A2(n_399),
.B(n_400),
.Y(n_397)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx4_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx6_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_408),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_410),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_412),
.Y(n_425)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_420),
.B(n_433),
.C(n_448),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_433),
.B1(n_434),
.B2(n_448),
.Y(n_421)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_422),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_423),
.B(n_424),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_436),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_435),
.B(n_437),
.C(n_442),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_442),
.Y(n_436)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

INVx5_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_444),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_450),
.B(n_451),
.Y(n_455)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_459),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_SL g459 ( 
.A1(n_460),
.A2(n_487),
.B1(n_488),
.B2(n_489),
.Y(n_459)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_460),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_466),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_461),
.Y(n_496)
);

OAI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_461)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_462),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_462),
.A2(n_465),
.B1(n_512),
.B2(n_519),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_462),
.B(n_464),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_487),
.C(n_496),
.Y(n_495)
);

XNOR2x1_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_486),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_480),
.Y(n_467)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_468),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g503 ( 
.A(n_470),
.Y(n_503)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_475),
.Y(n_479)
);

INVx4_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_486),
.C(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_482),
.Y(n_513)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

HB1xp67_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g493 ( 
.A(n_494),
.B(n_523),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_497),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_500),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_501),
.A2(n_510),
.B1(n_521),
.B2(n_522),
.Y(n_500)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

OAI21xp33_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_507),
.B(n_509),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_507),
.Y(n_509)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_510),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_511),
.B(n_520),
.Y(n_510)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

INVx5_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

INVx8_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);


endmodule