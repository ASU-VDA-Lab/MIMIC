module real_jpeg_23669_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_0),
.B(n_47),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_67),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_0),
.B(n_185),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_0),
.B(n_33),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_0),
.B(n_52),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_1),
.B(n_33),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_1),
.B(n_49),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_1),
.B(n_47),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_2),
.B(n_71),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_2),
.B(n_47),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_2),
.B(n_67),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_2),
.B(n_113),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_2),
.B(n_33),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_2),
.B(n_52),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_2),
.B(n_49),
.Y(n_281)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_4),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_4),
.B(n_27),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_4),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_4),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_4),
.B(n_33),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_4),
.B(n_52),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_5),
.B(n_47),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_5),
.B(n_67),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_5),
.B(n_49),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_5),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_5),
.B(n_33),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_5),
.B(n_27),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_9),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_9),
.B(n_27),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_52),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_9),
.B(n_49),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_9),
.B(n_33),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_9),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_9),
.B(n_47),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_9),
.B(n_67),
.Y(n_276)
);

INVx8_ASAP7_75t_SL g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_11),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_11),
.B(n_33),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_11),
.B(n_52),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_11),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_11),
.B(n_49),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_11),
.B(n_47),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_11),
.B(n_67),
.Y(n_297)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_14),
.B(n_71),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_14),
.B(n_49),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_14),
.B(n_47),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_14),
.B(n_52),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_14),
.B(n_33),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_14),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_14),
.B(n_67),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_14),
.B(n_27),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_15),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_47),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_15),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_15),
.B(n_52),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_15),
.B(n_67),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_15),
.B(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_16),
.B(n_52),
.Y(n_83)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_152),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_120),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_78),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_21),
.B(n_78),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_54),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_22),
.B(n_55),
.C(n_72),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_39),
.C(n_45),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_23),
.B(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_24),
.B(n_30),
.C(n_37),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_26),
.B(n_61),
.Y(n_127)
);

CKINVDCx5p33_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_30),
.A2(n_38),
.B1(n_82),
.B2(n_83),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_SL g134 ( 
.A(n_30),
.B(n_80),
.C(n_83),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_31),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_31),
.B(n_62),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_32),
.B(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_35),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_35),
.A2(n_37),
.B1(n_40),
.B2(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_36),
.Y(n_198)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_36),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_40),
.C(n_41),
.Y(n_39)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_39),
.B(n_45),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_40),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_41),
.A2(n_42),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_44),
.B(n_218),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g335 ( 
.A(n_45),
.Y(n_335)
);

FAx1_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.CI(n_51),
.CON(n_45),
.SN(n_45)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_46),
.B(n_48),
.C(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_52),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_66),
.C(n_70),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_56),
.A2(n_57),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_60),
.C(n_63),
.Y(n_57)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_58),
.B(n_63),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_65),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_66),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_66),
.B(n_75),
.C(n_77),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_70),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_77),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_74),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_84),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_79),
.B(n_85),
.C(n_86),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_81),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_82),
.A2(n_83),
.B1(n_129),
.B2(n_130),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_86),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_88),
.CI(n_89),
.CON(n_86),
.SN(n_86)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_87),
.B(n_88),
.C(n_89),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_90),
.B(n_334),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.C(n_108),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_91),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_92),
.B(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_94),
.B(n_100),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_97),
.B(n_292),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_104),
.B(n_108),
.Y(n_330)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.C(n_119),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_109),
.B(n_319),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_116),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_110),
.B(n_116),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_115),
.B(n_306),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_118),
.B(n_119),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_122),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_135),
.B2(n_136),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_131),
.B2(n_132),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_129),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_138),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_147),
.Y(n_142)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_332),
.C(n_333),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_322),
.C(n_323),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_308),
.C(n_309),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_285),
.C(n_286),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_255),
.C(n_256),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_230),
.C(n_231),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_188),
.C(n_200),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_173),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_161),
.B(n_168),
.C(n_173),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_163),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_169),
.B(n_171),
.C(n_172),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_174),
.B(n_180),
.C(n_181),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_199)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_183),
.B(n_187),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_199),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_189),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_192),
.A2(n_193),
.B1(n_199),
.B2(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_226),
.C(n_227),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_215),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_244),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_232),
.B(n_245),
.C(n_254),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_240),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_239),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_235),
.A2(n_236),
.B1(n_237),
.B2(n_238),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_235),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_236),
.B(n_238),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_240),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.CI(n_243),
.CON(n_240),
.SN(n_240)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_254),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_252),
.B2(n_253),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_250),
.B2(n_251),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_248),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_249),
.B(n_251),
.C(n_253),
.Y(n_272)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_252),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_271),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_260),
.B2(n_261),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_259),
.B(n_260),
.C(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_266),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_262),
.B(n_267),
.C(n_270),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_262),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_264),
.CI(n_265),
.CON(n_262),
.SN(n_262)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_264),
.C(n_265),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_272),
.B(n_278),
.C(n_283),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_278),
.B1(n_283),
.B2(n_284),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_274),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B(n_277),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_277),
.B(n_304),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_277),
.B(n_304),
.C(n_305),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_278),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_281),
.C(n_282),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_300),
.B2(n_307),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_301),
.C(n_302),
.Y(n_308)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g288 ( 
.A(n_289),
.B(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_291),
.C(n_293),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_293),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_299),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_298),
.C(n_299),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_297),
.Y(n_298)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_311),
.B1(n_320),
.B2(n_321),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_310),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_311),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_312),
.B(n_314),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_314),
.C(n_320),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_317),
.C(n_318),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_324),
.B(n_326),
.C(n_331),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_329),
.B2(n_331),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);


endmodule