module fake_jpeg_10567_n_36 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_36);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_36;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_6),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

INVx4_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_SL g19 ( 
.A1(n_17),
.A2(n_11),
.B1(n_8),
.B2(n_7),
.Y(n_19)
);

OA22x2_ASAP7_75t_L g22 ( 
.A1(n_19),
.A2(n_10),
.B1(n_8),
.B2(n_17),
.Y(n_22)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_20),
.Y(n_21)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_22),
.B(n_17),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_7),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_15),
.C(n_13),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_24),
.A2(n_22),
.B1(n_14),
.B2(n_18),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_25),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_30),
.A2(n_22),
.B(n_18),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_26),
.B(n_21),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_32),
.C(n_16),
.Y(n_33)
);

AO21x1_ASAP7_75t_L g34 ( 
.A1(n_33),
.A2(n_16),
.B(n_1),
.Y(n_34)
);

A2O1A1O1Ixp25_ASAP7_75t_L g35 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.C(n_2),
.D(n_5),
.Y(n_35)
);

BUFx24_ASAP7_75t_SL g36 ( 
.A(n_35),
.Y(n_36)
);


endmodule