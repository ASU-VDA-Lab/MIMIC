module fake_jpeg_15203_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_SL g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_41),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx4f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_21),
.B1(n_26),
.B2(n_30),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_51),
.A2(n_59),
.B1(n_64),
.B2(n_45),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_23),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_52),
.Y(n_77)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_60),
.Y(n_67)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_24),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_16),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_22),
.Y(n_79)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_62),
.Y(n_81)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

OA22x2_ASAP7_75t_SL g65 ( 
.A1(n_62),
.A2(n_37),
.B1(n_34),
.B2(n_30),
.Y(n_65)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_40),
.B1(n_30),
.B2(n_26),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_68),
.A2(n_69),
.B1(n_86),
.B2(n_50),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_30),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_25),
.Y(n_116)
);

OAI22xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_30),
.B1(n_17),
.B2(n_20),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_84),
.B1(n_22),
.B2(n_29),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_49),
.A2(n_30),
.B1(n_26),
.B2(n_20),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_76),
.B1(n_80),
.B2(n_87),
.Y(n_93)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_90),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_75),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_44),
.A2(n_26),
.B1(n_17),
.B2(n_32),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_79),
.B(n_27),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_55),
.B1(n_63),
.B2(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_59),
.A2(n_33),
.B1(n_18),
.B2(n_23),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_82),
.A2(n_85),
.B1(n_27),
.B2(n_19),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_33),
.B1(n_18),
.B2(n_22),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_64),
.A2(n_33),
.B1(n_23),
.B2(n_28),
.Y(n_85)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_32),
.Y(n_86)
);

OR2x6_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_32),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_44),
.A2(n_16),
.B1(n_29),
.B2(n_24),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_22),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_29),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_46),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_94),
.A2(n_101),
.B1(n_102),
.B2(n_115),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_97),
.A2(n_83),
.B1(n_72),
.B2(n_89),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_65),
.B(n_66),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_99),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_46),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_107),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_67),
.A2(n_48),
.B1(n_57),
.B2(n_47),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_48),
.B1(n_50),
.B2(n_47),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_67),
.B(n_16),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_105),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_28),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_19),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_69),
.B(n_28),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_112),
.Y(n_140)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_19),
.Y(n_113)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_78),
.A2(n_43),
.B1(n_25),
.B2(n_31),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_65),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_103),
.B(n_77),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_91),
.A2(n_87),
.B(n_71),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_119),
.A2(n_121),
.B(n_128),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_68),
.C(n_80),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_122),
.B(n_125),
.C(n_130),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_98),
.A2(n_84),
.B(n_65),
.C(n_71),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_81),
.C(n_73),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_96),
.A2(n_83),
.B1(n_72),
.B2(n_74),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_97),
.B(n_81),
.C(n_31),
.Y(n_130)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_131),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_101),
.B1(n_115),
.B2(n_94),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g136 ( 
.A(n_98),
.B(n_76),
.C(n_83),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_136),
.B(n_98),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_98),
.B(n_0),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_137),
.A2(n_139),
.B(n_121),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_98),
.A2(n_74),
.B(n_31),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g143 ( 
.A(n_92),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_98),
.B(n_31),
.C(n_25),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_146),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_131),
.B(n_95),
.Y(n_147)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_124),
.Y(n_150)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_135),
.A2(n_96),
.B(n_111),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_151),
.A2(n_173),
.B(n_123),
.Y(n_183)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_153),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_154),
.B(n_156),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_134),
.B(n_109),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_158),
.B(n_163),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_141),
.Y(n_159)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_125),
.A2(n_91),
.B1(n_93),
.B2(n_104),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_161),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_141),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_137),
.B1(n_132),
.B2(n_130),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_168),
.A2(n_170),
.B1(n_172),
.B2(n_114),
.Y(n_195)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_118),
.A2(n_93),
.B1(n_108),
.B2(n_112),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_174),
.B1(n_137),
.B2(n_128),
.Y(n_177)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_119),
.Y(n_172)
);

AO22x1_ASAP7_75t_SL g174 ( 
.A1(n_136),
.A2(n_102),
.B1(n_100),
.B2(n_105),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_144),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_175),
.B(n_178),
.C(n_179),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_177),
.A2(n_184),
.B1(n_188),
.B2(n_192),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_139),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_122),
.C(n_140),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_140),
.C(n_134),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_180),
.B(n_187),
.C(n_191),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_158),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_161),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_195),
.B(n_168),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_172),
.A2(n_118),
.B1(n_142),
.B2(n_120),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_165),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_186),
.B(n_162),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_160),
.B(n_95),
.C(n_99),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_149),
.A2(n_110),
.B1(n_107),
.B2(n_106),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_113),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_167),
.A2(n_110),
.B1(n_114),
.B2(n_2),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_169),
.B(n_25),
.C(n_14),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_14),
.C(n_13),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_171),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_201),
.A2(n_148),
.B1(n_151),
.B2(n_164),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_159),
.C(n_163),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_202),
.B(n_219),
.Y(n_226)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_203),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_205),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_173),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_206),
.B(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_146),
.Y(n_207)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_207),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_175),
.B(n_174),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_182),
.A2(n_157),
.B1(n_153),
.B2(n_150),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_209),
.A2(n_210),
.B1(n_217),
.B2(n_220),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_200),
.A2(n_162),
.B1(n_174),
.B2(n_154),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g211 ( 
.A(n_179),
.B(n_156),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_211),
.B(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_194),
.B(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_214),
.A2(n_224),
.B1(n_192),
.B2(n_188),
.Y(n_236)
);

AOI21x1_ASAP7_75t_SL g215 ( 
.A1(n_183),
.A2(n_152),
.B(n_170),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_215),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_199),
.C(n_201),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_152),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_193),
.A2(n_152),
.B1(n_13),
.B2(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_176),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_221),
.B(n_225),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_184),
.A2(n_197),
.B1(n_180),
.B2(n_187),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_222),
.A2(n_223),
.B1(n_2),
.B2(n_3),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_177),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_195),
.A2(n_11),
.B(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_176),
.B(n_0),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_209),
.B(n_198),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_227),
.B(n_230),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_207),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_235),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_236),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_216),
.A2(n_198),
.B1(n_190),
.B2(n_189),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_239),
.B1(n_222),
.B2(n_204),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_215),
.A2(n_190),
.B1(n_189),
.B2(n_181),
.Y(n_239)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_220),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_4),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_1),
.Y(n_242)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_242),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_243),
.A2(n_223),
.B1(n_224),
.B2(n_210),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_221),
.B(n_3),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_244),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_245),
.A2(n_218),
.B1(n_5),
.B2(n_6),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_232),
.A2(n_233),
.B1(n_228),
.B2(n_240),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_246),
.A2(n_259),
.B1(n_244),
.B2(n_245),
.Y(n_268)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_232),
.A2(n_206),
.B1(n_217),
.B2(n_205),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_252),
.Y(n_270)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_253),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_239),
.A2(n_208),
.B(n_204),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_226),
.A2(n_211),
.B(n_213),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_256),
.B(n_237),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g257 ( 
.A1(n_228),
.A2(n_213),
.B(n_5),
.C(n_6),
.Y(n_257)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_257),
.B(n_260),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_234),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_261),
.B(n_264),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_258),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_237),
.C(n_231),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_266),
.C(n_272),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_250),
.A2(n_229),
.B1(n_235),
.B2(n_242),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_238),
.C(n_229),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_243),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_267),
.B(n_268),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_241),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_246),
.B(n_248),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_276),
.Y(n_291)
);

INVx3_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

OAI21x1_ASAP7_75t_L g277 ( 
.A1(n_272),
.A2(n_257),
.B(n_256),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_277),
.B(n_278),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_265),
.A2(n_251),
.B1(n_255),
.B2(n_247),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_271),
.A2(n_259),
.B(n_247),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_252),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_12),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_284),
.B(n_9),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_285),
.B(n_289),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_276),
.A2(n_273),
.B(n_270),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_288),
.A2(n_290),
.B(n_9),
.Y(n_296)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_280),
.B(n_263),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_281),
.A2(n_10),
.B(n_8),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_292),
.B(n_279),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_274),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_294),
.B(n_295),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_280),
.B(n_9),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_298),
.B1(n_9),
.B2(n_10),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_287),
.B(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_300),
.B(n_10),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_301),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_303),
.B(n_293),
.Y(n_304)
);

INVxp33_ASAP7_75t_L g305 ( 
.A(n_304),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_305),
.B(n_289),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_299),
.C(n_10),
.Y(n_307)
);


endmodule