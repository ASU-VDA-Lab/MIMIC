module real_jpeg_25530_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_249;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_262;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_202;
wire n_213;
wire n_244;
wire n_167;
wire n_179;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_283;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_0),
.A2(n_25),
.B1(n_26),
.B2(n_42),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_0),
.A2(n_42),
.B1(n_56),
.B2(n_57),
.Y(n_123)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx8_ASAP7_75t_SL g59 ( 
.A(n_4),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_5),
.A2(n_28),
.B1(n_52),
.B2(n_54),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_28),
.B1(n_56),
.B2(n_57),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_5),
.A2(n_28),
.B1(n_39),
.B2(n_40),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_5),
.A2(n_60),
.B(n_159),
.C(n_160),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_5),
.B(n_55),
.Y(n_174)
);

O2A1O1Ixp33_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_57),
.B(n_72),
.C(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_5),
.B(n_26),
.C(n_37),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_5),
.B(n_124),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_5),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_5),
.B(n_35),
.Y(n_232)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_6),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_7),
.A2(n_53),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_7),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_7),
.A2(n_56),
.B1(n_57),
.B2(n_64),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_64),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_64),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_8),
.A2(n_31),
.B1(n_39),
.B2(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_8),
.A2(n_31),
.B1(n_56),
.B2(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_8),
.A2(n_31),
.B1(n_52),
.B2(n_53),
.Y(n_104)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_11),
.Y(n_163)
);

INVx6_ASAP7_75t_L g228 ( 
.A(n_11),
.Y(n_228)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_SL g13 ( 
.A1(n_14),
.A2(n_273),
.B1(n_286),
.B2(n_287),
.Y(n_13)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_14),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_128),
.B(n_272),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_105),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_16),
.B(n_105),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_80),
.C(n_87),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_17),
.B(n_80),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_47),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_18),
.B(n_48),
.C(n_68),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_33),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_19),
.B(n_33),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_20),
.B(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_23),
.Y(n_20)
);

INVx3_ASAP7_75t_SL g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_22),
.B(n_26),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_22),
.A2(n_24),
.B(n_32),
.Y(n_81)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_24),
.B(n_32),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_25),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_26),
.B(n_226),
.Y(n_225)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_28),
.A2(n_57),
.B(n_59),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g185 ( 
.A1(n_28),
.A2(n_39),
.B(n_73),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_29),
.A2(n_91),
.B(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_29),
.B(n_219),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_30),
.B(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_32),
.A2(n_91),
.B(n_92),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_32),
.B(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_38),
.B(n_43),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_34),
.B(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_34),
.A2(n_84),
.B(n_120),
.Y(n_140)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_35),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_35),
.B(n_46),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_35),
.B(n_189),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_84),
.B(n_85),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_39),
.A2(n_40),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_40),
.B(n_202),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp33_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_43),
.B(n_199),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_46),
.Y(n_43)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_44),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_44),
.B(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_67),
.B2(n_68),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_51),
.B(n_55),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_51),
.B(n_65),
.Y(n_138)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_52),
.Y(n_54)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_53),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_62),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_55),
.B(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_56),
.A2(n_57),
.B1(n_72),
.B2(n_73),
.Y(n_78)
);

INVx3_ASAP7_75t_SL g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_61),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_65),
.B(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_65),
.Y(n_113)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_74),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_69),
.B(n_150),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_69),
.A2(n_76),
.B(n_123),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_70),
.B(n_77),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_78),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_77),
.B(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_71),
.B(n_100),
.Y(n_152)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_75),
.B(n_143),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_79),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_77),
.B(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_86),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_81),
.B(n_83),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_81),
.A2(n_86),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_81),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_81),
.A2(n_86),
.B1(n_184),
.B2(n_244),
.Y(n_243)
);

AOI21xp33_ASAP7_75t_L g283 ( 
.A1(n_81),
.A2(n_109),
.B(n_111),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_85),
.B(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_85),
.B(n_188),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_87),
.B(n_270),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_99),
.C(n_101),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_88),
.A2(n_89),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_96),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_96),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_93),
.B(n_176),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_93),
.B(n_212),
.Y(n_233)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_97),
.B(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_98),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_99),
.A2(n_101),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_99),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_101),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_127),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_116),
.B2(n_117),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_107),
.B(n_117),
.C(n_127),
.Y(n_284)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_113),
.A2(n_114),
.B(n_115),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_122),
.B(n_126),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_122),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B(n_125),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_124),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_125),
.B(n_142),
.Y(n_141)
);

FAx1_ASAP7_75t_L g275 ( 
.A(n_126),
.B(n_276),
.CI(n_283),
.CON(n_275),
.SN(n_275)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_267),
.B(n_271),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_177),
.B(n_253),
.C(n_266),
.Y(n_129)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_165),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_131),
.B(n_165),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_132),
.A2(n_133),
.B1(n_147),
.B2(n_164),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_145),
.B2(n_146),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_134),
.B(n_146),
.C(n_164),
.Y(n_254)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_139),
.C(n_141),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_137),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_138),
.B(n_154),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_140),
.B1(n_141),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_139),
.A2(n_140),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_141),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

INVxp67_ASAP7_75t_SL g151 ( 
.A(n_144),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_157),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_149),
.A2(n_153),
.B1(n_155),
.B2(n_156),
.Y(n_148)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_149),
.B(n_156),
.C(n_157),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_150),
.B(n_152),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_153),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_162),
.Y(n_171)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_163),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_171),
.C(n_172),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_167),
.B1(n_191),
.B2(n_192),
.Y(n_190)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_172),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_174),
.C(n_175),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_173),
.B(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_174),
.B(n_175),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_176),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_178),
.B(n_252),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_193),
.B(n_251),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_190),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_180),
.B(n_190),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.C(n_186),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_181),
.B(n_249),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_183),
.B(n_186),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_184),
.Y(n_244)
);

INVxp33_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_246),
.B(n_250),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_195),
.A2(n_237),
.B(n_245),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_216),
.B(n_236),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_203),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_197),
.B(n_203),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_198),
.B(n_200),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_198),
.A2(n_200),
.B1(n_201),
.B2(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_205),
.B1(n_210),
.B2(n_215),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_206),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_209),
.C(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_210),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_214),
.B(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_217),
.A2(n_223),
.B(n_235),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_218),
.B(n_221),
.Y(n_235)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_219),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_231),
.B(n_234),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

INVx5_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_232),
.B(n_233),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_239),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_241),
.B(n_242),
.C(n_243),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_255),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_255),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_263),
.B2(n_264),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_264),
.C(n_265),
.Y(n_268)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g271 ( 
.A(n_268),
.B(n_269),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_273),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_285),
.Y(n_273)
);

OR2x2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_284),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_284),
.Y(n_285)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_275),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_281),
.B2(n_282),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);


endmodule