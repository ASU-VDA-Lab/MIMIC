module real_aes_7257_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_509, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_509;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_453;
wire n_379;
wire n_374;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_330;
wire n_388;
wire n_395;
wire n_332;
wire n_292;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_174;
wire n_104;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_178;
wire n_409;
wire n_298;
wire n_439;
wire n_506;
wire n_297;
wire n_383;
wire n_310;
wire n_119;
wire n_504;
wire n_455;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_484;
wire n_326;
wire n_492;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_313;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_507;
wire n_270;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_0), .A2(n_71), .B1(n_139), .B2(n_144), .Y(n_138) );
A2O1A1Ixp33_ASAP7_75t_SL g244 ( .A1(n_1), .A2(n_245), .B(n_246), .C(n_250), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_2), .B(n_239), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_3), .B(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_4), .A2(n_233), .B(n_335), .Y(n_334) );
AO21x2_ASAP7_75t_L g291 ( .A1(n_5), .A2(n_206), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g196 ( .A(n_6), .Y(n_196) );
AND2x6_ASAP7_75t_L g231 ( .A(n_6), .B(n_194), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_6), .B(n_497), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g309 ( .A1(n_7), .A2(n_214), .B(n_231), .C(n_310), .Y(n_309) );
AO22x2_ASAP7_75t_L g88 ( .A1(n_8), .A2(n_19), .B1(n_89), .B2(n_90), .Y(n_88) );
INVx1_ASAP7_75t_L g211 ( .A(n_9), .Y(n_211) );
NAND2xp5_ASAP7_75t_SL g298 ( .A(n_10), .B(n_225), .Y(n_298) );
AO22x2_ASAP7_75t_L g92 ( .A1(n_11), .A2(n_21), .B1(n_89), .B2(n_93), .Y(n_92) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_12), .A2(n_176), .B1(n_182), .B2(n_183), .Y(n_175) );
INVx1_ASAP7_75t_L g182 ( .A(n_12), .Y(n_182) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_12), .A2(n_214), .B(n_276), .C(n_281), .Y(n_275) );
A2O1A1Ixp33_ASAP7_75t_L g294 ( .A1(n_13), .A2(n_214), .B(n_281), .C(n_295), .Y(n_294) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_14), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g99 ( .A(n_15), .Y(n_99) );
AOI22xp33_ASAP7_75t_SL g148 ( .A1(n_16), .A2(n_65), .B1(n_149), .B2(n_154), .Y(n_148) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_17), .A2(n_233), .B(n_241), .Y(n_240) );
INVx2_ASAP7_75t_L g216 ( .A(n_18), .Y(n_216) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_20), .A2(n_229), .B(n_260), .C(n_261), .Y(n_259) );
OAI221xp5_ASAP7_75t_L g187 ( .A1(n_21), .A2(n_36), .B1(n_47), .B2(n_188), .C(n_189), .Y(n_187) );
INVxp67_ASAP7_75t_L g190 ( .A(n_21), .Y(n_190) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_22), .A2(n_80), .B1(n_173), .B2(n_174), .Y(n_79) );
INVx1_ASAP7_75t_L g173 ( .A(n_22), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_23), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_24), .B(n_274), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g314 ( .A(n_25), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_26), .Y(n_83) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_27), .B(n_225), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_28), .B(n_233), .Y(n_293) );
A2O1A1Ixp33_ASAP7_75t_L g320 ( .A1(n_29), .A2(n_229), .B(n_260), .C(n_321), .Y(n_320) );
AOI22xp33_ASAP7_75t_L g111 ( .A1(n_30), .A2(n_52), .B1(n_112), .B2(n_118), .Y(n_111) );
INVx1_ASAP7_75t_L g247 ( .A(n_31), .Y(n_247) );
INVx1_ASAP7_75t_L g322 ( .A(n_32), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_33), .B(n_233), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g166 ( .A1(n_34), .A2(n_59), .B1(n_167), .B2(n_171), .Y(n_166) );
CKINVDCx20_ASAP7_75t_R g285 ( .A(n_35), .Y(n_285) );
AO22x2_ASAP7_75t_L g98 ( .A1(n_36), .A2(n_58), .B1(n_89), .B2(n_93), .Y(n_98) );
INVxp67_ASAP7_75t_L g191 ( .A(n_36), .Y(n_191) );
INVx1_ASAP7_75t_L g194 ( .A(n_37), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_38), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_39), .B(n_239), .Y(n_340) );
A2O1A1Ixp33_ASAP7_75t_L g337 ( .A1(n_40), .A2(n_221), .B(n_280), .C(n_338), .Y(n_337) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_41), .Y(n_123) );
INVx1_ASAP7_75t_L g210 ( .A(n_42), .Y(n_210) );
CKINVDCx20_ASAP7_75t_R g188 ( .A(n_43), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g265 ( .A(n_44), .B(n_225), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_45), .B(n_226), .Y(n_311) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_46), .Y(n_110) );
AO22x2_ASAP7_75t_L g96 ( .A1(n_47), .A2(n_67), .B1(n_89), .B2(n_90), .Y(n_96) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_48), .Y(n_242) );
AOI22xp5_ASAP7_75t_SL g493 ( .A1(n_48), .A2(n_80), .B1(n_174), .B2(n_242), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_49), .B(n_264), .Y(n_277) );
A2O1A1Ixp33_ASAP7_75t_L g213 ( .A1(n_50), .A2(n_214), .B(n_219), .C(n_229), .Y(n_213) );
CKINVDCx16_ASAP7_75t_R g336 ( .A(n_51), .Y(n_336) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_53), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g278 ( .A(n_54), .B(n_263), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g176 ( .A1(n_55), .A2(n_177), .B1(n_178), .B2(n_181), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_55), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_56), .Y(n_269) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_57), .A2(n_73), .B1(n_179), .B2(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_57), .Y(n_179) );
INVx2_ASAP7_75t_L g208 ( .A(n_60), .Y(n_208) );
AOI22xp33_ASAP7_75t_SL g159 ( .A1(n_61), .A2(n_64), .B1(n_160), .B2(n_162), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_62), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g312 ( .A(n_63), .B(n_249), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_66), .B(n_233), .Y(n_258) );
INVx1_ASAP7_75t_L g262 ( .A(n_68), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g502 ( .A1(n_69), .A2(n_80), .B1(n_174), .B2(n_503), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g503 ( .A(n_69), .Y(n_503) );
INVxp67_ASAP7_75t_L g339 ( .A(n_70), .Y(n_339) );
INVx1_ASAP7_75t_L g89 ( .A(n_72), .Y(n_89) );
INVx1_ASAP7_75t_L g91 ( .A(n_72), .Y(n_91) );
INVx1_ASAP7_75t_L g180 ( .A(n_73), .Y(n_180) );
INVx1_ASAP7_75t_L g220 ( .A(n_74), .Y(n_220) );
INVx1_ASAP7_75t_L g307 ( .A(n_75), .Y(n_307) );
AND2x2_ASAP7_75t_L g324 ( .A(n_76), .B(n_267), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_184), .B1(n_197), .B2(n_489), .C(n_492), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_175), .Y(n_78) );
INVx1_ASAP7_75t_L g174 ( .A(n_80), .Y(n_174) );
AND2x2_ASAP7_75t_L g80 ( .A(n_81), .B(n_136), .Y(n_80) );
NOR3xp33_ASAP7_75t_L g81 ( .A(n_82), .B(n_104), .C(n_122), .Y(n_81) );
OAI22xp5_ASAP7_75t_L g82 ( .A1(n_83), .A2(n_84), .B1(n_99), .B2(n_100), .Y(n_82) );
BUFx3_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
OR2x2_ASAP7_75t_L g85 ( .A(n_86), .B(n_94), .Y(n_85) );
INVx2_ASAP7_75t_L g170 ( .A(n_86), .Y(n_170) );
OR2x2_ASAP7_75t_L g86 ( .A(n_87), .B(n_92), .Y(n_86) );
AND2x2_ASAP7_75t_L g103 ( .A(n_87), .B(n_92), .Y(n_103) );
AND2x2_ASAP7_75t_L g143 ( .A(n_87), .B(n_116), .Y(n_143) );
INVx2_ASAP7_75t_L g87 ( .A(n_88), .Y(n_87) );
AND2x2_ASAP7_75t_L g107 ( .A(n_88), .B(n_92), .Y(n_107) );
AND2x2_ASAP7_75t_L g117 ( .A(n_88), .B(n_98), .Y(n_117) );
INVx1_ASAP7_75t_L g90 ( .A(n_91), .Y(n_90) );
INVx1_ASAP7_75t_L g93 ( .A(n_91), .Y(n_93) );
INVx2_ASAP7_75t_L g116 ( .A(n_92), .Y(n_116) );
INVx1_ASAP7_75t_L g156 ( .A(n_92), .Y(n_156) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
NAND2x1p5_ASAP7_75t_L g102 ( .A(n_95), .B(n_103), .Y(n_102) );
AND2x4_ASAP7_75t_L g147 ( .A(n_95), .B(n_143), .Y(n_147) );
AND2x2_ASAP7_75t_L g95 ( .A(n_96), .B(n_97), .Y(n_95) );
INVx1_ASAP7_75t_L g109 ( .A(n_96), .Y(n_109) );
INVx1_ASAP7_75t_L g115 ( .A(n_96), .Y(n_115) );
INVx1_ASAP7_75t_L g135 ( .A(n_96), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_96), .B(n_98), .Y(n_157) );
AND2x2_ASAP7_75t_L g108 ( .A(n_97), .B(n_109), .Y(n_108) );
INVx2_ASAP7_75t_L g97 ( .A(n_98), .Y(n_97) );
AND2x2_ASAP7_75t_L g153 ( .A(n_98), .B(n_135), .Y(n_153) );
BUFx3_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
BUFx3_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_L g152 ( .A(n_103), .B(n_153), .Y(n_152) );
AND2x4_ASAP7_75t_L g172 ( .A(n_103), .B(n_108), .Y(n_172) );
OAI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_110), .B(n_111), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
AND2x2_ASAP7_75t_L g142 ( .A(n_108), .B(n_143), .Y(n_142) );
AND2x6_ASAP7_75t_L g169 ( .A(n_108), .B(n_170), .Y(n_169) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
AND2x4_ASAP7_75t_L g113 ( .A(n_114), .B(n_117), .Y(n_113) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
INVx1_ASAP7_75t_L g121 ( .A(n_115), .Y(n_121) );
INVx1_ASAP7_75t_L g127 ( .A(n_116), .Y(n_127) );
AND2x4_ASAP7_75t_L g120 ( .A(n_117), .B(n_121), .Y(n_120) );
NAND2x1p5_ASAP7_75t_L g126 ( .A(n_117), .B(n_127), .Y(n_126) );
BUFx4f_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI22xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_124), .B1(n_128), .B2(n_129), .Y(n_122) );
INVx3_ASAP7_75t_SL g124 ( .A(n_125), .Y(n_124) );
INVx4_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_131), .Y(n_130) );
OR2x6_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
NOR2xp33_ASAP7_75t_L g136 ( .A(n_137), .B(n_158), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_148), .Y(n_137) );
INVx2_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx3_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
AND2x2_ASAP7_75t_L g161 ( .A(n_143), .B(n_153), .Y(n_161) );
AND2x4_ASAP7_75t_L g164 ( .A(n_143), .B(n_165), .Y(n_164) );
INVx4_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx3_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx8_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_SL g154 ( .A(n_155), .Y(n_154) );
OR2x6_ASAP7_75t_L g155 ( .A(n_156), .B(n_157), .Y(n_155) );
INVx1_ASAP7_75t_L g165 ( .A(n_157), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_159), .B(n_166), .Y(n_158) );
BUFx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx4_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx11_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
BUFx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
CKINVDCx20_ASAP7_75t_R g183 ( .A(n_176), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_178), .Y(n_181) );
CKINVDCx16_ASAP7_75t_R g184 ( .A(n_185), .Y(n_184) );
CKINVDCx20_ASAP7_75t_R g185 ( .A(n_186), .Y(n_185) );
AND3x1_ASAP7_75t_SL g186 ( .A(n_187), .B(n_192), .C(n_195), .Y(n_186) );
INVxp67_ASAP7_75t_L g497 ( .A(n_187), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_191), .Y(n_189) );
INVx1_ASAP7_75t_SL g498 ( .A(n_192), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g500 ( .A1(n_192), .A2(n_214), .B(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g507 ( .A(n_192), .Y(n_507) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_193), .B(n_196), .Y(n_501) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
OR2x2_ASAP7_75t_SL g506 ( .A(n_195), .B(n_507), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NAND2x1p5_ASAP7_75t_L g199 ( .A(n_200), .B(n_432), .Y(n_199) );
AND4x1_ASAP7_75t_L g200 ( .A(n_201), .B(n_372), .C(n_387), .D(n_412), .Y(n_200) );
NOR2xp33_ASAP7_75t_SL g201 ( .A(n_202), .B(n_345), .Y(n_201) );
OAI21xp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_253), .B(n_325), .Y(n_202) );
AND2x2_ASAP7_75t_L g375 ( .A(n_203), .B(n_271), .Y(n_375) );
AND2x2_ASAP7_75t_L g388 ( .A(n_203), .B(n_270), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_203), .B(n_254), .Y(n_438) );
INVx1_ASAP7_75t_L g442 ( .A(n_203), .Y(n_442) );
AND2x2_ASAP7_75t_L g203 ( .A(n_204), .B(n_238), .Y(n_203) );
INVx2_ASAP7_75t_L g359 ( .A(n_204), .Y(n_359) );
BUFx2_ASAP7_75t_L g386 ( .A(n_204), .Y(n_386) );
AO21x2_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_212), .B(n_236), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_205), .B(n_237), .Y(n_236) );
INVx3_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_205), .B(n_269), .Y(n_268) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_205), .A2(n_306), .B(n_313), .Y(n_305) );
INVx4_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_206), .A2(n_293), .B(n_294), .Y(n_292) );
HB1xp67_ASAP7_75t_L g333 ( .A(n_206), .Y(n_333) );
BUFx6f_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g315 ( .A(n_207), .Y(n_315) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
AND2x2_ASAP7_75t_SL g267 ( .A(n_208), .B(n_209), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_232), .Y(n_212) );
INVx5_ASAP7_75t_L g243 ( .A(n_214), .Y(n_243) );
AND2x2_ASAP7_75t_L g491 ( .A(n_214), .B(n_281), .Y(n_491) );
AND2x6_ASAP7_75t_L g214 ( .A(n_215), .B(n_217), .Y(n_214) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_215), .Y(n_228) );
BUFx3_ASAP7_75t_L g251 ( .A(n_215), .Y(n_251) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g235 ( .A(n_216), .Y(n_235) );
INVx1_ASAP7_75t_L g301 ( .A(n_216), .Y(n_301) );
INVx1_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
BUFx6f_ASAP7_75t_L g223 ( .A(n_218), .Y(n_223) );
INVx3_ASAP7_75t_L g226 ( .A(n_218), .Y(n_226) );
AND2x2_ASAP7_75t_L g234 ( .A(n_218), .B(n_235), .Y(n_234) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_218), .Y(n_249) );
INVx1_ASAP7_75t_L g297 ( .A(n_218), .Y(n_297) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_224), .C(n_227), .Y(n_219) );
INVx1_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g264 ( .A(n_223), .Y(n_264) );
INVx2_ASAP7_75t_L g245 ( .A(n_225), .Y(n_245) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_225), .B(n_339), .Y(n_338) );
INVx5_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
O2A1O1Ixp33_ASAP7_75t_SL g241 ( .A1(n_230), .A2(n_242), .B(n_243), .C(n_244), .Y(n_241) );
O2A1O1Ixp33_ASAP7_75t_L g335 ( .A1(n_230), .A2(n_243), .B(n_336), .C(n_337), .Y(n_335) );
INVx4_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x4_ASAP7_75t_L g233 ( .A(n_231), .B(n_234), .Y(n_233) );
BUFx3_ASAP7_75t_L g281 ( .A(n_231), .Y(n_281) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_231), .B(n_234), .Y(n_308) );
BUFx2_ASAP7_75t_L g274 ( .A(n_233), .Y(n_274) );
INVx1_ASAP7_75t_L g280 ( .A(n_235), .Y(n_280) );
AND2x2_ASAP7_75t_L g326 ( .A(n_238), .B(n_271), .Y(n_326) );
INVx2_ASAP7_75t_L g342 ( .A(n_238), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_238), .B(n_270), .Y(n_351) );
AND2x2_ASAP7_75t_L g430 ( .A(n_238), .B(n_359), .Y(n_430) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_252), .Y(n_238) );
OAI322xp33_ASAP7_75t_L g492 ( .A1(n_242), .A2(n_493), .A3(n_494), .B1(n_498), .B2(n_499), .C1(n_502), .C2(n_504), .Y(n_492) );
INVx2_ASAP7_75t_L g260 ( .A(n_243), .Y(n_260) );
NOR2xp33_ASAP7_75t_L g246 ( .A(n_247), .B(n_248), .Y(n_246) );
INVx4_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
HB1xp67_ASAP7_75t_L g266 ( .A(n_251), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_254), .B(n_287), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_254), .B(n_357), .Y(n_395) );
INVx1_ASAP7_75t_L g483 ( .A(n_254), .Y(n_483) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_270), .Y(n_254) );
AND2x2_ASAP7_75t_L g341 ( .A(n_255), .B(n_342), .Y(n_341) );
OR2x2_ASAP7_75t_L g355 ( .A(n_255), .B(n_356), .Y(n_355) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_255), .Y(n_384) );
OR2x2_ASAP7_75t_L g416 ( .A(n_255), .B(n_358), .Y(n_416) );
AND2x2_ASAP7_75t_L g424 ( .A(n_255), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g457 ( .A(n_255), .B(n_426), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_255), .B(n_326), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_255), .B(n_386), .Y(n_482) );
AND2x2_ASAP7_75t_L g488 ( .A(n_255), .B(n_375), .Y(n_488) );
INVx5_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
BUFx2_ASAP7_75t_L g348 ( .A(n_256), .Y(n_348) );
AND2x2_ASAP7_75t_L g378 ( .A(n_256), .B(n_358), .Y(n_378) );
AND2x2_ASAP7_75t_L g411 ( .A(n_256), .B(n_371), .Y(n_411) );
AND2x2_ASAP7_75t_L g431 ( .A(n_256), .B(n_271), .Y(n_431) );
AND2x2_ASAP7_75t_L g465 ( .A(n_256), .B(n_331), .Y(n_465) );
OR2x6_ASAP7_75t_L g256 ( .A(n_257), .B(n_268), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_258), .A2(n_259), .B(n_267), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_263), .B(n_265), .C(n_266), .Y(n_261) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_263), .A2(n_266), .B(n_322), .C(n_323), .Y(n_321) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx2_ASAP7_75t_L g283 ( .A(n_267), .Y(n_283) );
INVx1_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g318 ( .A1(n_267), .A2(n_319), .B(n_320), .Y(n_318) );
AND2x4_ASAP7_75t_L g371 ( .A(n_270), .B(n_342), .Y(n_371) );
AND2x2_ASAP7_75t_L g382 ( .A(n_270), .B(n_378), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_270), .B(n_358), .Y(n_421) );
INVx2_ASAP7_75t_L g436 ( .A(n_270), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g459 ( .A(n_270), .B(n_370), .Y(n_459) );
AND2x2_ASAP7_75t_L g478 ( .A(n_270), .B(n_430), .Y(n_478) );
INVx5_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_271), .Y(n_377) );
AND2x2_ASAP7_75t_L g385 ( .A(n_271), .B(n_386), .Y(n_385) );
AND2x4_ASAP7_75t_L g426 ( .A(n_271), .B(n_342), .Y(n_426) );
OR2x6_ASAP7_75t_L g271 ( .A(n_272), .B(n_284), .Y(n_271) );
AOI21xp5_ASAP7_75t_SL g272 ( .A1(n_273), .A2(n_275), .B(n_282), .Y(n_272) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_277), .A2(n_278), .B(n_279), .Y(n_276) );
INVx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
NOR2xp33_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_302), .Y(n_288) );
AND2x2_ASAP7_75t_L g349 ( .A(n_289), .B(n_332), .Y(n_349) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_SL g329 ( .A(n_290), .B(n_305), .Y(n_329) );
OR2x2_ASAP7_75t_L g362 ( .A(n_290), .B(n_332), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_290), .B(n_332), .Y(n_367) );
AND2x2_ASAP7_75t_L g394 ( .A(n_290), .B(n_331), .Y(n_394) );
AND2x2_ASAP7_75t_L g446 ( .A(n_290), .B(n_304), .Y(n_446) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_291), .B(n_316), .Y(n_354) );
AND2x2_ASAP7_75t_L g390 ( .A(n_291), .B(n_305), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_298), .B(n_299), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_299), .A2(n_311), .B(n_312), .Y(n_310) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_302), .B(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
OR2x2_ASAP7_75t_L g380 ( .A(n_303), .B(n_362), .Y(n_380) );
OR2x2_ASAP7_75t_L g303 ( .A(n_304), .B(n_316), .Y(n_303) );
OAI322xp33_ASAP7_75t_L g345 ( .A1(n_304), .A2(n_346), .A3(n_350), .B1(n_352), .B2(n_355), .C1(n_360), .C2(n_368), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_304), .B(n_331), .Y(n_353) );
OR2x2_ASAP7_75t_L g363 ( .A(n_304), .B(n_317), .Y(n_363) );
AND2x2_ASAP7_75t_L g365 ( .A(n_304), .B(n_317), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_304), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_304), .B(n_332), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_304), .B(n_461), .Y(n_460) );
INVx5_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_305), .B(n_349), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_308), .B(n_309), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_316), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g343 ( .A(n_316), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_316), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g405 ( .A(n_316), .B(n_332), .Y(n_405) );
AOI211xp5_ASAP7_75t_SL g433 ( .A1(n_316), .A2(n_434), .B(n_437), .C(n_449), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_316), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g471 ( .A(n_316), .B(n_446), .Y(n_471) );
INVx5_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g399 ( .A(n_317), .B(n_332), .Y(n_399) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_317), .Y(n_408) );
AND2x2_ASAP7_75t_L g448 ( .A(n_317), .B(n_446), .Y(n_448) );
AND2x2_ASAP7_75t_SL g479 ( .A(n_317), .B(n_349), .Y(n_479) );
AND2x2_ASAP7_75t_L g486 ( .A(n_317), .B(n_445), .Y(n_486) );
OR2x6_ASAP7_75t_L g317 ( .A(n_318), .B(n_324), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_341), .B2(n_343), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_326), .B(n_348), .Y(n_396) );
INVx2_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g344 ( .A(n_329), .Y(n_344) );
OR2x2_ASAP7_75t_L g404 ( .A(n_329), .B(n_405), .Y(n_404) );
OAI221xp5_ASAP7_75t_SL g452 ( .A1(n_329), .A2(n_453), .B1(n_455), .B2(n_456), .C(n_458), .Y(n_452) );
INVx2_ASAP7_75t_L g391 ( .A(n_330), .Y(n_391) );
AND2x2_ASAP7_75t_L g364 ( .A(n_331), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g454 ( .A(n_331), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_331), .B(n_446), .Y(n_467) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVxp67_ASAP7_75t_L g409 ( .A(n_332), .Y(n_409) );
AND2x2_ASAP7_75t_L g445 ( .A(n_332), .B(n_446), .Y(n_445) );
OA21x2_ASAP7_75t_L g332 ( .A1(n_333), .A2(n_334), .B(n_340), .Y(n_332) );
AND2x2_ASAP7_75t_L g447 ( .A(n_341), .B(n_386), .Y(n_447) );
AND2x2_ASAP7_75t_L g357 ( .A(n_342), .B(n_358), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_342), .B(n_415), .Y(n_414) );
NOR2xp33_ASAP7_75t_SL g428 ( .A(n_344), .B(n_391), .Y(n_428) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
AND2x2_ASAP7_75t_L g434 ( .A(n_347), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g347 ( .A(n_348), .B(n_349), .Y(n_347) );
OR2x2_ASAP7_75t_L g420 ( .A(n_348), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g485 ( .A(n_348), .B(n_430), .Y(n_485) );
INVx2_ASAP7_75t_L g418 ( .A(n_349), .Y(n_418) );
NAND4xp25_ASAP7_75t_SL g481 ( .A(n_350), .B(n_482), .C(n_483), .D(n_484), .Y(n_481) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_351), .B(n_415), .Y(n_450) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_SL g487 ( .A(n_354), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_SL g449 ( .A1(n_355), .A2(n_418), .B(n_422), .C(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
AND2x2_ASAP7_75t_L g444 ( .A(n_357), .B(n_436), .Y(n_444) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_358), .Y(n_370) );
INVx1_ASAP7_75t_L g425 ( .A(n_358), .Y(n_425) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_359), .Y(n_402) );
AOI211xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_363), .B(n_364), .C(n_366), .Y(n_360) );
AND2x2_ASAP7_75t_L g381 ( .A(n_361), .B(n_365), .Y(n_381) );
OAI322xp33_ASAP7_75t_SL g419 ( .A1(n_361), .A2(n_420), .A3(n_422), .B1(n_423), .B2(n_427), .C1(n_428), .C2(n_429), .Y(n_419) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OR2x2_ASAP7_75t_L g441 ( .A(n_363), .B(n_367), .Y(n_441) );
INVx1_ASAP7_75t_L g422 ( .A(n_365), .Y(n_422) );
INVx1_ASAP7_75t_SL g440 ( .A(n_367), .Y(n_440) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
AOI222xp33_ASAP7_75t_L g372 ( .A1(n_373), .A2(n_379), .B1(n_381), .B2(n_382), .C1(n_383), .C2(n_509), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_374), .B(n_376), .Y(n_373) );
OAI322xp33_ASAP7_75t_L g462 ( .A1(n_374), .A2(n_436), .A3(n_441), .B1(n_463), .B2(n_464), .C1(n_466), .C2(n_467), .Y(n_462) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
AOI221xp5_ASAP7_75t_L g412 ( .A1(n_375), .A2(n_389), .B1(n_413), .B2(n_417), .C(n_419), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_377), .B(n_378), .Y(n_376) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OAI222xp33_ASAP7_75t_L g392 ( .A1(n_380), .A2(n_393), .B1(n_395), .B2(n_396), .C1(n_397), .C2(n_400), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_382), .A2(n_389), .B1(n_459), .B2(n_460), .Y(n_458) );
AND2x2_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
AOI211xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_389), .B(n_392), .C(n_403), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_389), .A2(n_426), .B(n_469), .C(n_472), .Y(n_468) );
AND2x4_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
AND2x2_ASAP7_75t_L g398 ( .A(n_390), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g461 ( .A(n_394), .Y(n_461) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_401), .B(n_426), .Y(n_455) );
BUFx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B(n_410), .Y(n_403) );
OAI221xp5_ASAP7_75t_SL g472 ( .A1(n_404), .A2(n_473), .B1(n_474), .B2(n_475), .C(n_476), .Y(n_472) );
INVxp33_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_408), .B(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_415), .B(n_426), .Y(n_466) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_426), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_430), .B(n_431), .Y(n_429) );
AND2x2_ASAP7_75t_L g477 ( .A(n_430), .B(n_436), .Y(n_477) );
AND4x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_451), .C(n_468), .D(n_480), .Y(n_432) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
OAI221xp5_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_439), .B1(n_441), .B2(n_442), .C(n_443), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_443) );
INVx1_ASAP7_75t_L g473 ( .A(n_444), .Y(n_473) );
INVx1_ASAP7_75t_SL g463 ( .A(n_448), .Y(n_463) );
NOR2xp33_ASAP7_75t_SL g451 ( .A(n_452), .B(n_462), .Y(n_451) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_464), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g476 ( .A1(n_471), .A2(n_477), .B1(n_478), .B2(n_479), .Y(n_476) );
AOI22xp5_ASAP7_75t_L g480 ( .A1(n_481), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_480) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_490), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g494 ( .A(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_496), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_500), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_505), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g505 ( .A(n_506), .Y(n_505) );
endmodule