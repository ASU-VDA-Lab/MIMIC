module fake_jpeg_703_n_217 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_217);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_217;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_184;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_28),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_45),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx12_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_7),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_8),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_14),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_19),
.Y(n_71)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_13),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_70),
.Y(n_76)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_77),
.B(n_83),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_49),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_79),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_55),
.B(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_80),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

INVx13_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_77),
.A2(n_62),
.B1(n_69),
.B2(n_71),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_84),
.A2(n_61),
.B1(n_71),
.B2(n_72),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_75),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_79),
.A2(n_62),
.B1(n_57),
.B2(n_71),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_88),
.A2(n_91),
.B1(n_56),
.B2(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_76),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_56),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_53),
.C(n_60),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_80),
.A2(n_57),
.B1(n_56),
.B2(n_61),
.Y(n_91)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_93),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_99),
.Y(n_116)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_93),
.Y(n_98)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_98),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_86),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_82),
.B1(n_81),
.B2(n_73),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_100),
.A2(n_59),
.B1(n_1),
.B2(n_2),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_108),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_103),
.B(n_104),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_89),
.B(n_58),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_105),
.B(n_97),
.Y(n_129)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_92),
.Y(n_106)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_106),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_107),
.A2(n_84),
.B1(n_64),
.B2(n_66),
.Y(n_114)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_95),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_85),
.B(n_66),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_63),
.B1(n_72),
.B2(n_73),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_74),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_74),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_121),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_105),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_118),
.B(n_125),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_101),
.A2(n_87),
.B(n_83),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_119),
.A2(n_0),
.B(n_3),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_102),
.B(n_68),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_0),
.C(n_1),
.Y(n_137)
);

AND2x6_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_47),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_126),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_106),
.A2(n_64),
.B1(n_65),
.B2(n_59),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_124),
.A2(n_126),
.B1(n_3),
.B2(n_4),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_59),
.B1(n_54),
.B2(n_2),
.Y(n_126)
);

NOR2x1_ASAP7_75t_R g128 ( 
.A(n_108),
.B(n_46),
.Y(n_128)
);

AO21x1_ASAP7_75t_L g156 ( 
.A1(n_128),
.A2(n_135),
.B(n_5),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_131),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_99),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_99),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_134),
.B(n_37),
.Y(n_155)
);

AO21x1_ASAP7_75t_SL g135 ( 
.A1(n_112),
.A2(n_96),
.B(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_138),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_150),
.Y(n_166)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_42),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_139),
.B(n_149),
.C(n_128),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_140),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_142),
.B(n_148),
.Y(n_171)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_144),
.B(n_152),
.Y(n_173)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_145),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_133),
.B(n_4),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_41),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_115),
.Y(n_151)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_114),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_154),
.A2(n_155),
.B(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_5),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_157),
.B(n_6),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_161),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_121),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_170),
.C(n_176),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_153),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_167),
.B(n_172),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_139),
.B(n_32),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_150),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_31),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_146),
.A2(n_30),
.B1(n_27),
.B2(n_24),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_10),
.B(n_11),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_147),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_137),
.B(n_23),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_177),
.B(n_179),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_182),
.Y(n_195)
);

CKINVDCx11_ASAP7_75t_R g182 ( 
.A(n_168),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_146),
.C(n_142),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_188),
.Y(n_192)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_175),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_186),
.B1(n_165),
.B2(n_173),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_164),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_158),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_187),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_163),
.B(n_152),
.C(n_156),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_196),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_171),
.B1(n_162),
.B2(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_197),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_181),
.B(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_198),
.C(n_177),
.Y(n_201)
);

OAI22x1_ASAP7_75t_L g196 ( 
.A1(n_178),
.A2(n_172),
.B1(n_162),
.B2(n_183),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_166),
.B1(n_176),
.B2(n_13),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_185),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_195),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_201),
.Y(n_208)
);

XNOR2x1_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_12),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_203),
.B(n_194),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_192),
.B(n_15),
.C(n_16),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_16),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_206),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_202),
.A2(n_189),
.B1(n_193),
.B2(n_196),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g209 ( 
.A(n_207),
.B(n_202),
.CI(n_18),
.CON(n_209),
.SN(n_209)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_209),
.A2(n_208),
.B1(n_200),
.B2(n_205),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_210),
.B1(n_209),
.B2(n_19),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_212),
.Y(n_213)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_213),
.A2(n_209),
.A3(n_18),
.B1(n_20),
.B2(n_21),
.C1(n_22),
.C2(n_23),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_214),
.A2(n_22),
.B(n_17),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_17),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_20),
.Y(n_217)
);


endmodule