module fake_jpeg_28257_n_305 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_305);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_305;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_303;
wire n_90;
wire n_304;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVxp67_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_4),
.B(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_3),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_33),
.Y(n_51)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_0),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_13),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_22),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_22),
.B1(n_26),
.B2(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

AND2x4_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_33),
.A2(n_29),
.B1(n_26),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_39),
.B1(n_38),
.B2(n_35),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_41),
.A2(n_29),
.B1(n_28),
.B2(n_19),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_53),
.A2(n_55),
.B1(n_17),
.B2(n_19),
.Y(n_65)
);

AOI21xp33_ASAP7_75t_SL g54 ( 
.A1(n_33),
.A2(n_23),
.B(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_18),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_22),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx2_ASAP7_75t_SL g71 ( 
.A(n_57),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_59),
.A2(n_46),
.B1(n_53),
.B2(n_55),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_60),
.B(n_61),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_37),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_35),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_63),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_66),
.B(n_77),
.Y(n_87)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_31),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_68),
.B(n_72),
.Y(n_95)
);

AND2x4_ASAP7_75t_L g69 ( 
.A(n_45),
.B(n_32),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_69),
.B(n_80),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_45),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_75),
.B(n_82),
.Y(n_104)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_54),
.A2(n_45),
.B(n_15),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_45),
.B(n_39),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_50),
.Y(n_94)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_64),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_84),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_70),
.A2(n_45),
.B1(n_57),
.B2(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_86),
.A2(n_89),
.B1(n_96),
.B2(n_83),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_57),
.B1(n_48),
.B2(n_47),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_92),
.B(n_99),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_94),
.B(n_59),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_60),
.A2(n_48),
.B1(n_47),
.B2(n_44),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_71),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_64),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_100),
.A2(n_102),
.B1(n_60),
.B2(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_74),
.B1(n_81),
.B2(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_68),
.B(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_64),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_105),
.B(n_79),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_76),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_80),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_128),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_129),
.B1(n_131),
.B2(n_92),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_117),
.B(n_118),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_69),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_119),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_90),
.C(n_98),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_132),
.C(n_89),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_98),
.A2(n_69),
.B(n_74),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_125),
.B(n_104),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_123),
.B(n_127),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_102),
.B(n_85),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_104),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_86),
.B(n_75),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_61),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_85),
.B(n_87),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_88),
.A2(n_72),
.B1(n_63),
.B2(n_66),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_63),
.B1(n_73),
.B2(n_48),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_88),
.C(n_96),
.Y(n_132)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_134),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_112),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_135),
.B(n_140),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_136),
.B(n_144),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_142),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_150),
.B1(n_153),
.B2(n_159),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_111),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_128),
.B(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_114),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_145),
.B(n_147),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_97),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_97),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_131),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_133),
.Y(n_148)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_99),
.B1(n_105),
.B2(n_82),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_154),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_116),
.A2(n_25),
.B1(n_16),
.B2(n_107),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_109),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_157),
.B(n_108),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_107),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_158),
.A2(n_150),
.B(n_154),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_126),
.A2(n_108),
.B1(n_49),
.B2(n_56),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_121),
.B(n_101),
.C(n_91),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_160),
.B(n_110),
.C(n_58),
.Y(n_169)
);

OAI22x1_ASAP7_75t_SL g161 ( 
.A1(n_139),
.A2(n_132),
.B1(n_125),
.B2(n_123),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_161),
.A2(n_167),
.B1(n_174),
.B2(n_25),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_146),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_162),
.B(n_185),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_SL g198 ( 
.A1(n_163),
.A2(n_178),
.B(n_183),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_125),
.B1(n_118),
.B2(n_122),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_168),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_169),
.B(n_177),
.C(n_181),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_143),
.B(n_16),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_170),
.B(n_172),
.Y(n_210)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_78),
.B1(n_101),
.B2(n_62),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_175),
.B(n_23),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_137),
.A2(n_56),
.B1(n_44),
.B2(n_62),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_49),
.B1(n_17),
.B2(n_16),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_58),
.C(n_79),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_141),
.A2(n_0),
.B(n_1),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_138),
.C(n_141),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_155),
.A2(n_0),
.B(n_1),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_158),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_184),
.B(n_24),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_136),
.B(n_40),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_140),
.B(n_79),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_186),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_142),
.B(n_149),
.C(n_151),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_188),
.B(n_175),
.C(n_169),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_162),
.B(n_149),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_190),
.B(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_187),
.A2(n_135),
.B1(n_145),
.B2(n_157),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_192),
.A2(n_195),
.B1(n_208),
.B2(n_174),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_153),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_156),
.B1(n_134),
.B2(n_49),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_200),
.C(n_202),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_188),
.Y(n_197)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_197),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_181),
.B(n_58),
.C(n_79),
.Y(n_200)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_201),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_18),
.C(n_40),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_20),
.C(n_23),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_204),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_185),
.B(n_167),
.C(n_180),
.Y(n_204)
);

XOR2x2_ASAP7_75t_L g205 ( 
.A(n_184),
.B(n_30),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_205),
.B(n_206),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_171),
.B(n_24),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_20),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_182),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_209),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_166),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_211),
.B(n_212),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_173),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_213),
.A2(n_165),
.B1(n_179),
.B2(n_183),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g214 ( 
.A(n_210),
.B(n_180),
.C(n_178),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_214),
.B(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_216),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_163),
.B(n_173),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_225),
.Y(n_248)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_209),
.Y(n_225)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_205),
.A2(n_179),
.B1(n_23),
.B2(n_21),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_227),
.A2(n_216),
.B1(n_217),
.B2(n_224),
.Y(n_235)
);

NAND3xp33_ASAP7_75t_L g230 ( 
.A(n_191),
.B(n_14),
.C(n_12),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_230),
.A2(n_232),
.B(n_233),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_199),
.Y(n_244)
);

NAND3xp33_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_14),
.C(n_12),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_204),
.B(n_14),
.Y(n_233)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_220),
.A2(n_194),
.B1(n_196),
.B2(n_206),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_243),
.Y(n_251)
);

BUFx4f_ASAP7_75t_SL g237 ( 
.A(n_219),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_237),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_245),
.C(n_247),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_215),
.A2(n_194),
.B1(n_200),
.B2(n_199),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_244),
.B(n_218),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_221),
.B(n_207),
.C(n_203),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_23),
.B1(n_21),
.B2(n_20),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_249),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_20),
.C(n_21),
.Y(n_247)
);

BUFx2_ASAP7_75t_L g249 ( 
.A(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_239),
.B(n_228),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_259),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_238),
.A2(n_229),
.B1(n_218),
.B2(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_254),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_261),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_229),
.C(n_20),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_256),
.B(n_260),
.C(n_245),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_241),
.A2(n_12),
.B1(n_11),
.B2(n_23),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_258),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_2),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_23),
.C(n_21),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_21),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_264),
.B(n_255),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_265),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_277)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_235),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_270),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_247),
.C(n_240),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_267),
.B(n_272),
.C(n_5),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_250),
.A2(n_242),
.B(n_248),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_268),
.A2(n_271),
.B(n_256),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_237),
.C(n_240),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_257),
.A2(n_237),
.B(n_249),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_246),
.C(n_21),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_3),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_273),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_258),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_277),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_276),
.A2(n_10),
.B(n_7),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_266),
.B(n_261),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_264),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_279),
.A2(n_284),
.B(n_263),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_283),
.C(n_272),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_5),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_5),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_286),
.Y(n_293)
);

INVxp33_ASAP7_75t_L g297 ( 
.A(n_287),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_288),
.B(n_289),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_282),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_281),
.B(n_269),
.C(n_7),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_290),
.A2(n_292),
.B(n_283),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_6),
.B(n_7),
.Y(n_291)
);

NAND3xp33_ASAP7_75t_SL g295 ( 
.A(n_291),
.B(n_6),
.C(n_7),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_294),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_298),
.B(n_293),
.C(n_8),
.Y(n_301)
);

AOI31xp33_ASAP7_75t_L g300 ( 
.A1(n_297),
.A2(n_285),
.A3(n_292),
.B(n_9),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_300),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_301),
.Y(n_303)
);

AO21x1_ASAP7_75t_L g304 ( 
.A1(n_303),
.A2(n_299),
.B(n_302),
.Y(n_304)
);

OAI21xp33_ASAP7_75t_L g305 ( 
.A1(n_304),
.A2(n_9),
.B(n_10),
.Y(n_305)
);


endmodule