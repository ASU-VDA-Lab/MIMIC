module fake_jpeg_16639_n_353 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_353);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_353;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_SL g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx13_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_20),
.B(n_15),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_42),
.Y(n_56)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_24),
.Y(n_40)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_22),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_41),
.B(n_45),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_23),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_47),
.B(n_48),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_18),
.A2(n_24),
.B(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_49),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_51),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_41),
.B(n_25),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g81 ( 
.A(n_53),
.B(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_48),
.A2(n_18),
.B1(n_30),
.B2(n_29),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_55),
.A2(n_29),
.B1(n_16),
.B2(n_20),
.Y(n_82)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_60),
.Y(n_85)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_40),
.A2(n_30),
.B1(n_18),
.B2(n_29),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_68),
.A2(n_16),
.B1(n_35),
.B2(n_26),
.Y(n_87)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_74),
.Y(n_84)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_77),
.Y(n_99)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_50),
.Y(n_76)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_76),
.Y(n_114)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

OAI22x1_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_16),
.B1(n_48),
.B2(n_30),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_94),
.B1(n_108),
.B2(n_19),
.Y(n_127)
);

OA22x2_ASAP7_75t_L g79 ( 
.A1(n_71),
.A2(n_51),
.B1(n_44),
.B2(n_38),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_79),
.A2(n_92),
.B1(n_112),
.B2(n_34),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_47),
.C(n_24),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_80),
.B(n_32),
.C(n_34),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_83),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_87),
.B1(n_90),
.B2(n_59),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_42),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_63),
.B(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_95),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_46),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_88),
.B(n_93),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_89),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_16),
.B1(n_25),
.B2(n_35),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_51),
.B1(n_44),
.B2(n_38),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_36),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_64),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_27),
.B1(n_36),
.B2(n_21),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_97),
.A2(n_19),
.B1(n_21),
.B2(n_33),
.Y(n_123)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_100),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_103),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_64),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_74),
.Y(n_105)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_105),
.Y(n_143)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_65),
.Y(n_107)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_0),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_21),
.B1(n_31),
.B2(n_13),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_78),
.B1(n_39),
.B2(n_109),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_73),
.A2(n_27),
.B1(n_31),
.B2(n_21),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_66),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_113),
.B(n_57),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_60),
.B(n_32),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_34),
.B(n_28),
.Y(n_135)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_119),
.Y(n_162)
);

OAI22xp33_ASAP7_75t_L g158 ( 
.A1(n_120),
.A2(n_123),
.B1(n_130),
.B2(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_122),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_88),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_125),
.B(n_133),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_92),
.B1(n_85),
.B2(n_105),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_127),
.A2(n_135),
.B(n_136),
.Y(n_177)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_106),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_94),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_80),
.B(n_32),
.C(n_34),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_136),
.C(n_115),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_94),
.Y(n_133)
);

CKINVDCx14_ASAP7_75t_R g147 ( 
.A(n_134),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_135),
.A2(n_137),
.B(n_108),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_28),
.C(n_17),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_140),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_104),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_104),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_141),
.B(n_145),
.Y(n_167)
);

BUFx12f_ASAP7_75t_L g142 ( 
.A(n_96),
.Y(n_142)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_142),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_148),
.B(n_164),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_149),
.A2(n_17),
.B(n_142),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_83),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_154),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_79),
.B1(n_108),
.B2(n_82),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_153),
.A2(n_166),
.B(n_168),
.Y(n_206)
);

NAND3xp33_ASAP7_75t_SL g154 ( 
.A(n_117),
.B(n_79),
.C(n_81),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_117),
.B(n_79),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_157),
.B(n_159),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_158),
.A2(n_177),
.B1(n_139),
.B2(n_146),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_112),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_110),
.B1(n_107),
.B2(n_114),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_160),
.A2(n_169),
.B1(n_122),
.B2(n_144),
.Y(n_182)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_119),
.Y(n_161)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_161),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_163),
.B(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g164 ( 
.A(n_127),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_132),
.B(n_92),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_133),
.B(n_92),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_130),
.B(n_99),
.Y(n_170)
);

OAI21xp33_ASAP7_75t_L g201 ( 
.A1(n_170),
.A2(n_11),
.B(n_13),
.Y(n_201)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_118),
.B(n_126),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_173),
.B(n_175),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_124),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_118),
.B(n_106),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_98),
.Y(n_190)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_134),
.A2(n_85),
.B1(n_114),
.B2(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_179),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_98),
.Y(n_180)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_182),
.A2(n_183),
.B(n_196),
.Y(n_234)
);

XNOR2x1_ASAP7_75t_SL g183 ( 
.A(n_177),
.B(n_131),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_129),
.B1(n_141),
.B2(n_143),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_184),
.A2(n_192),
.B1(n_197),
.B2(n_214),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_172),
.B(n_121),
.C(n_143),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_185),
.B(n_165),
.Y(n_235)
);

MAJx2_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_116),
.C(n_33),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_187),
.B(n_175),
.Y(n_227)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_190),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_160),
.A2(n_164),
.B1(n_166),
.B2(n_168),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_116),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_199),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_142),
.B(n_139),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_155),
.B(n_167),
.Y(n_199)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_201),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_204),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_155),
.B(n_144),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_162),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_146),
.B1(n_33),
.B2(n_28),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_207),
.A2(n_165),
.B1(n_96),
.B2(n_4),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_148),
.Y(n_220)
);

XNOR2x2_ASAP7_75t_L g209 ( 
.A(n_157),
.B(n_17),
.Y(n_209)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_209),
.A2(n_211),
.B(n_151),
.Y(n_217)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_210),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_170),
.A2(n_142),
.B(n_1),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_213),
.A2(n_0),
.B(n_2),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_169),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_198),
.A2(n_188),
.B1(n_194),
.B2(n_183),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_223),
.B1(n_228),
.B2(n_237),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_217),
.A2(n_239),
.B(n_207),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_200),
.Y(n_218)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_218),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_150),
.Y(n_219)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_219),
.Y(n_257)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_198),
.A2(n_163),
.B1(n_179),
.B2(n_153),
.Y(n_223)
);

BUFx24_ASAP7_75t_SL g224 ( 
.A(n_210),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_233),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_159),
.Y(n_225)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_225),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_191),
.Y(n_226)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_226),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_227),
.B(n_230),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_171),
.B1(n_152),
.B2(n_162),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_174),
.Y(n_229)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_229),
.Y(n_268)
);

OAI32xp33_ASAP7_75t_L g230 ( 
.A1(n_209),
.A2(n_174),
.A3(n_152),
.B1(n_3),
.B2(n_4),
.Y(n_230)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_212),
.C(n_185),
.Y(n_251)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_208),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_209),
.A2(n_96),
.B1(n_2),
.B2(n_4),
.Y(n_237)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_186),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_191),
.B(n_165),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_242),
.B(n_233),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_243),
.A2(n_213),
.B1(n_211),
.B2(n_187),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_244),
.A2(n_5),
.B(n_6),
.Y(n_289)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_252),
.B1(n_259),
.B2(n_264),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_253),
.C(n_258),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_218),
.A2(n_182),
.B1(n_206),
.B2(n_192),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_212),
.C(n_206),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_222),
.B(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_261),
.Y(n_271)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_234),
.B(n_184),
.C(n_196),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_240),
.A2(n_181),
.B1(n_189),
.B2(n_186),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_238),
.B(n_181),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_189),
.C(n_96),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_263),
.C(n_231),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_0),
.C(n_2),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_219),
.B1(n_225),
.B2(n_223),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_266)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_228),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_281),
.C(n_286),
.Y(n_292)
);

NAND2x1_ASAP7_75t_L g273 ( 
.A(n_244),
.B(n_230),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_273),
.B(n_280),
.Y(n_301)
);

XOR2x1_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_237),
.Y(n_275)
);

OAI311xp33_ASAP7_75t_L g306 ( 
.A1(n_275),
.A2(n_266),
.A3(n_263),
.B1(n_9),
.C1(n_10),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_236),
.Y(n_276)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_276),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_259),
.A2(n_215),
.B(n_232),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_278),
.A2(n_279),
.B(n_289),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_256),
.A2(n_241),
.B(n_238),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_221),
.C(n_239),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_243),
.Y(n_281)
);

NOR3xp33_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_221),
.C(n_11),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_289),
.Y(n_297)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_255),
.Y(n_285)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_285),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_251),
.B(n_256),
.C(n_264),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.C(n_247),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_252),
.B(n_231),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_277),
.A2(n_268),
.B1(n_260),
.B2(n_257),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_295),
.B(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx13_ASAP7_75t_L g298 ( 
.A(n_273),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_269),
.B(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_299),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_287),
.A2(n_257),
.B1(n_268),
.B2(n_246),
.Y(n_300)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_300),
.Y(n_320)
);

BUFx12_ASAP7_75t_L g302 ( 
.A(n_275),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_271),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_288),
.B(n_247),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_303),
.B(n_305),
.C(n_286),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_270),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_9),
.Y(n_321)
);

OAI21x1_ASAP7_75t_SL g307 ( 
.A1(n_306),
.A2(n_284),
.B(n_8),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_307),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_302),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_282),
.C(n_281),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_282),
.C(n_272),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_291),
.A2(n_283),
.B1(n_272),
.B2(n_280),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_314),
.B1(n_298),
.B2(n_290),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_248),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_315),
.A2(n_316),
.B(n_321),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_304),
.A2(n_6),
.B(n_8),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_9),
.C(n_10),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_9),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_308),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g339 ( 
.A(n_322),
.B(n_294),
.Y(n_339)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_323),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_317),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_324),
.B(n_325),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_313),
.A2(n_290),
.B1(n_291),
.B2(n_296),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_303),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_330),
.B(n_309),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_328),
.B(n_329),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_315),
.B(n_293),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_326),
.B(n_310),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g345 ( 
.A(n_334),
.B(n_311),
.Y(n_345)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_336),
.Y(n_341)
);

OAI21xp5_ASAP7_75t_SL g338 ( 
.A1(n_327),
.A2(n_331),
.B(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_338),
.B(n_339),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g340 ( 
.A(n_325),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_SL g342 ( 
.A(n_340),
.B(n_323),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_343),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g343 ( 
.A(n_335),
.B(n_332),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_345),
.B(n_312),
.C(n_344),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_346),
.A2(n_347),
.B(n_320),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_341),
.B(n_333),
.C(n_337),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_349),
.A2(n_348),
.B(n_340),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_339),
.B(n_319),
.Y(n_351)
);

AOI31xp67_ASAP7_75t_L g352 ( 
.A1(n_351),
.A2(n_301),
.A3(n_302),
.B(n_10),
.Y(n_352)
);

FAx1_ASAP7_75t_SL g353 ( 
.A(n_352),
.B(n_301),
.CI(n_307),
.CON(n_353),
.SN(n_353)
);


endmodule