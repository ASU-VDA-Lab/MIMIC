module fake_jpeg_11318_n_581 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_581);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_581;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_548;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_8),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_14),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_6),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_0),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_11),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_7),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_58),
.Y(n_161)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_60),
.Y(n_183)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

INVx4_ASAP7_75t_SL g62 ( 
.A(n_20),
.Y(n_62)
);

INVx4_ASAP7_75t_SL g150 ( 
.A(n_62),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_20),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g178 ( 
.A(n_63),
.Y(n_178)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_64),
.Y(n_126)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_65),
.Y(n_187)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_66),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_67),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_47),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_68),
.A2(n_18),
.B1(n_32),
.B2(n_29),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_69),
.Y(n_140)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_72),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_45),
.Y(n_77)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_77),
.Y(n_154)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_7),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_79),
.B(n_106),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

BUFx4f_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_83),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_84),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_87),
.Y(n_193)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_40),
.Y(n_89)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_56),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_90),
.Y(n_166)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_91),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_92),
.Y(n_157)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_93),
.Y(n_172)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_22),
.Y(n_94)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_95),
.Y(n_184)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_40),
.Y(n_96)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_96),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_40),
.Y(n_97)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_97),
.Y(n_177)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_98),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_99),
.B(n_105),
.Y(n_164)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_33),
.Y(n_101)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_101),
.Y(n_159)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_102),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_19),
.B(n_8),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_50),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_48),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g162 ( 
.A(n_104),
.Y(n_162)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_18),
.B(n_13),
.Y(n_106)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_107),
.Y(n_180)
);

INVx5_ASAP7_75t_SL g108 ( 
.A(n_41),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_113),
.Y(n_176)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_109),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_110),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_48),
.Y(n_111)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_111),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_112),
.Y(n_192)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_22),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_23),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_116),
.Y(n_131)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_33),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_115),
.B(n_117),
.Y(n_130)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_21),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_31),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_120),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_21),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_121),
.A2(n_133),
.B1(n_146),
.B2(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_122),
.B(n_123),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_79),
.B(n_50),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_106),
.B(n_17),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_127),
.B(n_144),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_21),
.B1(n_72),
.B2(n_65),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_96),
.A2(n_31),
.B1(n_36),
.B2(n_34),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_136),
.A2(n_170),
.B1(n_35),
.B2(n_51),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_138),
.B(n_128),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_108),
.A2(n_38),
.B1(n_42),
.B2(n_41),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_143),
.A2(n_175),
.B1(n_37),
.B2(n_46),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_17),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_117),
.A2(n_26),
.B1(n_27),
.B2(n_44),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_86),
.B(n_26),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_151),
.B(n_171),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_87),
.A2(n_44),
.B1(n_27),
.B2(n_42),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_89),
.B(n_34),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_168),
.B(n_174),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_58),
.A2(n_77),
.B1(n_67),
.B2(n_73),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_86),
.B(n_49),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_60),
.B(n_49),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_114),
.A2(n_38),
.B1(n_119),
.B2(n_41),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_75),
.B(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_179),
.B(n_181),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_80),
.B(n_39),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_84),
.B(n_54),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_194),
.B(n_0),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_92),
.B(n_39),
.C(n_32),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_39),
.C(n_54),
.Y(n_241)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_161),
.Y(n_197)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_135),
.Y(n_198)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_198),
.Y(n_281)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_148),
.Y(n_199)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_199),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_124),
.B(n_37),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_200),
.B(n_206),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_164),
.A2(n_112),
.B1(n_111),
.B2(n_110),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_202),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g203 ( 
.A(n_150),
.Y(n_203)
);

INVx4_ASAP7_75t_SL g266 ( 
.A(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_176),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_204),
.B(n_225),
.Y(n_294)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g284 ( 
.A(n_205),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_35),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_130),
.B(n_43),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_204),
.C(n_241),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_184),
.Y(n_209)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_209),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_210),
.A2(n_218),
.B1(n_224),
.B2(n_1),
.Y(n_310)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_128),
.Y(n_211)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_211),
.Y(n_288)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_212),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_166),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_213),
.B(n_253),
.Y(n_285)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_180),
.Y(n_214)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_214),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_166),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_215),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_140),
.Y(n_216)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_216),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_176),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_217),
.B(n_227),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_175),
.A2(n_104),
.B1(n_97),
.B2(n_43),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_156),
.B(n_32),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_220),
.B(n_221),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_159),
.B(n_29),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g222 ( 
.A(n_164),
.B(n_131),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_222),
.A2(n_145),
.B(n_126),
.Y(n_297)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_170),
.A2(n_43),
.B1(n_29),
.B2(n_54),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_141),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_185),
.Y(n_226)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_226),
.Y(n_304)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_135),
.Y(n_228)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_228),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_161),
.Y(n_229)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_229),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_231),
.B(n_233),
.Y(n_289)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_162),
.Y(n_232)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_232),
.Y(n_317)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_190),
.Y(n_233)
);

INVx4_ASAP7_75t_L g234 ( 
.A(n_162),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_234),
.B(n_240),
.Y(n_293)
);

BUFx8_ASAP7_75t_L g235 ( 
.A(n_150),
.Y(n_235)
);

INVx5_ASAP7_75t_SL g298 ( 
.A(n_235),
.Y(n_298)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_165),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_236),
.B(n_237),
.Y(n_295)
);

INVx3_ASAP7_75t_SL g237 ( 
.A(n_134),
.Y(n_237)
);

INVxp67_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

AOI21xp33_ASAP7_75t_SL g268 ( 
.A1(n_238),
.A2(n_178),
.B(n_12),
.Y(n_268)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_239),
.Y(n_267)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_192),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_241),
.B(n_248),
.Y(n_319)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_242),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_129),
.B(n_51),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_L g244 ( 
.A1(n_136),
.A2(n_51),
.B1(n_37),
.B2(n_35),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g314 ( 
.A1(n_244),
.A2(n_199),
.B1(n_214),
.B2(n_207),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_245),
.A2(n_246),
.B1(n_247),
.B2(n_249),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_172),
.A2(n_46),
.B1(n_62),
.B2(n_69),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_172),
.A2(n_46),
.B1(n_83),
.B2(n_10),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_183),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_191),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_251),
.A2(n_255),
.B1(n_261),
.B2(n_265),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_158),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_252),
.B(n_257),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_137),
.B(n_15),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_139),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_256),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_189),
.A2(n_46),
.B1(n_15),
.B2(n_12),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_142),
.B(n_0),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_177),
.B(n_1),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_1),
.Y(n_292)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_167),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_260),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_178),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_152),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_261)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_188),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_262),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_152),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_263),
.B(n_178),
.Y(n_305)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_191),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_268),
.B(n_273),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_208),
.B(n_182),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_270),
.B(n_274),
.C(n_279),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_195),
.C(n_187),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_201),
.A2(n_153),
.B1(n_173),
.B2(n_160),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_278),
.A2(n_282),
.B1(n_308),
.B2(n_309),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_200),
.B(n_132),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_201),
.A2(n_157),
.B1(n_187),
.B2(n_195),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_230),
.B(n_157),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_286),
.B(n_292),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_219),
.B(n_256),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_254),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_297),
.A2(n_225),
.B(n_260),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_222),
.B(n_145),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_302),
.B(n_235),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_305),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_250),
.B(n_193),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_306),
.B(n_197),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_231),
.A2(n_134),
.B(n_173),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_307),
.A2(n_228),
.B(n_198),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_202),
.A2(n_160),
.B1(n_154),
.B2(n_153),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_206),
.A2(n_154),
.B1(n_193),
.B2(n_3),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_310),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_224),
.B1(n_226),
.B2(n_248),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_210),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_320),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_298),
.A2(n_209),
.B1(n_242),
.B2(n_232),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_322),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_326),
.Y(n_376)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_324),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_258),
.Y(n_326)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_277),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_327),
.B(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_283),
.Y(n_328)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_328),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g331 ( 
.A(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_331),
.B(n_334),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_332),
.A2(n_335),
.B1(n_364),
.B2(n_310),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_298),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_277),
.B(n_223),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_278),
.A2(n_248),
.B1(n_264),
.B2(n_237),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_336),
.A2(n_339),
.B(n_343),
.Y(n_367)
);

AO22x1_ASAP7_75t_L g338 ( 
.A1(n_315),
.A2(n_234),
.B1(n_212),
.B2(n_236),
.Y(n_338)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_287),
.Y(n_340)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_341),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_290),
.B(n_262),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_342),
.B(n_350),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_289),
.A2(n_203),
.B(n_235),
.Y(n_343)
);

BUFx24_ASAP7_75t_L g344 ( 
.A(n_298),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_291),
.Y(n_345)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_345),
.Y(n_389)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_291),
.Y(n_346)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_346),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_347),
.B(n_302),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_293),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_349),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_275),
.B(n_216),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_284),
.Y(n_351)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_351),
.Y(n_395)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_271),
.Y(n_352)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_352),
.A2(n_356),
.B1(n_358),
.B2(n_359),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_294),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g400 ( 
.A(n_353),
.B(n_357),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_SL g355 ( 
.A1(n_289),
.A2(n_211),
.B(n_265),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_355),
.A2(n_297),
.B(n_307),
.Y(n_378)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_284),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_286),
.B(n_239),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_304),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_304),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_284),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_360),
.B(n_361),
.Y(n_375)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_271),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_272),
.A2(n_229),
.B1(n_249),
.B2(n_251),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_363),
.A2(n_308),
.B1(n_316),
.B2(n_309),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_366),
.A2(n_399),
.B1(n_361),
.B2(n_352),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_388),
.B1(n_396),
.B2(n_398),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g406 ( 
.A(n_370),
.B(n_383),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_273),
.C(n_319),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_371),
.B(n_381),
.C(n_390),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_378),
.A2(n_380),
.B(n_384),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_343),
.A2(n_268),
.B(n_300),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_319),
.C(n_270),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_323),
.B(n_319),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_347),
.A2(n_285),
.B(n_275),
.Y(n_384)
);

FAx1_ASAP7_75t_SL g386 ( 
.A(n_326),
.B(n_296),
.CI(n_279),
.CON(n_386),
.SN(n_386)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_386),
.B(n_345),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_342),
.A2(n_272),
.B1(n_274),
.B2(n_294),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_354),
.B(n_276),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_276),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_334),
.C(n_340),
.Y(n_421)
);

AO22x1_ASAP7_75t_SL g392 ( 
.A1(n_330),
.A2(n_311),
.B1(n_317),
.B2(n_318),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_332),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_292),
.B1(n_299),
.B2(n_316),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_347),
.A2(n_299),
.B1(n_295),
.B2(n_267),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_330),
.A2(n_303),
.B1(n_313),
.B2(n_293),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_350),
.A2(n_295),
.B1(n_303),
.B2(n_311),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_401),
.A2(n_357),
.B1(n_335),
.B2(n_337),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g402 ( 
.A1(n_336),
.A2(n_312),
.B(n_317),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_402),
.A2(n_324),
.B(n_341),
.Y(n_419)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_403),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_404),
.A2(n_408),
.B1(n_415),
.B2(n_418),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_383),
.B(n_337),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_412),
.C(n_416),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_376),
.B(n_348),
.Y(n_407)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_407),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_368),
.A2(n_339),
.B1(n_329),
.B2(n_349),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_372),
.Y(n_409)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_376),
.B(n_346),
.Y(n_410)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_410),
.Y(n_460)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_381),
.B(n_355),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_SL g413 ( 
.A(n_369),
.B(n_397),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_413),
.B(n_417),
.Y(n_443)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_372),
.Y(n_414)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_414),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_377),
.A2(n_385),
.B1(n_388),
.B2(n_378),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_325),
.Y(n_416)
);

CKINVDCx14_ASAP7_75t_R g417 ( 
.A(n_400),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_377),
.A2(n_328),
.B1(n_359),
.B2(n_358),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_419),
.A2(n_429),
.B(n_344),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_421),
.B(n_428),
.C(n_433),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_338),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g424 ( 
.A1(n_385),
.A2(n_333),
.B1(n_363),
.B2(n_360),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_424),
.A2(n_387),
.B1(n_394),
.B2(n_389),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_401),
.B(n_356),
.Y(n_425)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_425),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_374),
.B(n_280),
.Y(n_426)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_398),
.Y(n_427)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_427),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_371),
.B(n_391),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g429 ( 
.A1(n_367),
.A2(n_344),
.B(n_312),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_430),
.A2(n_435),
.B1(n_365),
.B2(n_402),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g431 ( 
.A(n_373),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_431),
.B(n_434),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_373),
.B(n_351),
.Y(n_432)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_432),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_390),
.B(n_280),
.C(n_295),
.Y(n_433)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_379),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_399),
.A2(n_344),
.B1(n_338),
.B2(n_321),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_384),
.B(n_288),
.C(n_301),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_436),
.B(n_367),
.C(n_396),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_418),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_439),
.B(n_449),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_446),
.A2(n_408),
.B1(n_415),
.B2(n_404),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_450),
.C(n_455),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g474 ( 
.A1(n_448),
.A2(n_452),
.B1(n_459),
.B2(n_461),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_432),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_428),
.B(n_386),
.C(n_380),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_411),
.A2(n_382),
.B1(n_392),
.B2(n_394),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_453),
.Y(n_475)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_435),
.Y(n_454)
);

INVxp33_ASAP7_75t_L g485 ( 
.A(n_454),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_386),
.C(n_379),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_406),
.B(n_387),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_456),
.B(n_406),
.Y(n_473)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_458),
.Y(n_472)
);

AOI22xp33_ASAP7_75t_L g459 ( 
.A1(n_424),
.A2(n_382),
.B1(n_393),
.B2(n_392),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_SL g461 ( 
.A1(n_427),
.A2(n_393),
.B1(n_375),
.B2(n_395),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_462),
.B(n_412),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_420),
.B(n_389),
.C(n_395),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_464),
.B(n_436),
.C(n_433),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_407),
.B(n_318),
.Y(n_466)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_466),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_451),
.B(n_410),
.Y(n_468)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_468),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_469),
.A2(n_477),
.B1(n_489),
.B2(n_452),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g503 ( 
.A(n_473),
.B(n_479),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_437),
.A2(n_429),
.B(n_423),
.Y(n_476)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_476),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_454),
.A2(n_403),
.B1(n_423),
.B2(n_425),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_451),
.B(n_434),
.Y(n_480)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_480),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_440),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_481),
.B(n_443),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_482),
.B(n_491),
.C(n_493),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g483 ( 
.A(n_442),
.B(n_416),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_483),
.B(n_484),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_444),
.B(n_421),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_440),
.Y(n_486)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_486),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_442),
.B(n_405),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_488),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_444),
.B(n_419),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_446),
.A2(n_430),
.B1(n_413),
.B2(n_431),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_414),
.Y(n_490)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_490),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_288),
.C(n_321),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_438),
.Y(n_492)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_492),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_455),
.B(n_269),
.C(n_281),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_474),
.Y(n_518)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_496),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_460),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_499),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_480),
.B(n_466),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_488),
.B(n_447),
.C(n_450),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_SL g522 ( 
.A(n_500),
.B(n_504),
.Y(n_522)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_489),
.A2(n_457),
.B1(n_437),
.B2(n_441),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_490),
.B(n_463),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_506),
.B(n_448),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_471),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_508),
.B(n_509),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_456),
.C(n_453),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_487),
.B(n_467),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_512),
.B(n_493),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g513 ( 
.A(n_475),
.B(n_462),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_513),
.A2(n_515),
.B1(n_477),
.B2(n_476),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_469),
.A2(n_445),
.B1(n_463),
.B2(n_441),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_509),
.B(n_473),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_517),
.B(n_503),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_518),
.A2(n_494),
.B1(n_515),
.B2(n_514),
.Y(n_533)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_519),
.Y(n_535)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_520),
.Y(n_540)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_498),
.B(n_482),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g534 ( 
.A(n_523),
.B(n_525),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_498),
.B(n_491),
.C(n_483),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_524),
.B(n_529),
.C(n_503),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_501),
.B(n_470),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_507),
.B(n_479),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_526),
.B(n_531),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_505),
.B(n_511),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_528),
.A2(n_532),
.B(n_506),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_501),
.B(n_470),
.C(n_485),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_507),
.B(n_445),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g532 ( 
.A1(n_513),
.A2(n_485),
.B(n_478),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g555 ( 
.A(n_533),
.B(n_536),
.Y(n_555)
);

FAx1_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_510),
.CI(n_514),
.CON(n_537),
.SN(n_537)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_537),
.B(n_546),
.Y(n_551)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_538),
.Y(n_556)
);

AOI21xp5_ASAP7_75t_L g539 ( 
.A1(n_530),
.A2(n_500),
.B(n_511),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_539),
.B(n_543),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_541),
.B(n_545),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_523),
.B(n_510),
.C(n_502),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_524),
.B(n_502),
.C(n_497),
.Y(n_545)
);

NOR2xp67_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_465),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_534),
.B(n_522),
.C(n_518),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_547),
.B(n_557),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_542),
.A2(n_527),
.B1(n_499),
.B2(n_465),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_549),
.A2(n_535),
.B1(n_540),
.B2(n_537),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_543),
.B(n_519),
.Y(n_552)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_552),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g553 ( 
.A(n_534),
.B(n_526),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_553),
.B(n_554),
.Y(n_565)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_533),
.A2(n_545),
.B(n_537),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_541),
.B(n_531),
.C(n_517),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_558),
.B(n_566),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_548),
.B(n_544),
.C(n_536),
.Y(n_560)
);

AOI21xp5_ASAP7_75t_L g571 ( 
.A1(n_560),
.A2(n_561),
.B(n_562),
.Y(n_571)
);

OAI21xp5_ASAP7_75t_SL g561 ( 
.A1(n_551),
.A2(n_544),
.B(n_495),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g562 ( 
.A1(n_551),
.A2(n_495),
.B(n_472),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_SL g563 ( 
.A1(n_554),
.A2(n_266),
.B(n_281),
.Y(n_563)
);

OAI21xp5_ASAP7_75t_SL g568 ( 
.A1(n_563),
.A2(n_549),
.B(n_266),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_550),
.A2(n_556),
.B(n_547),
.Y(n_566)
);

NAND3xp33_ASAP7_75t_SL g574 ( 
.A(n_568),
.B(n_569),
.C(n_555),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_552),
.Y(n_569)
);

NOR2x1_ASAP7_75t_L g570 ( 
.A(n_564),
.B(n_557),
.Y(n_570)
);

AO21x1_ASAP7_75t_L g573 ( 
.A1(n_570),
.A2(n_565),
.B(n_567),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_565),
.B(n_555),
.C(n_269),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_572),
.B(n_266),
.C(n_3),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g577 ( 
.A1(n_573),
.A2(n_574),
.B(n_567),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_575),
.B(n_2),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_577),
.C(n_571),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g579 ( 
.A1(n_578),
.A2(n_2),
.B(n_4),
.Y(n_579)
);

AOI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_4),
.B(n_6),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_580),
.B(n_4),
.Y(n_581)
);


endmodule