module fake_ariane_297_n_2861 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_197, n_463, n_176, n_34, n_404, n_172, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_416, n_283, n_50, n_187, n_525, n_367, n_598, n_345, n_374, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_339, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_222, n_478, n_510, n_256, n_326, n_227, n_48, n_188, n_323, n_550, n_330, n_400, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_293, n_228, n_325, n_276, n_93, n_427, n_108, n_587, n_497, n_303, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_588, n_136, n_334, n_192, n_488, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_16, n_440, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_565, n_281, n_24, n_7, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_464, n_575, n_546, n_297, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_217, n_452, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_513, n_288, n_179, n_395, n_195, n_606, n_213, n_110, n_304, n_67, n_509, n_583, n_306, n_313, n_92, n_430, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_337, n_437, n_111, n_21, n_274, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_184, n_177, n_477, n_364, n_258, n_425, n_431, n_508, n_118, n_121, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_359, n_155, n_573, n_127, n_531, n_2861);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_197;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_330;
input n_400;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_588;
input n_136;
input n_334;
input n_192;
input n_488;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_16;
input n_440;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_565;
input n_281;
input n_24;
input n_7;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_464;
input n_575;
input n_546;
input n_297;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_217;
input n_452;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_513;
input n_288;
input n_179;
input n_395;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_67;
input n_509;
input n_583;
input n_306;
input n_313;
input n_92;
input n_430;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_425;
input n_431;
input n_508;
input n_118;
input n_121;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;

output n_2861;

wire n_2752;
wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_2484;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_2679;
wire n_1355;
wire n_2131;
wire n_2559;
wire n_2500;
wire n_2509;
wire n_1383;
wire n_2182;
wire n_2135;
wire n_2334;
wire n_2680;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_1713;
wire n_1436;
wire n_2407;
wire n_690;
wire n_2818;
wire n_1109;
wire n_1430;
wire n_2537;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2694;
wire n_2011;
wire n_2729;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_2786;
wire n_1566;
wire n_2837;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_2446;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_2671;
wire n_2790;
wire n_1706;
wire n_2207;
wire n_2461;
wire n_2702;
wire n_2731;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2529;
wire n_2374;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_2646;
wire n_737;
wire n_1298;
wire n_2653;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_2482;
wire n_1682;
wire n_2750;
wire n_1836;
wire n_870;
wire n_2547;
wire n_1453;
wire n_945;
wire n_958;
wire n_2554;
wire n_2248;
wire n_813;
wire n_1985;
wire n_2288;
wire n_2621;
wire n_995;
wire n_2579;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_754;
wire n_665;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_2844;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_738;
wire n_1690;
wire n_2221;
wire n_2807;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_2735;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2634;
wire n_2709;
wire n_625;
wire n_2322;
wire n_2746;
wire n_1107;
wire n_2832;
wire n_1688;
wire n_989;
wire n_645;
wire n_1944;
wire n_2370;
wire n_2233;
wire n_2663;
wire n_1988;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_770;
wire n_1514;
wire n_2539;
wire n_1528;
wire n_901;
wire n_2782;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_2458;
wire n_2779;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_2859;
wire n_2847;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_1636;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_1977;
wire n_693;
wire n_863;
wire n_2650;
wire n_1254;
wire n_929;
wire n_2433;
wire n_1703;
wire n_899;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_2571;
wire n_2427;
wire n_661;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_1917;
wire n_2456;
wire n_2769;
wire n_1924;
wire n_1560;
wire n_1654;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_2575;
wire n_2722;
wire n_1396;
wire n_1230;
wire n_1840;
wire n_2739;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2685;
wire n_2094;
wire n_2512;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_2788;
wire n_1021;
wire n_1443;
wire n_2595;
wire n_1465;
wire n_2686;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_2727;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_1121;
wire n_1416;
wire n_1461;
wire n_2717;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_2527;
wire n_1112;
wire n_1159;
wire n_700;
wire n_772;
wire n_1216;
wire n_2759;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_1675;
wire n_2466;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2800;
wire n_2568;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_2326;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_2806;
wire n_1716;
wire n_1872;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_1108;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_2426;
wire n_652;
wire n_1819;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_2703;
wire n_696;
wire n_1442;
wire n_2620;
wire n_798;
wire n_1833;
wire n_1691;
wire n_916;
wire n_1386;
wire n_2810;
wire n_912;
wire n_1884;
wire n_1555;
wire n_1842;
wire n_2499;
wire n_2549;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_762;
wire n_2791;
wire n_2683;
wire n_804;
wire n_1656;
wire n_1382;
wire n_992;
wire n_966;
wire n_955;
wire n_1182;
wire n_794;
wire n_2855;
wire n_2166;
wire n_2848;
wire n_1692;
wire n_2611;
wire n_1562;
wire n_2748;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_1292;
wire n_1178;
wire n_1972;
wire n_2015;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_2415;
wire n_2693;
wire n_2745;
wire n_2087;
wire n_931;
wire n_669;
wire n_1491;
wire n_2628;
wire n_619;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1787;
wire n_2462;
wire n_1389;
wire n_2155;
wire n_2659;
wire n_615;
wire n_1139;
wire n_2836;
wire n_2439;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_2172;
wire n_2601;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_2167;
wire n_2293;
wire n_2753;
wire n_1340;
wire n_2668;
wire n_1240;
wire n_1087;
wire n_2701;
wire n_2400;
wire n_632;
wire n_650;
wire n_2388;
wire n_2273;
wire n_2712;
wire n_1433;
wire n_1911;
wire n_2567;
wire n_2557;
wire n_2695;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_2598;
wire n_1071;
wire n_2755;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_2795;
wire n_2682;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_2762;
wire n_964;
wire n_1627;
wire n_2220;
wire n_2294;
wire n_2274;
wire n_974;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2829;
wire n_2378;
wire n_2467;
wire n_2768;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_2019;
wire n_698;
wire n_2728;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2507;
wire n_2142;
wire n_1633;
wire n_2625;
wire n_1913;
wire n_2069;
wire n_2495;
wire n_1058;
wire n_2328;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2473;
wire n_2144;
wire n_2511;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_760;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_2681;
wire n_1111;
wire n_970;
wire n_1689;
wire n_2535;
wire n_713;
wire n_1255;
wire n_2632;
wire n_1646;
wire n_2262;
wire n_2565;
wire n_1237;
wire n_927;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_706;
wire n_2120;
wire n_2631;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_2860;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_2697;
wire n_1387;
wire n_1263;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_2312;
wire n_670;
wire n_2677;
wire n_1826;
wire n_2834;
wire n_2483;
wire n_1951;
wire n_2490;
wire n_1032;
wire n_1217;
wire n_2558;
wire n_1496;
wire n_637;
wire n_1592;
wire n_2812;
wire n_2662;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_2655;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_2718;
wire n_720;
wire n_926;
wire n_1943;
wire n_2687;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_2765;
wire n_1163;
wire n_2640;
wire n_2811;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_2531;
wire n_1570;
wire n_2099;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2617;
wire n_2481;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_2476;
wire n_2814;
wire n_2059;
wire n_2437;
wire n_2636;
wire n_1439;
wire n_814;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_2841;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_1609;
wire n_1053;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_1899;
wire n_2195;
wire n_2194;
wire n_1467;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_677;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_2783;
wire n_2599;
wire n_699;
wire n_727;
wire n_2075;
wire n_1726;
wire n_2523;
wire n_1945;
wire n_1015;
wire n_2418;
wire n_2496;
wire n_1377;
wire n_1162;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_2853;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_2802;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2125;
wire n_2716;
wire n_1132;
wire n_1156;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_1823;
wire n_2780;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_2618;
wire n_957;
wire n_1402;
wire n_1242;
wire n_2754;
wire n_2707;
wire n_2774;
wire n_2849;
wire n_1607;
wire n_1489;
wire n_2799;
wire n_1218;
wire n_2756;
wire n_2217;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2763;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_1859;
wire n_2660;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_2732;
wire n_1883;
wire n_2516;
wire n_2776;
wire n_2555;
wire n_1969;
wire n_2708;
wire n_735;
wire n_1005;
wire n_2379;
wire n_1294;
wire n_2661;
wire n_1667;
wire n_888;
wire n_845;
wire n_2300;
wire n_1649;
wire n_2452;
wire n_1677;
wire n_2470;
wire n_1927;
wire n_1297;
wire n_2827;
wire n_1708;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_2526;
wire n_1957;
wire n_1953;
wire n_2643;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_2508;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_2594;
wire n_2266;
wire n_2449;
wire n_890;
wire n_842;
wire n_1898;
wire n_1741;
wire n_745;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1373;
wire n_1081;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_2742;
wire n_769;
wire n_1797;
wire n_2366;
wire n_2493;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_832;
wire n_744;
wire n_1895;
wire n_2821;
wire n_2690;
wire n_2474;
wire n_2623;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_2785;
wire n_2460;
wire n_2840;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2448;
wire n_2211;
wire n_2292;
wire n_2480;
wire n_951;
wire n_2772;
wire n_862;
wire n_1700;
wire n_2637;
wire n_659;
wire n_1332;
wire n_2306;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_2737;
wire n_1867;
wire n_852;
wire n_1394;
wire n_2576;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_2696;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_2468;
wire n_1400;
wire n_2035;
wire n_2614;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_2581;
wire n_1783;
wire n_2494;
wire n_1538;
wire n_2831;
wire n_2457;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_2629;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_2540;
wire n_1605;
wire n_1078;
wire n_2486;
wire n_1897;
wire n_2520;
wire n_2137;
wire n_1161;
wire n_2489;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_2492;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_1406;
wire n_1405;
wire n_2684;
wire n_2726;
wire n_2622;
wire n_2272;
wire n_1757;
wire n_1499;
wire n_1318;
wire n_854;
wire n_2091;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_2691;
wire n_805;
wire n_2032;
wire n_2090;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_1596;
wire n_2348;
wire n_2656;
wire n_1281;
wire n_2364;
wire n_1997;
wire n_2574;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_1733;
wire n_1524;
wire n_1476;
wire n_1856;
wire n_2016;
wire n_2667;
wire n_2723;
wire n_2725;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_2850;
wire n_1874;
wire n_1293;
wire n_961;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_2857;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_2730;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_2720;
wire n_1352;
wire n_2405;
wire n_2815;
wire n_1824;
wire n_643;
wire n_2606;
wire n_2700;
wire n_1492;
wire n_2383;
wire n_2764;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2633;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1776;
wire n_686;
wire n_1154;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2698;
wire n_2320;
wire n_979;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2417;
wire n_2789;
wire n_2525;
wire n_1815;
wire n_2813;
wire n_897;
wire n_2546;
wire n_949;
wire n_2454;
wire n_1493;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_2760;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_2368;
wire n_802;
wire n_1151;
wire n_960;
wire n_2352;
wire n_2502;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_2652;
wire n_1133;
wire n_883;
wire n_1852;
wire n_801;
wire n_1286;
wire n_2612;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2477;
wire n_2279;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2497;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_2001;
wire n_1047;
wire n_2506;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_2610;
wire n_1050;
wire n_2626;
wire n_2158;
wire n_2578;
wire n_2607;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_2605;
wire n_858;
wire n_2804;
wire n_1185;
wire n_2475;
wire n_2796;
wire n_2173;
wire n_2715;
wire n_1035;
wire n_1143;
wire n_2665;
wire n_2070;
wire n_2136;
wire n_2771;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_928;
wire n_1153;
wire n_1103;
wire n_825;
wire n_732;
wire n_2619;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_1291;
wire n_2020;
wire n_748;
wire n_2310;
wire n_1045;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_2711;
wire n_1881;
wire n_2635;
wire n_988;
wire n_914;
wire n_689;
wire n_1116;
wire n_1958;
wire n_2747;
wire n_1511;
wire n_2177;
wire n_2713;
wire n_1422;
wire n_2766;
wire n_1965;
wire n_644;
wire n_1197;
wire n_2820;
wire n_2613;
wire n_1165;
wire n_1641;
wire n_2845;
wire n_1517;
wire n_2036;
wire n_843;
wire n_2647;
wire n_638;
wire n_2003;
wire n_2533;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2777;
wire n_2450;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2431;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_2666;
wire n_1370;
wire n_1603;
wire n_728;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2588;
wire n_2331;
wire n_935;
wire n_2478;
wire n_685;
wire n_911;
wire n_2658;
wire n_623;
wire n_2608;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_1534;
wire n_1948;
wire n_2767;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_2692;
wire n_683;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_2553;
wire n_2645;
wire n_907;
wire n_2749;
wire n_1454;
wire n_2592;
wire n_660;
wire n_2459;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_2566;
wire n_2751;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_673;
wire n_2842;
wire n_2833;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_1695;
wire n_2560;
wire n_1164;
wire n_2313;
wire n_1193;
wire n_1345;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_2609;
wire n_2561;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_2303;
wire n_2669;
wire n_1157;
wire n_1584;
wire n_848;
wire n_1664;
wire n_629;
wire n_1739;
wire n_2642;
wire n_1814;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_2688;
wire n_692;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_2498;
wire n_800;
wire n_2638;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_2803;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_621;
wire n_2648;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_2672;
wire n_1772;
wire n_2444;
wire n_2602;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_875;
wire n_1617;
wire n_2455;
wire n_827;
wire n_2600;
wire n_2231;
wire n_697;
wire n_2828;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2530;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_1785;
wire n_1262;
wire n_792;
wire n_1942;
wire n_2180;
wire n_1579;
wire n_2809;
wire n_2181;
wire n_2014;
wire n_975;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2503;
wire n_2270;
wire n_2443;
wire n_1407;
wire n_2465;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_2586;
wire n_1360;
wire n_973;
wire n_2858;
wire n_972;
wire n_2251;
wire n_2843;
wire n_856;
wire n_2572;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_2487;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_2534;
wire n_2488;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_1721;
wire n_2564;
wire n_2591;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_2550;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_1024;
wire n_830;
wire n_2291;
wire n_2816;
wire n_1980;
wire n_2518;
wire n_987;
wire n_936;
wire n_2510;
wire n_1620;
wire n_2501;
wire n_2542;
wire n_1385;
wire n_1525;
wire n_2793;
wire n_1998;
wire n_2165;
wire n_2675;
wire n_2604;
wire n_1775;
wire n_908;
wire n_788;
wire n_2639;
wire n_1036;
wire n_2169;
wire n_2603;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_2630;
wire n_2794;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_2773;
wire n_2817;
wire n_1926;
wire n_2402;
wire n_1458;
wire n_679;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_2808;
wire n_2453;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_1930;
wire n_765;
wire n_1809;
wire n_2787;
wire n_1843;
wire n_1904;
wire n_2000;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2758;
wire n_2395;
wire n_917;
wire n_1271;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_2770;
wire n_631;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_1261;
wire n_2471;
wire n_702;
wire n_898;
wire n_857;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_2584;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_1813;
wire n_2268;
wire n_1452;
wire n_2835;
wire n_1573;
wire n_2734;
wire n_668;
wire n_2569;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_2583;
wire n_1473;
wire n_835;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2445;
wire n_2733;
wire n_1770;
wire n_701;
wire n_1003;
wire n_2469;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_2522;
wire n_2641;
wire n_2463;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_2580;
wire n_2699;
wire n_1792;
wire n_2062;
wire n_1141;
wire n_1629;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2710;
wire n_2505;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_2397;
wire n_2521;
wire n_1727;
wire n_2740;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_2721;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_2615;
wire n_2775;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_2784;
wire n_2541;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_1152;
wire n_2657;
wire n_2447;
wire n_2034;
wire n_1845;
wire n_2538;
wire n_1934;
wire n_2101;
wire n_2577;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_2552;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_2704;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2856;
wire n_2088;
wire n_1275;
wire n_904;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_2736;
wire n_1039;
wire n_2246;
wire n_1150;
wire n_977;
wire n_2339;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2532;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2472;
wire n_2664;
wire n_2705;
wire n_2056;
wire n_2852;
wire n_1136;
wire n_2515;
wire n_1782;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_2519;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_1393;
wire n_723;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_2846;
wire n_1781;
wire n_709;
wire n_2544;
wire n_809;
wire n_2432;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_2504;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_1223;
wire n_2545;
wire n_1768;
wire n_2513;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2451;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_2587;
wire n_1347;
wire n_2839;
wire n_860;
wire n_1043;
wire n_1923;
wire n_2670;
wire n_1764;
wire n_2674;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_2644;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_2562;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_2673;
wire n_664;
wire n_1591;
wire n_2585;
wire n_1229;
wire n_1683;
wire n_2582;
wire n_2548;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2384;
wire n_2678;
wire n_2179;
wire n_1280;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_768;
wire n_1091;
wire n_2052;
wire n_2485;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_2275;
wire n_2563;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2761;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_1639;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_626;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_2792;
wire n_1634;
wire n_2596;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_937;
wire n_1474;
wire n_2081;
wire n_2536;
wire n_2524;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_2318;
wire n_1827;
wire n_866;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_2819;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_2551;
wire n_1102;
wire n_719;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2798;
wire n_2316;
wire n_2464;
wire n_1010;
wire n_2830;
wire n_882;
wire n_2706;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_2514;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_2573;
wire n_2336;
wire n_1662;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_2654;
wire n_2491;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_2517;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_2259;
wire n_849;
wire n_2095;
wire n_2719;
wire n_2738;
wire n_1820;
wire n_2590;
wire n_2797;
wire n_1251;
wire n_1989;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_2689;
wire n_2778;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_2479;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2824;
wire n_2037;
wire n_1308;
wire n_796;
wire n_2851;
wire n_2823;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx14_ASAP7_75t_R g615 ( 
.A(n_614),
.Y(n_615)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_456),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_443),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_12),
.Y(n_618)
);

INVx1_ASAP7_75t_SL g619 ( 
.A(n_459),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_118),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_252),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_126),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_569),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_110),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_413),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_176),
.Y(n_626)
);

CKINVDCx14_ASAP7_75t_R g627 ( 
.A(n_608),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_461),
.Y(n_628)
);

BUFx6f_ASAP7_75t_L g629 ( 
.A(n_156),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_157),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_388),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_104),
.Y(n_632)
);

CKINVDCx5p33_ASAP7_75t_R g633 ( 
.A(n_97),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_6),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_426),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_237),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_136),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_227),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_597),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_570),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_433),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_590),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_42),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_271),
.Y(n_644)
);

INVx1_ASAP7_75t_SL g645 ( 
.A(n_249),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_182),
.Y(n_646)
);

CKINVDCx20_ASAP7_75t_R g647 ( 
.A(n_272),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_17),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_96),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_236),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_500),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_314),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_445),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_250),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_187),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_213),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_160),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_566),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_313),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_231),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_208),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_477),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_565),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_473),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_564),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_11),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_578),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_602),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_562),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_55),
.Y(n_670)
);

CKINVDCx5p33_ASAP7_75t_R g671 ( 
.A(n_516),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_389),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_106),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_29),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_125),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_66),
.Y(n_676)
);

CKINVDCx20_ASAP7_75t_R g677 ( 
.A(n_239),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_295),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_107),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_391),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_292),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_66),
.Y(n_682)
);

CKINVDCx16_ASAP7_75t_R g683 ( 
.A(n_180),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_490),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_317),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_182),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_52),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_557),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_156),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_329),
.Y(n_690)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_11),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_463),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_311),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_101),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_563),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_296),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_474),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_327),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_370),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_551),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_176),
.Y(n_701)
);

CKINVDCx16_ASAP7_75t_R g702 ( 
.A(n_270),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_5),
.Y(n_703)
);

INVx2_ASAP7_75t_SL g704 ( 
.A(n_212),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_143),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_288),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_228),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_38),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_538),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_250),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_256),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_382),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_547),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_33),
.Y(n_714)
);

BUFx10_ASAP7_75t_L g715 ( 
.A(n_72),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_466),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_175),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_412),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_378),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_475),
.Y(n_720)
);

BUFx2_ASAP7_75t_L g721 ( 
.A(n_45),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_21),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_235),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_15),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_190),
.Y(n_725)
);

CKINVDCx16_ASAP7_75t_R g726 ( 
.A(n_204),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_49),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_310),
.Y(n_728)
);

CKINVDCx16_ASAP7_75t_R g729 ( 
.A(n_92),
.Y(n_729)
);

INVx1_ASAP7_75t_SL g730 ( 
.A(n_613),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_543),
.Y(n_731)
);

BUFx6f_ASAP7_75t_L g732 ( 
.A(n_168),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_588),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_267),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_472),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_65),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_88),
.Y(n_737)
);

INVxp67_ASAP7_75t_L g738 ( 
.A(n_228),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_324),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_505),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_436),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_141),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_355),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_190),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_434),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_315),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_317),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_272),
.Y(n_748)
);

INVx1_ASAP7_75t_SL g749 ( 
.A(n_85),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_506),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_81),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_417),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_586),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_48),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_434),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_436),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_31),
.Y(n_757)
);

INVxp67_ASAP7_75t_L g758 ( 
.A(n_558),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_271),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_559),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_307),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_481),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_321),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_281),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_172),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_26),
.Y(n_766)
);

INVxp33_ASAP7_75t_R g767 ( 
.A(n_335),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_524),
.Y(n_768)
);

CKINVDCx20_ASAP7_75t_R g769 ( 
.A(n_557),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_567),
.Y(n_770)
);

BUFx6f_ASAP7_75t_L g771 ( 
.A(n_536),
.Y(n_771)
);

BUFx6f_ASAP7_75t_L g772 ( 
.A(n_267),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_245),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_345),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_392),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_339),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_41),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_165),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_522),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_208),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_397),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_473),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_457),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_422),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_483),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_506),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_220),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_236),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_65),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_564),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_606),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_232),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_256),
.Y(n_793)
);

CKINVDCx16_ASAP7_75t_R g794 ( 
.A(n_371),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_59),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_155),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_544),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_311),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_398),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_265),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_119),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_309),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_425),
.Y(n_803)
);

CKINVDCx20_ASAP7_75t_R g804 ( 
.A(n_523),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_612),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_257),
.Y(n_806)
);

CKINVDCx16_ASAP7_75t_R g807 ( 
.A(n_394),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_153),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_276),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_375),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_221),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_456),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_411),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_458),
.Y(n_814)
);

CKINVDCx16_ASAP7_75t_R g815 ( 
.A(n_22),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_217),
.Y(n_816)
);

INVx3_ASAP7_75t_L g817 ( 
.A(n_258),
.Y(n_817)
);

BUFx2_ASAP7_75t_L g818 ( 
.A(n_555),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_561),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_483),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_85),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_16),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_274),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_422),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_263),
.Y(n_825)
);

CKINVDCx16_ASAP7_75t_R g826 ( 
.A(n_398),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_449),
.Y(n_827)
);

HB1xp67_ASAP7_75t_L g828 ( 
.A(n_550),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_293),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_531),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_544),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_443),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_22),
.Y(n_833)
);

CKINVDCx16_ASAP7_75t_R g834 ( 
.A(n_30),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_497),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_247),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_44),
.Y(n_837)
);

BUFx3_ASAP7_75t_L g838 ( 
.A(n_146),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_560),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_297),
.Y(n_840)
);

BUFx2_ASAP7_75t_SL g841 ( 
.A(n_293),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_30),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_240),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_556),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_418),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_121),
.Y(n_846)
);

BUFx10_ASAP7_75t_L g847 ( 
.A(n_259),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_532),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_147),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_87),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_611),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_173),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_343),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_472),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_129),
.Y(n_855)
);

BUFx10_ASAP7_75t_L g856 ( 
.A(n_391),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_122),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_351),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_411),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_394),
.Y(n_860)
);

CKINVDCx5p33_ASAP7_75t_R g861 ( 
.A(n_128),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_142),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_576),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_92),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_817),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_623),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_817),
.B(n_1),
.Y(n_867)
);

CKINVDCx16_ASAP7_75t_R g868 ( 
.A(n_622),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_639),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_639),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_640),
.Y(n_872)
);

INVxp67_ASAP7_75t_L g873 ( 
.A(n_721),
.Y(n_873)
);

INVxp33_ASAP7_75t_L g874 ( 
.A(n_617),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_754),
.Y(n_875)
);

CKINVDCx16_ASAP7_75t_R g876 ( 
.A(n_683),
.Y(n_876)
);

INVx2_ASAP7_75t_L g877 ( 
.A(n_629),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_629),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_629),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_629),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_629),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_732),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_732),
.Y(n_883)
);

BUFx3_ASAP7_75t_L g884 ( 
.A(n_623),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_732),
.Y(n_885)
);

INVxp67_ASAP7_75t_SL g886 ( 
.A(n_754),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_732),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_647),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_771),
.Y(n_889)
);

INVxp33_ASAP7_75t_L g890 ( 
.A(n_709),
.Y(n_890)
);

BUFx6f_ASAP7_75t_L g891 ( 
.A(n_771),
.Y(n_891)
);

INVxp33_ASAP7_75t_L g892 ( 
.A(n_828),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_771),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_818),
.Y(n_894)
);

CKINVDCx20_ASAP7_75t_R g895 ( 
.A(n_677),
.Y(n_895)
);

CKINVDCx20_ASAP7_75t_R g896 ( 
.A(n_695),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_771),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_772),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_640),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_733),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_838),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_838),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_772),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_621),
.Y(n_904)
);

INVxp67_ASAP7_75t_SL g905 ( 
.A(n_772),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_772),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_772),
.Y(n_907)
);

INVxp33_ASAP7_75t_L g908 ( 
.A(n_644),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_649),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_791),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_651),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_652),
.Y(n_912)
);

BUFx3_ASAP7_75t_L g913 ( 
.A(n_805),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_642),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_641),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_654),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_657),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_851),
.Y(n_918)
);

INVxp33_ASAP7_75t_L g919 ( 
.A(n_659),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_662),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_863),
.Y(n_921)
);

BUFx5_ASAP7_75t_L g922 ( 
.A(n_665),
.Y(n_922)
);

CKINVDCx20_ASAP7_75t_R g923 ( 
.A(n_701),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_641),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_666),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_670),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_642),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_643),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_643),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_667),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_681),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_685),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_702),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_688),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_694),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_696),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_697),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_726),
.Y(n_938)
);

INVxp67_ASAP7_75t_SL g939 ( 
.A(n_658),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_703),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_769),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_705),
.Y(n_942)
);

INVxp67_ASAP7_75t_SL g943 ( 
.A(n_658),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_841),
.Y(n_944)
);

HB1xp67_ASAP7_75t_L g945 ( 
.A(n_729),
.Y(n_945)
);

BUFx3_ASAP7_75t_L g946 ( 
.A(n_668),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_706),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_711),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_712),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_708),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_708),
.Y(n_951)
);

BUFx2_ASAP7_75t_L g952 ( 
.A(n_775),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_722),
.Y(n_953)
);

CKINVDCx20_ASAP7_75t_R g954 ( 
.A(n_787),
.Y(n_954)
);

INVxp67_ASAP7_75t_L g955 ( 
.A(n_636),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_722),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_794),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_807),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_782),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_782),
.Y(n_960)
);

INVxp67_ASAP7_75t_SL g961 ( 
.A(n_821),
.Y(n_961)
);

INVx2_ASAP7_75t_L g962 ( 
.A(n_821),
.Y(n_962)
);

BUFx3_ASAP7_75t_L g963 ( 
.A(n_753),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_840),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_840),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_843),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_891),
.Y(n_967)
);

INVxp67_ASAP7_75t_L g968 ( 
.A(n_945),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_884),
.B(n_636),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_891),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_952),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_933),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_884),
.B(n_678),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_878),
.Y(n_974)
);

NOR2xp33_ASAP7_75t_L g975 ( 
.A(n_930),
.B(n_615),
.Y(n_975)
);

NOR2xp33_ASAP7_75t_L g976 ( 
.A(n_930),
.B(n_627),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_891),
.Y(n_977)
);

INVx2_ASAP7_75t_SL g978 ( 
.A(n_869),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_878),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_939),
.B(n_715),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_879),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_946),
.B(n_730),
.Y(n_982)
);

INVx4_ASAP7_75t_L g983 ( 
.A(n_866),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_869),
.Y(n_984)
);

INVxp67_ASAP7_75t_L g985 ( 
.A(n_952),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_946),
.B(n_815),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_943),
.B(n_715),
.Y(n_987)
);

INVx3_ASAP7_75t_L g988 ( 
.A(n_891),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_871),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_891),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_963),
.B(n_678),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_871),
.Y(n_992)
);

HB1xp67_ASAP7_75t_L g993 ( 
.A(n_933),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_877),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_963),
.B(n_704),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_872),
.B(n_826),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_879),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_877),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_L g999 ( 
.A(n_872),
.B(n_834),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_961),
.B(n_715),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_880),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_881),
.Y(n_1002)
);

NOR2xp33_ASAP7_75t_L g1003 ( 
.A(n_899),
.B(n_704),
.Y(n_1003)
);

BUFx6f_ASAP7_75t_L g1004 ( 
.A(n_881),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_887),
.Y(n_1005)
);

BUFx8_ASAP7_75t_L g1006 ( 
.A(n_866),
.Y(n_1006)
);

INVx4_ASAP7_75t_L g1007 ( 
.A(n_866),
.Y(n_1007)
);

BUFx3_ASAP7_75t_L g1008 ( 
.A(n_866),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_868),
.B(n_847),
.Y(n_1009)
);

INVx6_ASAP7_75t_L g1010 ( 
.A(n_866),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_870),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_887),
.Y(n_1012)
);

BUFx6f_ASAP7_75t_L g1013 ( 
.A(n_907),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_880),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_907),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_882),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_899),
.B(n_839),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_914),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_886),
.B(n_839),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_905),
.B(n_660),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_906),
.B(n_661),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_865),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_900),
.B(n_843),
.Y(n_1023)
);

INVx3_ASAP7_75t_L g1024 ( 
.A(n_865),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_938),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_900),
.B(n_716),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_914),
.B(n_663),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_927),
.B(n_664),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_922),
.Y(n_1029)
);

INVx3_ASAP7_75t_L g1030 ( 
.A(n_882),
.Y(n_1030)
);

BUFx3_ASAP7_75t_L g1031 ( 
.A(n_875),
.Y(n_1031)
);

INVx4_ASAP7_75t_L g1032 ( 
.A(n_913),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_883),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_974),
.Y(n_1034)
);

AND2x2_ASAP7_75t_L g1035 ( 
.A(n_980),
.B(n_913),
.Y(n_1035)
);

AND2x4_ASAP7_75t_L g1036 ( 
.A(n_1026),
.B(n_921),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_974),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_968),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_980),
.B(n_987),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_979),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_979),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_981),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_981),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_1029),
.B(n_922),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_997),
.Y(n_1045)
);

AND2x2_ASAP7_75t_L g1046 ( 
.A(n_987),
.B(n_921),
.Y(n_1046)
);

BUFx6f_ASAP7_75t_L g1047 ( 
.A(n_994),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_1030),
.Y(n_1048)
);

AND2x2_ASAP7_75t_SL g1049 ( 
.A(n_996),
.B(n_867),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_1030),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_1000),
.B(n_910),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_997),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_1030),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_1001),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_1030),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_1002),
.Y(n_1056)
);

NOR2xp33_ASAP7_75t_L g1057 ( 
.A(n_1027),
.B(n_927),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_1026),
.B(n_910),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1001),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_1014),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1014),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_1002),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_1015),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_994),
.Y(n_1064)
);

HB1xp67_ASAP7_75t_L g1065 ( 
.A(n_971),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1015),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_1024),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1024),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_1024),
.Y(n_1069)
);

INVx3_ASAP7_75t_L g1070 ( 
.A(n_1016),
.Y(n_1070)
);

INVx2_ASAP7_75t_L g1071 ( 
.A(n_1016),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_985),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_1024),
.Y(n_1073)
);

AND2x2_ASAP7_75t_L g1074 ( 
.A(n_1000),
.B(n_918),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1023),
.B(n_918),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1016),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_1016),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_1016),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_1033),
.Y(n_1079)
);

CKINVDCx20_ASAP7_75t_R g1080 ( 
.A(n_984),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1033),
.Y(n_1081)
);

INVx4_ASAP7_75t_L g1082 ( 
.A(n_1029),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_1033),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_1033),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_1033),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_1029),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_999),
.B(n_804),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_967),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_1023),
.B(n_908),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_967),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_970),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_967),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_1032),
.B(n_922),
.Y(n_1093)
);

AND2x2_ASAP7_75t_L g1094 ( 
.A(n_1023),
.B(n_919),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_967),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_988),
.Y(n_1096)
);

INVx3_ASAP7_75t_L g1097 ( 
.A(n_994),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_988),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_1026),
.B(n_901),
.Y(n_1099)
);

NAND3xp33_ASAP7_75t_L g1100 ( 
.A(n_1003),
.B(n_944),
.C(n_885),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_988),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_970),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_977),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_988),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_994),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_994),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_998),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_998),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_998),
.Y(n_1109)
);

BUFx2_ASAP7_75t_L g1110 ( 
.A(n_1025),
.Y(n_1110)
);

NOR2x1_ASAP7_75t_L g1111 ( 
.A(n_982),
.B(n_904),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1023),
.B(n_874),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_977),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_998),
.Y(n_1114)
);

OR2x6_ASAP7_75t_L g1115 ( 
.A(n_972),
.B(n_924),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_998),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1004),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1011),
.B(n_890),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1004),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1004),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1032),
.B(n_922),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1004),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1038),
.B(n_876),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_1056),
.Y(n_1124)
);

CKINVDCx6p67_ASAP7_75t_R g1125 ( 
.A(n_1080),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_1056),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1034),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_1110),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_SL g1129 ( 
.A(n_1049),
.B(n_978),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_1056),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1038),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_1063),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_1063),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1057),
.B(n_984),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1063),
.Y(n_1135)
);

NAND2xp33_ASAP7_75t_SL g1136 ( 
.A(n_1039),
.B(n_978),
.Y(n_1136)
);

INVx3_ASAP7_75t_L g1137 ( 
.A(n_1070),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1034),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_1066),
.Y(n_1139)
);

INVx2_ASAP7_75t_L g1140 ( 
.A(n_1066),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_1049),
.Y(n_1141)
);

INVx2_ASAP7_75t_SL g1142 ( 
.A(n_1118),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1066),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_1048),
.Y(n_1144)
);

NOR2x1p5_ASAP7_75t_L g1145 ( 
.A(n_1039),
.B(n_972),
.Y(n_1145)
);

INVx3_ASAP7_75t_L g1146 ( 
.A(n_1070),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_1049),
.B(n_992),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_1072),
.B(n_989),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1048),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1051),
.B(n_1017),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1048),
.Y(n_1151)
);

NOR2xp33_ASAP7_75t_L g1152 ( 
.A(n_1072),
.B(n_989),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1050),
.Y(n_1153)
);

HB1xp67_ASAP7_75t_L g1154 ( 
.A(n_1065),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1037),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1050),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_1087),
.B(n_992),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1050),
.Y(n_1158)
);

INVx8_ASAP7_75t_L g1159 ( 
.A(n_1115),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1087),
.B(n_1018),
.Y(n_1160)
);

INVx3_ASAP7_75t_L g1161 ( 
.A(n_1070),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1110),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1053),
.Y(n_1163)
);

AOI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1093),
.A2(n_995),
.B(n_991),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1037),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1053),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1053),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1055),
.Y(n_1168)
);

AND2x6_ASAP7_75t_L g1169 ( 
.A(n_1051),
.B(n_969),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1074),
.B(n_975),
.Y(n_1170)
);

AOI22xp5_ASAP7_75t_L g1171 ( 
.A1(n_1074),
.A2(n_836),
.B1(n_1018),
.B2(n_986),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1040),
.Y(n_1172)
);

NOR2xp33_ASAP7_75t_L g1173 ( 
.A(n_1065),
.B(n_1025),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_1055),
.Y(n_1174)
);

BUFx6f_ASAP7_75t_L g1175 ( 
.A(n_1047),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_1047),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1112),
.B(n_993),
.Y(n_1177)
);

OAI21xp33_ASAP7_75t_SL g1178 ( 
.A1(n_1040),
.A2(n_1019),
.B(n_1028),
.Y(n_1178)
);

INVx8_ASAP7_75t_L g1179 ( 
.A(n_1115),
.Y(n_1179)
);

NAND3xp33_ASAP7_75t_L g1180 ( 
.A(n_1100),
.B(n_1007),
.C(n_983),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1041),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1055),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1070),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1035),
.B(n_976),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_1062),
.Y(n_1185)
);

INVxp67_ASAP7_75t_SL g1186 ( 
.A(n_1086),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1041),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_1097),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_1036),
.B(n_1032),
.Y(n_1189)
);

OAI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1100),
.A2(n_957),
.B1(n_958),
.B2(n_938),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1062),
.Y(n_1191)
);

AOI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1093),
.A2(n_1021),
.B(n_1020),
.Y(n_1192)
);

NOR2xp33_ASAP7_75t_L g1193 ( 
.A(n_1118),
.B(n_1009),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1035),
.B(n_1032),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_1042),
.Y(n_1195)
);

INVxp67_ASAP7_75t_L g1196 ( 
.A(n_1089),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1042),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1043),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1043),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1045),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1046),
.B(n_1111),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_SL g1202 ( 
.A(n_1036),
.B(n_958),
.Y(n_1202)
);

AND2x2_ASAP7_75t_L g1203 ( 
.A(n_1046),
.B(n_1026),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1089),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1045),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_1036),
.B(n_957),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1111),
.B(n_969),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1058),
.B(n_969),
.Y(n_1208)
);

INVx2_ASAP7_75t_L g1209 ( 
.A(n_1052),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1052),
.Y(n_1210)
);

INVx2_ASAP7_75t_L g1211 ( 
.A(n_1054),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1054),
.Y(n_1212)
);

OAI21xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1059),
.A2(n_718),
.B(n_717),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1059),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1060),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1060),
.Y(n_1216)
);

INVxp33_ASAP7_75t_SL g1217 ( 
.A(n_1112),
.Y(n_1217)
);

OR2x6_ASAP7_75t_L g1218 ( 
.A(n_1115),
.B(n_969),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_SL g1219 ( 
.A(n_1036),
.B(n_973),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1094),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1061),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1061),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1067),
.Y(n_1223)
);

HB1xp67_ASAP7_75t_L g1224 ( 
.A(n_1094),
.Y(n_1224)
);

BUFx6f_ASAP7_75t_SL g1225 ( 
.A(n_1115),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1067),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1068),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1058),
.B(n_973),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1068),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_1069),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1069),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1058),
.B(n_973),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1073),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1073),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1088),
.Y(n_1235)
);

BUFx6f_ASAP7_75t_L g1236 ( 
.A(n_1122),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1088),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1099),
.B(n_888),
.Y(n_1238)
);

INVx2_ASAP7_75t_SL g1239 ( 
.A(n_1075),
.Y(n_1239)
);

AO21x2_ASAP7_75t_L g1240 ( 
.A1(n_1044),
.A2(n_885),
.B(n_883),
.Y(n_1240)
);

INVxp67_ASAP7_75t_SL g1241 ( 
.A(n_1086),
.Y(n_1241)
);

INVx3_ASAP7_75t_L g1242 ( 
.A(n_1097),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1058),
.B(n_973),
.Y(n_1243)
);

NAND3xp33_ASAP7_75t_L g1244 ( 
.A(n_1121),
.B(n_1007),
.C(n_983),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_1091),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1090),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1091),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1091),
.Y(n_1248)
);

INVx2_ASAP7_75t_L g1249 ( 
.A(n_1102),
.Y(n_1249)
);

OAI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1115),
.A2(n_873),
.B1(n_626),
.B2(n_645),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1102),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1102),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1103),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1075),
.B(n_1031),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1099),
.B(n_895),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1090),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1092),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_SL g1258 ( 
.A(n_1099),
.B(n_618),
.Y(n_1258)
);

NOR2xp33_ASAP7_75t_L g1259 ( 
.A(n_1099),
.B(n_896),
.Y(n_1259)
);

BUFx10_ASAP7_75t_L g1260 ( 
.A(n_1115),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_1175),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1195),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1195),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1175),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1197),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1217),
.B(n_1121),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1124),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1124),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1126),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1197),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1126),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1148),
.B(n_892),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1198),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1152),
.B(n_923),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1175),
.Y(n_1275)
);

INVx2_ASAP7_75t_L g1276 ( 
.A(n_1130),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1130),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1198),
.Y(n_1278)
);

NAND2xp33_ASAP7_75t_R g1279 ( 
.A(n_1217),
.B(n_941),
.Y(n_1279)
);

INVxp33_ASAP7_75t_L g1280 ( 
.A(n_1123),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1199),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1125),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1128),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1186),
.A2(n_1044),
.B(n_1241),
.Y(n_1284)
);

INVxp67_ASAP7_75t_SL g1285 ( 
.A(n_1127),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1199),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1205),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1205),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_SL g1289 ( 
.A(n_1141),
.B(n_1082),
.Y(n_1289)
);

AND2x4_ASAP7_75t_L g1290 ( 
.A(n_1145),
.B(n_1011),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1127),
.B(n_1086),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1134),
.B(n_1082),
.Y(n_1292)
);

CKINVDCx20_ASAP7_75t_R g1293 ( 
.A(n_1125),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1131),
.B(n_954),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1132),
.Y(n_1295)
);

XOR2xp5_ASAP7_75t_L g1296 ( 
.A(n_1123),
.B(n_894),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1128),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1209),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1209),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1210),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1210),
.Y(n_1301)
);

OAI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1178),
.A2(n_1086),
.B(n_1092),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1211),
.Y(n_1303)
);

INVx3_ASAP7_75t_R g1304 ( 
.A(n_1177),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1138),
.B(n_1082),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1211),
.Y(n_1306)
);

AND2x6_ASAP7_75t_L g1307 ( 
.A(n_1138),
.B(n_1071),
.Y(n_1307)
);

INVxp67_ASAP7_75t_L g1308 ( 
.A(n_1154),
.Y(n_1308)
);

CKINVDCx20_ASAP7_75t_R g1309 ( 
.A(n_1162),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1162),
.B(n_1031),
.Y(n_1310)
);

XNOR2x2_ASAP7_75t_L g1311 ( 
.A(n_1171),
.B(n_767),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1214),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1173),
.B(n_1177),
.Y(n_1313)
);

CKINVDCx20_ASAP7_75t_R g1314 ( 
.A(n_1171),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1214),
.Y(n_1315)
);

AOI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1164),
.A2(n_1192),
.B(n_1165),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1132),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1155),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1155),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1133),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1165),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1172),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1172),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1220),
.B(n_1224),
.Y(n_1324)
);

XNOR2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1145),
.B(n_618),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1133),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1181),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1181),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1203),
.B(n_955),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1187),
.Y(n_1330)
);

CKINVDCx20_ASAP7_75t_R g1331 ( 
.A(n_1238),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1187),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1200),
.Y(n_1333)
);

INVx4_ASAP7_75t_L g1334 ( 
.A(n_1179),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1200),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1212),
.Y(n_1336)
);

CKINVDCx20_ASAP7_75t_R g1337 ( 
.A(n_1255),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1212),
.Y(n_1338)
);

CKINVDCx20_ASAP7_75t_R g1339 ( 
.A(n_1259),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1215),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1215),
.Y(n_1341)
);

CKINVDCx5p33_ASAP7_75t_R g1342 ( 
.A(n_1142),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_1193),
.Y(n_1343)
);

INVxp33_ASAP7_75t_L g1344 ( 
.A(n_1203),
.Y(n_1344)
);

XOR2xp5_ASAP7_75t_L g1345 ( 
.A(n_1160),
.B(n_902),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1216),
.B(n_1082),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1178),
.A2(n_1222),
.B(n_1221),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1221),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1222),
.Y(n_1349)
);

CKINVDCx14_ASAP7_75t_R g1350 ( 
.A(n_1218),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1235),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1235),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1135),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1239),
.B(n_1097),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_L g1355 ( 
.A(n_1129),
.B(n_1095),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1237),
.Y(n_1356)
);

NOR2xp33_ASAP7_75t_L g1357 ( 
.A(n_1147),
.B(n_1095),
.Y(n_1357)
);

XOR2x2_ASAP7_75t_L g1358 ( 
.A(n_1157),
.B(n_619),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1237),
.Y(n_1359)
);

XOR2xp5_ASAP7_75t_L g1360 ( 
.A(n_1190),
.B(n_620),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1204),
.B(n_1097),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1135),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1246),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1246),
.Y(n_1364)
);

XNOR2xp5_ASAP7_75t_L g1365 ( 
.A(n_1250),
.B(n_909),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1256),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1139),
.Y(n_1367)
);

OAI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1244),
.A2(n_1098),
.B(n_1096),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1256),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1257),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1196),
.B(n_911),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1257),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1142),
.B(n_912),
.Y(n_1373)
);

NOR2xp33_ASAP7_75t_L g1374 ( 
.A(n_1150),
.B(n_1184),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_SL g1375 ( 
.A(n_1141),
.B(n_1047),
.Y(n_1375)
);

BUFx2_ASAP7_75t_R g1376 ( 
.A(n_1202),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1223),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1204),
.B(n_916),
.Y(n_1378)
);

XOR2xp5_ASAP7_75t_L g1379 ( 
.A(n_1206),
.B(n_620),
.Y(n_1379)
);

NAND2xp33_ASAP7_75t_SL g1380 ( 
.A(n_1170),
.B(n_1096),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1239),
.B(n_917),
.Y(n_1381)
);

INVxp33_ASAP7_75t_SL g1382 ( 
.A(n_1194),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1223),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1230),
.Y(n_1384)
);

NOR2xp33_ASAP7_75t_L g1385 ( 
.A(n_1141),
.B(n_1098),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1234),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1201),
.B(n_920),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1219),
.B(n_925),
.Y(n_1388)
);

INVxp67_ASAP7_75t_SL g1389 ( 
.A(n_1175),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1139),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1218),
.B(n_1101),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1140),
.Y(n_1392)
);

AND2x2_ASAP7_75t_L g1393 ( 
.A(n_1218),
.B(n_926),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1226),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1218),
.B(n_931),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1228),
.B(n_932),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1169),
.B(n_1101),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1226),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1227),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1227),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1140),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1229),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_1258),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1229),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_1225),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1143),
.Y(n_1406)
);

INVxp67_ASAP7_75t_SL g1407 ( 
.A(n_1175),
.Y(n_1407)
);

NOR2xp33_ASAP7_75t_L g1408 ( 
.A(n_1254),
.B(n_1207),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_1225),
.Y(n_1409)
);

AND2x2_ASAP7_75t_L g1410 ( 
.A(n_1208),
.B(n_1232),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1231),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1231),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1233),
.Y(n_1413)
);

NOR2xp33_ASAP7_75t_L g1414 ( 
.A(n_1243),
.B(n_1104),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1136),
.B(n_934),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1233),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1185),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1185),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1191),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1191),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1159),
.Y(n_1421)
);

OR2x6_ASAP7_75t_L g1422 ( 
.A(n_1179),
.B(n_924),
.Y(n_1422)
);

XNOR2xp5_ASAP7_75t_L g1423 ( 
.A(n_1189),
.B(n_1180),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1144),
.Y(n_1424)
);

NOR2xp33_ASAP7_75t_L g1425 ( 
.A(n_1137),
.B(n_1104),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1137),
.B(n_1076),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1159),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1144),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1143),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1149),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1149),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1159),
.Y(n_1432)
);

XNOR2xp5_ASAP7_75t_L g1433 ( 
.A(n_1180),
.B(n_935),
.Y(n_1433)
);

NAND2x1p5_ASAP7_75t_L g1434 ( 
.A(n_1176),
.B(n_1084),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1151),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1151),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1153),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1153),
.Y(n_1438)
);

NOR2xp67_ASAP7_75t_L g1439 ( 
.A(n_1213),
.B(n_983),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1169),
.B(n_936),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1156),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1156),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1158),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1158),
.Y(n_1444)
);

CKINVDCx5p33_ASAP7_75t_R g1445 ( 
.A(n_1225),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1163),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1163),
.Y(n_1447)
);

INVx4_ASAP7_75t_SL g1448 ( 
.A(n_1169),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_SL g1449 ( 
.A(n_1179),
.B(n_749),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1166),
.Y(n_1450)
);

AND2x2_ASAP7_75t_L g1451 ( 
.A(n_1169),
.B(n_937),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_SL g1452 ( 
.A(n_1260),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1166),
.Y(n_1453)
);

OR2x2_ASAP7_75t_SL g1454 ( 
.A(n_1159),
.B(n_940),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1167),
.Y(n_1455)
);

NAND2xp33_ASAP7_75t_R g1456 ( 
.A(n_1188),
.B(n_1105),
.Y(n_1456)
);

XOR2xp5_ASAP7_75t_L g1457 ( 
.A(n_1164),
.B(n_624),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1167),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1168),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1168),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1374),
.B(n_1169),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1313),
.B(n_847),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1274),
.B(n_1213),
.C(n_738),
.Y(n_1463)
);

NOR2xp33_ASAP7_75t_L g1464 ( 
.A(n_1343),
.B(n_1179),
.Y(n_1464)
);

OR2x2_ASAP7_75t_L g1465 ( 
.A(n_1272),
.B(n_1294),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1373),
.Y(n_1466)
);

NAND2xp33_ASAP7_75t_L g1467 ( 
.A(n_1307),
.B(n_1169),
.Y(n_1467)
);

AOI21xp5_ASAP7_75t_L g1468 ( 
.A1(n_1292),
.A2(n_1244),
.B(n_1236),
.Y(n_1468)
);

AOI22xp5_ASAP7_75t_L g1469 ( 
.A1(n_1314),
.A2(n_1169),
.B1(n_1179),
.B2(n_1260),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1374),
.B(n_1174),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1394),
.Y(n_1471)
);

INVx2_ASAP7_75t_L g1472 ( 
.A(n_1398),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1381),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1378),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1318),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1285),
.B(n_1174),
.Y(n_1476)
);

BUFx4_ASAP7_75t_L g1477 ( 
.A(n_1304),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1285),
.B(n_1182),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1309),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1399),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1319),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1400),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1408),
.B(n_1182),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1408),
.B(n_1137),
.Y(n_1484)
);

NOR2xp33_ASAP7_75t_L g1485 ( 
.A(n_1343),
.B(n_1260),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1292),
.A2(n_1161),
.B1(n_1183),
.B2(n_1146),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1321),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1410),
.B(n_1146),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1322),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1266),
.B(n_1146),
.Y(n_1490)
);

NOR2xp33_ASAP7_75t_SL g1491 ( 
.A(n_1282),
.B(n_847),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1421),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1266),
.B(n_1161),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_SL g1494 ( 
.A(n_1382),
.B(n_1176),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_SL g1495 ( 
.A(n_1342),
.B(n_1176),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1323),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1327),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1329),
.B(n_1161),
.Y(n_1498)
);

OR2x2_ASAP7_75t_L g1499 ( 
.A(n_1296),
.B(n_1183),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1280),
.B(n_856),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1328),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1387),
.B(n_1183),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_L g1503 ( 
.A(n_1280),
.B(n_1188),
.Y(n_1503)
);

AO221x1_ASAP7_75t_L g1504 ( 
.A1(n_1360),
.A2(n_758),
.B1(n_616),
.B2(n_1236),
.C(n_1176),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1396),
.B(n_1188),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1371),
.B(n_1242),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1344),
.B(n_1331),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_SL g1508 ( 
.A(n_1283),
.B(n_1176),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1402),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1404),
.Y(n_1510)
);

INVx4_ASAP7_75t_L g1511 ( 
.A(n_1448),
.Y(n_1511)
);

NAND3xp33_ASAP7_75t_L g1512 ( 
.A(n_1347),
.B(n_672),
.C(n_671),
.Y(n_1512)
);

NOR2xp33_ASAP7_75t_L g1513 ( 
.A(n_1344),
.B(n_1331),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1330),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1411),
.Y(n_1515)
);

NAND3xp33_ASAP7_75t_L g1516 ( 
.A(n_1347),
.B(n_674),
.C(n_673),
.Y(n_1516)
);

BUFx3_ASAP7_75t_L g1517 ( 
.A(n_1297),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1332),
.Y(n_1518)
);

BUFx5_ASAP7_75t_L g1519 ( 
.A(n_1307),
.Y(n_1519)
);

AND2x6_ASAP7_75t_L g1520 ( 
.A(n_1391),
.B(n_1242),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1333),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1308),
.B(n_1236),
.Y(n_1522)
);

BUFx3_ASAP7_75t_L g1523 ( 
.A(n_1297),
.Y(n_1523)
);

NOR2xp33_ASAP7_75t_L g1524 ( 
.A(n_1337),
.B(n_1242),
.Y(n_1524)
);

AOI22xp5_ASAP7_75t_L g1525 ( 
.A1(n_1337),
.A2(n_852),
.B1(n_766),
.B2(n_675),
.Y(n_1525)
);

NAND3xp33_ASAP7_75t_L g1526 ( 
.A(n_1380),
.B(n_679),
.C(n_676),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1412),
.Y(n_1527)
);

NAND2xp5_ASAP7_75t_L g1528 ( 
.A(n_1324),
.B(n_1245),
.Y(n_1528)
);

O2A1O1Ixp5_ASAP7_75t_L g1529 ( 
.A1(n_1380),
.A2(n_1192),
.B(n_1076),
.C(n_1078),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1335),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1388),
.B(n_1247),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1336),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1339),
.B(n_1245),
.Y(n_1533)
);

NOR2xp33_ASAP7_75t_L g1534 ( 
.A(n_1339),
.B(n_1247),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1440),
.B(n_1249),
.Y(n_1535)
);

NAND2xp5_ASAP7_75t_L g1536 ( 
.A(n_1451),
.B(n_1249),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1393),
.B(n_1251),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1395),
.B(n_1251),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1311),
.A2(n_1248),
.B1(n_1253),
.B2(n_1252),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1413),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1279),
.A2(n_628),
.B1(n_630),
.B2(n_624),
.Y(n_1541)
);

INVx2_ASAP7_75t_SL g1542 ( 
.A(n_1310),
.Y(n_1542)
);

NOR2xp67_ASAP7_75t_L g1543 ( 
.A(n_1415),
.B(n_1071),
.Y(n_1543)
);

NAND3xp33_ASAP7_75t_L g1544 ( 
.A(n_1365),
.B(n_682),
.C(n_669),
.Y(n_1544)
);

INVx8_ASAP7_75t_L g1545 ( 
.A(n_1422),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1379),
.B(n_1248),
.Y(n_1546)
);

AOI221xp5_ASAP7_75t_L g1547 ( 
.A1(n_1457),
.A2(n_948),
.B1(n_949),
.B2(n_947),
.C(n_942),
.Y(n_1547)
);

NAND2xp33_ASAP7_75t_L g1548 ( 
.A(n_1307),
.B(n_1236),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_SL g1549 ( 
.A(n_1290),
.B(n_1047),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1416),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1433),
.B(n_1252),
.Y(n_1551)
);

INVx3_ASAP7_75t_L g1552 ( 
.A(n_1334),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1262),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1338),
.Y(n_1554)
);

BUFx3_ASAP7_75t_L g1555 ( 
.A(n_1293),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1340),
.A2(n_725),
.B1(n_728),
.B2(n_720),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1263),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1265),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1279),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_SL g1560 ( 
.A(n_1290),
.B(n_1047),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1341),
.B(n_1253),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1350),
.B(n_856),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1345),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1270),
.Y(n_1564)
);

OR2x2_ASAP7_75t_L g1565 ( 
.A(n_1454),
.B(n_962),
.Y(n_1565)
);

AO22x1_ASAP7_75t_L g1566 ( 
.A1(n_1405),
.A2(n_630),
.B1(n_631),
.B2(n_625),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_SL g1567 ( 
.A(n_1448),
.B(n_1449),
.Y(n_1567)
);

BUFx6f_ASAP7_75t_SL g1568 ( 
.A(n_1391),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1348),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1349),
.B(n_1240),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1273),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1278),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1448),
.B(n_1385),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1351),
.B(n_1240),
.Y(n_1574)
);

INVx2_ASAP7_75t_L g1575 ( 
.A(n_1281),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1352),
.B(n_922),
.Y(n_1576)
);

NOR2xp33_ASAP7_75t_L g1577 ( 
.A(n_1403),
.B(n_1376),
.Y(n_1577)
);

OR2x2_ASAP7_75t_L g1578 ( 
.A(n_1358),
.B(n_962),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1356),
.B(n_922),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1359),
.B(n_922),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1286),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1287),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1363),
.A2(n_737),
.B1(n_743),
.B2(n_736),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1350),
.B(n_856),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1288),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1364),
.B(n_922),
.Y(n_1586)
);

INVx2_ASAP7_75t_L g1587 ( 
.A(n_1298),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1403),
.B(n_1077),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1366),
.A2(n_1370),
.B1(n_1372),
.B2(n_1369),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1377),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_SL g1591 ( 
.A(n_1423),
.B(n_1334),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1383),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1384),
.B(n_1077),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1386),
.B(n_1079),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1299),
.B(n_1081),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1376),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_L g1597 ( 
.A(n_1361),
.B(n_1081),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1427),
.A2(n_631),
.B1(n_632),
.B2(n_625),
.Y(n_1598)
);

INVx2_ASAP7_75t_L g1599 ( 
.A(n_1300),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1301),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1303),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1306),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1312),
.B(n_1083),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1315),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1417),
.B(n_1083),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1418),
.B(n_1419),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_SL g1607 ( 
.A(n_1261),
.B(n_1064),
.Y(n_1607)
);

NAND2xp33_ASAP7_75t_L g1608 ( 
.A(n_1307),
.B(n_1085),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1432),
.B(n_915),
.Y(n_1609)
);

OAI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1414),
.A2(n_1291),
.B1(n_1346),
.B2(n_1305),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1409),
.B(n_915),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1422),
.B(n_1361),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1355),
.B(n_1085),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1420),
.B(n_1071),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1414),
.B(n_1084),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1291),
.B(n_1084),
.Y(n_1616)
);

NOR2xp33_ASAP7_75t_L g1617 ( 
.A(n_1355),
.B(n_1357),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1424),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1261),
.B(n_1064),
.Y(n_1619)
);

INVx3_ASAP7_75t_L g1620 ( 
.A(n_1261),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1428),
.B(n_1430),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1431),
.B(n_1105),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1435),
.B(n_1106),
.Y(n_1623)
);

OR2x6_ASAP7_75t_L g1624 ( 
.A(n_1422),
.B(n_1116),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1436),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1437),
.B(n_1106),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1267),
.A2(n_632),
.B1(n_633),
.B2(n_628),
.Y(n_1627)
);

INVx2_ASAP7_75t_L g1628 ( 
.A(n_1268),
.Y(n_1628)
);

BUFx8_ASAP7_75t_L g1629 ( 
.A(n_1452),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1438),
.B(n_1107),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1441),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1445),
.B(n_928),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1442),
.B(n_1107),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1357),
.B(n_1108),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1443),
.B(n_1108),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1444),
.B(n_1109),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1446),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1452),
.Y(n_1638)
);

AOI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1269),
.A2(n_634),
.B1(n_635),
.B2(n_633),
.Y(n_1639)
);

INVx2_ASAP7_75t_SL g1640 ( 
.A(n_1354),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1447),
.Y(n_1641)
);

NOR2xp33_ASAP7_75t_L g1642 ( 
.A(n_1375),
.B(n_1109),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1450),
.B(n_1114),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1271),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1375),
.B(n_1114),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1453),
.B(n_1117),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1455),
.B(n_928),
.Y(n_1647)
);

CKINVDCx5p33_ASAP7_75t_R g1648 ( 
.A(n_1456),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1276),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1354),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1277),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1458),
.Y(n_1652)
);

AOI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1295),
.A2(n_635),
.B1(n_637),
.B2(n_634),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1459),
.B(n_1117),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_SL g1655 ( 
.A(n_1325),
.B(n_637),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1460),
.B(n_638),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1317),
.Y(n_1657)
);

INVxp67_ASAP7_75t_SL g1658 ( 
.A(n_1456),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1261),
.B(n_1064),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1389),
.B(n_638),
.Y(n_1660)
);

INVx8_ASAP7_75t_L g1661 ( 
.A(n_1307),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1305),
.A2(n_745),
.B1(n_760),
.B2(n_744),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1320),
.Y(n_1663)
);

INVxp67_ASAP7_75t_L g1664 ( 
.A(n_1439),
.Y(n_1664)
);

INVx4_ASAP7_75t_L g1665 ( 
.A(n_1520),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1617),
.B(n_1326),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1466),
.B(n_1353),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1475),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1473),
.B(n_1474),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1471),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1533),
.B(n_1362),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1534),
.A2(n_1289),
.B1(n_1397),
.B2(n_1426),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1477),
.Y(n_1673)
);

NOR2xp33_ASAP7_75t_SL g1674 ( 
.A(n_1648),
.B(n_1407),
.Y(n_1674)
);

OR2x6_ASAP7_75t_L g1675 ( 
.A(n_1545),
.B(n_1397),
.Y(n_1675)
);

OAI22xp5_ASAP7_75t_L g1676 ( 
.A1(n_1461),
.A2(n_1346),
.B1(n_1426),
.B2(n_1302),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1609),
.B(n_646),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1472),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_SL g1679 ( 
.A(n_1524),
.B(n_1264),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1610),
.A2(n_1284),
.B(n_1302),
.Y(n_1680)
);

NOR2xp33_ASAP7_75t_L g1681 ( 
.A(n_1507),
.B(n_1275),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1546),
.B(n_646),
.Y(n_1682)
);

OAI21xp33_ASAP7_75t_L g1683 ( 
.A1(n_1463),
.A2(n_650),
.B(n_648),
.Y(n_1683)
);

AO21x1_ASAP7_75t_L g1684 ( 
.A1(n_1658),
.A2(n_1289),
.B(n_1316),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1551),
.B(n_1367),
.Y(n_1685)
);

OAI22xp5_ASAP7_75t_L g1686 ( 
.A1(n_1490),
.A2(n_1425),
.B1(n_1284),
.B2(n_1264),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1588),
.B(n_1264),
.Y(n_1687)
);

NOR2xp67_ASAP7_75t_L g1688 ( 
.A(n_1559),
.B(n_1513),
.Y(n_1688)
);

AOI21xp5_ASAP7_75t_L g1689 ( 
.A1(n_1608),
.A2(n_1548),
.B(n_1467),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1462),
.B(n_648),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1468),
.A2(n_1425),
.B(n_1275),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1484),
.A2(n_1368),
.B(n_1434),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1520),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1465),
.B(n_1390),
.Y(n_1694)
);

AOI21xp5_ASAP7_75t_L g1695 ( 
.A1(n_1484),
.A2(n_1368),
.B(n_1434),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1499),
.Y(n_1696)
);

OAI21xp33_ASAP7_75t_L g1697 ( 
.A1(n_1512),
.A2(n_653),
.B(n_650),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1517),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1516),
.A2(n_1401),
.B(n_1406),
.C(n_1392),
.Y(n_1699)
);

AOI21xp5_ASAP7_75t_L g1700 ( 
.A1(n_1476),
.A2(n_1429),
.B(n_1119),
.Y(n_1700)
);

INVxp67_ASAP7_75t_L g1701 ( 
.A(n_1632),
.Y(n_1701)
);

AND2x2_ASAP7_75t_SL g1702 ( 
.A(n_1655),
.B(n_761),
.Y(n_1702)
);

OAI21xp33_ASAP7_75t_L g1703 ( 
.A1(n_1662),
.A2(n_655),
.B(n_653),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1470),
.B(n_655),
.Y(n_1704)
);

AOI22xp5_ASAP7_75t_L g1705 ( 
.A1(n_1544),
.A2(n_740),
.B1(n_748),
.B2(n_656),
.Y(n_1705)
);

A2O1A1Ixp33_ASAP7_75t_L g1706 ( 
.A1(n_1613),
.A2(n_1119),
.B(n_1120),
.C(n_1116),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1577),
.B(n_765),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1500),
.B(n_656),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1470),
.B(n_1528),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1476),
.A2(n_1119),
.B(n_1116),
.Y(n_1710)
);

AOI33xp33_ASAP7_75t_L g1711 ( 
.A1(n_1541),
.A2(n_773),
.A3(n_790),
.B1(n_798),
.B2(n_797),
.B3(n_768),
.Y(n_1711)
);

INVx4_ASAP7_75t_L g1712 ( 
.A(n_1520),
.Y(n_1712)
);

AOI21xp33_ASAP7_75t_L g1713 ( 
.A1(n_1662),
.A2(n_1120),
.B(n_1113),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1542),
.B(n_1498),
.Y(n_1714)
);

BUFx3_ASAP7_75t_L g1715 ( 
.A(n_1629),
.Y(n_1715)
);

AOI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1478),
.A2(n_1120),
.B(n_1064),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1478),
.A2(n_1486),
.B(n_1615),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1486),
.A2(n_1122),
.B(n_1064),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_SL g1719 ( 
.A(n_1490),
.B(n_1122),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1503),
.B(n_740),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1615),
.A2(n_1122),
.B(n_1113),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1523),
.B(n_748),
.Y(n_1722)
);

A2O1A1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1634),
.A2(n_819),
.B(n_820),
.C(n_811),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1483),
.A2(n_1493),
.B(n_1616),
.Y(n_1724)
);

NOR3xp33_ASAP7_75t_L g1725 ( 
.A(n_1566),
.B(n_864),
.C(n_845),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_SL g1726 ( 
.A(n_1464),
.B(n_1122),
.Y(n_1726)
);

AOI21xp5_ASAP7_75t_L g1727 ( 
.A1(n_1483),
.A2(n_1122),
.B(n_1113),
.Y(n_1727)
);

AOI21xp5_ASAP7_75t_L g1728 ( 
.A1(n_1616),
.A2(n_1103),
.B(n_1007),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1479),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1563),
.B(n_929),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1480),
.Y(n_1731)
);

A2O1A1Ixp33_ASAP7_75t_L g1732 ( 
.A1(n_1526),
.A2(n_849),
.B(n_855),
.C(n_831),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1481),
.B(n_827),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1482),
.Y(n_1734)
);

A2O1A1Ixp33_ASAP7_75t_L g1735 ( 
.A1(n_1502),
.A2(n_1506),
.B(n_1664),
.C(n_1485),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1487),
.B(n_827),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1509),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1489),
.B(n_829),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1496),
.B(n_829),
.Y(n_1739)
);

AOI21xp5_ASAP7_75t_L g1740 ( 
.A1(n_1661),
.A2(n_1488),
.B(n_1607),
.Y(n_1740)
);

BUFx2_ASAP7_75t_L g1741 ( 
.A(n_1555),
.Y(n_1741)
);

O2A1O1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1556),
.A2(n_860),
.B(n_858),
.C(n_929),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_SL g1743 ( 
.A(n_1494),
.B(n_983),
.Y(n_1743)
);

OAI21xp5_ASAP7_75t_L g1744 ( 
.A1(n_1529),
.A2(n_1103),
.B(n_1007),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1510),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_SL g1746 ( 
.A(n_1552),
.B(n_830),
.Y(n_1746)
);

O2A1O1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1556),
.A2(n_951),
.B(n_953),
.C(n_950),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1497),
.B(n_830),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1515),
.Y(n_1749)
);

NAND2x1p5_ASAP7_75t_L g1750 ( 
.A(n_1511),
.B(n_1008),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1598),
.B(n_832),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1501),
.B(n_832),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1514),
.B(n_1518),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1521),
.Y(n_1754)
);

A2O1A1Ixp33_ASAP7_75t_L g1755 ( 
.A1(n_1505),
.A2(n_1008),
.B(n_951),
.C(n_953),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_SL g1756 ( 
.A(n_1552),
.B(n_1488),
.Y(n_1756)
);

AND2x4_ASAP7_75t_L g1757 ( 
.A(n_1612),
.B(n_1008),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1527),
.Y(n_1758)
);

INVx11_ASAP7_75t_L g1759 ( 
.A(n_1629),
.Y(n_1759)
);

A2O1A1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1597),
.A2(n_956),
.B(n_959),
.C(n_950),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1583),
.A2(n_959),
.B(n_960),
.C(n_956),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1530),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_SL g1763 ( 
.A(n_1591),
.B(n_1537),
.Y(n_1763)
);

AOI21xp5_ASAP7_75t_L g1764 ( 
.A1(n_1661),
.A2(n_893),
.B(n_889),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1661),
.A2(n_893),
.B(n_889),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1504),
.A2(n_835),
.B1(n_837),
.B2(n_833),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_L g1767 ( 
.A(n_1532),
.B(n_833),
.Y(n_1767)
);

A2O1A1Ixp33_ASAP7_75t_L g1768 ( 
.A1(n_1642),
.A2(n_964),
.B(n_965),
.C(n_960),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1492),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1589),
.A2(n_854),
.B1(n_835),
.B2(n_842),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1554),
.B(n_837),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1569),
.B(n_842),
.Y(n_1772)
);

BUFx6f_ASAP7_75t_L g1773 ( 
.A(n_1492),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1619),
.A2(n_898),
.B(n_897),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1538),
.B(n_844),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1469),
.B(n_844),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1659),
.A2(n_898),
.B(n_897),
.Y(n_1777)
);

AOI21xp5_ASAP7_75t_L g1778 ( 
.A1(n_1589),
.A2(n_903),
.B(n_990),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1594),
.A2(n_990),
.B(n_1004),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1525),
.B(n_1491),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1590),
.B(n_846),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1568),
.B(n_846),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1592),
.B(n_1647),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_L g1784 ( 
.A(n_1611),
.Y(n_1784)
);

AOI22xp5_ASAP7_75t_L g1785 ( 
.A1(n_1520),
.A2(n_850),
.B1(n_853),
.B2(n_848),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1535),
.B(n_848),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1565),
.Y(n_1787)
);

NAND2xp5_ASAP7_75t_L g1788 ( 
.A(n_1562),
.B(n_850),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_SL g1789 ( 
.A(n_1536),
.B(n_853),
.Y(n_1789)
);

AOI21xp5_ASAP7_75t_L g1790 ( 
.A1(n_1594),
.A2(n_1574),
.B(n_1570),
.Y(n_1790)
);

O2A1O1Ixp5_ASAP7_75t_L g1791 ( 
.A1(n_1495),
.A2(n_965),
.B(n_966),
.C(n_964),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1584),
.B(n_854),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1600),
.Y(n_1793)
);

OAI21x1_ASAP7_75t_SL g1794 ( 
.A1(n_1640),
.A2(n_966),
.B(n_2),
.Y(n_1794)
);

AOI21xp5_ASAP7_75t_L g1795 ( 
.A1(n_1561),
.A2(n_990),
.B(n_1005),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1568),
.B(n_857),
.Y(n_1796)
);

AND2x2_ASAP7_75t_SL g1797 ( 
.A(n_1511),
.B(n_1005),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1547),
.B(n_857),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_L g1799 ( 
.A1(n_1576),
.A2(n_1022),
.B(n_684),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1579),
.A2(n_990),
.B(n_1005),
.Y(n_1800)
);

AOI21xp5_ASAP7_75t_L g1801 ( 
.A1(n_1580),
.A2(n_1013),
.B(n_1005),
.Y(n_1801)
);

O2A1O1Ixp33_ASAP7_75t_SL g1802 ( 
.A1(n_1522),
.A2(n_2),
.B(n_0),
.C(n_1),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1601),
.B(n_859),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_SL g1804 ( 
.A(n_1492),
.B(n_859),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1604),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_SL g1806 ( 
.A(n_1650),
.B(n_861),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_SL g1807 ( 
.A(n_1543),
.B(n_861),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_SL g1808 ( 
.A(n_1519),
.B(n_1573),
.Y(n_1808)
);

AOI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1586),
.A2(n_1013),
.B(n_1005),
.Y(n_1809)
);

INVx3_ASAP7_75t_L g1810 ( 
.A(n_1624),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1618),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1593),
.A2(n_1013),
.B(n_1022),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1578),
.A2(n_862),
.B1(n_686),
.B2(n_687),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1625),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1596),
.B(n_862),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1540),
.B(n_680),
.Y(n_1816)
);

AND2x6_ASAP7_75t_L g1817 ( 
.A(n_1620),
.B(n_1006),
.Y(n_1817)
);

NOR2xp33_ASAP7_75t_SL g1818 ( 
.A(n_1545),
.B(n_1006),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1595),
.A2(n_1022),
.B(n_1006),
.Y(n_1819)
);

AOI21xp33_ASAP7_75t_L g1820 ( 
.A1(n_1660),
.A2(n_1006),
.B(n_1022),
.Y(n_1820)
);

NOR2xp33_ASAP7_75t_L g1821 ( 
.A(n_1549),
.B(n_689),
.Y(n_1821)
);

OAI21xp5_ASAP7_75t_L g1822 ( 
.A1(n_1645),
.A2(n_691),
.B(n_690),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1595),
.A2(n_693),
.B(n_692),
.Y(n_1823)
);

BUFx4f_ASAP7_75t_L g1824 ( 
.A(n_1545),
.Y(n_1824)
);

INVx3_ASAP7_75t_L g1825 ( 
.A(n_1624),
.Y(n_1825)
);

INVx3_ASAP7_75t_L g1826 ( 
.A(n_1624),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1550),
.B(n_698),
.Y(n_1827)
);

INVx1_ASAP7_75t_SL g1828 ( 
.A(n_1560),
.Y(n_1828)
);

OAI21xp33_ASAP7_75t_L g1829 ( 
.A1(n_1627),
.A2(n_822),
.B(n_734),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1553),
.B(n_699),
.Y(n_1830)
);

HB1xp67_ASAP7_75t_L g1831 ( 
.A(n_1612),
.Y(n_1831)
);

NOR2xp33_ASAP7_75t_L g1832 ( 
.A(n_1638),
.B(n_700),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1557),
.B(n_707),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1603),
.A2(n_1605),
.B(n_1622),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1558),
.B(n_710),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1656),
.A2(n_714),
.B1(n_719),
.B2(n_713),
.Y(n_1836)
);

AOI21xp5_ASAP7_75t_L g1837 ( 
.A1(n_1603),
.A2(n_724),
.B(n_723),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1564),
.B(n_727),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1583),
.B(n_731),
.Y(n_1839)
);

AOI21xp5_ASAP7_75t_L g1840 ( 
.A1(n_1605),
.A2(n_739),
.B(n_735),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1571),
.B(n_741),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1606),
.A2(n_746),
.B(n_742),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1631),
.Y(n_1843)
);

O2A1O1Ixp33_ASAP7_75t_L g1844 ( 
.A1(n_1508),
.A2(n_750),
.B(n_751),
.C(n_747),
.Y(n_1844)
);

AO21x1_ASAP7_75t_L g1845 ( 
.A1(n_1606),
.A2(n_1010),
.B(n_0),
.Y(n_1845)
);

AOI21xp5_ASAP7_75t_L g1846 ( 
.A1(n_1622),
.A2(n_755),
.B(n_752),
.Y(n_1846)
);

OAI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1623),
.A2(n_757),
.B(n_756),
.Y(n_1847)
);

OAI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1623),
.A2(n_762),
.B(n_759),
.Y(n_1848)
);

AOI21xp5_ASAP7_75t_L g1849 ( 
.A1(n_1626),
.A2(n_764),
.B(n_763),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1626),
.A2(n_774),
.B(n_770),
.Y(n_1850)
);

AOI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1630),
.A2(n_777),
.B(n_776),
.Y(n_1851)
);

INVx2_ASAP7_75t_SL g1852 ( 
.A(n_1612),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1572),
.B(n_778),
.Y(n_1853)
);

A2O1A1Ixp33_ASAP7_75t_L g1854 ( 
.A1(n_1531),
.A2(n_780),
.B(n_781),
.C(n_779),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1567),
.A2(n_784),
.B1(n_785),
.B2(n_783),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1680),
.A2(n_1621),
.B(n_1630),
.Y(n_1856)
);

NOR2xp33_ASAP7_75t_L g1857 ( 
.A(n_1701),
.B(n_786),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1784),
.B(n_1575),
.Y(n_1858)
);

AOI21xp5_ASAP7_75t_L g1859 ( 
.A1(n_1689),
.A2(n_1621),
.B(n_1633),
.Y(n_1859)
);

NOR2xp33_ASAP7_75t_SL g1860 ( 
.A(n_1702),
.B(n_1581),
.Y(n_1860)
);

A2O1A1Ixp33_ASAP7_75t_SL g1861 ( 
.A1(n_1832),
.A2(n_1620),
.B(n_1653),
.C(n_1639),
.Y(n_1861)
);

OAI21xp33_ASAP7_75t_L g1862 ( 
.A1(n_1839),
.A2(n_789),
.B(n_788),
.Y(n_1862)
);

OAI21xp5_ASAP7_75t_L g1863 ( 
.A1(n_1735),
.A2(n_1635),
.B(n_1633),
.Y(n_1863)
);

CKINVDCx8_ASAP7_75t_R g1864 ( 
.A(n_1769),
.Y(n_1864)
);

AOI22xp33_ASAP7_75t_L g1865 ( 
.A1(n_1707),
.A2(n_1539),
.B1(n_1644),
.B2(n_1628),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1670),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1847),
.A2(n_1641),
.B(n_1652),
.C(n_1637),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1666),
.B(n_1582),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1753),
.Y(n_1869)
);

AO22x1_ASAP7_75t_L g1870 ( 
.A1(n_1780),
.A2(n_1673),
.B1(n_1751),
.B2(n_1725),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1717),
.A2(n_1636),
.B(n_1635),
.Y(n_1871)
);

O2A1O1Ixp33_ASAP7_75t_L g1872 ( 
.A1(n_1723),
.A2(n_1636),
.B(n_1646),
.C(n_1643),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1783),
.B(n_1585),
.Y(n_1873)
);

INVx3_ASAP7_75t_L g1874 ( 
.A(n_1665),
.Y(n_1874)
);

AOI21xp33_ASAP7_75t_L g1875 ( 
.A1(n_1822),
.A2(n_1646),
.B(n_1643),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1694),
.B(n_1587),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_SL g1877 ( 
.A(n_1674),
.B(n_1519),
.Y(n_1877)
);

A2O1A1Ixp33_ASAP7_75t_SL g1878 ( 
.A1(n_1847),
.A2(n_1602),
.B(n_1599),
.C(n_1649),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1709),
.B(n_1651),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1671),
.B(n_1657),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1682),
.B(n_792),
.Y(n_1881)
);

AOI21xp5_ASAP7_75t_L g1882 ( 
.A1(n_1724),
.A2(n_1654),
.B(n_1614),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1676),
.A2(n_1519),
.B(n_1663),
.Y(n_1883)
);

AOI21xp5_ASAP7_75t_L g1884 ( 
.A1(n_1686),
.A2(n_1519),
.B(n_795),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1669),
.B(n_793),
.Y(n_1885)
);

OR2x2_ASAP7_75t_L g1886 ( 
.A(n_1696),
.B(n_796),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1678),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1698),
.Y(n_1888)
);

AOI21xp5_ASAP7_75t_L g1889 ( 
.A1(n_1718),
.A2(n_1519),
.B(n_800),
.Y(n_1889)
);

OAI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1848),
.A2(n_801),
.B1(n_802),
.B2(n_799),
.Y(n_1890)
);

AOI21xp5_ASAP7_75t_L g1891 ( 
.A1(n_1834),
.A2(n_1519),
.B(n_806),
.Y(n_1891)
);

NOR3xp33_ASAP7_75t_L g1892 ( 
.A(n_1683),
.B(n_808),
.C(n_803),
.Y(n_1892)
);

INVx3_ASAP7_75t_L g1893 ( 
.A(n_1665),
.Y(n_1893)
);

CKINVDCx20_ASAP7_75t_R g1894 ( 
.A(n_1715),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1685),
.B(n_809),
.Y(n_1895)
);

NAND2x1p5_ASAP7_75t_L g1896 ( 
.A(n_1824),
.B(n_1693),
.Y(n_1896)
);

INVx2_ASAP7_75t_SL g1897 ( 
.A(n_1769),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1731),
.Y(n_1898)
);

NOR2xp33_ASAP7_75t_L g1899 ( 
.A(n_1741),
.B(n_810),
.Y(n_1899)
);

NOR2xp67_ASAP7_75t_L g1900 ( 
.A(n_1681),
.B(n_1012),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1677),
.B(n_812),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1852),
.B(n_1810),
.Y(n_1902)
);

AOI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1834),
.A2(n_814),
.B(n_813),
.Y(n_1903)
);

NOR2xp33_ASAP7_75t_L g1904 ( 
.A(n_1788),
.B(n_1792),
.Y(n_1904)
);

OAI22xp33_ASAP7_75t_L g1905 ( 
.A1(n_1766),
.A2(n_823),
.B1(n_824),
.B2(n_816),
.Y(n_1905)
);

AOI21xp5_ASAP7_75t_L g1906 ( 
.A1(n_1691),
.A2(n_825),
.B(n_1012),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1704),
.B(n_1010),
.Y(n_1907)
);

BUFx12f_ASAP7_75t_L g1908 ( 
.A(n_1769),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1692),
.A2(n_1012),
.B(n_3),
.Y(n_1909)
);

AOI22xp5_ASAP7_75t_L g1910 ( 
.A1(n_1703),
.A2(n_1010),
.B1(n_1012),
.B2(n_5),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1695),
.A2(n_1012),
.B(n_3),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1790),
.A2(n_4),
.B(n_6),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1696),
.B(n_4),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1787),
.B(n_7),
.Y(n_1914)
);

AOI21xp5_ASAP7_75t_L g1915 ( 
.A1(n_1740),
.A2(n_7),
.B(n_8),
.Y(n_1915)
);

OA22x2_ASAP7_75t_L g1916 ( 
.A1(n_1848),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1668),
.Y(n_1917)
);

INVx3_ASAP7_75t_SL g1918 ( 
.A(n_1773),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1798),
.A2(n_12),
.B1(n_9),
.B2(n_10),
.Y(n_1919)
);

BUFx6f_ASAP7_75t_L g1920 ( 
.A(n_1824),
.Y(n_1920)
);

NOR2xp33_ASAP7_75t_L g1921 ( 
.A(n_1782),
.B(n_13),
.Y(n_1921)
);

BUFx8_ASAP7_75t_L g1922 ( 
.A(n_1722),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1714),
.B(n_13),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1754),
.B(n_14),
.Y(n_1924)
);

BUFx6f_ASAP7_75t_L g1925 ( 
.A(n_1773),
.Y(n_1925)
);

INVx3_ASAP7_75t_L g1926 ( 
.A(n_1693),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1716),
.A2(n_14),
.B(n_15),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1810),
.B(n_16),
.Y(n_1928)
);

BUFx3_ASAP7_75t_L g1929 ( 
.A(n_1773),
.Y(n_1929)
);

OAI22xp5_ASAP7_75t_L g1930 ( 
.A1(n_1785),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1779),
.A2(n_18),
.B(n_19),
.Y(n_1931)
);

OA22x2_ASAP7_75t_L g1932 ( 
.A1(n_1855),
.A2(n_23),
.B1(n_20),
.B2(n_21),
.Y(n_1932)
);

AO32x1_ASAP7_75t_L g1933 ( 
.A1(n_1770),
.A2(n_24),
.A3(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1762),
.B(n_24),
.Y(n_1934)
);

OAI21xp5_ASAP7_75t_L g1935 ( 
.A1(n_1822),
.A2(n_25),
.B(n_26),
.Y(n_1935)
);

A2O1A1Ixp33_ASAP7_75t_L g1936 ( 
.A1(n_1697),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_1936)
);

OAI22xp5_ASAP7_75t_L g1937 ( 
.A1(n_1672),
.A2(n_31),
.B1(n_27),
.B2(n_28),
.Y(n_1937)
);

BUFx12f_ASAP7_75t_L g1938 ( 
.A(n_1730),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1734),
.Y(n_1939)
);

O2A1O1Ixp33_ASAP7_75t_L g1940 ( 
.A1(n_1732),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1721),
.A2(n_32),
.B(n_34),
.Y(n_1941)
);

AOI21xp5_ASAP7_75t_L g1942 ( 
.A1(n_1800),
.A2(n_35),
.B(n_36),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1711),
.B(n_35),
.Y(n_1943)
);

CKINVDCx8_ASAP7_75t_R g1944 ( 
.A(n_1796),
.Y(n_1944)
);

O2A1O1Ixp5_ASAP7_75t_L g1945 ( 
.A1(n_1845),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1667),
.B(n_37),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1829),
.B(n_39),
.C(n_40),
.Y(n_1947)
);

NOR2x1p5_ASAP7_75t_L g1948 ( 
.A(n_1712),
.B(n_39),
.Y(n_1948)
);

INVx1_ASAP7_75t_SL g1949 ( 
.A(n_1729),
.Y(n_1949)
);

OA22x2_ASAP7_75t_L g1950 ( 
.A1(n_1763),
.A2(n_42),
.B1(n_40),
.B2(n_41),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_L g1951 ( 
.A(n_1690),
.B(n_43),
.Y(n_1951)
);

OR2x6_ASAP7_75t_L g1952 ( 
.A(n_1712),
.B(n_568),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1801),
.A2(n_1809),
.B(n_1819),
.Y(n_1953)
);

OAI21xp33_ASAP7_75t_L g1954 ( 
.A1(n_1705),
.A2(n_43),
.B(n_44),
.Y(n_1954)
);

AOI21xp5_ASAP7_75t_L g1955 ( 
.A1(n_1719),
.A2(n_45),
.B(n_46),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1793),
.B(n_46),
.Y(n_1956)
);

O2A1O1Ixp33_ASAP7_75t_L g1957 ( 
.A1(n_1854),
.A2(n_49),
.B(n_47),
.C(n_48),
.Y(n_1957)
);

AOI22x1_ASAP7_75t_L g1958 ( 
.A1(n_1823),
.A2(n_51),
.B1(n_47),
.B2(n_50),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1708),
.B(n_50),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1805),
.B(n_51),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1811),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1675),
.Y(n_1962)
);

AOI21xp5_ASAP7_75t_L g1963 ( 
.A1(n_1727),
.A2(n_52),
.B(n_53),
.Y(n_1963)
);

OAI22xp5_ASAP7_75t_L g1964 ( 
.A1(n_1720),
.A2(n_55),
.B1(n_53),
.B2(n_54),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_SL g1965 ( 
.A(n_1674),
.B(n_54),
.Y(n_1965)
);

BUFx3_ASAP7_75t_L g1966 ( 
.A(n_1815),
.Y(n_1966)
);

AOI21xp5_ASAP7_75t_L g1967 ( 
.A1(n_1799),
.A2(n_56),
.B(n_57),
.Y(n_1967)
);

O2A1O1Ixp5_ASAP7_75t_L g1968 ( 
.A1(n_1726),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1968)
);

BUFx4f_ASAP7_75t_L g1969 ( 
.A(n_1675),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1814),
.Y(n_1970)
);

INVxp67_ASAP7_75t_SL g1971 ( 
.A(n_1687),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1843),
.B(n_58),
.Y(n_1972)
);

AOI21xp5_ASAP7_75t_L g1973 ( 
.A1(n_1799),
.A2(n_59),
.B(n_60),
.Y(n_1973)
);

INVx5_ASAP7_75t_L g1974 ( 
.A(n_1817),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1737),
.Y(n_1975)
);

NOR3xp33_ASAP7_75t_L g1976 ( 
.A(n_1679),
.B(n_1836),
.C(n_1804),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1744),
.A2(n_60),
.B(n_61),
.Y(n_1977)
);

AOI21xp5_ASAP7_75t_L g1978 ( 
.A1(n_1744),
.A2(n_61),
.B(n_62),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1688),
.B(n_62),
.Y(n_1979)
);

A2O1A1Ixp33_ASAP7_75t_L g1980 ( 
.A1(n_1742),
.A2(n_67),
.B(n_63),
.C(n_64),
.Y(n_1980)
);

AOI21xp5_ASAP7_75t_L g1981 ( 
.A1(n_1795),
.A2(n_63),
.B(n_64),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1733),
.A2(n_69),
.B1(n_67),
.B2(n_68),
.Y(n_1982)
);

O2A1O1Ixp33_ASAP7_75t_L g1983 ( 
.A1(n_1786),
.A2(n_70),
.B(n_68),
.C(n_69),
.Y(n_1983)
);

BUFx2_ASAP7_75t_L g1984 ( 
.A(n_1675),
.Y(n_1984)
);

OAI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1736),
.A2(n_72),
.B1(n_70),
.B2(n_71),
.Y(n_1985)
);

AOI22xp5_ASAP7_75t_L g1986 ( 
.A1(n_1776),
.A2(n_1821),
.B1(n_1813),
.B2(n_1789),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_L g1987 ( 
.A1(n_1797),
.A2(n_71),
.B(n_73),
.Y(n_1987)
);

AOI21xp5_ASAP7_75t_L g1988 ( 
.A1(n_1710),
.A2(n_73),
.B(n_74),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1745),
.B(n_74),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1749),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1828),
.B(n_75),
.Y(n_1991)
);

OAI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1738),
.A2(n_1739),
.B1(n_1752),
.B2(n_1748),
.Y(n_1992)
);

AO32x1_ASAP7_75t_L g1993 ( 
.A1(n_1758),
.A2(n_77),
.A3(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_1993)
);

BUFx4f_ASAP7_75t_SL g1994 ( 
.A(n_1759),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_SL g1995 ( 
.A(n_1828),
.B(n_76),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1757),
.B(n_77),
.Y(n_1996)
);

AOI21xp5_ASAP7_75t_L g1997 ( 
.A1(n_1706),
.A2(n_78),
.B(n_79),
.Y(n_1997)
);

AOI21xp5_ASAP7_75t_L g1998 ( 
.A1(n_1756),
.A2(n_79),
.B(n_80),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1768),
.Y(n_1999)
);

O2A1O1Ixp33_ASAP7_75t_L g2000 ( 
.A1(n_1775),
.A2(n_82),
.B(n_80),
.C(n_81),
.Y(n_2000)
);

O2A1O1Ixp33_ASAP7_75t_L g2001 ( 
.A1(n_1802),
.A2(n_84),
.B(n_82),
.C(n_83),
.Y(n_2001)
);

AOI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1728),
.A2(n_83),
.B(n_84),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_L g2003 ( 
.A(n_1760),
.B(n_86),
.Y(n_2003)
);

INVx1_ASAP7_75t_SL g2004 ( 
.A(n_1831),
.Y(n_2004)
);

INVx4_ASAP7_75t_L g2005 ( 
.A(n_1757),
.Y(n_2005)
);

O2A1O1Ixp33_ASAP7_75t_L g2006 ( 
.A1(n_1746),
.A2(n_88),
.B(n_86),
.C(n_87),
.Y(n_2006)
);

INVx3_ASAP7_75t_L g2007 ( 
.A(n_1825),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1767),
.B(n_1771),
.Y(n_2008)
);

OAI21xp33_ASAP7_75t_SL g2009 ( 
.A1(n_1743),
.A2(n_89),
.B(n_90),
.Y(n_2009)
);

AOI21xp5_ASAP7_75t_L g2010 ( 
.A1(n_1700),
.A2(n_89),
.B(n_90),
.Y(n_2010)
);

NOR3xp33_ASAP7_75t_L g2011 ( 
.A(n_1806),
.B(n_1844),
.C(n_1807),
.Y(n_2011)
);

AND2x4_ASAP7_75t_L g2012 ( 
.A(n_1825),
.B(n_91),
.Y(n_2012)
);

HB1xp67_ASAP7_75t_L g2013 ( 
.A(n_1826),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1772),
.B(n_91),
.Y(n_2014)
);

A2O1A1Ixp33_ASAP7_75t_L g2015 ( 
.A1(n_1842),
.A2(n_95),
.B(n_93),
.C(n_94),
.Y(n_2015)
);

NOR2xp67_ASAP7_75t_L g2016 ( 
.A(n_1803),
.B(n_571),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_L g2017 ( 
.A(n_1781),
.B(n_93),
.Y(n_2017)
);

HB1xp67_ASAP7_75t_L g2018 ( 
.A(n_1826),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1837),
.A2(n_96),
.B1(n_94),
.B2(n_95),
.Y(n_2019)
);

INVx5_ASAP7_75t_L g2020 ( 
.A(n_1817),
.Y(n_2020)
);

OAI21xp33_ASAP7_75t_L g2021 ( 
.A1(n_1840),
.A2(n_97),
.B(n_98),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1853),
.B(n_98),
.Y(n_2022)
);

OAI21xp33_ASAP7_75t_L g2023 ( 
.A1(n_1846),
.A2(n_1850),
.B(n_1849),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_L g2024 ( 
.A(n_1816),
.B(n_99),
.Y(n_2024)
);

CKINVDCx5p33_ASAP7_75t_R g2025 ( 
.A(n_1827),
.Y(n_2025)
);

OAI22xp5_ASAP7_75t_L g2026 ( 
.A1(n_1851),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_2026)
);

INVx3_ASAP7_75t_L g2027 ( 
.A(n_1750),
.Y(n_2027)
);

OAI22xp5_ASAP7_75t_L g2028 ( 
.A1(n_1830),
.A2(n_103),
.B1(n_100),
.B2(n_102),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1818),
.B(n_572),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1917),
.Y(n_2030)
);

OAI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1860),
.A2(n_1818),
.B1(n_1835),
.B2(n_1833),
.Y(n_2031)
);

OAI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1967),
.A2(n_1778),
.B(n_1791),
.Y(n_2032)
);

INVxp67_ASAP7_75t_SL g2033 ( 
.A(n_2013),
.Y(n_2033)
);

AOI21x1_ASAP7_75t_L g2034 ( 
.A1(n_1900),
.A2(n_1684),
.B(n_1808),
.Y(n_2034)
);

BUFx12f_ASAP7_75t_L g2035 ( 
.A(n_1922),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1908),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1904),
.B(n_102),
.Y(n_2037)
);

A2O1A1Ixp33_ASAP7_75t_L g2038 ( 
.A1(n_1921),
.A2(n_1747),
.B(n_1761),
.C(n_1838),
.Y(n_2038)
);

NOR2xp33_ASAP7_75t_L g2039 ( 
.A(n_1922),
.B(n_103),
.Y(n_2039)
);

AO22x2_ASAP7_75t_L g2040 ( 
.A1(n_1975),
.A2(n_1794),
.B1(n_1841),
.B2(n_1764),
.Y(n_2040)
);

AOI211x1_ASAP7_75t_L g2041 ( 
.A1(n_1862),
.A2(n_1765),
.B(n_1777),
.C(n_1774),
.Y(n_2041)
);

OA21x2_ASAP7_75t_L g2042 ( 
.A1(n_1953),
.A2(n_1755),
.B(n_1820),
.Y(n_2042)
);

A2O1A1Ixp33_ASAP7_75t_L g2043 ( 
.A1(n_1954),
.A2(n_1699),
.B(n_1713),
.C(n_1812),
.Y(n_2043)
);

BUFx6f_ASAP7_75t_L g2044 ( 
.A(n_1920),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1859),
.A2(n_1817),
.B(n_574),
.Y(n_2045)
);

AOI21x1_ASAP7_75t_L g2046 ( 
.A1(n_1977),
.A2(n_1817),
.B(n_104),
.Y(n_2046)
);

OAI21xp5_ASAP7_75t_SL g2047 ( 
.A1(n_1919),
.A2(n_105),
.B(n_106),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1961),
.Y(n_2048)
);

AO31x2_ASAP7_75t_L g2049 ( 
.A1(n_1882),
.A2(n_575),
.A3(n_577),
.B(n_573),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1869),
.B(n_105),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_L g2051 ( 
.A(n_1949),
.B(n_1858),
.Y(n_2051)
);

OAI21xp5_ASAP7_75t_L g2052 ( 
.A1(n_1973),
.A2(n_107),
.B(n_108),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1873),
.B(n_108),
.Y(n_2053)
);

AND2x2_ASAP7_75t_L g2054 ( 
.A(n_1888),
.B(n_1970),
.Y(n_2054)
);

A2O1A1Ixp33_ASAP7_75t_L g2055 ( 
.A1(n_1935),
.A2(n_1957),
.B(n_1947),
.C(n_1940),
.Y(n_2055)
);

INVx6_ASAP7_75t_L g2056 ( 
.A(n_1920),
.Y(n_2056)
);

AOI21xp5_ASAP7_75t_L g2057 ( 
.A1(n_1871),
.A2(n_109),
.B(n_110),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_L g2058 ( 
.A(n_1868),
.B(n_109),
.Y(n_2058)
);

OAI21x1_ASAP7_75t_SL g2059 ( 
.A1(n_1863),
.A2(n_111),
.B(n_112),
.Y(n_2059)
);

NOR2xp33_ASAP7_75t_L g2060 ( 
.A(n_2025),
.B(n_1944),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1994),
.Y(n_2061)
);

AO22x2_ASAP7_75t_L g2062 ( 
.A1(n_1990),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1876),
.B(n_113),
.Y(n_2063)
);

OAI21x1_ASAP7_75t_SL g2064 ( 
.A1(n_1978),
.A2(n_114),
.B(n_115),
.Y(n_2064)
);

INVx2_ASAP7_75t_L g2065 ( 
.A(n_1866),
.Y(n_2065)
);

OAI21x1_ASAP7_75t_SL g2066 ( 
.A1(n_1891),
.A2(n_114),
.B(n_115),
.Y(n_2066)
);

AOI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_1856),
.A2(n_116),
.B(n_117),
.Y(n_2067)
);

OAI21x1_ASAP7_75t_L g2068 ( 
.A1(n_1883),
.A2(n_580),
.B(n_579),
.Y(n_2068)
);

OAI21x1_ASAP7_75t_L g2069 ( 
.A1(n_1909),
.A2(n_582),
.B(n_581),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1879),
.B(n_116),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1877),
.A2(n_117),
.B(n_118),
.Y(n_2071)
);

OR2x2_ASAP7_75t_L g2072 ( 
.A(n_2004),
.B(n_119),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_1928),
.B(n_120),
.Y(n_2073)
);

A2O1A1Ixp33_ASAP7_75t_L g2074 ( 
.A1(n_2023),
.A2(n_122),
.B(n_120),
.C(n_121),
.Y(n_2074)
);

INVx5_ASAP7_75t_L g2075 ( 
.A(n_1952),
.Y(n_2075)
);

AOI21xp5_ASAP7_75t_L g2076 ( 
.A1(n_1872),
.A2(n_123),
.B(n_124),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_1884),
.A2(n_123),
.B(n_124),
.Y(n_2077)
);

BUFx2_ASAP7_75t_L g2078 ( 
.A(n_1918),
.Y(n_2078)
);

AOI21xp5_ASAP7_75t_L g2079 ( 
.A1(n_1911),
.A2(n_125),
.B(n_126),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1880),
.B(n_127),
.Y(n_2080)
);

OAI22xp5_ASAP7_75t_L g2081 ( 
.A1(n_1986),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2081)
);

AOI21xp5_ASAP7_75t_L g2082 ( 
.A1(n_1969),
.A2(n_130),
.B(n_131),
.Y(n_2082)
);

OAI21x1_ASAP7_75t_L g2083 ( 
.A1(n_1981),
.A2(n_584),
.B(n_583),
.Y(n_2083)
);

AOI211x1_ASAP7_75t_L g2084 ( 
.A1(n_1951),
.A2(n_132),
.B(n_130),
.C(n_131),
.Y(n_2084)
);

OAI21x1_ASAP7_75t_L g2085 ( 
.A1(n_1963),
.A2(n_587),
.B(n_585),
.Y(n_2085)
);

A2O1A1Ixp33_ASAP7_75t_L g2086 ( 
.A1(n_2021),
.A2(n_134),
.B(n_132),
.C(n_133),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1929),
.Y(n_2087)
);

NOR2xp33_ASAP7_75t_L g2088 ( 
.A(n_2008),
.B(n_133),
.Y(n_2088)
);

INVx2_ASAP7_75t_SL g2089 ( 
.A(n_1925),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_1923),
.B(n_134),
.Y(n_2090)
);

OAI21xp33_ASAP7_75t_L g2091 ( 
.A1(n_1916),
.A2(n_1950),
.B(n_1936),
.Y(n_2091)
);

OAI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_1937),
.A2(n_135),
.B(n_136),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1928),
.B(n_2012),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2012),
.B(n_135),
.Y(n_2094)
);

AND2x4_ASAP7_75t_L g2095 ( 
.A(n_1962),
.B(n_589),
.Y(n_2095)
);

NOR2xp67_ASAP7_75t_L g2096 ( 
.A(n_1938),
.B(n_137),
.Y(n_2096)
);

INVx4_ASAP7_75t_L g2097 ( 
.A(n_1920),
.Y(n_2097)
);

OAI21x1_ASAP7_75t_L g2098 ( 
.A1(n_1931),
.A2(n_592),
.B(n_591),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_1946),
.B(n_137),
.Y(n_2099)
);

AOI21xp5_ASAP7_75t_L g2100 ( 
.A1(n_1969),
.A2(n_138),
.B(n_139),
.Y(n_2100)
);

NAND3x1_ASAP7_75t_L g2101 ( 
.A(n_1913),
.B(n_138),
.C(n_139),
.Y(n_2101)
);

INVx2_ASAP7_75t_L g2102 ( 
.A(n_1887),
.Y(n_2102)
);

OAI21x1_ASAP7_75t_L g2103 ( 
.A1(n_1941),
.A2(n_594),
.B(n_593),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_1992),
.B(n_140),
.Y(n_2104)
);

OAI21x1_ASAP7_75t_SL g2105 ( 
.A1(n_2001),
.A2(n_140),
.B(n_141),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1924),
.B(n_142),
.Y(n_2106)
);

NAND2x1p5_ASAP7_75t_L g2107 ( 
.A(n_1974),
.B(n_595),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_1959),
.B(n_143),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2018),
.Y(n_2109)
);

AO31x2_ASAP7_75t_L g2110 ( 
.A1(n_1867),
.A2(n_598),
.A3(n_599),
.B(n_596),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_1934),
.B(n_144),
.Y(n_2111)
);

OAI21x1_ASAP7_75t_L g2112 ( 
.A1(n_1942),
.A2(n_1889),
.B(n_1927),
.Y(n_2112)
);

AOI21xp33_ASAP7_75t_L g2113 ( 
.A1(n_1878),
.A2(n_144),
.B(n_145),
.Y(n_2113)
);

OAI21x1_ASAP7_75t_L g2114 ( 
.A1(n_2010),
.A2(n_601),
.B(n_600),
.Y(n_2114)
);

BUFx3_ASAP7_75t_L g2115 ( 
.A(n_1894),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_1966),
.B(n_145),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_1898),
.Y(n_2117)
);

OAI21xp5_ASAP7_75t_L g2118 ( 
.A1(n_1912),
.A2(n_146),
.B(n_147),
.Y(n_2118)
);

CKINVDCx8_ASAP7_75t_R g2119 ( 
.A(n_1925),
.Y(n_2119)
);

AOI22xp5_ASAP7_75t_L g2120 ( 
.A1(n_1870),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1984),
.B(n_1902),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1939),
.Y(n_2122)
);

OAI21x1_ASAP7_75t_L g2123 ( 
.A1(n_1988),
.A2(n_2002),
.B(n_1915),
.Y(n_2123)
);

OAI21x1_ASAP7_75t_L g2124 ( 
.A1(n_1906),
.A2(n_604),
.B(n_603),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1971),
.Y(n_2125)
);

NAND2xp5_ASAP7_75t_L g2126 ( 
.A(n_1956),
.B(n_148),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1881),
.B(n_149),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_1902),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_1874),
.B(n_605),
.Y(n_2129)
);

OAI22x1_ASAP7_75t_L g2130 ( 
.A1(n_1948),
.A2(n_152),
.B1(n_150),
.B2(n_151),
.Y(n_2130)
);

AOI21xp5_ASAP7_75t_L g2131 ( 
.A1(n_1875),
.A2(n_151),
.B(n_152),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_1965),
.A2(n_1993),
.B(n_1952),
.Y(n_2132)
);

OAI21xp5_ASAP7_75t_L g2133 ( 
.A1(n_1980),
.A2(n_153),
.B(n_154),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2007),
.Y(n_2134)
);

BUFx4f_ASAP7_75t_L g2135 ( 
.A(n_1896),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_1989),
.Y(n_2136)
);

OR2x2_ASAP7_75t_L g2137 ( 
.A(n_1886),
.B(n_154),
.Y(n_2137)
);

BUFx2_ASAP7_75t_L g2138 ( 
.A(n_1925),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1960),
.B(n_1972),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2005),
.B(n_155),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_L g2141 ( 
.A(n_1976),
.B(n_157),
.Y(n_2141)
);

OAI21x1_ASAP7_75t_L g2142 ( 
.A1(n_1997),
.A2(n_609),
.B(n_607),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2007),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_2005),
.B(n_610),
.Y(n_2144)
);

OA21x2_ASAP7_75t_L g2145 ( 
.A1(n_1945),
.A2(n_158),
.B(n_159),
.Y(n_2145)
);

INVx2_ASAP7_75t_SL g2146 ( 
.A(n_1897),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_1914),
.B(n_158),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_1864),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_1895),
.B(n_1885),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_2125),
.B(n_2014),
.Y(n_2150)
);

INVx4_ASAP7_75t_L g2151 ( 
.A(n_2075),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2054),
.B(n_1899),
.Y(n_2152)
);

XNOR2xp5_ASAP7_75t_L g2153 ( 
.A(n_2061),
.B(n_1901),
.Y(n_2153)
);

AOI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2141),
.A2(n_2029),
.B(n_1933),
.Y(n_2154)
);

AND2x4_ASAP7_75t_L g2155 ( 
.A(n_2033),
.B(n_1974),
.Y(n_2155)
);

INVx1_ASAP7_75t_L g2156 ( 
.A(n_2030),
.Y(n_2156)
);

BUFx6f_ASAP7_75t_L g2157 ( 
.A(n_2135),
.Y(n_2157)
);

AOI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_2091),
.A2(n_1932),
.B1(n_1865),
.B2(n_1958),
.Y(n_2158)
);

INVx2_ASAP7_75t_SL g2159 ( 
.A(n_2078),
.Y(n_2159)
);

AND2x4_ASAP7_75t_L g2160 ( 
.A(n_2121),
.B(n_1974),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2030),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2048),
.Y(n_2162)
);

AOI22xp5_ASAP7_75t_L g2163 ( 
.A1(n_2037),
.A2(n_1930),
.B1(n_1964),
.B2(n_1982),
.Y(n_2163)
);

AND2x2_ASAP7_75t_SL g2164 ( 
.A(n_2148),
.B(n_1874),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_2055),
.A2(n_1933),
.B(n_1993),
.Y(n_2165)
);

OR2x2_ASAP7_75t_L g2166 ( 
.A(n_2051),
.B(n_2017),
.Y(n_2166)
);

INVx2_ASAP7_75t_L g2167 ( 
.A(n_2065),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_SL g2168 ( 
.A(n_2075),
.B(n_1893),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2087),
.B(n_2121),
.Y(n_2169)
);

NAND2xp33_ASAP7_75t_L g2170 ( 
.A(n_2092),
.B(n_2011),
.Y(n_2170)
);

OAI22xp5_ASAP7_75t_L g2171 ( 
.A1(n_2104),
.A2(n_1943),
.B1(n_2003),
.B2(n_1910),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_2048),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2102),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_2119),
.Y(n_2174)
);

BUFx6f_ASAP7_75t_SL g2175 ( 
.A(n_2115),
.Y(n_2175)
);

BUFx3_ASAP7_75t_L g2176 ( 
.A(n_2035),
.Y(n_2176)
);

NAND2x1p5_ASAP7_75t_L g2177 ( 
.A(n_2075),
.B(n_2020),
.Y(n_2177)
);

BUFx6f_ASAP7_75t_L g2178 ( 
.A(n_2135),
.Y(n_2178)
);

AOI21xp5_ASAP7_75t_SL g2179 ( 
.A1(n_2074),
.A2(n_1979),
.B(n_2015),
.Y(n_2179)
);

INVx1_ASAP7_75t_SL g2180 ( 
.A(n_2138),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2139),
.B(n_2022),
.Y(n_2181)
);

AND2x4_ASAP7_75t_L g2182 ( 
.A(n_2125),
.B(n_2020),
.Y(n_2182)
);

AOI222xp33_ASAP7_75t_L g2183 ( 
.A1(n_2088),
.A2(n_2047),
.B1(n_2127),
.B2(n_2133),
.C1(n_2130),
.C2(n_2039),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2109),
.B(n_2024),
.Y(n_2184)
);

NOR2xp67_ASAP7_75t_SL g2185 ( 
.A(n_2148),
.B(n_2020),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2109),
.B(n_1903),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2117),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2093),
.B(n_1893),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2122),
.Y(n_2189)
);

BUFx2_ASAP7_75t_L g2190 ( 
.A(n_2146),
.Y(n_2190)
);

INVxp67_ASAP7_75t_SL g2191 ( 
.A(n_2134),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_2134),
.Y(n_2192)
);

A2O1A1Ixp33_ASAP7_75t_L g2193 ( 
.A1(n_2082),
.A2(n_2016),
.B(n_1861),
.C(n_2000),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_2143),
.Y(n_2194)
);

INVx1_ASAP7_75t_L g2195 ( 
.A(n_2143),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2128),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_2136),
.B(n_1857),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2050),
.Y(n_2198)
);

AND2x2_ASAP7_75t_L g2199 ( 
.A(n_2108),
.B(n_1926),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_2120),
.A2(n_1985),
.B1(n_2028),
.B2(n_1987),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2062),
.Y(n_2201)
);

A2O1A1Ixp33_ASAP7_75t_L g2202 ( 
.A1(n_2100),
.A2(n_1983),
.B(n_2006),
.C(n_1892),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2084),
.A2(n_1999),
.B1(n_1995),
.B2(n_1991),
.Y(n_2203)
);

INVx2_ASAP7_75t_L g2204 ( 
.A(n_2062),
.Y(n_2204)
);

AND2x4_ASAP7_75t_L g2205 ( 
.A(n_2148),
.B(n_1926),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2060),
.B(n_159),
.Y(n_2206)
);

NAND2x1p5_ASAP7_75t_L g2207 ( 
.A(n_2095),
.B(n_2027),
.Y(n_2207)
);

INVx1_ASAP7_75t_L g2208 ( 
.A(n_2070),
.Y(n_2208)
);

INVx2_ASAP7_75t_SL g2209 ( 
.A(n_2036),
.Y(n_2209)
);

NAND2xp5_ASAP7_75t_L g2210 ( 
.A(n_2058),
.B(n_1907),
.Y(n_2210)
);

INVx2_ASAP7_75t_SL g2211 ( 
.A(n_2056),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2034),
.Y(n_2212)
);

OA21x2_ASAP7_75t_L g2213 ( 
.A1(n_2132),
.A2(n_1968),
.B(n_1955),
.Y(n_2213)
);

BUFx6f_ASAP7_75t_L g2214 ( 
.A(n_2044),
.Y(n_2214)
);

BUFx6f_ASAP7_75t_L g2215 ( 
.A(n_2044),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2080),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_2076),
.A2(n_1933),
.B(n_1993),
.Y(n_2217)
);

INVx1_ASAP7_75t_SL g2218 ( 
.A(n_2089),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2063),
.Y(n_2219)
);

AOI21xp5_ASAP7_75t_L g2220 ( 
.A1(n_2043),
.A2(n_1996),
.B(n_1998),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2053),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_SL g2222 ( 
.A(n_2031),
.B(n_2027),
.Y(n_2222)
);

INVx1_ASAP7_75t_SL g2223 ( 
.A(n_2056),
.Y(n_2223)
);

BUFx3_ASAP7_75t_L g2224 ( 
.A(n_2176),
.Y(n_2224)
);

BUFx2_ASAP7_75t_L g2225 ( 
.A(n_2190),
.Y(n_2225)
);

OR2x2_ASAP7_75t_L g2226 ( 
.A(n_2150),
.B(n_2072),
.Y(n_2226)
);

INVx2_ASAP7_75t_SL g2227 ( 
.A(n_2159),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2156),
.Y(n_2228)
);

OAI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2163),
.A2(n_2154),
.B1(n_2204),
.B2(n_2201),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2161),
.Y(n_2230)
);

AOI22xp33_ASAP7_75t_SL g2231 ( 
.A1(n_2170),
.A2(n_2040),
.B1(n_2052),
.B2(n_2081),
.Y(n_2231)
);

AOI22xp33_ASAP7_75t_SL g2232 ( 
.A1(n_2200),
.A2(n_2171),
.B1(n_2165),
.B2(n_2040),
.Y(n_2232)
);

INVx6_ASAP7_75t_L g2233 ( 
.A(n_2157),
.Y(n_2233)
);

AOI22xp33_ASAP7_75t_SL g2234 ( 
.A1(n_2200),
.A2(n_2171),
.B1(n_2213),
.B2(n_2203),
.Y(n_2234)
);

AOI22xp33_ASAP7_75t_L g2235 ( 
.A1(n_2183),
.A2(n_2158),
.B1(n_2163),
.B2(n_2118),
.Y(n_2235)
);

INVxp67_ASAP7_75t_L g2236 ( 
.A(n_2184),
.Y(n_2236)
);

OAI21xp33_ASAP7_75t_L g2237 ( 
.A1(n_2183),
.A2(n_2099),
.B(n_2090),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2162),
.Y(n_2238)
);

INVx6_ASAP7_75t_L g2239 ( 
.A(n_2157),
.Y(n_2239)
);

BUFx12f_ASAP7_75t_L g2240 ( 
.A(n_2157),
.Y(n_2240)
);

AOI22xp33_ASAP7_75t_L g2241 ( 
.A1(n_2203),
.A2(n_2105),
.B1(n_2149),
.B2(n_2137),
.Y(n_2241)
);

BUFx10_ASAP7_75t_L g2242 ( 
.A(n_2178),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_2189),
.Y(n_2243)
);

BUFx12f_ASAP7_75t_L g2244 ( 
.A(n_2178),
.Y(n_2244)
);

OAI22xp5_ASAP7_75t_SL g2245 ( 
.A1(n_2206),
.A2(n_2147),
.B1(n_2094),
.B2(n_2111),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_2167),
.Y(n_2246)
);

CKINVDCx20_ASAP7_75t_R g2247 ( 
.A(n_2153),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2172),
.Y(n_2248)
);

INVx6_ASAP7_75t_L g2249 ( 
.A(n_2178),
.Y(n_2249)
);

OAI21xp33_ASAP7_75t_SL g2250 ( 
.A1(n_2164),
.A2(n_2126),
.B(n_2106),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2192),
.Y(n_2251)
);

BUFx8_ASAP7_75t_L g2252 ( 
.A(n_2175),
.Y(n_2252)
);

INVx2_ASAP7_75t_L g2253 ( 
.A(n_2173),
.Y(n_2253)
);

AOI22xp33_ASAP7_75t_SL g2254 ( 
.A1(n_2213),
.A2(n_2059),
.B1(n_2066),
.B2(n_2145),
.Y(n_2254)
);

INVx2_ASAP7_75t_L g2255 ( 
.A(n_2187),
.Y(n_2255)
);

BUFx3_ASAP7_75t_L g2256 ( 
.A(n_2174),
.Y(n_2256)
);

INVx2_ASAP7_75t_L g2257 ( 
.A(n_2194),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2195),
.Y(n_2258)
);

INVx6_ASAP7_75t_L g2259 ( 
.A(n_2151),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2150),
.B(n_2116),
.Y(n_2260)
);

INVx1_ASAP7_75t_SL g2261 ( 
.A(n_2152),
.Y(n_2261)
);

BUFx3_ASAP7_75t_L g2262 ( 
.A(n_2174),
.Y(n_2262)
);

OAI22xp33_ASAP7_75t_L g2263 ( 
.A1(n_2207),
.A2(n_2057),
.B1(n_2067),
.B2(n_2131),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2196),
.Y(n_2264)
);

BUFx12f_ASAP7_75t_SL g2265 ( 
.A(n_2199),
.Y(n_2265)
);

CKINVDCx5p33_ASAP7_75t_R g2266 ( 
.A(n_2175),
.Y(n_2266)
);

INVx1_ASAP7_75t_L g2267 ( 
.A(n_2191),
.Y(n_2267)
);

OAI22xp33_ASAP7_75t_L g2268 ( 
.A1(n_2207),
.A2(n_2077),
.B1(n_2079),
.B2(n_2046),
.Y(n_2268)
);

OAI22xp5_ASAP7_75t_L g2269 ( 
.A1(n_2202),
.A2(n_2086),
.B1(n_2101),
.B2(n_2038),
.Y(n_2269)
);

AOI22xp33_ASAP7_75t_L g2270 ( 
.A1(n_2220),
.A2(n_2064),
.B1(n_2026),
.B2(n_2019),
.Y(n_2270)
);

AOI22xp33_ASAP7_75t_L g2271 ( 
.A1(n_2208),
.A2(n_2145),
.B1(n_1905),
.B2(n_1890),
.Y(n_2271)
);

AND2x2_ASAP7_75t_SL g2272 ( 
.A(n_2235),
.B(n_2151),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2225),
.B(n_2169),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_SL g2274 ( 
.A1(n_2235),
.A2(n_2209),
.B1(n_2181),
.B2(n_2198),
.Y(n_2274)
);

HB1xp67_ASAP7_75t_L g2275 ( 
.A(n_2251),
.Y(n_2275)
);

AND2x2_ASAP7_75t_L g2276 ( 
.A(n_2227),
.B(n_2180),
.Y(n_2276)
);

HB1xp67_ASAP7_75t_L g2277 ( 
.A(n_2251),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2257),
.Y(n_2278)
);

AOI21xp5_ASAP7_75t_L g2279 ( 
.A1(n_2269),
.A2(n_2179),
.B(n_2168),
.Y(n_2279)
);

INVx4_ASAP7_75t_L g2280 ( 
.A(n_2266),
.Y(n_2280)
);

A2O1A1Ixp33_ASAP7_75t_L g2281 ( 
.A1(n_2237),
.A2(n_2193),
.B(n_2096),
.C(n_2217),
.Y(n_2281)
);

HB1xp67_ASAP7_75t_L g2282 ( 
.A(n_2267),
.Y(n_2282)
);

NOR2xp67_ASAP7_75t_L g2283 ( 
.A(n_2250),
.B(n_2212),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2236),
.B(n_2216),
.Y(n_2284)
);

OAI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2231),
.A2(n_2186),
.B1(n_2180),
.B2(n_2210),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2261),
.B(n_2219),
.Y(n_2286)
);

A2O1A1Ixp33_ASAP7_75t_L g2287 ( 
.A1(n_2232),
.A2(n_2166),
.B(n_2221),
.C(n_2197),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2257),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2255),
.Y(n_2289)
);

OAI22xp5_ASAP7_75t_L g2290 ( 
.A1(n_2234),
.A2(n_2186),
.B1(n_2210),
.B2(n_2218),
.Y(n_2290)
);

OAI22xp5_ASAP7_75t_L g2291 ( 
.A1(n_2241),
.A2(n_2218),
.B1(n_2223),
.B2(n_2155),
.Y(n_2291)
);

OAI22xp5_ASAP7_75t_L g2292 ( 
.A1(n_2241),
.A2(n_2223),
.B1(n_2155),
.B2(n_2205),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2271),
.A2(n_2205),
.B1(n_2211),
.B2(n_2222),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_2256),
.B(n_2188),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2256),
.B(n_2182),
.Y(n_2295)
);

O2A1O1Ixp5_ASAP7_75t_L g2296 ( 
.A1(n_2229),
.A2(n_2182),
.B(n_2071),
.C(n_2129),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2262),
.B(n_2160),
.Y(n_2297)
);

INVx4_ASAP7_75t_SL g2298 ( 
.A(n_2274),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2290),
.B(n_2258),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2282),
.B(n_2260),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2275),
.Y(n_2301)
);

NAND2xp33_ASAP7_75t_R g2302 ( 
.A(n_2279),
.B(n_2226),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_SL g2303 ( 
.A1(n_2281),
.A2(n_2270),
.B(n_2229),
.Y(n_2303)
);

BUFx4f_ASAP7_75t_L g2304 ( 
.A(n_2272),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_L g2305 ( 
.A(n_2285),
.B(n_2228),
.Y(n_2305)
);

CKINVDCx16_ASAP7_75t_R g2306 ( 
.A(n_2280),
.Y(n_2306)
);

AND2x2_ASAP7_75t_L g2307 ( 
.A(n_2295),
.B(n_2262),
.Y(n_2307)
);

OAI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2303),
.A2(n_2287),
.B(n_2272),
.Y(n_2308)
);

HB1xp67_ASAP7_75t_L g2309 ( 
.A(n_2301),
.Y(n_2309)
);

INVx2_ASAP7_75t_L g2310 ( 
.A(n_2298),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2300),
.Y(n_2311)
);

OAI21xp5_ASAP7_75t_L g2312 ( 
.A1(n_2304),
.A2(n_2283),
.B(n_2296),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2299),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_2307),
.B(n_2294),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_2298),
.Y(n_2315)
);

BUFx2_ASAP7_75t_L g2316 ( 
.A(n_2310),
.Y(n_2316)
);

NOR2xp33_ASAP7_75t_L g2317 ( 
.A(n_2310),
.B(n_2306),
.Y(n_2317)
);

NAND2xp5_ASAP7_75t_L g2318 ( 
.A(n_2313),
.B(n_2305),
.Y(n_2318)
);

INVx1_ASAP7_75t_L g2319 ( 
.A(n_2309),
.Y(n_2319)
);

NOR2xp67_ASAP7_75t_L g2320 ( 
.A(n_2315),
.B(n_2280),
.Y(n_2320)
);

HB1xp67_ASAP7_75t_L g2321 ( 
.A(n_2313),
.Y(n_2321)
);

NAND2xp5_ASAP7_75t_L g2322 ( 
.A(n_2311),
.B(n_2277),
.Y(n_2322)
);

AND2x2_ASAP7_75t_L g2323 ( 
.A(n_2314),
.B(n_2276),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2314),
.B(n_2312),
.Y(n_2324)
);

NOR2xp33_ASAP7_75t_L g2325 ( 
.A(n_2315),
.B(n_2280),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_2319),
.Y(n_2326)
);

AND2x4_ASAP7_75t_SL g2327 ( 
.A(n_2317),
.B(n_2247),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2324),
.A2(n_2308),
.B1(n_2304),
.B2(n_2293),
.Y(n_2328)
);

AND2x2_ASAP7_75t_L g2329 ( 
.A(n_2323),
.B(n_2276),
.Y(n_2329)
);

OAI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2318),
.A2(n_2291),
.B1(n_2283),
.B2(n_2292),
.Y(n_2330)
);

AOI22xp33_ASAP7_75t_L g2331 ( 
.A1(n_2317),
.A2(n_2245),
.B1(n_2271),
.B2(n_2254),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_2316),
.Y(n_2332)
);

OAI221xp5_ASAP7_75t_SL g2333 ( 
.A1(n_2321),
.A2(n_2270),
.B1(n_2302),
.B2(n_2263),
.C(n_2268),
.Y(n_2333)
);

OAI22xp5_ASAP7_75t_L g2334 ( 
.A1(n_2321),
.A2(n_2263),
.B1(n_2224),
.B2(n_2284),
.Y(n_2334)
);

AOI22xp33_ASAP7_75t_L g2335 ( 
.A1(n_2325),
.A2(n_2268),
.B1(n_2286),
.B2(n_2255),
.Y(n_2335)
);

OAI221xp5_ASAP7_75t_L g2336 ( 
.A1(n_2320),
.A2(n_2289),
.B1(n_2288),
.B2(n_2278),
.C(n_2224),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2326),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2327),
.B(n_2322),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2332),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2329),
.Y(n_2340)
);

AND2x2_ASAP7_75t_L g2341 ( 
.A(n_2328),
.B(n_2273),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2335),
.B(n_2273),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_2330),
.Y(n_2343)
);

INVx2_ASAP7_75t_L g2344 ( 
.A(n_2334),
.Y(n_2344)
);

AND2x4_ASAP7_75t_L g2345 ( 
.A(n_2331),
.B(n_2297),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2338),
.Y(n_2346)
);

OR2x2_ASAP7_75t_L g2347 ( 
.A(n_2340),
.B(n_2333),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2340),
.B(n_2334),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2339),
.Y(n_2349)
);

INVx2_ASAP7_75t_L g2350 ( 
.A(n_2346),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2349),
.Y(n_2351)
);

OA21x2_ASAP7_75t_L g2352 ( 
.A1(n_2348),
.A2(n_2344),
.B(n_2343),
.Y(n_2352)
);

O2A1O1Ixp5_ASAP7_75t_L g2353 ( 
.A1(n_2347),
.A2(n_2344),
.B(n_2339),
.C(n_2337),
.Y(n_2353)
);

OAI211xp5_ASAP7_75t_SL g2354 ( 
.A1(n_2353),
.A2(n_2336),
.B(n_2341),
.C(n_2345),
.Y(n_2354)
);

INVx1_ASAP7_75t_L g2355 ( 
.A(n_2352),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2352),
.Y(n_2356)
);

AND2x4_ASAP7_75t_L g2357 ( 
.A(n_2350),
.B(n_2342),
.Y(n_2357)
);

INVx1_ASAP7_75t_L g2358 ( 
.A(n_2352),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2350),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2357),
.B(n_2351),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2355),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_2356),
.B(n_2351),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2358),
.Y(n_2363)
);

CKINVDCx16_ASAP7_75t_R g2364 ( 
.A(n_2359),
.Y(n_2364)
);

NAND2xp5_ASAP7_75t_L g2365 ( 
.A(n_2354),
.B(n_2345),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2357),
.B(n_2345),
.Y(n_2366)
);

INVx4_ASAP7_75t_L g2367 ( 
.A(n_2359),
.Y(n_2367)
);

INVxp67_ASAP7_75t_L g2368 ( 
.A(n_2357),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2357),
.B(n_2252),
.Y(n_2369)
);

OAI21xp33_ASAP7_75t_L g2370 ( 
.A1(n_2365),
.A2(n_2140),
.B(n_2073),
.Y(n_2370)
);

OR2x6_ASAP7_75t_L g2371 ( 
.A(n_2367),
.B(n_2240),
.Y(n_2371)
);

AOI21xp33_ASAP7_75t_L g2372 ( 
.A1(n_2367),
.A2(n_2362),
.B(n_2369),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_2366),
.B(n_2294),
.Y(n_2373)
);

INVx2_ASAP7_75t_L g2374 ( 
.A(n_2364),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2360),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2368),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2361),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2363),
.Y(n_2378)
);

INVxp67_ASAP7_75t_L g2379 ( 
.A(n_2369),
.Y(n_2379)
);

AOI22xp5_ASAP7_75t_L g2380 ( 
.A1(n_2364),
.A2(n_2252),
.B1(n_2244),
.B2(n_2233),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2364),
.B(n_2278),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2365),
.A2(n_2113),
.B(n_2295),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2374),
.Y(n_2383)
);

INVx1_ASAP7_75t_L g2384 ( 
.A(n_2377),
.Y(n_2384)
);

AOI211xp5_ASAP7_75t_L g2385 ( 
.A1(n_2372),
.A2(n_2009),
.B(n_2144),
.C(n_2297),
.Y(n_2385)
);

AOI21xp5_ASAP7_75t_L g2386 ( 
.A1(n_2371),
.A2(n_2144),
.B(n_160),
.Y(n_2386)
);

OR2x2_ASAP7_75t_L g2387 ( 
.A(n_2375),
.B(n_2230),
.Y(n_2387)
);

NOR2xp33_ASAP7_75t_R g2388 ( 
.A(n_2376),
.B(n_161),
.Y(n_2388)
);

INVxp67_ASAP7_75t_L g2389 ( 
.A(n_2371),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_2378),
.Y(n_2390)
);

AND2x2_ASAP7_75t_L g2391 ( 
.A(n_2373),
.B(n_2242),
.Y(n_2391)
);

NAND3xp33_ASAP7_75t_L g2392 ( 
.A(n_2379),
.B(n_2095),
.C(n_2041),
.Y(n_2392)
);

NAND2xp5_ASAP7_75t_L g2393 ( 
.A(n_2370),
.B(n_2288),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2380),
.B(n_2233),
.Y(n_2394)
);

CKINVDCx16_ASAP7_75t_R g2395 ( 
.A(n_2381),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_SL g2396 ( 
.A(n_2382),
.B(n_2242),
.Y(n_2396)
);

OAI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2374),
.A2(n_2233),
.B1(n_2249),
.B2(n_2239),
.Y(n_2397)
);

INVx1_ASAP7_75t_SL g2398 ( 
.A(n_2388),
.Y(n_2398)
);

AOI22xp33_ASAP7_75t_L g2399 ( 
.A1(n_2395),
.A2(n_2239),
.B1(n_2249),
.B2(n_2044),
.Y(n_2399)
);

AND2x2_ASAP7_75t_L g2400 ( 
.A(n_2383),
.B(n_2239),
.Y(n_2400)
);

INVx2_ASAP7_75t_L g2401 ( 
.A(n_2384),
.Y(n_2401)
);

INVx1_ASAP7_75t_SL g2402 ( 
.A(n_2390),
.Y(n_2402)
);

NOR2xp67_ASAP7_75t_SL g2403 ( 
.A(n_2386),
.B(n_2249),
.Y(n_2403)
);

AOI22xp33_ASAP7_75t_L g2404 ( 
.A1(n_2393),
.A2(n_2289),
.B1(n_2215),
.B2(n_2214),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2387),
.Y(n_2405)
);

INVx1_ASAP7_75t_SL g2406 ( 
.A(n_2391),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2389),
.Y(n_2407)
);

NOR3xp33_ASAP7_75t_SL g2408 ( 
.A(n_2396),
.B(n_161),
.C(n_162),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_L g2409 ( 
.A(n_2394),
.B(n_2097),
.Y(n_2409)
);

AOI221xp5_ASAP7_75t_L g2410 ( 
.A1(n_2385),
.A2(n_2032),
.B1(n_2248),
.B2(n_2238),
.C(n_164),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2397),
.B(n_2392),
.Y(n_2411)
);

OAI211xp5_ASAP7_75t_SL g2412 ( 
.A1(n_2402),
.A2(n_164),
.B(n_162),
.C(n_163),
.Y(n_2412)
);

NAND4xp25_ASAP7_75t_L g2413 ( 
.A(n_2401),
.B(n_2097),
.C(n_166),
.D(n_163),
.Y(n_2413)
);

INVx1_ASAP7_75t_L g2414 ( 
.A(n_2398),
.Y(n_2414)
);

NOR2xp33_ASAP7_75t_L g2415 ( 
.A(n_2398),
.B(n_165),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2405),
.A2(n_2259),
.B1(n_2185),
.B2(n_2107),
.Y(n_2416)
);

NAND3xp33_ASAP7_75t_SL g2417 ( 
.A(n_2407),
.B(n_2177),
.C(n_166),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2408),
.B(n_167),
.Y(n_2418)
);

NAND3xp33_ASAP7_75t_L g2419 ( 
.A(n_2400),
.B(n_167),
.C(n_168),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2406),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2403),
.B(n_169),
.Y(n_2421)
);

AOI22xp33_ASAP7_75t_L g2422 ( 
.A1(n_2411),
.A2(n_2215),
.B1(n_2214),
.B2(n_2243),
.Y(n_2422)
);

INVx1_ASAP7_75t_L g2423 ( 
.A(n_2410),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2409),
.B(n_169),
.Y(n_2424)
);

NAND2xp33_ASAP7_75t_L g2425 ( 
.A(n_2399),
.B(n_2214),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_L g2426 ( 
.A(n_2404),
.B(n_170),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2402),
.B(n_170),
.Y(n_2427)
);

NAND2xp5_ASAP7_75t_L g2428 ( 
.A(n_2402),
.B(n_171),
.Y(n_2428)
);

O2A1O1Ixp33_ASAP7_75t_SL g2429 ( 
.A1(n_2402),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2429)
);

AOI221x1_ASAP7_75t_L g2430 ( 
.A1(n_2407),
.A2(n_177),
.B1(n_174),
.B2(n_175),
.C(n_178),
.Y(n_2430)
);

OA22x2_ASAP7_75t_L g2431 ( 
.A1(n_2402),
.A2(n_2069),
.B1(n_2142),
.B2(n_2098),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2402),
.Y(n_2432)
);

NOR2xp33_ASAP7_75t_L g2433 ( 
.A(n_2402),
.B(n_174),
.Y(n_2433)
);

AOI21xp5_ASAP7_75t_L g2434 ( 
.A1(n_2429),
.A2(n_177),
.B(n_178),
.Y(n_2434)
);

NOR3xp33_ASAP7_75t_L g2435 ( 
.A(n_2432),
.B(n_179),
.C(n_180),
.Y(n_2435)
);

AOI211xp5_ASAP7_75t_L g2436 ( 
.A1(n_2433),
.A2(n_183),
.B(n_179),
.C(n_181),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2420),
.Y(n_2437)
);

CKINVDCx20_ASAP7_75t_L g2438 ( 
.A(n_2414),
.Y(n_2438)
);

NAND3xp33_ASAP7_75t_L g2439 ( 
.A(n_2415),
.B(n_181),
.C(n_183),
.Y(n_2439)
);

NAND2x1_ASAP7_75t_L g2440 ( 
.A(n_2427),
.B(n_2259),
.Y(n_2440)
);

HB1xp67_ASAP7_75t_L g2441 ( 
.A(n_2418),
.Y(n_2441)
);

NOR2xp33_ASAP7_75t_L g2442 ( 
.A(n_2412),
.B(n_184),
.Y(n_2442)
);

NOR4xp25_ASAP7_75t_L g2443 ( 
.A(n_2428),
.B(n_186),
.C(n_184),
.D(n_185),
.Y(n_2443)
);

NOR3xp33_ASAP7_75t_L g2444 ( 
.A(n_2421),
.B(n_185),
.C(n_186),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2413),
.B(n_187),
.Y(n_2445)
);

NAND2xp5_ASAP7_75t_L g2446 ( 
.A(n_2430),
.B(n_188),
.Y(n_2446)
);

NAND4xp25_ASAP7_75t_L g2447 ( 
.A(n_2424),
.B(n_191),
.C(n_188),
.D(n_189),
.Y(n_2447)
);

AND2x2_ASAP7_75t_L g2448 ( 
.A(n_2423),
.B(n_2259),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2419),
.B(n_189),
.Y(n_2449)
);

NAND2xp5_ASAP7_75t_L g2450 ( 
.A(n_2417),
.B(n_191),
.Y(n_2450)
);

AOI221xp5_ASAP7_75t_L g2451 ( 
.A1(n_2426),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_2451)
);

NOR2xp33_ASAP7_75t_L g2452 ( 
.A(n_2425),
.B(n_192),
.Y(n_2452)
);

NOR2xp33_ASAP7_75t_L g2453 ( 
.A(n_2422),
.B(n_193),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2416),
.B(n_194),
.Y(n_2454)
);

AOI21xp5_ASAP7_75t_L g2455 ( 
.A1(n_2431),
.A2(n_195),
.B(n_196),
.Y(n_2455)
);

NAND3xp33_ASAP7_75t_L g2456 ( 
.A(n_2432),
.B(n_196),
.C(n_197),
.Y(n_2456)
);

AND2x2_ASAP7_75t_L g2457 ( 
.A(n_2420),
.B(n_197),
.Y(n_2457)
);

AOI221xp5_ASAP7_75t_L g2458 ( 
.A1(n_2432),
.A2(n_200),
.B1(n_198),
.B2(n_199),
.C(n_201),
.Y(n_2458)
);

NAND4xp25_ASAP7_75t_SL g2459 ( 
.A(n_2420),
.B(n_200),
.C(n_198),
.D(n_199),
.Y(n_2459)
);

INVxp67_ASAP7_75t_L g2460 ( 
.A(n_2415),
.Y(n_2460)
);

NAND3xp33_ASAP7_75t_L g2461 ( 
.A(n_2432),
.B(n_201),
.C(n_202),
.Y(n_2461)
);

INVxp67_ASAP7_75t_L g2462 ( 
.A(n_2415),
.Y(n_2462)
);

O2A1O1Ixp5_ASAP7_75t_SL g2463 ( 
.A1(n_2420),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2429),
.Y(n_2464)
);

OAI21xp5_ASAP7_75t_L g2465 ( 
.A1(n_2427),
.A2(n_2103),
.B(n_2085),
.Y(n_2465)
);

NAND2xp5_ASAP7_75t_L g2466 ( 
.A(n_2430),
.B(n_203),
.Y(n_2466)
);

AO22x2_ASAP7_75t_L g2467 ( 
.A1(n_2432),
.A2(n_207),
.B1(n_205),
.B2(n_206),
.Y(n_2467)
);

INVxp67_ASAP7_75t_SL g2468 ( 
.A(n_2418),
.Y(n_2468)
);

NOR2xp33_ASAP7_75t_L g2469 ( 
.A(n_2412),
.B(n_205),
.Y(n_2469)
);

NAND4xp25_ASAP7_75t_L g2470 ( 
.A(n_2432),
.B(n_209),
.C(n_206),
.D(n_207),
.Y(n_2470)
);

AOI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2437),
.A2(n_211),
.B(n_209),
.C(n_210),
.Y(n_2471)
);

NOR3xp33_ASAP7_75t_L g2472 ( 
.A(n_2460),
.B(n_210),
.C(n_211),
.Y(n_2472)
);

NOR2xp33_ASAP7_75t_SL g2473 ( 
.A(n_2464),
.B(n_2470),
.Y(n_2473)
);

AOI21xp5_ASAP7_75t_L g2474 ( 
.A1(n_2434),
.A2(n_212),
.B(n_213),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2468),
.A2(n_2441),
.B1(n_2469),
.B2(n_2442),
.Y(n_2475)
);

OAI22xp5_ASAP7_75t_L g2476 ( 
.A1(n_2456),
.A2(n_2177),
.B1(n_2215),
.B2(n_2243),
.Y(n_2476)
);

NOR3xp33_ASAP7_75t_SL g2477 ( 
.A(n_2446),
.B(n_214),
.C(n_215),
.Y(n_2477)
);

NOR3xp33_ASAP7_75t_SL g2478 ( 
.A(n_2466),
.B(n_214),
.C(n_215),
.Y(n_2478)
);

AOI211xp5_ASAP7_75t_L g2479 ( 
.A1(n_2459),
.A2(n_218),
.B(n_216),
.C(n_217),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2443),
.B(n_2049),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2467),
.B(n_2049),
.Y(n_2481)
);

OA211x2_ASAP7_75t_L g2482 ( 
.A1(n_2458),
.A2(n_219),
.B(n_216),
.C(n_218),
.Y(n_2482)
);

NAND4xp25_ASAP7_75t_L g2483 ( 
.A(n_2452),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2483)
);

AND2x2_ASAP7_75t_L g2484 ( 
.A(n_2457),
.B(n_222),
.Y(n_2484)
);

NOR2x1_ASAP7_75t_L g2485 ( 
.A(n_2461),
.B(n_222),
.Y(n_2485)
);

AOI211xp5_ASAP7_75t_L g2486 ( 
.A1(n_2450),
.A2(n_225),
.B(n_223),
.C(n_224),
.Y(n_2486)
);

NOR4xp25_ASAP7_75t_L g2487 ( 
.A(n_2462),
.B(n_225),
.C(n_223),
.D(n_224),
.Y(n_2487)
);

NOR4xp75_ASAP7_75t_L g2488 ( 
.A(n_2454),
.B(n_229),
.C(n_226),
.D(n_227),
.Y(n_2488)
);

NAND2xp5_ASAP7_75t_L g2489 ( 
.A(n_2467),
.B(n_2049),
.Y(n_2489)
);

NOR3xp33_ASAP7_75t_L g2490 ( 
.A(n_2439),
.B(n_226),
.C(n_229),
.Y(n_2490)
);

INVx1_ASAP7_75t_L g2491 ( 
.A(n_2445),
.Y(n_2491)
);

NOR3xp33_ASAP7_75t_L g2492 ( 
.A(n_2435),
.B(n_230),
.C(n_231),
.Y(n_2492)
);

AOI222xp33_ASAP7_75t_L g2493 ( 
.A1(n_2453),
.A2(n_2448),
.B1(n_2449),
.B2(n_2451),
.C1(n_2465),
.C2(n_2438),
.Y(n_2493)
);

NOR2xp33_ASAP7_75t_L g2494 ( 
.A(n_2447),
.B(n_2440),
.Y(n_2494)
);

OAI211xp5_ASAP7_75t_L g2495 ( 
.A1(n_2436),
.A2(n_233),
.B(n_230),
.C(n_232),
.Y(n_2495)
);

NAND3xp33_ASAP7_75t_SL g2496 ( 
.A(n_2463),
.B(n_233),
.C(n_234),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2444),
.Y(n_2497)
);

AOI221xp5_ASAP7_75t_L g2498 ( 
.A1(n_2455),
.A2(n_237),
.B1(n_234),
.B2(n_235),
.C(n_238),
.Y(n_2498)
);

INVx2_ASAP7_75t_L g2499 ( 
.A(n_2467),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2434),
.A2(n_238),
.B(n_239),
.Y(n_2500)
);

OAI32xp33_ASAP7_75t_L g2501 ( 
.A1(n_2437),
.A2(n_242),
.A3(n_240),
.B1(n_241),
.B2(n_243),
.Y(n_2501)
);

OAI211xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2464),
.A2(n_243),
.B(n_241),
.C(n_242),
.Y(n_2502)
);

NAND4xp25_ASAP7_75t_L g2503 ( 
.A(n_2442),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2503)
);

NAND2xp5_ASAP7_75t_L g2504 ( 
.A(n_2464),
.B(n_2110),
.Y(n_2504)
);

NOR2xp33_ASAP7_75t_L g2505 ( 
.A(n_2464),
.B(n_244),
.Y(n_2505)
);

NAND2xp5_ASAP7_75t_L g2506 ( 
.A(n_2464),
.B(n_2110),
.Y(n_2506)
);

NOR2x1_ASAP7_75t_L g2507 ( 
.A(n_2437),
.B(n_246),
.Y(n_2507)
);

A2O1A1Ixp33_ASAP7_75t_SL g2508 ( 
.A1(n_2437),
.A2(n_249),
.B(n_247),
.C(n_248),
.Y(n_2508)
);

OAI21xp5_ASAP7_75t_L g2509 ( 
.A1(n_2474),
.A2(n_2083),
.B(n_2114),
.Y(n_2509)
);

AOI221xp5_ASAP7_75t_L g2510 ( 
.A1(n_2505),
.A2(n_252),
.B1(n_248),
.B2(n_251),
.C(n_253),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2499),
.B(n_251),
.Y(n_2511)
);

OA211x2_ASAP7_75t_L g2512 ( 
.A1(n_2473),
.A2(n_2498),
.B(n_2494),
.C(n_2496),
.Y(n_2512)
);

NOR2xp67_ASAP7_75t_SL g2513 ( 
.A(n_2491),
.B(n_253),
.Y(n_2513)
);

NOR2xp67_ASAP7_75t_L g2514 ( 
.A(n_2483),
.B(n_254),
.Y(n_2514)
);

NAND3xp33_ASAP7_75t_L g2515 ( 
.A(n_2507),
.B(n_254),
.C(n_255),
.Y(n_2515)
);

OAI221xp5_ASAP7_75t_L g2516 ( 
.A1(n_2508),
.A2(n_258),
.B1(n_255),
.B2(n_257),
.C(n_259),
.Y(n_2516)
);

NAND4xp25_ASAP7_75t_L g2517 ( 
.A(n_2475),
.B(n_262),
.C(n_260),
.D(n_261),
.Y(n_2517)
);

NAND3xp33_ASAP7_75t_SL g2518 ( 
.A(n_2486),
.B(n_2487),
.C(n_2478),
.Y(n_2518)
);

INVx1_ASAP7_75t_L g2519 ( 
.A(n_2484),
.Y(n_2519)
);

AND4x1_ASAP7_75t_L g2520 ( 
.A(n_2477),
.B(n_262),
.C(n_260),
.D(n_261),
.Y(n_2520)
);

NAND2xp5_ASAP7_75t_L g2521 ( 
.A(n_2500),
.B(n_263),
.Y(n_2521)
);

NAND3xp33_ASAP7_75t_L g2522 ( 
.A(n_2472),
.B(n_264),
.C(n_265),
.Y(n_2522)
);

AND2x2_ASAP7_75t_L g2523 ( 
.A(n_2479),
.B(n_264),
.Y(n_2523)
);

NAND4xp25_ASAP7_75t_L g2524 ( 
.A(n_2482),
.B(n_269),
.C(n_266),
.D(n_268),
.Y(n_2524)
);

NOR2x1_ASAP7_75t_L g2525 ( 
.A(n_2502),
.B(n_266),
.Y(n_2525)
);

NOR2x1_ASAP7_75t_L g2526 ( 
.A(n_2503),
.B(n_268),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2480),
.B(n_269),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2488),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2485),
.Y(n_2529)
);

NAND4xp75_ASAP7_75t_L g2530 ( 
.A(n_2497),
.B(n_274),
.C(n_270),
.D(n_273),
.Y(n_2530)
);

OR2x2_ASAP7_75t_L g2531 ( 
.A(n_2481),
.B(n_273),
.Y(n_2531)
);

NOR3x1_ASAP7_75t_L g2532 ( 
.A(n_2495),
.B(n_275),
.C(n_276),
.Y(n_2532)
);

NOR4xp75_ASAP7_75t_L g2533 ( 
.A(n_2504),
.B(n_278),
.C(n_275),
.D(n_277),
.Y(n_2533)
);

NAND4xp25_ASAP7_75t_L g2534 ( 
.A(n_2493),
.B(n_2492),
.C(n_2490),
.D(n_2471),
.Y(n_2534)
);

AOI211xp5_ASAP7_75t_L g2535 ( 
.A1(n_2501),
.A2(n_279),
.B(n_277),
.C(n_278),
.Y(n_2535)
);

O2A1O1Ixp33_ASAP7_75t_L g2536 ( 
.A1(n_2506),
.A2(n_281),
.B(n_279),
.C(n_280),
.Y(n_2536)
);

NAND5xp2_ASAP7_75t_L g2537 ( 
.A(n_2489),
.B(n_283),
.C(n_280),
.D(n_282),
.E(n_284),
.Y(n_2537)
);

AOI211xp5_ASAP7_75t_L g2538 ( 
.A1(n_2476),
.A2(n_284),
.B(n_282),
.C(n_283),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2499),
.B(n_285),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2499),
.B(n_285),
.Y(n_2540)
);

NOR2xp67_ASAP7_75t_L g2541 ( 
.A(n_2483),
.B(n_286),
.Y(n_2541)
);

NOR4xp75_ASAP7_75t_L g2542 ( 
.A(n_2496),
.B(n_288),
.C(n_286),
.D(n_287),
.Y(n_2542)
);

AOI211xp5_ASAP7_75t_L g2543 ( 
.A1(n_2505),
.A2(n_290),
.B(n_287),
.C(n_289),
.Y(n_2543)
);

NOR5xp2_ASAP7_75t_L g2544 ( 
.A(n_2502),
.B(n_291),
.C(n_289),
.D(n_290),
.E(n_292),
.Y(n_2544)
);

AOI221xp5_ASAP7_75t_L g2545 ( 
.A1(n_2505),
.A2(n_295),
.B1(n_291),
.B2(n_294),
.C(n_296),
.Y(n_2545)
);

NAND3xp33_ASAP7_75t_SL g2546 ( 
.A(n_2475),
.B(n_294),
.C(n_297),
.Y(n_2546)
);

AND2x4_ASAP7_75t_L g2547 ( 
.A(n_2507),
.B(n_298),
.Y(n_2547)
);

NAND4xp25_ASAP7_75t_SL g2548 ( 
.A(n_2493),
.B(n_300),
.C(n_298),
.D(n_299),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_SL g2549 ( 
.A(n_2484),
.B(n_2265),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_L g2550 ( 
.A(n_2499),
.B(n_299),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2473),
.B(n_300),
.C(n_301),
.Y(n_2551)
);

NOR2x1_ASAP7_75t_L g2552 ( 
.A(n_2505),
.B(n_301),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2487),
.B(n_302),
.Y(n_2553)
);

NOR3xp33_ASAP7_75t_L g2554 ( 
.A(n_2491),
.B(n_302),
.C(n_303),
.Y(n_2554)
);

AOI221xp5_ASAP7_75t_L g2555 ( 
.A1(n_2505),
.A2(n_305),
.B1(n_303),
.B2(n_304),
.C(n_306),
.Y(n_2555)
);

NOR3xp33_ASAP7_75t_L g2556 ( 
.A(n_2491),
.B(n_304),
.C(n_305),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_2484),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2507),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_2499),
.B(n_306),
.Y(n_2559)
);

OAI211xp5_ASAP7_75t_SL g2560 ( 
.A1(n_2475),
.A2(n_309),
.B(n_307),
.C(n_308),
.Y(n_2560)
);

NAND2xp5_ASAP7_75t_SL g2561 ( 
.A(n_2487),
.B(n_308),
.Y(n_2561)
);

AOI221x1_ASAP7_75t_L g2562 ( 
.A1(n_2505),
.A2(n_313),
.B1(n_310),
.B2(n_312),
.C(n_314),
.Y(n_2562)
);

NAND3xp33_ASAP7_75t_SL g2563 ( 
.A(n_2475),
.B(n_312),
.C(n_315),
.Y(n_2563)
);

NOR3xp33_ASAP7_75t_SL g2564 ( 
.A(n_2496),
.B(n_316),
.C(n_318),
.Y(n_2564)
);

AOI322xp5_ASAP7_75t_L g2565 ( 
.A1(n_2494),
.A2(n_2110),
.A3(n_2253),
.B1(n_2246),
.B2(n_2264),
.C1(n_2160),
.C2(n_322),
.Y(n_2565)
);

HB1xp67_ASAP7_75t_L g2566 ( 
.A(n_2488),
.Y(n_2566)
);

INVx1_ASAP7_75t_SL g2567 ( 
.A(n_2484),
.Y(n_2567)
);

NAND4xp25_ASAP7_75t_L g2568 ( 
.A(n_2473),
.B(n_319),
.C(n_316),
.D(n_318),
.Y(n_2568)
);

OAI22xp5_ASAP7_75t_L g2569 ( 
.A1(n_2505),
.A2(n_2042),
.B1(n_2246),
.B2(n_2264),
.Y(n_2569)
);

NAND3xp33_ASAP7_75t_SL g2570 ( 
.A(n_2475),
.B(n_319),
.C(n_320),
.Y(n_2570)
);

OAI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2515),
.A2(n_2124),
.B(n_2045),
.Y(n_2571)
);

OAI22xp5_ASAP7_75t_L g2572 ( 
.A1(n_2516),
.A2(n_2042),
.B1(n_322),
.B2(n_320),
.Y(n_2572)
);

NOR2x1_ASAP7_75t_L g2573 ( 
.A(n_2548),
.B(n_321),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_SL g2574 ( 
.A(n_2528),
.B(n_323),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2566),
.Y(n_2575)
);

AOI221xp5_ASAP7_75t_L g2576 ( 
.A1(n_2540),
.A2(n_325),
.B1(n_323),
.B2(n_324),
.C(n_326),
.Y(n_2576)
);

AND2x2_ASAP7_75t_SL g2577 ( 
.A(n_2544),
.B(n_325),
.Y(n_2577)
);

INVx1_ASAP7_75t_SL g2578 ( 
.A(n_2567),
.Y(n_2578)
);

AOI221x1_ASAP7_75t_L g2579 ( 
.A1(n_2550),
.A2(n_328),
.B1(n_326),
.B2(n_327),
.C(n_329),
.Y(n_2579)
);

OAI21xp33_ASAP7_75t_L g2580 ( 
.A1(n_2537),
.A2(n_328),
.B(n_330),
.Y(n_2580)
);

AO22x2_ASAP7_75t_L g2581 ( 
.A1(n_2558),
.A2(n_332),
.B1(n_330),
.B2(n_331),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2547),
.B(n_331),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2547),
.Y(n_2583)
);

OAI22xp33_ASAP7_75t_L g2584 ( 
.A1(n_2511),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2584)
);

AOI22x1_ASAP7_75t_L g2585 ( 
.A1(n_2529),
.A2(n_2523),
.B1(n_2557),
.B2(n_2519),
.Y(n_2585)
);

INVxp67_ASAP7_75t_L g2586 ( 
.A(n_2552),
.Y(n_2586)
);

A2O1A1Ixp33_ASAP7_75t_SL g2587 ( 
.A1(n_2559),
.A2(n_335),
.B(n_333),
.C(n_334),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_SL g2588 ( 
.A(n_2543),
.B(n_336),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2520),
.Y(n_2589)
);

NAND2xp33_ASAP7_75t_R g2590 ( 
.A(n_2564),
.B(n_336),
.Y(n_2590)
);

NOR3xp33_ASAP7_75t_L g2591 ( 
.A(n_2539),
.B(n_337),
.C(n_338),
.Y(n_2591)
);

INVx1_ASAP7_75t_SL g2592 ( 
.A(n_2542),
.Y(n_2592)
);

NAND2xp5_ASAP7_75t_L g2593 ( 
.A(n_2549),
.B(n_337),
.Y(n_2593)
);

A2O1A1Ixp33_ASAP7_75t_L g2594 ( 
.A1(n_2536),
.A2(n_340),
.B(n_338),
.C(n_339),
.Y(n_2594)
);

XNOR2x1_ASAP7_75t_L g2595 ( 
.A(n_2512),
.B(n_340),
.Y(n_2595)
);

INVx5_ASAP7_75t_L g2596 ( 
.A(n_2513),
.Y(n_2596)
);

AOI221xp5_ASAP7_75t_L g2597 ( 
.A1(n_2534),
.A2(n_343),
.B1(n_341),
.B2(n_342),
.C(n_344),
.Y(n_2597)
);

NAND4xp25_ASAP7_75t_L g2598 ( 
.A(n_2532),
.B(n_344),
.C(n_341),
.D(n_342),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2525),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_L g2600 ( 
.A(n_2514),
.B(n_345),
.Y(n_2600)
);

NOR2xp33_ASAP7_75t_R g2601 ( 
.A(n_2546),
.B(n_346),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2551),
.A2(n_348),
.B1(n_346),
.B2(n_347),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2553),
.Y(n_2603)
);

AOI221xp5_ASAP7_75t_L g2604 ( 
.A1(n_2563),
.A2(n_349),
.B1(n_347),
.B2(n_348),
.C(n_350),
.Y(n_2604)
);

OAI21xp5_ASAP7_75t_L g2605 ( 
.A1(n_2527),
.A2(n_2068),
.B(n_2123),
.Y(n_2605)
);

NAND2xp5_ASAP7_75t_L g2606 ( 
.A(n_2541),
.B(n_349),
.Y(n_2606)
);

AOI21xp5_ASAP7_75t_L g2607 ( 
.A1(n_2561),
.A2(n_350),
.B(n_351),
.Y(n_2607)
);

INVx1_ASAP7_75t_SL g2608 ( 
.A(n_2530),
.Y(n_2608)
);

AOI22xp5_ASAP7_75t_L g2609 ( 
.A1(n_2518),
.A2(n_2112),
.B1(n_354),
.B2(n_352),
.Y(n_2609)
);

INVx1_ASAP7_75t_SL g2610 ( 
.A(n_2521),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2533),
.Y(n_2611)
);

INVx1_ASAP7_75t_L g2612 ( 
.A(n_2526),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2524),
.Y(n_2613)
);

OAI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2535),
.A2(n_354),
.B1(n_352),
.B2(n_353),
.Y(n_2614)
);

INVx1_ASAP7_75t_SL g2615 ( 
.A(n_2531),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2562),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2554),
.B(n_353),
.Y(n_2617)
);

OAI221xp5_ASAP7_75t_L g2618 ( 
.A1(n_2538),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.C(n_358),
.Y(n_2618)
);

NOR2x1_ASAP7_75t_L g2619 ( 
.A(n_2568),
.B(n_356),
.Y(n_2619)
);

OR2x2_ASAP7_75t_L g2620 ( 
.A(n_2517),
.B(n_357),
.Y(n_2620)
);

NAND2xp5_ASAP7_75t_L g2621 ( 
.A(n_2556),
.B(n_358),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2522),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2570),
.Y(n_2623)
);

OAI21xp5_ASAP7_75t_SL g2624 ( 
.A1(n_2560),
.A2(n_359),
.B(n_360),
.Y(n_2624)
);

INVxp67_ASAP7_75t_L g2625 ( 
.A(n_2510),
.Y(n_2625)
);

INVx1_ASAP7_75t_L g2626 ( 
.A(n_2545),
.Y(n_2626)
);

NOR2xp33_ASAP7_75t_R g2627 ( 
.A(n_2555),
.B(n_359),
.Y(n_2627)
);

AND2x2_ASAP7_75t_L g2628 ( 
.A(n_2509),
.B(n_360),
.Y(n_2628)
);

AOI22xp5_ASAP7_75t_L g2629 ( 
.A1(n_2569),
.A2(n_363),
.B1(n_361),
.B2(n_362),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2565),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2566),
.Y(n_2631)
);

INVx1_ASAP7_75t_SL g2632 ( 
.A(n_2567),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_L g2633 ( 
.A(n_2547),
.B(n_361),
.Y(n_2633)
);

NAND2xp5_ASAP7_75t_SL g2634 ( 
.A(n_2528),
.B(n_362),
.Y(n_2634)
);

OAI22xp33_ASAP7_75t_SL g2635 ( 
.A1(n_2558),
.A2(n_365),
.B1(n_363),
.B2(n_364),
.Y(n_2635)
);

BUFx6f_ASAP7_75t_L g2636 ( 
.A(n_2511),
.Y(n_2636)
);

AOI322xp5_ASAP7_75t_L g2637 ( 
.A1(n_2566),
.A2(n_364),
.A3(n_365),
.B1(n_366),
.B2(n_367),
.C1(n_368),
.C2(n_369),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2577),
.B(n_366),
.Y(n_2638)
);

XNOR2xp5_ASAP7_75t_L g2639 ( 
.A(n_2595),
.B(n_2578),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2611),
.Y(n_2640)
);

OR2x2_ASAP7_75t_L g2641 ( 
.A(n_2632),
.B(n_367),
.Y(n_2641)
);

NOR2x1_ASAP7_75t_L g2642 ( 
.A(n_2575),
.B(n_368),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2596),
.B(n_369),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2616),
.Y(n_2644)
);

XNOR2x1_ASAP7_75t_L g2645 ( 
.A(n_2585),
.B(n_370),
.Y(n_2645)
);

INVx2_ASAP7_75t_L g2646 ( 
.A(n_2581),
.Y(n_2646)
);

NAND4xp75_ASAP7_75t_L g2647 ( 
.A(n_2631),
.B(n_373),
.C(n_371),
.D(n_372),
.Y(n_2647)
);

INVx1_ASAP7_75t_L g2648 ( 
.A(n_2582),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2596),
.B(n_372),
.Y(n_2649)
);

AOI22xp5_ASAP7_75t_L g2650 ( 
.A1(n_2613),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_2650)
);

AND2x2_ASAP7_75t_SL g2651 ( 
.A(n_2600),
.B(n_374),
.Y(n_2651)
);

NOR2x1_ASAP7_75t_SL g2652 ( 
.A(n_2574),
.B(n_2634),
.Y(n_2652)
);

NOR2xp67_ASAP7_75t_L g2653 ( 
.A(n_2598),
.B(n_376),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2633),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2583),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2596),
.Y(n_2656)
);

NOR2x1_ASAP7_75t_L g2657 ( 
.A(n_2603),
.B(n_376),
.Y(n_2657)
);

AND3x4_ASAP7_75t_L g2658 ( 
.A(n_2573),
.B(n_377),
.C(n_378),
.Y(n_2658)
);

AND2x2_ASAP7_75t_L g2659 ( 
.A(n_2592),
.B(n_377),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2581),
.Y(n_2660)
);

AOI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2590),
.A2(n_381),
.B1(n_379),
.B2(n_380),
.Y(n_2661)
);

HB1xp67_ASAP7_75t_L g2662 ( 
.A(n_2586),
.Y(n_2662)
);

NOR2x1_ASAP7_75t_L g2663 ( 
.A(n_2612),
.B(n_379),
.Y(n_2663)
);

NOR3xp33_ASAP7_75t_L g2664 ( 
.A(n_2615),
.B(n_380),
.C(n_381),
.Y(n_2664)
);

NAND4xp75_ASAP7_75t_L g2665 ( 
.A(n_2599),
.B(n_384),
.C(n_382),
.D(n_383),
.Y(n_2665)
);

NAND4xp75_ASAP7_75t_L g2666 ( 
.A(n_2606),
.B(n_385),
.C(n_383),
.D(n_384),
.Y(n_2666)
);

NAND4xp75_ASAP7_75t_L g2667 ( 
.A(n_2619),
.B(n_387),
.C(n_385),
.D(n_386),
.Y(n_2667)
);

OR2x2_ASAP7_75t_L g2668 ( 
.A(n_2589),
.B(n_386),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2580),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2636),
.Y(n_2670)
);

NAND4xp75_ASAP7_75t_L g2671 ( 
.A(n_2607),
.B(n_389),
.C(n_387),
.D(n_388),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2636),
.Y(n_2672)
);

NAND4xp75_ASAP7_75t_L g2673 ( 
.A(n_2579),
.B(n_2623),
.C(n_2593),
.D(n_2621),
.Y(n_2673)
);

NAND4xp75_ASAP7_75t_L g2674 ( 
.A(n_2617),
.B(n_393),
.C(n_390),
.D(n_392),
.Y(n_2674)
);

INVx2_ASAP7_75t_L g2675 ( 
.A(n_2620),
.Y(n_2675)
);

NOR3xp33_ASAP7_75t_L g2676 ( 
.A(n_2610),
.B(n_390),
.C(n_393),
.Y(n_2676)
);

OAI22x1_ASAP7_75t_L g2677 ( 
.A1(n_2608),
.A2(n_397),
.B1(n_395),
.B2(n_396),
.Y(n_2677)
);

INVx2_ASAP7_75t_L g2678 ( 
.A(n_2628),
.Y(n_2678)
);

NOR2xp33_ASAP7_75t_L g2679 ( 
.A(n_2624),
.B(n_395),
.Y(n_2679)
);

NOR2x1_ASAP7_75t_L g2680 ( 
.A(n_2584),
.B(n_396),
.Y(n_2680)
);

NAND4xp75_ASAP7_75t_L g2681 ( 
.A(n_2626),
.B(n_401),
.C(n_399),
.D(n_400),
.Y(n_2681)
);

NOR2x1_ASAP7_75t_L g2682 ( 
.A(n_2622),
.B(n_399),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2635),
.Y(n_2683)
);

NOR3xp33_ASAP7_75t_L g2684 ( 
.A(n_2591),
.B(n_400),
.C(n_401),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2588),
.Y(n_2685)
);

XNOR2xp5_ASAP7_75t_L g2686 ( 
.A(n_2614),
.B(n_402),
.Y(n_2686)
);

INVx2_ASAP7_75t_L g2687 ( 
.A(n_2630),
.Y(n_2687)
);

XOR2xp5_ASAP7_75t_L g2688 ( 
.A(n_2602),
.B(n_402),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_L g2689 ( 
.A(n_2587),
.B(n_403),
.Y(n_2689)
);

INVx2_ASAP7_75t_SL g2690 ( 
.A(n_2601),
.Y(n_2690)
);

NAND4xp75_ASAP7_75t_L g2691 ( 
.A(n_2604),
.B(n_405),
.C(n_403),
.D(n_404),
.Y(n_2691)
);

INVxp67_ASAP7_75t_L g2692 ( 
.A(n_2618),
.Y(n_2692)
);

NOR2x1_ASAP7_75t_L g2693 ( 
.A(n_2594),
.B(n_404),
.Y(n_2693)
);

NAND2x1p5_ASAP7_75t_L g2694 ( 
.A(n_2629),
.B(n_405),
.Y(n_2694)
);

HB1xp67_ASAP7_75t_L g2695 ( 
.A(n_2627),
.Y(n_2695)
);

AND2x4_ASAP7_75t_L g2696 ( 
.A(n_2625),
.B(n_2609),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2572),
.Y(n_2697)
);

XNOR2xp5_ASAP7_75t_L g2698 ( 
.A(n_2576),
.B(n_406),
.Y(n_2698)
);

HB1xp67_ASAP7_75t_L g2699 ( 
.A(n_2597),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2571),
.A2(n_408),
.B1(n_406),
.B2(n_407),
.Y(n_2700)
);

XOR2xp5_ASAP7_75t_L g2701 ( 
.A(n_2639),
.B(n_2637),
.Y(n_2701)
);

NOR4xp25_ASAP7_75t_L g2702 ( 
.A(n_2656),
.B(n_2605),
.C(n_409),
.D(n_407),
.Y(n_2702)
);

XNOR2x1_ASAP7_75t_L g2703 ( 
.A(n_2662),
.B(n_408),
.Y(n_2703)
);

NAND2xp5_ASAP7_75t_L g2704 ( 
.A(n_2660),
.B(n_2646),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2644),
.B(n_409),
.Y(n_2705)
);

AND3x4_ASAP7_75t_L g2706 ( 
.A(n_2653),
.B(n_410),
.C(n_412),
.Y(n_2706)
);

INVx3_ASAP7_75t_L g2707 ( 
.A(n_2658),
.Y(n_2707)
);

NOR2x1_ASAP7_75t_L g2708 ( 
.A(n_2643),
.B(n_410),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_L g2709 ( 
.A(n_2640),
.B(n_413),
.Y(n_2709)
);

NOR5xp2_ASAP7_75t_L g2710 ( 
.A(n_2699),
.B(n_414),
.C(n_415),
.D(n_416),
.E(n_417),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_SL g2711 ( 
.A(n_2638),
.B(n_2687),
.Y(n_2711)
);

OR2x2_ASAP7_75t_L g2712 ( 
.A(n_2649),
.B(n_414),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2663),
.Y(n_2713)
);

NOR3xp33_ASAP7_75t_SL g2714 ( 
.A(n_2655),
.B(n_415),
.C(n_416),
.Y(n_2714)
);

OAI211xp5_ASAP7_75t_SL g2715 ( 
.A1(n_2670),
.A2(n_2672),
.B(n_2683),
.C(n_2654),
.Y(n_2715)
);

XNOR2xp5_ASAP7_75t_L g2716 ( 
.A(n_2645),
.B(n_418),
.Y(n_2716)
);

NAND4xp75_ASAP7_75t_L g2717 ( 
.A(n_2642),
.B(n_421),
.C(n_419),
.D(n_420),
.Y(n_2717)
);

NOR2x1_ASAP7_75t_L g2718 ( 
.A(n_2641),
.B(n_2673),
.Y(n_2718)
);

BUFx2_ASAP7_75t_L g2719 ( 
.A(n_2657),
.Y(n_2719)
);

NOR3xp33_ASAP7_75t_L g2720 ( 
.A(n_2648),
.B(n_419),
.C(n_420),
.Y(n_2720)
);

AOI32xp33_ASAP7_75t_L g2721 ( 
.A1(n_2679),
.A2(n_421),
.A3(n_423),
.B1(n_424),
.B2(n_425),
.Y(n_2721)
);

INVx1_ASAP7_75t_L g2722 ( 
.A(n_2682),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2689),
.Y(n_2723)
);

NAND4xp75_ASAP7_75t_L g2724 ( 
.A(n_2651),
.B(n_423),
.C(n_424),
.D(n_426),
.Y(n_2724)
);

AND2x4_ASAP7_75t_L g2725 ( 
.A(n_2652),
.B(n_427),
.Y(n_2725)
);

INVx1_ASAP7_75t_SL g2726 ( 
.A(n_2668),
.Y(n_2726)
);

NAND2xp5_ASAP7_75t_SL g2727 ( 
.A(n_2661),
.B(n_427),
.Y(n_2727)
);

AND2x2_ASAP7_75t_L g2728 ( 
.A(n_2652),
.B(n_428),
.Y(n_2728)
);

NAND5xp2_ASAP7_75t_L g2729 ( 
.A(n_2694),
.B(n_2669),
.C(n_2685),
.D(n_2697),
.E(n_2684),
.Y(n_2729)
);

NAND4xp25_ASAP7_75t_L g2730 ( 
.A(n_2664),
.B(n_428),
.C(n_429),
.D(n_430),
.Y(n_2730)
);

NOR5xp2_ASAP7_75t_L g2731 ( 
.A(n_2692),
.B(n_429),
.C(n_430),
.D(n_431),
.E(n_432),
.Y(n_2731)
);

NOR2xp33_ASAP7_75t_L g2732 ( 
.A(n_2690),
.B(n_431),
.Y(n_2732)
);

AOI211x1_ASAP7_75t_L g2733 ( 
.A1(n_2659),
.A2(n_432),
.B(n_433),
.C(n_435),
.Y(n_2733)
);

NOR3xp33_ASAP7_75t_L g2734 ( 
.A(n_2675),
.B(n_435),
.C(n_437),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2667),
.Y(n_2735)
);

AOI21xp5_ASAP7_75t_L g2736 ( 
.A1(n_2677),
.A2(n_437),
.B(n_438),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2678),
.B(n_438),
.Y(n_2737)
);

NOR4xp25_ASAP7_75t_L g2738 ( 
.A(n_2695),
.B(n_439),
.C(n_440),
.D(n_441),
.Y(n_2738)
);

NOR3xp33_ASAP7_75t_L g2739 ( 
.A(n_2696),
.B(n_439),
.C(n_440),
.Y(n_2739)
);

O2A1O1Ixp33_ASAP7_75t_L g2740 ( 
.A1(n_2696),
.A2(n_441),
.B(n_442),
.C(n_444),
.Y(n_2740)
);

HB1xp67_ASAP7_75t_L g2741 ( 
.A(n_2666),
.Y(n_2741)
);

NOR3xp33_ASAP7_75t_L g2742 ( 
.A(n_2676),
.B(n_442),
.C(n_444),
.Y(n_2742)
);

OAI211xp5_ASAP7_75t_SL g2743 ( 
.A1(n_2680),
.A2(n_445),
.B(n_446),
.C(n_447),
.Y(n_2743)
);

NAND4xp75_ASAP7_75t_L g2744 ( 
.A(n_2693),
.B(n_2700),
.C(n_2650),
.D(n_2674),
.Y(n_2744)
);

NAND5xp2_ASAP7_75t_L g2745 ( 
.A(n_2686),
.B(n_446),
.C(n_447),
.D(n_448),
.E(n_449),
.Y(n_2745)
);

NAND2xp33_ASAP7_75t_SL g2746 ( 
.A(n_2714),
.B(n_2698),
.Y(n_2746)
);

INVx1_ASAP7_75t_L g2747 ( 
.A(n_2719),
.Y(n_2747)
);

AOI322xp5_ASAP7_75t_L g2748 ( 
.A1(n_2718),
.A2(n_2688),
.A3(n_2671),
.B1(n_2691),
.B2(n_2681),
.C1(n_2647),
.C2(n_2665),
.Y(n_2748)
);

AOI22xp5_ASAP7_75t_L g2749 ( 
.A1(n_2715),
.A2(n_2704),
.B1(n_2707),
.B2(n_2711),
.Y(n_2749)
);

CKINVDCx5p33_ASAP7_75t_R g2750 ( 
.A(n_2726),
.Y(n_2750)
);

INVx2_ASAP7_75t_SL g2751 ( 
.A(n_2708),
.Y(n_2751)
);

INVx1_ASAP7_75t_SL g2752 ( 
.A(n_2728),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2707),
.B(n_448),
.Y(n_2753)
);

CKINVDCx5p33_ASAP7_75t_R g2754 ( 
.A(n_2723),
.Y(n_2754)
);

NOR2xp33_ASAP7_75t_R g2755 ( 
.A(n_2716),
.B(n_450),
.Y(n_2755)
);

NAND2xp5_ASAP7_75t_L g2756 ( 
.A(n_2713),
.B(n_450),
.Y(n_2756)
);

CKINVDCx20_ASAP7_75t_R g2757 ( 
.A(n_2701),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2725),
.Y(n_2758)
);

CKINVDCx5p33_ASAP7_75t_R g2759 ( 
.A(n_2722),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2725),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2706),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2703),
.Y(n_2762)
);

HB1xp67_ASAP7_75t_L g2763 ( 
.A(n_2712),
.Y(n_2763)
);

AND2x4_ASAP7_75t_L g2764 ( 
.A(n_2735),
.B(n_451),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_2741),
.Y(n_2765)
);

INVx1_ASAP7_75t_SL g2766 ( 
.A(n_2705),
.Y(n_2766)
);

CKINVDCx16_ASAP7_75t_R g2767 ( 
.A(n_2737),
.Y(n_2767)
);

CKINVDCx16_ASAP7_75t_R g2768 ( 
.A(n_2709),
.Y(n_2768)
);

INVx1_ASAP7_75t_SL g2769 ( 
.A(n_2724),
.Y(n_2769)
);

BUFx2_ASAP7_75t_L g2770 ( 
.A(n_2717),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2738),
.B(n_451),
.Y(n_2771)
);

CKINVDCx5p33_ASAP7_75t_R g2772 ( 
.A(n_2727),
.Y(n_2772)
);

INVx1_ASAP7_75t_L g2773 ( 
.A(n_2733),
.Y(n_2773)
);

CKINVDCx5p33_ASAP7_75t_R g2774 ( 
.A(n_2732),
.Y(n_2774)
);

CKINVDCx5p33_ASAP7_75t_R g2775 ( 
.A(n_2736),
.Y(n_2775)
);

AND2x2_ASAP7_75t_L g2776 ( 
.A(n_2734),
.B(n_452),
.Y(n_2776)
);

NOR2x1p5_ASAP7_75t_L g2777 ( 
.A(n_2744),
.B(n_452),
.Y(n_2777)
);

AND3x4_ASAP7_75t_L g2778 ( 
.A(n_2742),
.B(n_453),
.C(n_454),
.Y(n_2778)
);

HB1xp67_ASAP7_75t_L g2779 ( 
.A(n_2730),
.Y(n_2779)
);

INVx1_ASAP7_75t_SL g2780 ( 
.A(n_2729),
.Y(n_2780)
);

OAI211xp5_ASAP7_75t_L g2781 ( 
.A1(n_2749),
.A2(n_2721),
.B(n_2702),
.C(n_2740),
.Y(n_2781)
);

OAI22xp5_ASAP7_75t_L g2782 ( 
.A1(n_2757),
.A2(n_2720),
.B1(n_2739),
.B2(n_2745),
.Y(n_2782)
);

AOI22xp5_ASAP7_75t_L g2783 ( 
.A1(n_2750),
.A2(n_2743),
.B1(n_2731),
.B2(n_2710),
.Y(n_2783)
);

AOI32xp33_ASAP7_75t_L g2784 ( 
.A1(n_2780),
.A2(n_453),
.A3(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_2784)
);

INVx1_ASAP7_75t_L g2785 ( 
.A(n_2763),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2758),
.Y(n_2786)
);

O2A1O1Ixp33_ASAP7_75t_L g2787 ( 
.A1(n_2747),
.A2(n_455),
.B(n_458),
.C(n_459),
.Y(n_2787)
);

AOI221xp5_ASAP7_75t_L g2788 ( 
.A1(n_2765),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.C(n_463),
.Y(n_2788)
);

OAI221xp5_ASAP7_75t_L g2789 ( 
.A1(n_2752),
.A2(n_460),
.B1(n_462),
.B2(n_464),
.C(n_465),
.Y(n_2789)
);

HB1xp67_ASAP7_75t_L g2790 ( 
.A(n_2760),
.Y(n_2790)
);

AOI322xp5_ASAP7_75t_L g2791 ( 
.A1(n_2751),
.A2(n_464),
.A3(n_465),
.B1(n_466),
.B2(n_467),
.C1(n_468),
.C2(n_469),
.Y(n_2791)
);

OAI211xp5_ASAP7_75t_L g2792 ( 
.A1(n_2759),
.A2(n_467),
.B(n_468),
.C(n_469),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2768),
.B(n_470),
.Y(n_2793)
);

O2A1O1Ixp33_ASAP7_75t_L g2794 ( 
.A1(n_2761),
.A2(n_470),
.B(n_471),
.C(n_474),
.Y(n_2794)
);

AOI322xp5_ASAP7_75t_L g2795 ( 
.A1(n_2746),
.A2(n_471),
.A3(n_475),
.B1(n_476),
.B2(n_477),
.C1(n_478),
.C2(n_479),
.Y(n_2795)
);

OAI211xp5_ASAP7_75t_SL g2796 ( 
.A1(n_2766),
.A2(n_476),
.B(n_478),
.C(n_479),
.Y(n_2796)
);

OAI211xp5_ASAP7_75t_L g2797 ( 
.A1(n_2754),
.A2(n_480),
.B(n_481),
.C(n_482),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2773),
.Y(n_2798)
);

OAI221xp5_ASAP7_75t_L g2799 ( 
.A1(n_2769),
.A2(n_480),
.B1(n_482),
.B2(n_484),
.C(n_485),
.Y(n_2799)
);

AOI322xp5_ASAP7_75t_L g2800 ( 
.A1(n_2771),
.A2(n_484),
.A3(n_485),
.B1(n_486),
.B2(n_487),
.C1(n_488),
.C2(n_489),
.Y(n_2800)
);

AOI221xp5_ASAP7_75t_SL g2801 ( 
.A1(n_2762),
.A2(n_486),
.B1(n_487),
.B2(n_488),
.C(n_489),
.Y(n_2801)
);

AOI322xp5_ASAP7_75t_L g2802 ( 
.A1(n_2767),
.A2(n_490),
.A3(n_491),
.B1(n_492),
.B2(n_493),
.C1(n_494),
.C2(n_495),
.Y(n_2802)
);

OAI322xp33_ASAP7_75t_L g2803 ( 
.A1(n_2775),
.A2(n_491),
.A3(n_492),
.B1(n_493),
.B2(n_494),
.C1(n_495),
.C2(n_496),
.Y(n_2803)
);

INVx2_ASAP7_75t_L g2804 ( 
.A(n_2777),
.Y(n_2804)
);

OAI22xp5_ASAP7_75t_L g2805 ( 
.A1(n_2779),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2805)
);

OAI211xp5_ASAP7_75t_L g2806 ( 
.A1(n_2755),
.A2(n_498),
.B(n_499),
.C(n_500),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2790),
.Y(n_2807)
);

AOI22xp5_ASAP7_75t_L g2808 ( 
.A1(n_2785),
.A2(n_2774),
.B1(n_2770),
.B2(n_2778),
.Y(n_2808)
);

BUFx2_ASAP7_75t_L g2809 ( 
.A(n_2798),
.Y(n_2809)
);

AOI22xp33_ASAP7_75t_L g2810 ( 
.A1(n_2786),
.A2(n_2772),
.B1(n_2776),
.B2(n_2753),
.Y(n_2810)
);

AOI22xp5_ASAP7_75t_L g2811 ( 
.A1(n_2783),
.A2(n_2756),
.B1(n_2764),
.B2(n_2748),
.Y(n_2811)
);

INVx2_ASAP7_75t_L g2812 ( 
.A(n_2804),
.Y(n_2812)
);

AOI31xp33_ASAP7_75t_L g2813 ( 
.A1(n_2782),
.A2(n_2764),
.A3(n_501),
.B(n_502),
.Y(n_2813)
);

AO22x2_ASAP7_75t_SL g2814 ( 
.A1(n_2781),
.A2(n_499),
.B1(n_501),
.B2(n_502),
.Y(n_2814)
);

AOI31xp33_ASAP7_75t_L g2815 ( 
.A1(n_2806),
.A2(n_503),
.A3(n_504),
.B(n_505),
.Y(n_2815)
);

NAND4xp75_ASAP7_75t_L g2816 ( 
.A(n_2801),
.B(n_503),
.C(n_504),
.D(n_507),
.Y(n_2816)
);

OAI22xp5_ASAP7_75t_SL g2817 ( 
.A1(n_2793),
.A2(n_507),
.B1(n_508),
.B2(n_509),
.Y(n_2817)
);

OA22x2_ASAP7_75t_L g2818 ( 
.A1(n_2792),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.Y(n_2818)
);

OAI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2789),
.A2(n_510),
.B1(n_511),
.B2(n_512),
.Y(n_2819)
);

AO22x2_ASAP7_75t_L g2820 ( 
.A1(n_2805),
.A2(n_511),
.B1(n_512),
.B2(n_513),
.Y(n_2820)
);

INVx1_ASAP7_75t_SL g2821 ( 
.A(n_2800),
.Y(n_2821)
);

AOI22xp5_ASAP7_75t_L g2822 ( 
.A1(n_2796),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_2822)
);

AOI22xp5_ASAP7_75t_L g2823 ( 
.A1(n_2797),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_2823)
);

NAND5xp2_ASAP7_75t_L g2824 ( 
.A(n_2807),
.B(n_2784),
.C(n_2787),
.D(n_2794),
.E(n_2788),
.Y(n_2824)
);

OA22x2_ASAP7_75t_L g2825 ( 
.A1(n_2809),
.A2(n_2799),
.B1(n_2803),
.B2(n_2795),
.Y(n_2825)
);

AOI221xp5_ASAP7_75t_L g2826 ( 
.A1(n_2813),
.A2(n_2802),
.B1(n_2791),
.B2(n_519),
.C(n_520),
.Y(n_2826)
);

INVx2_ASAP7_75t_L g2827 ( 
.A(n_2812),
.Y(n_2827)
);

AOI22xp5_ASAP7_75t_L g2828 ( 
.A1(n_2808),
.A2(n_517),
.B1(n_518),
.B2(n_519),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_L g2829 ( 
.A(n_2811),
.B(n_517),
.Y(n_2829)
);

NOR3xp33_ASAP7_75t_L g2830 ( 
.A(n_2821),
.B(n_518),
.C(n_520),
.Y(n_2830)
);

NAND3xp33_ASAP7_75t_L g2831 ( 
.A(n_2810),
.B(n_2823),
.C(n_2815),
.Y(n_2831)
);

NAND3xp33_ASAP7_75t_L g2832 ( 
.A(n_2819),
.B(n_2822),
.C(n_2814),
.Y(n_2832)
);

OR3x1_ASAP7_75t_L g2833 ( 
.A(n_2818),
.B(n_521),
.C(n_522),
.Y(n_2833)
);

AND3x2_ASAP7_75t_L g2834 ( 
.A(n_2817),
.B(n_521),
.C(n_523),
.Y(n_2834)
);

AOI221xp5_ASAP7_75t_L g2835 ( 
.A1(n_2820),
.A2(n_524),
.B1(n_525),
.B2(n_526),
.C(n_527),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_SL g2836 ( 
.A1(n_2827),
.A2(n_2816),
.B(n_526),
.Y(n_2836)
);

NAND3xp33_ASAP7_75t_L g2837 ( 
.A(n_2831),
.B(n_525),
.C(n_527),
.Y(n_2837)
);

OAI22xp5_ASAP7_75t_SL g2838 ( 
.A1(n_2833),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_2838)
);

AO21x2_ASAP7_75t_L g2839 ( 
.A1(n_2829),
.A2(n_528),
.B(n_529),
.Y(n_2839)
);

XNOR2xp5_ASAP7_75t_L g2840 ( 
.A(n_2825),
.B(n_530),
.Y(n_2840)
);

AOI221xp5_ASAP7_75t_L g2841 ( 
.A1(n_2830),
.A2(n_531),
.B1(n_532),
.B2(n_533),
.C(n_534),
.Y(n_2841)
);

AOI22xp5_ASAP7_75t_L g2842 ( 
.A1(n_2835),
.A2(n_533),
.B1(n_534),
.B2(n_535),
.Y(n_2842)
);

OAI21xp5_ASAP7_75t_SL g2843 ( 
.A1(n_2840),
.A2(n_2832),
.B(n_2834),
.Y(n_2843)
);

OAI22xp5_ASAP7_75t_L g2844 ( 
.A1(n_2838),
.A2(n_2828),
.B1(n_2826),
.B2(n_2824),
.Y(n_2844)
);

XNOR2x1_ASAP7_75t_L g2845 ( 
.A(n_2842),
.B(n_2837),
.Y(n_2845)
);

OAI22xp5_ASAP7_75t_L g2846 ( 
.A1(n_2836),
.A2(n_535),
.B1(n_536),
.B2(n_537),
.Y(n_2846)
);

INVxp67_ASAP7_75t_L g2847 ( 
.A(n_2839),
.Y(n_2847)
);

OAI22xp5_ASAP7_75t_L g2848 ( 
.A1(n_2841),
.A2(n_537),
.B1(n_538),
.B2(n_539),
.Y(n_2848)
);

AOI22xp5_ASAP7_75t_L g2849 ( 
.A1(n_2847),
.A2(n_539),
.B1(n_540),
.B2(n_541),
.Y(n_2849)
);

OAI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2843),
.A2(n_540),
.B(n_541),
.Y(n_2850)
);

OAI21xp33_ASAP7_75t_L g2851 ( 
.A1(n_2845),
.A2(n_542),
.B(n_543),
.Y(n_2851)
);

NOR2xp33_ASAP7_75t_R g2852 ( 
.A(n_2850),
.B(n_2844),
.Y(n_2852)
);

OA21x2_ASAP7_75t_L g2853 ( 
.A1(n_2851),
.A2(n_2846),
.B(n_2848),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2849),
.B(n_542),
.Y(n_2854)
);

AOI21xp5_ASAP7_75t_L g2855 ( 
.A1(n_2854),
.A2(n_545),
.B(n_546),
.Y(n_2855)
);

AOI22xp5_ASAP7_75t_SL g2856 ( 
.A1(n_2853),
.A2(n_545),
.B1(n_546),
.B2(n_547),
.Y(n_2856)
);

OA21x2_ASAP7_75t_L g2857 ( 
.A1(n_2855),
.A2(n_2852),
.B(n_549),
.Y(n_2857)
);

XNOR2xp5_ASAP7_75t_L g2858 ( 
.A(n_2857),
.B(n_2856),
.Y(n_2858)
);

AOI221xp5_ASAP7_75t_L g2859 ( 
.A1(n_2858),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.C(n_551),
.Y(n_2859)
);

AOI22xp5_ASAP7_75t_L g2860 ( 
.A1(n_2859),
.A2(n_548),
.B1(n_552),
.B2(n_553),
.Y(n_2860)
);

AOI211xp5_ASAP7_75t_L g2861 ( 
.A1(n_2860),
.A2(n_552),
.B(n_553),
.C(n_554),
.Y(n_2861)
);


endmodule