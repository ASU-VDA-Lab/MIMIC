module fake_jpeg_25051_n_330 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_330);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_330;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_14),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_14),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_43),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_7),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_39),
.B(n_26),
.Y(n_61)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_24),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_44),
.Y(n_56)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_49),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_20),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_53),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_46),
.A2(n_20),
.B1(n_25),
.B2(n_23),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_52),
.A2(n_48),
.B1(n_29),
.B2(n_30),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_31),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_45),
.A2(n_32),
.B1(n_29),
.B2(n_33),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_32),
.B1(n_31),
.B2(n_33),
.Y(n_77)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_57),
.B(n_61),
.Y(n_83)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_38),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_65),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_34),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g109 ( 
.A(n_66),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_46),
.B(n_25),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_23),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_22),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g75 ( 
.A(n_59),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_75),
.B(n_76),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_50),
.B(n_43),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_77),
.A2(n_101),
.B1(n_89),
.B2(n_67),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_78),
.A2(n_89),
.B1(n_91),
.B2(n_72),
.Y(n_127)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_41),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_79),
.B(n_90),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_45),
.Y(n_80)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_80),
.A2(n_104),
.B(n_106),
.C(n_79),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_84),
.B(n_85),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_63),
.B(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_65),
.B(n_16),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_86),
.B(n_92),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_59),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_87),
.Y(n_115)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_52),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_89)
);

OA22x2_ASAP7_75t_SL g90 ( 
.A1(n_51),
.A2(n_45),
.B1(n_42),
.B2(n_41),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_60),
.A2(n_37),
.B1(n_42),
.B2(n_28),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_28),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_93),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_58),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_53),
.B(n_15),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_95),
.B(n_96),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_64),
.B(n_37),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_37),
.B1(n_44),
.B2(n_47),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_60),
.A2(n_15),
.B1(n_34),
.B2(n_21),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_100),
.A2(n_18),
.B1(n_22),
.B2(n_36),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_68),
.A2(n_21),
.B1(n_36),
.B2(n_27),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_55),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_102),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_64),
.B(n_49),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_103),
.Y(n_117)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_55),
.B(n_44),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_105),
.Y(n_120)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_111),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_57),
.A2(n_71),
.B(n_1),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_112),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_114),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_18),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_119),
.B(n_145),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_125),
.A2(n_140),
.B(n_3),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_89),
.A2(n_72),
.B1(n_66),
.B2(n_11),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_127),
.A2(n_138),
.B1(n_99),
.B2(n_97),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_89),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_131),
.A2(n_93),
.B1(n_88),
.B2(n_112),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_136),
.B(n_74),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_79),
.A2(n_22),
.B1(n_18),
.B2(n_47),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_137),
.A2(n_78),
.B1(n_91),
.B2(n_107),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_73),
.A2(n_47),
.B1(n_49),
.B2(n_27),
.Y(n_138)
);

AOI22x1_ASAP7_75t_SL g140 ( 
.A1(n_90),
.A2(n_49),
.B1(n_47),
.B2(n_7),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_141),
.A2(n_150),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_0),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_80),
.B(n_0),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_146),
.B(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_80),
.B(n_0),
.Y(n_149)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_83),
.A2(n_47),
.B(n_8),
.C(n_9),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_110),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_151),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_152),
.A2(n_134),
.B1(n_147),
.B2(n_132),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_109),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_156),
.Y(n_198)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_158),
.Y(n_188)
);

O2A1O1Ixp33_ASAP7_75t_L g158 ( 
.A1(n_140),
.A2(n_90),
.B(n_111),
.C(n_99),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_160),
.B(n_161),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_119),
.B(n_113),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_121),
.B(n_104),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_162),
.B(n_164),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_117),
.B(n_109),
.Y(n_163)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_105),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_165),
.A2(n_175),
.B1(n_183),
.B2(n_134),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_141),
.B(n_102),
.C(n_98),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_166),
.B(n_167),
.C(n_142),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_121),
.B(n_148),
.C(n_115),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_171),
.B1(n_176),
.B2(n_147),
.Y(n_204)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_98),
.B1(n_99),
.B2(n_81),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_170),
.A2(n_172),
.B1(n_177),
.B2(n_136),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_148),
.A2(n_108),
.B1(n_94),
.B2(n_9),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_6),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_174),
.B(n_183),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_127),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_138),
.A2(n_117),
.B1(n_135),
.B2(n_139),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_150),
.B(n_145),
.Y(n_186)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_144),
.Y(n_180)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_135),
.B(n_12),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_181),
.Y(n_208)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_151),
.Y(n_182)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_182),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_125),
.A2(n_5),
.B1(n_13),
.B2(n_149),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_124),
.B(n_13),
.Y(n_185)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_185),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_190),
.B(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_167),
.B(n_166),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_193),
.Y(n_220)
);

AND2x4_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_142),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_170),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_192),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_172),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_164),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_199),
.A2(n_116),
.B1(n_123),
.B2(n_133),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_178),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_205),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_184),
.B1(n_154),
.B2(n_165),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_204),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_209),
.B(n_210),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g210 ( 
.A(n_180),
.Y(n_210)
);

NOR2x1_ASAP7_75t_L g212 ( 
.A(n_168),
.B(n_128),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_215),
.Y(n_231)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_156),
.Y(n_213)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_213),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_173),
.A2(n_124),
.B1(n_116),
.B2(n_123),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_214),
.A2(n_154),
.B1(n_169),
.B2(n_157),
.Y(n_230)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_162),
.B(n_120),
.C(n_133),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_217),
.B(n_189),
.Y(n_239)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_214),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_196),
.A2(n_184),
.B1(n_159),
.B2(n_160),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_226),
.A2(n_229),
.B1(n_230),
.B2(n_199),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_211),
.Y(n_227)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_227),
.Y(n_248)
);

XOR2x1_ASAP7_75t_L g228 ( 
.A(n_190),
.B(n_179),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_239),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_188),
.A2(n_155),
.B(n_175),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_235),
.B(n_192),
.Y(n_244)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_188),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_236),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g234 ( 
.A(n_206),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_216),
.Y(n_235)
);

AO22x1_ASAP7_75t_SL g236 ( 
.A1(n_190),
.A2(n_155),
.B1(n_144),
.B2(n_120),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_210),
.Y(n_237)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_194),
.B1(n_200),
.B2(n_203),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_130),
.B1(n_132),
.B2(n_174),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_243),
.A2(n_202),
.B1(n_195),
.B2(n_217),
.Y(n_256)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_244),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_225),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_245),
.B(n_246),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_252),
.A2(n_254),
.B1(n_257),
.B2(n_223),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_255),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_256),
.B(n_242),
.Y(n_279)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_235),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_219),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_259),
.B(n_226),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g266 ( 
.A1(n_260),
.A2(n_218),
.B1(n_228),
.B2(n_236),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_233),
.A2(n_207),
.B1(n_186),
.B2(n_187),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_261),
.A2(n_264),
.B1(n_232),
.B2(n_253),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_207),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_263),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_224),
.A2(n_212),
.B1(n_193),
.B2(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_266),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_239),
.C(n_221),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_275),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_268),
.A2(n_280),
.B1(n_252),
.B2(n_250),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NOR2xp67_ASAP7_75t_SL g272 ( 
.A(n_244),
.B(n_242),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_272),
.A2(n_248),
.B(n_257),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_273),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_255),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_220),
.C(n_236),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_278),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_220),
.C(n_231),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_279),
.B(n_247),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_254),
.A2(n_243),
.B1(n_231),
.B2(n_219),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_264),
.B(n_238),
.Y(n_281)
);

OA21x2_ASAP7_75t_SL g293 ( 
.A1(n_281),
.A2(n_246),
.B(n_258),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_286),
.B(n_288),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_247),
.B(n_261),
.Y(n_289)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_289),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_276),
.B(n_263),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_291),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_279),
.B(n_253),
.Y(n_292)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_292),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_293),
.A2(n_283),
.B1(n_287),
.B2(n_282),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_294),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_267),
.B(n_249),
.Y(n_296)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_296),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_297),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_274),
.B1(n_265),
.B2(n_268),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_301),
.B(n_302),
.Y(n_313)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_295),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_303),
.A2(n_274),
.B1(n_270),
.B2(n_292),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_290),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_310),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_308),
.A2(n_303),
.B1(n_266),
.B2(n_271),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_277),
.B1(n_270),
.B2(n_285),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_309),
.B(n_312),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_291),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_300),
.A2(n_296),
.B(n_294),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_311),
.A2(n_13),
.B(n_5),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_305),
.B(n_271),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_299),
.C(n_301),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_315),
.B(n_316),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_304),
.Y(n_316)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_319),
.A2(n_313),
.B(n_308),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_321),
.B(n_318),
.Y(n_324)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_324),
.B(n_323),
.C(n_317),
.Y(n_326)
);

INVxp33_ASAP7_75t_L g327 ( 
.A(n_326),
.Y(n_327)
);

A2O1A1Ixp33_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_325),
.B(n_310),
.C(n_320),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_328),
.B(n_320),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_130),
.Y(n_330)
);


endmodule