module fake_jpeg_29651_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_19),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_10),
.B(n_38),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_39),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_14),
.B(n_0),
.Y(n_64)
);

BUFx16f_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

INVx2_ASAP7_75t_R g69 ( 
.A(n_25),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_10),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_65),
.Y(n_73)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_73),
.Y(n_86)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_80),
.Y(n_82)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_77),
.Y(n_92)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_78),
.B(n_51),
.Y(n_95)
);

INVx4_ASAP7_75t_SL g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_79),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_69),
.B(n_0),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_60),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_81),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_80),
.B(n_70),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_94),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_56),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_85),
.B(n_87),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_64),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_75),
.A2(n_59),
.B1(n_68),
.B2(n_70),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_93),
.B1(n_62),
.B2(n_66),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_68),
.B1(n_63),
.B2(n_60),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_74),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_95),
.B(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_104),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_L g98 ( 
.A1(n_82),
.A2(n_71),
.B(n_67),
.C(n_52),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_98),
.B(n_103),
.Y(n_119)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_100),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_90),
.A2(n_51),
.B1(n_52),
.B2(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_101),
.A2(n_105),
.B1(n_106),
.B2(n_110),
.Y(n_117)
);

INVxp33_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_67),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_SL g105 ( 
.A1(n_91),
.A2(n_74),
.B(n_84),
.C(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_107),
.Y(n_122)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_86),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_109),
.Y(n_131)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_92),
.A2(n_62),
.B1(n_72),
.B2(n_61),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_84),
.A2(n_58),
.B1(n_55),
.B2(n_54),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_111),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_112),
.B(n_115),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g113 ( 
.A(n_94),
.B(n_1),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_113),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_87),
.B(n_2),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_114),
.B(n_27),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_2),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_26),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_132),
.C(n_29),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_97),
.B(n_3),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_135),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_125),
.Y(n_140)
);

NOR2x1_ASAP7_75t_L g124 ( 
.A(n_110),
.B(n_3),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_127),
.B(n_50),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_98),
.B(n_4),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_101),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_133),
.B1(n_12),
.B2(n_15),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_32),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_105),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_105),
.B(n_8),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_148),
.B1(n_124),
.B2(n_132),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_119),
.B(n_36),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_138),
.B(n_139),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_34),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_120),
.A2(n_12),
.B(n_16),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_141),
.A2(n_144),
.B(n_146),
.Y(n_154)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_143),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_18),
.B(n_20),
.C(n_22),
.D(n_23),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_131),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_136),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_142),
.A2(n_128),
.B(n_117),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_155),
.B(n_117),
.C(n_149),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_154),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_150),
.A2(n_140),
.B(n_141),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_150),
.B(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_160),
.B(n_153),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_146),
.B(n_144),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_162),
.A2(n_151),
.B1(n_41),
.B2(n_43),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_163),
.A2(n_33),
.A3(n_45),
.B1(n_46),
.B2(n_47),
.C1(n_48),
.C2(n_49),
.Y(n_164)
);


endmodule