module fake_jpeg_3066_n_653 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_653);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_653;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_19),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_12),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_0),
.Y(n_53)
);

INVx8_ASAP7_75t_SL g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_26),
.A2(n_10),
.B1(n_18),
.B2(n_17),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_58),
.A2(n_34),
.B1(n_44),
.B2(n_28),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_59),
.Y(n_158)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_60),
.Y(n_180)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_61),
.Y(n_141)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_10),
.Y(n_62)
);

OR2x2_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_132),
.Y(n_156)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx3_ASAP7_75t_SL g204 ( 
.A(n_63),
.Y(n_204)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_64),
.Y(n_160)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_65),
.Y(n_166)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_66),
.B(n_69),
.Y(n_133)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_67),
.Y(n_143)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_40),
.B(n_9),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_70),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_71),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_72),
.Y(n_150)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_20),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_73),
.B(n_93),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx4_ASAP7_75t_SL g164 ( 
.A(n_74),
.Y(n_164)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_76),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_37),
.B(n_19),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_77),
.B(n_83),
.Y(n_147)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_26),
.Y(n_78)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_78),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_79),
.Y(n_170)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_80),
.Y(n_157)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_26),
.Y(n_81)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_81),
.Y(n_222)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

INVx8_ASAP7_75t_L g163 ( 
.A(n_82),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_31),
.B(n_41),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_84),
.Y(n_174)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_85),
.Y(n_214)
);

INVx11_ASAP7_75t_L g86 ( 
.A(n_29),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g233 ( 
.A(n_86),
.Y(n_233)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_88),
.Y(n_182)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_89),
.Y(n_206)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_90),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_19),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_92),
.B(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_29),
.Y(n_94)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_94),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_54),
.Y(n_95)
);

CKINVDCx14_ASAP7_75t_R g161 ( 
.A(n_95),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_96),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_99),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g100 ( 
.A(n_47),
.Y(n_100)
);

BUFx4f_ASAP7_75t_L g196 ( 
.A(n_100),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_56),
.Y(n_101)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_101),
.Y(n_234)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_29),
.Y(n_102)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_102),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_41),
.B(n_49),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_9),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_106),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_21),
.Y(n_105)
);

INVx8_ASAP7_75t_L g201 ( 
.A(n_105),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_49),
.B(n_9),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_56),
.Y(n_107)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_107),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_27),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_108),
.Y(n_137)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_29),
.Y(n_109)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_109),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g171 ( 
.A(n_110),
.Y(n_171)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_29),
.Y(n_111)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_111),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_27),
.A2(n_9),
.B1(n_18),
.B2(n_17),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_112),
.A2(n_117),
.B1(n_53),
.B2(n_57),
.Y(n_134)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_36),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_118),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_23),
.B(n_8),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_116),
.Y(n_155)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_38),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_23),
.A2(n_8),
.B1(n_18),
.B2(n_16),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_38),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_50),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g194 ( 
.A(n_119),
.B(n_100),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_36),
.Y(n_120)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_38),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_121),
.B(n_124),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_36),
.Y(n_122)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_36),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_123),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_46),
.Y(n_124)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_46),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_125),
.Y(n_230)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_46),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g154 ( 
.A(n_126),
.Y(n_154)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_33),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_127),
.B(n_129),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_128),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_50),
.B(n_7),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_130),
.Y(n_183)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_33),
.Y(n_131)
);

CKINVDCx9p33_ASAP7_75t_R g178 ( 
.A(n_131),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_57),
.A2(n_7),
.B1(n_16),
.B2(n_15),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g315 ( 
.A1(n_134),
.A2(n_194),
.B(n_189),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_43),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_139),
.B(n_145),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_43),
.Y(n_145)
);

OA22x2_ASAP7_75t_L g254 ( 
.A1(n_146),
.A2(n_192),
.B1(n_154),
.B2(n_180),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_70),
.A2(n_76),
.B1(n_97),
.B2(n_91),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_149),
.A2(n_151),
.B1(n_153),
.B2(n_191),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_71),
.A2(n_24),
.B1(n_45),
.B2(n_44),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_72),
.A2(n_45),
.B1(n_34),
.B2(n_24),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_SL g168 ( 
.A1(n_79),
.A2(n_28),
.B(n_25),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_168),
.B(n_194),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_119),
.B(n_105),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_172),
.B(n_179),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_108),
.A2(n_25),
.B1(n_33),
.B2(n_48),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_176),
.A2(n_186),
.B1(n_191),
.B2(n_212),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g278 ( 
.A(n_177),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_74),
.B(n_15),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_74),
.B(n_15),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_181),
.B(n_185),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_98),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_184),
.B(n_193),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_105),
.B(n_14),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_82),
.A2(n_48),
.B1(n_33),
.B2(n_30),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_99),
.A2(n_48),
.B1(n_33),
.B2(n_30),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_187),
.A2(n_208),
.B1(n_3),
.B2(n_178),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_101),
.A2(n_48),
.B1(n_30),
.B2(n_21),
.Y(n_191)
);

BUFx16f_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_192),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_107),
.B(n_0),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_126),
.B(n_14),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_195),
.B(n_197),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_111),
.B(n_14),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_60),
.A2(n_48),
.B1(n_30),
.B2(n_21),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_198),
.A2(n_225),
.B1(n_212),
.B2(n_186),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_114),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_202),
.B(n_227),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_78),
.B(n_13),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_203),
.B(n_210),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_59),
.A2(n_30),
.B1(n_21),
.B2(n_13),
.Y(n_208)
);

CKINVDCx12_ASAP7_75t_R g209 ( 
.A(n_86),
.Y(n_209)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_209),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_120),
.B(n_130),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_19),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_211),
.B(n_218),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_63),
.A2(n_6),
.B1(n_16),
.B2(n_2),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_123),
.B(n_0),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_213),
.B(n_224),
.Y(n_283)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_125),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_216),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_0),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_131),
.B(n_0),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_219),
.B(n_231),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g220 ( 
.A(n_96),
.B(n_1),
.Y(n_220)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_220),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_65),
.B(n_1),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_58),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_64),
.A2(n_2),
.B1(n_3),
.B2(n_77),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_204),
.B1(n_141),
.B2(n_150),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_115),
.B(n_2),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_115),
.B(n_2),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_228),
.B(n_161),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_69),
.B(n_3),
.Y(n_231)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_236),
.Y(n_337)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_192),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g360 ( 
.A(n_237),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g330 ( 
.A1(n_238),
.A2(n_254),
.B1(n_302),
.B2(n_309),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_156),
.A2(n_193),
.B1(n_184),
.B2(n_139),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_239),
.A2(n_245),
.B1(n_292),
.B2(n_303),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_145),
.B1(n_168),
.B2(n_176),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_240),
.A2(n_249),
.B1(n_273),
.B2(n_280),
.Y(n_374)
);

A2O1A1Ixp33_ASAP7_75t_L g241 ( 
.A1(n_167),
.A2(n_165),
.B(n_147),
.C(n_156),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_241),
.B(n_320),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_164),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g340 ( 
.A(n_242),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_164),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_244),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_226),
.B1(n_148),
.B2(n_142),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_150),
.Y(n_247)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_247),
.Y(n_370)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_140),
.Y(n_248)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_248),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_182),
.A2(n_206),
.B1(n_217),
.B2(n_142),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_228),
.B1(n_135),
.B2(n_234),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_250),
.A2(n_260),
.B1(n_262),
.B2(n_271),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_289),
.Y(n_326)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_253),
.A2(n_321),
.B1(n_272),
.B2(n_270),
.Y(n_367)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_140),
.Y(n_257)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_154),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_261),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_135),
.A2(n_235),
.B1(n_234),
.B2(n_221),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_199),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_263),
.B(n_297),
.Y(n_339)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_175),
.Y(n_264)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_264),
.Y(n_343)
);

AOI22x1_ASAP7_75t_SL g266 ( 
.A1(n_170),
.A2(n_214),
.B1(n_162),
.B2(n_155),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_266),
.Y(n_329)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_175),
.Y(n_267)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_267),
.Y(n_365)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_182),
.Y(n_268)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_268),
.Y(n_375)
);

INVx11_ASAP7_75t_L g269 ( 
.A(n_233),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_144),
.B(n_133),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_270),
.B(n_274),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_173),
.A2(n_235),
.B1(n_207),
.B2(n_221),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_152),
.A2(n_199),
.B1(n_215),
.B2(n_170),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_272),
.A2(n_284),
.B(n_263),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_L g273 ( 
.A1(n_206),
.A2(n_217),
.B1(n_141),
.B2(n_204),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_157),
.B(n_223),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_196),
.Y(n_275)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_275),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_276),
.B(n_291),
.Y(n_331)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_169),
.Y(n_277)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_277),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_204),
.A2(n_190),
.B1(n_169),
.B2(n_150),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_199),
.A2(n_152),
.B(n_196),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g381 ( 
.A1(n_284),
.A2(n_278),
.B(n_285),
.Y(n_381)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_196),
.Y(n_286)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_286),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_157),
.B(n_223),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_287),
.B(n_288),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_152),
.B(n_183),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_162),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_188),
.B(n_232),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_173),
.A2(n_207),
.B1(n_160),
.B2(n_166),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_138),
.B(n_202),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_293),
.B(n_307),
.Y(n_348)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_200),
.Y(n_294)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_136),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g341 ( 
.A(n_295),
.Y(n_341)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_190),
.A2(n_229),
.B1(n_158),
.B2(n_138),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_296),
.A2(n_301),
.B1(n_304),
.B2(n_317),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g297 ( 
.A(n_162),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_200),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_298),
.B(n_300),
.Y(n_355)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_174),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_229),
.A2(n_158),
.B1(n_159),
.B2(n_183),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_180),
.A2(n_174),
.B1(n_164),
.B2(n_143),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_160),
.A2(n_166),
.B1(n_163),
.B2(n_229),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_163),
.A2(n_215),
.B1(n_159),
.B2(n_171),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_188),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_305),
.B(n_306),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_205),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_177),
.B(n_216),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_232),
.B(n_136),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_308),
.B(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_174),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_309),
.B(n_312),
.Y(n_377)
);

OA22x2_ASAP7_75t_L g310 ( 
.A1(n_214),
.A2(n_143),
.B1(n_233),
.B2(n_171),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g346 ( 
.A1(n_310),
.A2(n_238),
.B(n_304),
.C(n_319),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_137),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_311),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_233),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_230),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_313),
.B(n_314),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_233),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_315),
.A2(n_319),
.B1(n_300),
.B2(n_303),
.Y(n_349)
);

BUFx12f_ASAP7_75t_L g316 ( 
.A(n_201),
.Y(n_316)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_316),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_137),
.A2(n_171),
.B1(n_201),
.B2(n_222),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_137),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_318),
.B(n_325),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_137),
.A2(n_171),
.B1(n_222),
.B2(n_189),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_230),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_151),
.A2(n_153),
.B1(n_149),
.B2(n_92),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_139),
.B(n_193),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_323),
.B(n_290),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_147),
.B(n_167),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_182),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_328),
.A2(n_362),
.B(n_310),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_330),
.Y(n_417)
);

MAJx2_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_239),
.C(n_252),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_334),
.B(n_350),
.C(n_354),
.Y(n_401)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_346),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_349),
.B(n_381),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_259),
.B(n_243),
.C(n_241),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_259),
.B(n_283),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g403 ( 
.A(n_352),
.B(n_356),
.C(n_385),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_243),
.B(n_256),
.C(n_245),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_283),
.B(n_282),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_357),
.B(n_316),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_274),
.B(n_287),
.C(n_265),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_358),
.B(n_361),
.C(n_373),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_246),
.A2(n_260),
.B1(n_250),
.B2(n_299),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_359),
.A2(n_363),
.B1(n_317),
.B2(n_314),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_288),
.B(n_322),
.C(n_308),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_293),
.A2(n_281),
.B1(n_292),
.B2(n_271),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_246),
.A2(n_255),
.B1(n_253),
.B2(n_262),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_307),
.B(n_294),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_386),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_367),
.A2(n_376),
.B1(n_329),
.B2(n_363),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_268),
.B(n_325),
.C(n_254),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_266),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_310),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_306),
.B(n_254),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_379),
.B(n_380),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_254),
.B(n_312),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_279),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_248),
.B(n_298),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_257),
.B(n_267),
.C(n_264),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_387),
.B(n_326),
.Y(n_430)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_384),
.Y(n_388)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_388),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g389 ( 
.A1(n_380),
.A2(n_285),
.B(n_278),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_389),
.A2(n_392),
.B(n_393),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_390),
.A2(n_400),
.B1(n_421),
.B2(n_426),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_386),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_395),
.B(n_404),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_305),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_396),
.B(n_402),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_406),
.B1(n_407),
.B2(n_423),
.Y(n_456)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_359),
.A2(n_333),
.B1(n_329),
.B2(n_348),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_350),
.B(n_347),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_377),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_332),
.Y(n_405)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_405),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_333),
.A2(n_277),
.B1(n_247),
.B2(n_310),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_345),
.A2(n_247),
.B1(n_297),
.B2(n_289),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_348),
.B(n_236),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_408),
.B(n_411),
.Y(n_445)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_332),
.Y(n_409)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_409),
.Y(n_437)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_342),
.Y(n_410)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_331),
.B(n_286),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_242),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_412),
.B(n_413),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_331),
.B(n_358),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g414 ( 
.A(n_381),
.B(n_347),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_414),
.B(n_419),
.Y(n_466)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_342),
.Y(n_415)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_415),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_328),
.B(n_244),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_418),
.A2(n_340),
.B(n_344),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_352),
.B(n_318),
.Y(n_419)
);

FAx1_ASAP7_75t_SL g420 ( 
.A(n_334),
.B(n_269),
.CI(n_275),
.CON(n_420),
.SN(n_420)
);

FAx1_ASAP7_75t_SL g473 ( 
.A(n_420),
.B(n_353),
.CI(n_341),
.CON(n_473),
.SN(n_473)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_338),
.A2(n_313),
.B1(n_320),
.B2(n_311),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_361),
.B(n_237),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_422),
.B(n_424),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_345),
.A2(n_311),
.B1(n_316),
.B2(n_258),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_327),
.B(n_258),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_327),
.B(n_258),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_425),
.B(n_428),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_336),
.A2(n_258),
.B1(n_316),
.B2(n_326),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_377),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_432),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_326),
.B(n_339),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g463 ( 
.A(n_429),
.B(n_371),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_430),
.B(n_343),
.Y(n_459)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_343),
.Y(n_431)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_431),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_372),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_379),
.A2(n_336),
.B1(n_374),
.B2(n_373),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_433),
.A2(n_357),
.B1(n_356),
.B2(n_349),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_334),
.B(n_354),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_434),
.B(n_369),
.Y(n_452)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_394),
.A2(n_383),
.B(n_346),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_438),
.A2(n_455),
.B(n_414),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_439),
.A2(n_440),
.B1(n_476),
.B2(n_432),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_399),
.A2(n_398),
.B1(n_433),
.B2(n_395),
.Y(n_440)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_405),
.Y(n_442)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_442),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_401),
.B(n_387),
.C(n_339),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_449),
.B(n_453),
.C(n_458),
.Y(n_478)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_409),
.Y(n_451)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_451),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_452),
.B(n_454),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_434),
.C(n_416),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_416),
.B(n_369),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_394),
.A2(n_383),
.B(n_346),
.Y(n_455)
);

OAI22x1_ASAP7_75t_L g457 ( 
.A1(n_399),
.A2(n_355),
.B1(n_372),
.B2(n_365),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_457),
.A2(n_418),
.B1(n_404),
.B2(n_397),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_355),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_459),
.B(n_462),
.C(n_475),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_351),
.B1(n_365),
.B2(n_382),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g489 ( 
.A1(n_460),
.A2(n_461),
.B1(n_467),
.B2(n_431),
.Y(n_489)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_390),
.A2(n_351),
.B1(n_382),
.B2(n_368),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_429),
.C(n_413),
.Y(n_462)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_463),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_396),
.Y(n_465)
);

INVxp33_ASAP7_75t_SL g509 ( 
.A(n_465),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_406),
.A2(n_368),
.B1(n_344),
.B2(n_370),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_402),
.B(n_335),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_469),
.B(n_471),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_403),
.B(n_428),
.Y(n_471)
);

OAI21xp5_ASAP7_75t_SL g485 ( 
.A1(n_472),
.A2(n_473),
.B(n_418),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_341),
.C(n_353),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_391),
.A2(n_370),
.B1(n_337),
.B2(n_375),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_L g517 ( 
.A1(n_479),
.A2(n_482),
.B1(n_489),
.B2(n_493),
.Y(n_517)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_442),
.Y(n_480)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_480),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_436),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_481),
.B(n_487),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_440),
.A2(n_389),
.B1(n_417),
.B2(n_397),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_451),
.Y(n_483)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_483),
.Y(n_520)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_484),
.Y(n_525)
);

INVxp67_ASAP7_75t_L g549 ( 
.A(n_485),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_444),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_488),
.B(n_497),
.Y(n_534)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_437),
.Y(n_490)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_391),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_464),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_L g493 ( 
.A1(n_461),
.A2(n_408),
.B1(n_407),
.B2(n_423),
.Y(n_493)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_443),
.Y(n_496)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_496),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_445),
.B(n_427),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_SL g498 ( 
.A1(n_435),
.A2(n_418),
.B(n_397),
.Y(n_498)
);

CKINVDCx16_ASAP7_75t_R g499 ( 
.A(n_438),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_499),
.B(n_502),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_500),
.A2(n_506),
.B1(n_473),
.B2(n_463),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g501 ( 
.A1(n_435),
.A2(n_414),
.B(n_418),
.Y(n_501)
);

NOR2x1_ASAP7_75t_L g544 ( 
.A(n_501),
.B(n_510),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_476),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_455),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_503),
.B(n_504),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_445),
.B(n_412),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_446),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_505),
.B(n_511),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_447),
.A2(n_393),
.B1(n_426),
.B2(n_403),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_472),
.A2(n_392),
.B(n_420),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_SL g526 ( 
.A(n_508),
.B(n_513),
.C(n_473),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_460),
.B(n_425),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_466),
.A2(n_424),
.B(n_420),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_466),
.A2(n_420),
.B(n_419),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_447),
.A2(n_411),
.B(n_415),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_453),
.B(n_410),
.C(n_360),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_514),
.B(n_515),
.C(n_459),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_449),
.B(n_337),
.C(n_421),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_443),
.Y(n_516)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_516),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_439),
.B1(n_456),
.B2(n_457),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_521),
.A2(n_536),
.B1(n_482),
.B2(n_493),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_SL g572 ( 
.A(n_522),
.B(n_540),
.C(n_504),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_523),
.B(n_528),
.C(n_515),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_478),
.B(n_462),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_524),
.B(n_527),
.Y(n_558)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_526),
.B(n_477),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_478),
.B(n_452),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_458),
.C(n_474),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_529),
.B(n_527),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_497),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_531),
.B(n_532),
.Y(n_566)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_488),
.Y(n_532)
);

NAND3xp33_ASAP7_75t_L g533 ( 
.A(n_477),
.B(n_441),
.C(n_464),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_533),
.B(n_481),
.Y(n_571)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_495),
.Y(n_535)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_535),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g536 ( 
.A1(n_510),
.A2(n_474),
.B1(n_467),
.B2(n_463),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_486),
.B(n_448),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_546),
.Y(n_559)
);

INVx3_ASAP7_75t_SL g538 ( 
.A(n_495),
.Y(n_538)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_538),
.Y(n_553)
);

A2O1A1O1Ixp25_ASAP7_75t_L g540 ( 
.A1(n_512),
.A2(n_475),
.B(n_448),
.C(n_468),
.D(n_470),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g541 ( 
.A1(n_479),
.A2(n_470),
.B1(n_450),
.B2(n_446),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_541),
.A2(n_545),
.B1(n_550),
.B2(n_525),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_506),
.A2(n_450),
.B1(n_388),
.B2(n_384),
.Y(n_545)
);

XNOR2xp5_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_494),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_494),
.B(n_375),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g567 ( 
.A(n_547),
.B(n_487),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_552),
.B(n_562),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_554),
.A2(n_563),
.B1(n_577),
.B2(n_578),
.Y(n_590)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_534),
.Y(n_555)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

XOR2xp5_ASAP7_75t_L g592 ( 
.A(n_556),
.B(n_544),
.Y(n_592)
);

XNOR2xp5_ASAP7_75t_L g557 ( 
.A(n_524),
.B(n_537),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_557),
.B(n_560),
.Y(n_582)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_550),
.Y(n_561)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_561),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g562 ( 
.A(n_530),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_518),
.B(n_500),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_523),
.B(n_492),
.C(n_491),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_564),
.B(n_568),
.C(n_573),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_528),
.B(n_501),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_565),
.B(n_567),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_498),
.C(n_509),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_521),
.A2(n_503),
.B1(n_499),
.B2(n_508),
.Y(n_569)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_569),
.Y(n_585)
);

XNOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_529),
.B(n_511),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_571),
.B(n_544),
.Y(n_596)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_572),
.B(n_574),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_547),
.B(n_513),
.C(n_485),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_536),
.B(n_516),
.Y(n_574)
);

OAI22xp5_ASAP7_75t_SL g575 ( 
.A1(n_548),
.A2(n_502),
.B1(n_496),
.B2(n_490),
.Y(n_575)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_575),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_549),
.B(n_483),
.C(n_480),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_576),
.B(n_520),
.C(n_519),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g578 ( 
.A1(n_517),
.A2(n_484),
.B1(n_505),
.B2(n_507),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_542),
.Y(n_579)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_579),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_575),
.B(n_541),
.Y(n_580)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_580),
.Y(n_604)
);

CKINVDCx16_ASAP7_75t_R g583 ( 
.A(n_576),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_583),
.B(n_593),
.Y(n_609)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_566),
.Y(n_584)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_584),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_539),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_592),
.B(n_565),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_553),
.B(n_543),
.Y(n_594)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_594),
.Y(n_615)
);

NOR3xp33_ASAP7_75t_SL g610 ( 
.A(n_596),
.B(n_572),
.C(n_570),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g597 ( 
.A1(n_563),
.A2(n_549),
.B1(n_526),
.B2(n_540),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g611 ( 
.A1(n_597),
.A2(n_558),
.B1(n_577),
.B2(n_560),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_558),
.B(n_545),
.C(n_535),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_598),
.B(n_564),
.C(n_569),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_388),
.Y(n_599)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_599),
.Y(n_617)
);

FAx1_ASAP7_75t_SL g600 ( 
.A(n_552),
.B(n_507),
.CI(n_538),
.CON(n_600),
.SN(n_600)
);

MAJIxp5_ASAP7_75t_SL g613 ( 
.A(n_600),
.B(n_557),
.C(n_551),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_603),
.B(n_614),
.Y(n_622)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_585),
.A2(n_568),
.B(n_573),
.Y(n_606)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_606),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_L g607 ( 
.A1(n_585),
.A2(n_586),
.B(n_581),
.Y(n_607)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_607),
.Y(n_626)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_587),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_608),
.B(n_610),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_611),
.A2(n_592),
.B1(n_602),
.B2(n_597),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_613),
.B(n_616),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_582),
.B(n_559),
.C(n_340),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_595),
.A2(n_559),
.B1(n_384),
.B2(n_378),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_582),
.B(n_378),
.C(n_366),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_618),
.B(n_589),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_593),
.B(n_366),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_619),
.B(n_598),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_624),
.B(n_628),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_625),
.B(n_621),
.Y(n_633)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_627),
.A2(n_619),
.B(n_605),
.Y(n_638)
);

AOI22xp5_ASAP7_75t_L g628 ( 
.A1(n_604),
.A2(n_590),
.B1(n_586),
.B2(n_580),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_607),
.A2(n_588),
.B1(n_602),
.B2(n_594),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_629),
.B(n_630),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_609),
.B(n_591),
.C(n_589),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_612),
.B(n_601),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_631),
.B(n_619),
.Y(n_639)
);

OAI21xp5_ASAP7_75t_SL g632 ( 
.A1(n_620),
.A2(n_606),
.B(n_611),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_SL g641 ( 
.A1(n_632),
.A2(n_638),
.B(n_621),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_633),
.B(n_640),
.Y(n_644)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_630),
.B(n_603),
.C(n_614),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_634),
.B(n_639),
.Y(n_645)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_620),
.B(n_615),
.Y(n_636)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_636),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_623),
.B(n_617),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g648 ( 
.A(n_641),
.B(n_613),
.C(n_629),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_634),
.B(n_637),
.C(n_632),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_642),
.B(n_635),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g650 ( 
.A1(n_646),
.A2(n_647),
.B(n_648),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_645),
.B(n_626),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g649 ( 
.A(n_646),
.B(n_643),
.C(n_644),
.Y(n_649)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_649),
.B(n_645),
.C(n_622),
.Y(n_651)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_651),
.B(n_650),
.C(n_628),
.Y(n_652)
);

XOR2xp5_ASAP7_75t_L g653 ( 
.A(n_652),
.B(n_625),
.Y(n_653)
);


endmodule