module fake_jpeg_30409_n_411 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_411);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_411;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_7),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_21),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_45),
.B(n_54),
.Y(n_89)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_49),
.Y(n_109)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_20),
.B(n_0),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_50),
.B(n_38),
.C(n_40),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_17),
.B(n_28),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_83),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_20),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_85),
.Y(n_94)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_53),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_21),
.B(n_14),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_56),
.Y(n_106)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_57),
.Y(n_110)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_31),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_60),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_22),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_62),
.Y(n_138)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_63),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_17),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_67),
.Y(n_98)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_31),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_23),
.B(n_14),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_23),
.A2(n_41),
.B1(n_28),
.B2(n_24),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_68),
.A2(n_16),
.B1(n_19),
.B2(n_29),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_13),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_71),
.Y(n_101)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_70),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_26),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_26),
.B(n_1),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_77),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_32),
.Y(n_74)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_32),
.Y(n_75)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_75),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_22),
.Y(n_76)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_76),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_36),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g140 ( 
.A(n_78),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_36),
.B(n_2),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_2),
.Y(n_80)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_81),
.B(n_82),
.Y(n_131)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_37),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_84),
.B(n_39),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_2),
.Y(n_85)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_86),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_88),
.B(n_104),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_52),
.A2(n_16),
.B1(n_19),
.B2(n_29),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_91),
.A2(n_95),
.B1(n_114),
.B2(n_120),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_64),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_116),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_65),
.A2(n_39),
.B1(n_40),
.B2(n_35),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_85),
.B(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_115),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_50),
.A2(n_16),
.B1(n_19),
.B2(n_40),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_100),
.A2(n_112),
.B1(n_125),
.B2(n_135),
.Y(n_175)
);

AO22x1_ASAP7_75t_SL g112 ( 
.A1(n_50),
.A2(n_40),
.B1(n_35),
.B2(n_38),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_49),
.A2(n_39),
.B1(n_35),
.B2(n_31),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_46),
.B(n_34),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_77),
.B(n_25),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_83),
.A2(n_35),
.B1(n_39),
.B2(n_38),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_121),
.B(n_133),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_73),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_122),
.A2(n_127),
.B1(n_132),
.B2(n_62),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_84),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_86),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_57),
.B(n_6),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_130),
.B(n_135),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_47),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_51),
.B(n_7),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_59),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_48),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_81),
.B1(n_63),
.B2(n_55),
.Y(n_180)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_126),
.Y(n_141)
);

INVx13_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_126),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_142),
.Y(n_220)
);

OR2x2_ASAP7_75t_SL g144 ( 
.A(n_99),
.B(n_51),
.Y(n_144)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_147),
.Y(n_225)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_145),
.Y(n_201)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_146),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_88),
.A2(n_53),
.B1(n_43),
.B2(n_56),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g148 ( 
.A(n_111),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_148),
.B(n_153),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_149),
.B(n_164),
.Y(n_192)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx11_ASAP7_75t_L g152 ( 
.A(n_138),
.Y(n_152)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_152),
.Y(n_219)
);

OR2x4_ASAP7_75t_L g153 ( 
.A(n_112),
.B(n_75),
.Y(n_153)
);

AND2x2_ASAP7_75t_SL g154 ( 
.A(n_94),
.B(n_58),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_154),
.B(n_187),
.C(n_188),
.Y(n_230)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_97),
.Y(n_156)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_156),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_111),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_157),
.B(n_160),
.Y(n_215)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_159),
.A2(n_184),
.B(n_109),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_110),
.B1(n_112),
.B2(n_93),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_94),
.B(n_74),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_161),
.B(n_169),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_139),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_162),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_118),
.Y(n_164)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_140),
.Y(n_165)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx6_ASAP7_75t_SL g226 ( 
.A(n_166),
.Y(n_226)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_87),
.Y(n_167)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_167),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_104),
.B(n_66),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_170),
.B(n_183),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_137),
.A2(n_43),
.B1(n_53),
.B2(n_55),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_182),
.B1(n_10),
.B2(n_12),
.C(n_96),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_173),
.B(n_177),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_174),
.Y(n_197)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_140),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g177 ( 
.A(n_140),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_98),
.B(n_82),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_178),
.B(n_179),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_89),
.B(n_82),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_180),
.A2(n_181),
.B1(n_137),
.B2(n_108),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_100),
.A2(n_81),
.B1(n_56),
.B2(n_70),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_119),
.A2(n_10),
.B(n_12),
.Y(n_182)
);

A2O1A1Ixp33_ASAP7_75t_L g183 ( 
.A1(n_130),
.A2(n_60),
.B(n_44),
.C(n_78),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_124),
.A2(n_61),
.B1(n_62),
.B2(n_76),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_128),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_185),
.Y(n_205)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_87),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_186),
.B(n_189),
.Y(n_194)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_102),
.B(n_61),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_102),
.B(n_76),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_101),
.B(n_78),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_190),
.B(n_105),
.Y(n_208)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_129),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_191),
.B(n_128),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_131),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_193),
.B(n_144),
.C(n_154),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_195),
.A2(n_232),
.B1(n_187),
.B2(n_188),
.Y(n_250)
);

BUFx12_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_196),
.B(n_174),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_160),
.A2(n_170),
.B1(n_149),
.B2(n_153),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_203),
.A2(n_218),
.B1(n_224),
.B2(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_175),
.A2(n_117),
.B1(n_124),
.B2(n_106),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_207),
.A2(n_214),
.B1(n_232),
.B2(n_172),
.Y(n_240)
);

OAI21xp33_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_213),
.B(n_228),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_209),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g248 ( 
.A(n_211),
.B(n_157),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_171),
.A2(n_117),
.B1(n_109),
.B2(n_103),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_168),
.B(n_106),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_161),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_147),
.A2(n_103),
.B1(n_123),
.B2(n_90),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_168),
.A2(n_123),
.B1(n_90),
.B2(n_107),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_107),
.B1(n_96),
.B2(n_105),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_150),
.A2(n_180),
.B1(n_181),
.B2(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_203),
.B(n_150),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_233),
.B(n_235),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_SL g273 ( 
.A(n_234),
.B(n_230),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_236),
.Y(n_278)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_222),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_237),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_223),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_238),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_194),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_239),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_240),
.A2(n_250),
.B1(n_221),
.B2(n_195),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_241),
.Y(n_290)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_220),
.Y(n_242)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_243),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_143),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_245),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_207),
.A2(n_156),
.B1(n_158),
.B2(n_146),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_246),
.A2(n_256),
.B1(n_257),
.B2(n_259),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_193),
.B(n_169),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_253),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_248),
.B(n_251),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_164),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_249),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_216),
.B(n_150),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_192),
.B(n_163),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_252),
.B(n_264),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_221),
.B(n_169),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_148),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_255),
.Y(n_288)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_199),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_210),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_227),
.A2(n_212),
.B1(n_215),
.B2(n_224),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_258),
.A2(n_265),
.B1(n_244),
.B2(n_263),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_223),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_212),
.B(n_167),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_263),
.Y(n_286)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_225),
.A2(n_183),
.B(n_189),
.C(n_186),
.D(n_191),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_261),
.B(n_211),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_225),
.B(n_221),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_229),
.B(n_205),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_215),
.B(n_188),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_198),
.B(n_187),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_218),
.A2(n_155),
.B1(n_151),
.B2(n_177),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_206),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_209),
.B(n_197),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_271),
.A2(n_277),
.B1(n_176),
.B2(n_242),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_272),
.A2(n_283),
.B(n_248),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_273),
.B(n_279),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_244),
.A2(n_230),
.B1(n_217),
.B2(n_194),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_274),
.A2(n_275),
.B1(n_287),
.B2(n_291),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_250),
.A2(n_217),
.B1(n_226),
.B2(n_229),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g314 ( 
.A(n_282),
.B(n_226),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_262),
.A2(n_197),
.B(n_205),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_258),
.A2(n_201),
.B1(n_165),
.B2(n_220),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_233),
.A2(n_267),
.B1(n_239),
.B2(n_251),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_235),
.A2(n_201),
.B1(n_165),
.B2(n_202),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_292),
.B(n_295),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_260),
.A2(n_254),
.B(n_266),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_257),
.B(n_256),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_240),
.A2(n_202),
.B1(n_166),
.B2(n_162),
.Y(n_295)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_299),
.Y(n_344)
);

NOR3xp33_ASAP7_75t_SL g301 ( 
.A(n_278),
.B(n_261),
.C(n_248),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_301),
.B(n_309),
.Y(n_324)
);

AO21x1_ASAP7_75t_L g335 ( 
.A1(n_302),
.A2(n_310),
.B(n_320),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_289),
.Y(n_303)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_303),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_272),
.A2(n_253),
.B(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_304),
.B(n_307),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_273),
.B(n_247),
.C(n_234),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_316),
.C(n_286),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_269),
.B(n_255),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_308),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_269),
.B(n_259),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_268),
.B(n_243),
.Y(n_311)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_311),
.Y(n_328)
);

BUFx12_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_312),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_293),
.B(n_238),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_313),
.B(n_317),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_314),
.B(n_282),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_280),
.B(n_196),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_322),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_280),
.B(n_196),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_318),
.B(n_319),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_288),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_297),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_321),
.A2(n_287),
.B1(n_295),
.B2(n_275),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_297),
.B(n_268),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_237),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_279),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_298),
.A2(n_271),
.B1(n_277),
.B2(n_276),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_330),
.A2(n_333),
.B1(n_343),
.B2(n_321),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_331),
.B(n_332),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_316),
.B(n_291),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_298),
.A2(n_276),
.B1(n_281),
.B2(n_294),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_306),
.B(n_274),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_334),
.B(n_341),
.C(n_345),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_336),
.A2(n_270),
.B1(n_328),
.B2(n_342),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_281),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_340),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_300),
.A2(n_318),
.B1(n_319),
.B2(n_317),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_286),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_346),
.A2(n_350),
.B1(n_354),
.B2(n_344),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_329),
.A2(n_304),
.B(n_310),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_348),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_311),
.Y(n_349)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_349),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_330),
.A2(n_300),
.B1(n_302),
.B2(n_301),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_307),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_352),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_338),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_343),
.A2(n_292),
.B1(n_290),
.B2(n_303),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_341),
.B(n_314),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_355),
.B(n_345),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g357 ( 
.A(n_324),
.B(n_313),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_357),
.B(n_363),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_358),
.A2(n_336),
.B1(n_344),
.B2(n_331),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g359 ( 
.A1(n_335),
.A2(n_299),
.B(n_289),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g374 ( 
.A1(n_359),
.A2(n_360),
.B(n_348),
.Y(n_374)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_335),
.A2(n_305),
.B(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_325),
.Y(n_361)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_334),
.B(n_285),
.C(n_312),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_362),
.B(n_332),
.C(n_326),
.Y(n_369)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_327),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_364),
.B(n_367),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_326),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_369),
.B(n_374),
.Y(n_382)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_371),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_373),
.B(n_378),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_308),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_375),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_353),
.B(n_337),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_376),
.B(n_377),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_355),
.B(n_340),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g378 ( 
.A(n_347),
.B(n_312),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_372),
.B(n_360),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_381),
.Y(n_394)
);

BUFx24_ASAP7_75t_SL g381 ( 
.A(n_366),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_367),
.B(n_362),
.C(n_356),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_384),
.B(n_388),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_369),
.B(n_356),
.C(n_354),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_385),
.A2(n_368),
.B1(n_365),
.B2(n_346),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_390),
.B(n_392),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_387),
.A2(n_368),
.B1(n_358),
.B2(n_359),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_391),
.B(n_347),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_386),
.A2(n_350),
.B1(n_371),
.B2(n_370),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_382),
.B(n_378),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_393),
.B(n_395),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_388),
.B(n_364),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_377),
.B(n_376),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g401 ( 
.A1(n_396),
.A2(n_384),
.B(n_380),
.Y(n_401)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_394),
.Y(n_398)
);

AOI322xp5_ASAP7_75t_L g403 ( 
.A1(n_398),
.A2(n_399),
.A3(n_400),
.B1(n_393),
.B2(n_395),
.C1(n_380),
.C2(n_391),
.Y(n_403)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_389),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_401),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_404),
.B(n_405),
.Y(n_408)
);

AOI322xp5_ASAP7_75t_L g404 ( 
.A1(n_397),
.A2(n_303),
.A3(n_219),
.B1(n_200),
.B2(n_142),
.C1(n_141),
.C2(n_145),
.Y(n_404)
);

AOI322xp5_ASAP7_75t_L g405 ( 
.A1(n_400),
.A2(n_219),
.A3(n_200),
.B1(n_173),
.B2(n_222),
.C1(n_152),
.C2(n_204),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_406),
.B(n_402),
.C(n_204),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_407),
.B(n_113),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_409),
.B(n_408),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_410),
.B(n_113),
.Y(n_411)
);


endmodule