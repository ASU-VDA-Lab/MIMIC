module fake_netlist_6_3155_n_827 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_827);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_827;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_760;
wire n_741;
wire n_680;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_683;
wire n_420;
wire n_811;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_620;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_203;
wire n_254;
wire n_207;
wire n_242;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_106),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_41),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_167),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_90),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_173),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_89),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_172),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_168),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_176),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_5),
.Y(n_188)
);

BUFx10_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

BUFx10_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_92),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_101),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_147),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_117),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_58),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_126),
.Y(n_198)
);

INVx2_ASAP7_75t_SL g199 ( 
.A(n_51),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_86),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_127),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_77),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_94),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_63),
.B(n_44),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_140),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_19),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_129),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_153),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_75),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_103),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_29),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_28),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_121),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_27),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_31),
.Y(n_221)
);

NOR2xp67_ASAP7_75t_L g222 ( 
.A(n_124),
.B(n_116),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_170),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_82),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_46),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_62),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_95),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_146),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_109),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_93),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_5),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_25),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_72),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_166),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_163),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_26),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_10),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_111),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_69),
.Y(n_242)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_156),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_96),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_22),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_169),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_88),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_158),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_186),
.Y(n_250)
);

AOI22x1_ASAP7_75t_SL g251 ( 
.A1(n_188),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_240),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_209),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_0),
.Y(n_256)
);

INVx2_ASAP7_75t_SL g257 ( 
.A(n_246),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

AND2x4_ASAP7_75t_L g260 ( 
.A(n_193),
.B(n_23),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_1),
.Y(n_261)
);

INVx6_ASAP7_75t_L g262 ( 
.A(n_189),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g264 ( 
.A1(n_196),
.A2(n_2),
.B(n_3),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_189),
.B(n_190),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_199),
.B(n_4),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_180),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_196),
.B(n_4),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_227),
.B(n_6),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_186),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_182),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_183),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_220),
.B(n_6),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_184),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_220),
.B(n_7),
.Y(n_279)
);

BUFx12f_ASAP7_75t_L g280 ( 
.A(n_190),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_221),
.B(n_24),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_223),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_223),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_226),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_221),
.B(n_225),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_185),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_191),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g288 ( 
.A(n_249),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_225),
.B(n_7),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_194),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_226),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_195),
.B(n_32),
.Y(n_292)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_226),
.Y(n_293)
);

BUFx8_ASAP7_75t_SL g294 ( 
.A(n_248),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_200),
.B(n_33),
.Y(n_295)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_205),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g297 ( 
.A(n_206),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_208),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_216),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_261),
.B(n_248),
.Y(n_301)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_293),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_267),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_255),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_255),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_274),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_269),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_275),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_258),
.B(n_213),
.Y(n_311)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_215),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

NOR2x1p5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_207),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_273),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_256),
.B(n_8),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_265),
.B(n_217),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_257),
.B(n_224),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_257),
.B(n_228),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_292),
.B(n_230),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_261),
.B(n_222),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_231),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_260),
.B(n_178),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_262),
.B(n_233),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_292),
.B(n_235),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_260),
.B(n_179),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_250),
.Y(n_329)
);

NAND2xp33_ASAP7_75t_L g330 ( 
.A(n_266),
.B(n_187),
.Y(n_330)
);

INVx3_ASAP7_75t_L g331 ( 
.A(n_250),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_276),
.Y(n_332)
);

INVx2_ASAP7_75t_SL g333 ( 
.A(n_262),
.Y(n_333)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_286),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_276),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_284),
.Y(n_337)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_288),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_284),
.Y(n_339)
);

AND3x4_ASAP7_75t_L g340 ( 
.A(n_251),
.B(n_8),
.C(n_9),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_260),
.B(n_192),
.Y(n_341)
);

AND3x2_ASAP7_75t_L g342 ( 
.A(n_265),
.B(n_237),
.C(n_236),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

BUFx6f_ASAP7_75t_SL g344 ( 
.A(n_295),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_262),
.B(n_242),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_295),
.B(n_247),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_284),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_298),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_254),
.A2(n_245),
.B1(n_244),
.B2(n_241),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_321),
.B(n_281),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_303),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_338),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_318),
.B(n_254),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_323),
.B(n_281),
.Y(n_356)
);

OR2x6_ASAP7_75t_L g357 ( 
.A(n_301),
.B(n_315),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_329),
.Y(n_358)
);

INVx2_ASAP7_75t_SL g359 ( 
.A(n_312),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_327),
.B(n_347),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_318),
.B(n_280),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_337),
.Y(n_362)
);

OR2x6_ASAP7_75t_L g363 ( 
.A(n_301),
.B(n_282),
.Y(n_363)
);

AND2x4_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_295),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_322),
.B(n_262),
.Y(n_365)
);

BUFx8_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

OR2x2_ASAP7_75t_L g367 ( 
.A(n_311),
.B(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_305),
.Y(n_368)
);

O2A1O1Ixp33_ASAP7_75t_L g369 ( 
.A1(n_322),
.A2(n_268),
.B(n_289),
.C(n_277),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_293),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_311),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_307),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_313),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g374 ( 
.A(n_351),
.B(n_271),
.Y(n_374)
);

NAND2xp33_ASAP7_75t_L g375 ( 
.A(n_319),
.B(n_197),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_310),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_325),
.B(n_283),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_337),
.Y(n_378)
);

NOR3xp33_ASAP7_75t_SL g379 ( 
.A(n_317),
.B(n_256),
.C(n_279),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_328),
.B(n_293),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_328),
.B(n_283),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_239),
.B1(n_201),
.B2(n_203),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_341),
.B(n_293),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_304),
.B(n_285),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_L g385 ( 
.A1(n_341),
.A2(n_285),
.B1(n_253),
.B2(n_252),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_339),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_339),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_333),
.B(n_198),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_320),
.B(n_296),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_348),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_324),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_326),
.B(n_296),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_348),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_306),
.B(n_285),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_335),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_330),
.A2(n_238),
.B1(n_210),
.B2(n_211),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_349),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_346),
.B(n_204),
.Y(n_401)
);

NAND2x1_ASAP7_75t_L g402 ( 
.A(n_329),
.B(n_250),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_314),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_350),
.B(n_297),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_308),
.B(n_212),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_308),
.B(n_299),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_344),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_331),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_344),
.A2(n_218),
.B1(n_219),
.B2(n_229),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_309),
.B(n_297),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_331),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_331),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g414 ( 
.A1(n_340),
.A2(n_263),
.B1(n_299),
.B2(n_300),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_344),
.B(n_294),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_316),
.Y(n_416)
);

OAI221xp5_ASAP7_75t_L g417 ( 
.A1(n_316),
.A2(n_263),
.B1(n_300),
.B2(n_291),
.C(n_250),
.Y(n_417)
);

A2O1A1Ixp33_ASAP7_75t_L g418 ( 
.A1(n_369),
.A2(n_360),
.B(n_352),
.C(n_356),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_L g419 ( 
.A1(n_360),
.A2(n_264),
.B(n_336),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_352),
.B(n_332),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_356),
.B(n_332),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g422 ( 
.A1(n_384),
.A2(n_334),
.B(n_302),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_396),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_336),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_384),
.A2(n_334),
.B(n_302),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_389),
.B(n_300),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_403),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_362),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_364),
.B(n_263),
.Y(n_429)
);

AOI21x1_ASAP7_75t_L g430 ( 
.A1(n_394),
.A2(n_264),
.B(n_334),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_364),
.B(n_342),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_394),
.A2(n_380),
.B(n_370),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_383),
.A2(n_302),
.B(n_250),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_366),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_405),
.A2(n_291),
.B(n_340),
.Y(n_435)
);

OAI21xp33_ASAP7_75t_L g436 ( 
.A1(n_377),
.A2(n_291),
.B(n_294),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_358),
.Y(n_438)
);

NAND2xp33_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_359),
.Y(n_439)
);

O2A1O1Ixp5_ASAP7_75t_L g440 ( 
.A1(n_374),
.A2(n_401),
.B(n_358),
.C(n_355),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_365),
.B(n_291),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_368),
.B(n_34),
.Y(n_442)
);

OAI21xp33_ASAP7_75t_L g443 ( 
.A1(n_381),
.A2(n_9),
.B(n_10),
.Y(n_443)
);

AOI22x1_ASAP7_75t_L g444 ( 
.A1(n_372),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_444)
);

BUFx12f_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_376),
.B(n_35),
.Y(n_446)
);

NAND2x1p5_ASAP7_75t_L g447 ( 
.A(n_391),
.B(n_37),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_385),
.B(n_11),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_395),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_397),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_378),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g452 ( 
.A1(n_385),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_386),
.B(n_38),
.Y(n_453)
);

BUFx2_ASAP7_75t_L g454 ( 
.A(n_363),
.Y(n_454)
);

INVx3_ASAP7_75t_L g455 ( 
.A(n_387),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_407),
.A2(n_409),
.B(n_406),
.Y(n_456)
);

BUFx8_ASAP7_75t_L g457 ( 
.A(n_367),
.Y(n_457)
);

O2A1O1Ixp5_ASAP7_75t_L g458 ( 
.A1(n_390),
.A2(n_91),
.B(n_165),
.C(n_164),
.Y(n_458)
);

AOI33xp33_ASAP7_75t_L g459 ( 
.A1(n_373),
.A2(n_14),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.B3(n_18),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_407),
.A2(n_87),
.B(n_162),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_382),
.B(n_15),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_393),
.Y(n_462)
);

O2A1O1Ixp33_ASAP7_75t_L g463 ( 
.A1(n_375),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_463)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_412),
.A2(n_99),
.B(n_161),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_363),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_399),
.B(n_39),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_413),
.A2(n_98),
.B(n_160),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_411),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_402),
.A2(n_388),
.B(n_404),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_357),
.A2(n_85),
.B1(n_159),
.B2(n_157),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_410),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_L g473 ( 
.A1(n_357),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_408),
.A2(n_417),
.B(n_361),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_357),
.A2(n_84),
.B(n_155),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_415),
.B(n_174),
.Y(n_476)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_414),
.A2(n_20),
.B(n_21),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_363),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_354),
.A2(n_100),
.B(n_40),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_414),
.A2(n_102),
.B(n_42),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_379),
.B(n_104),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_359),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_443),
.A2(n_83),
.B1(n_43),
.B2(n_45),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_418),
.B(n_22),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_47),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_428),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_420),
.B(n_48),
.Y(n_487)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_420),
.A2(n_49),
.B(n_50),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g489 ( 
.A1(n_432),
.A2(n_52),
.B(n_53),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_437),
.B(n_54),
.Y(n_490)
);

OAI21x1_ASAP7_75t_L g491 ( 
.A1(n_456),
.A2(n_55),
.B(n_56),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_L g492 ( 
.A1(n_440),
.A2(n_57),
.B(n_59),
.Y(n_492)
);

AOI221x1_ASAP7_75t_L g493 ( 
.A1(n_419),
.A2(n_480),
.B1(n_475),
.B2(n_441),
.C(n_436),
.Y(n_493)
);

AO31x2_ASAP7_75t_L g494 ( 
.A1(n_477),
.A2(n_60),
.A3(n_64),
.B(n_65),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_472),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g496 ( 
.A(n_482),
.Y(n_496)
);

BUFx2_ASAP7_75t_L g497 ( 
.A(n_457),
.Y(n_497)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_421),
.A2(n_438),
.B(n_429),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_462),
.Y(n_499)
);

NAND2x1p5_ASAP7_75t_L g500 ( 
.A(n_423),
.B(n_70),
.Y(n_500)
);

AO31x2_ASAP7_75t_L g501 ( 
.A1(n_473),
.A2(n_71),
.A3(n_73),
.B(n_74),
.Y(n_501)
);

INVx2_ASAP7_75t_SL g502 ( 
.A(n_423),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_469),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_452),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_449),
.B(n_80),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_430),
.A2(n_81),
.B(n_105),
.Y(n_506)
);

INVx5_ASAP7_75t_L g507 ( 
.A(n_423),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g508 ( 
.A1(n_419),
.A2(n_108),
.B(n_110),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_450),
.B(n_112),
.Y(n_509)
);

O2A1O1Ixp5_ASAP7_75t_L g510 ( 
.A1(n_426),
.A2(n_113),
.B(n_114),
.C(n_118),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_468),
.B(n_119),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_439),
.B(n_122),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_470),
.A2(n_123),
.B(n_128),
.Y(n_513)
);

INVx4_ASAP7_75t_L g514 ( 
.A(n_455),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_451),
.B(n_130),
.Y(n_515)
);

OAI21x1_ASAP7_75t_L g516 ( 
.A1(n_453),
.A2(n_154),
.B(n_132),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_478),
.B(n_131),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_442),
.A2(n_133),
.B(n_134),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_455),
.B(n_135),
.Y(n_519)
);

INVx4_ASAP7_75t_L g520 ( 
.A(n_447),
.Y(n_520)
);

OAI21x1_ASAP7_75t_L g521 ( 
.A1(n_466),
.A2(n_152),
.B(n_138),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_454),
.B(n_137),
.Y(n_522)
);

AO31x2_ASAP7_75t_L g523 ( 
.A1(n_473),
.A2(n_139),
.A3(n_142),
.B(n_143),
.Y(n_523)
);

OAI21x1_ASAP7_75t_L g524 ( 
.A1(n_446),
.A2(n_433),
.B(n_458),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_474),
.B(n_461),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_448),
.B(n_476),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_431),
.B(n_435),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_463),
.A2(n_144),
.B(n_145),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_459),
.B(n_148),
.Y(n_529)
);

A2O1A1Ixp33_ASAP7_75t_L g530 ( 
.A1(n_471),
.A2(n_149),
.B(n_151),
.C(n_479),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_447),
.B(n_481),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_444),
.Y(n_532)
);

OAI21x1_ASAP7_75t_L g533 ( 
.A1(n_464),
.A2(n_467),
.B(n_460),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_465),
.B(n_427),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_422),
.B(n_425),
.Y(n_535)
);

AOI21xp5_ASAP7_75t_L g536 ( 
.A1(n_457),
.A2(n_434),
.B(n_445),
.Y(n_536)
);

INVx2_ASAP7_75t_SL g537 ( 
.A(n_482),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_418),
.B(n_360),
.Y(n_539)
);

AOI21xp5_ASAP7_75t_L g540 ( 
.A1(n_420),
.A2(n_421),
.B(n_418),
.Y(n_540)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_514),
.Y(n_541)
);

NAND2x1p5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_508),
.Y(n_542)
);

OAI22xp33_ASAP7_75t_L g543 ( 
.A1(n_483),
.A2(n_507),
.B1(n_539),
.B2(n_496),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_529),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_514),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_527),
.A2(n_504),
.B1(n_484),
.B2(n_528),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g547 ( 
.A1(n_493),
.A2(n_540),
.B(n_492),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_502),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_503),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_489),
.A2(n_528),
.B(n_525),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_483),
.A2(n_511),
.B1(n_517),
.B2(n_532),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_513),
.A2(n_533),
.B(n_524),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_532),
.B(n_486),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g554 ( 
.A(n_507),
.Y(n_554)
);

OA21x2_ASAP7_75t_L g555 ( 
.A1(n_506),
.A2(n_491),
.B(n_487),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_507),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_538),
.Y(n_558)
);

AOI21x1_ASAP7_75t_L g559 ( 
.A1(n_485),
.A2(n_531),
.B(n_498),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_522),
.Y(n_560)
);

AO31x2_ASAP7_75t_L g561 ( 
.A1(n_530),
.A2(n_495),
.A3(n_520),
.B(n_526),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_486),
.Y(n_562)
);

AO21x2_ASAP7_75t_L g563 ( 
.A1(n_535),
.A2(n_515),
.B(n_488),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_510),
.A2(n_516),
.B(n_521),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g565 ( 
.A1(n_490),
.A2(n_509),
.B1(n_505),
.B2(n_512),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_499),
.Y(n_566)
);

O2A1O1Ixp33_ASAP7_75t_SL g567 ( 
.A1(n_519),
.A2(n_518),
.B(n_499),
.C(n_494),
.Y(n_567)
);

O2A1O1Ixp33_ASAP7_75t_L g568 ( 
.A1(n_500),
.A2(n_534),
.B(n_536),
.C(n_497),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_501),
.B(n_523),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_494),
.A2(n_501),
.B(n_523),
.Y(n_570)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_501),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_494),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_523),
.B(n_367),
.Y(n_573)
);

INVx4_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_SL g575 ( 
.A1(n_530),
.A2(n_418),
.B(n_539),
.C(n_531),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_527),
.B(n_507),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_503),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g578 ( 
.A1(n_493),
.A2(n_540),
.B(n_419),
.Y(n_578)
);

BUFx2_ASAP7_75t_L g579 ( 
.A(n_496),
.Y(n_579)
);

NAND2x1p5_ASAP7_75t_L g580 ( 
.A(n_520),
.B(n_508),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_527),
.B(n_507),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_486),
.Y(n_582)
);

OA21x2_ASAP7_75t_L g583 ( 
.A1(n_493),
.A2(n_540),
.B(n_419),
.Y(n_583)
);

OAI211xp5_ASAP7_75t_L g584 ( 
.A1(n_483),
.A2(n_377),
.B(n_381),
.C(n_301),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_527),
.B(n_371),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_557),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_557),
.Y(n_587)
);

OR2x2_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_584),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_541),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_548),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_577),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_577),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_553),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_553),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_549),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_562),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_562),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_582),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_582),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_566),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_544),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_585),
.B(n_551),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_581),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_548),
.Y(n_605)
);

O2A1O1Ixp5_ASAP7_75t_L g606 ( 
.A1(n_565),
.A2(n_559),
.B(n_543),
.C(n_569),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_546),
.A2(n_560),
.B1(n_581),
.B2(n_576),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_579),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_579),
.Y(n_609)
);

OA21x2_ASAP7_75t_L g610 ( 
.A1(n_570),
.A2(n_572),
.B(n_552),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_541),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_576),
.B(n_581),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_576),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_541),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_558),
.A2(n_554),
.B1(n_556),
.B2(n_574),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g616 ( 
.A(n_569),
.B(n_550),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_556),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_545),
.Y(n_618)
);

AOI22xp5_ASAP7_75t_SL g619 ( 
.A1(n_558),
.A2(n_574),
.B1(n_550),
.B2(n_569),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_545),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_545),
.Y(n_621)
);

INVx3_ASAP7_75t_L g622 ( 
.A(n_574),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_572),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_575),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_568),
.B(n_542),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_626),
.B(n_542),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_595),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_603),
.B(n_550),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_595),
.Y(n_630)
);

HB1xp67_ASAP7_75t_L g631 ( 
.A(n_608),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_590),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_591),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_609),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_612),
.Y(n_637)
);

INVx2_ASAP7_75t_SL g638 ( 
.A(n_609),
.Y(n_638)
);

INVxp67_ASAP7_75t_L g639 ( 
.A(n_605),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_603),
.B(n_561),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_612),
.B(n_561),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_604),
.B(n_561),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_592),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_604),
.B(n_561),
.Y(n_644)
);

NAND2x1_ASAP7_75t_L g645 ( 
.A(n_626),
.B(n_555),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_593),
.B(n_561),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_592),
.Y(n_647)
);

INVx2_ASAP7_75t_R g648 ( 
.A(n_624),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_593),
.B(n_583),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_594),
.B(n_583),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_623),
.Y(n_652)
);

OR2x2_ASAP7_75t_L g653 ( 
.A(n_588),
.B(n_578),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_594),
.B(n_571),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_596),
.B(n_571),
.Y(n_655)
);

HB1xp67_ASAP7_75t_L g656 ( 
.A(n_617),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_601),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_613),
.B(n_567),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_586),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_600),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_622),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_615),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_601),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_L g664 ( 
.A1(n_607),
.A2(n_547),
.B1(n_580),
.B2(n_542),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_599),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_597),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_597),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_598),
.Y(n_669)
);

OR2x2_ASAP7_75t_L g670 ( 
.A(n_653),
.B(n_588),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_642),
.B(n_602),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_653),
.B(n_629),
.Y(n_672)
);

INVxp67_ASAP7_75t_L g673 ( 
.A(n_631),
.Y(n_673)
);

NOR2x1_ASAP7_75t_L g674 ( 
.A(n_636),
.B(n_626),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_639),
.B(n_632),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_633),
.B(n_602),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_628),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_652),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_656),
.B(n_598),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_659),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_634),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_636),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_637),
.B(n_625),
.Y(n_684)
);

AND2x2_ASAP7_75t_L g685 ( 
.A(n_640),
.B(n_616),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_640),
.B(n_616),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_644),
.B(n_629),
.Y(n_687)
);

AND2x4_ASAP7_75t_SL g688 ( 
.A(n_637),
.B(n_626),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_635),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_662),
.A2(n_619),
.B1(n_622),
.B2(n_589),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_637),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_644),
.B(n_646),
.Y(n_692)
);

INVxp67_ASAP7_75t_SL g693 ( 
.A(n_665),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_643),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_646),
.B(n_641),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_647),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_659),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_637),
.B(n_614),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_666),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_637),
.B(n_614),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_627),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_652),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_657),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_657),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_641),
.B(n_610),
.Y(n_705)
);

HB1xp67_ASAP7_75t_L g706 ( 
.A(n_638),
.Y(n_706)
);

BUFx3_ASAP7_75t_L g707 ( 
.A(n_638),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_649),
.B(n_610),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_673),
.B(n_663),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_678),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_675),
.B(n_663),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_706),
.Y(n_712)
);

HB1xp67_ASAP7_75t_L g713 ( 
.A(n_683),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_687),
.B(n_650),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_687),
.B(n_650),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_692),
.B(n_649),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_678),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_671),
.B(n_651),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_692),
.B(n_648),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_695),
.B(n_648),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_702),
.Y(n_721)
);

BUFx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_682),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_689),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_685),
.B(n_654),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_701),
.B(n_627),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_694),
.Y(n_727)
);

INVxp67_ASAP7_75t_SL g728 ( 
.A(n_693),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_696),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_677),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_685),
.B(n_654),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_681),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_707),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_686),
.B(n_627),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_672),
.B(n_670),
.Y(n_735)
);

NOR3xp33_ASAP7_75t_L g736 ( 
.A(n_690),
.B(n_658),
.C(n_606),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_672),
.B(n_670),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_699),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_703),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_704),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_679),
.B(n_660),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_710),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_717),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_721),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_719),
.B(n_705),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_723),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_724),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_719),
.B(n_705),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_713),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_727),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_729),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_735),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_730),
.Y(n_753)
);

INVx3_ASAP7_75t_L g754 ( 
.A(n_726),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_726),
.B(n_701),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_732),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_726),
.Y(n_757)
);

AOI21xp33_ASAP7_75t_L g758 ( 
.A1(n_718),
.A2(n_684),
.B(n_676),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_720),
.B(n_708),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_728),
.B(n_686),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_738),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_711),
.B(n_707),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_735),
.Y(n_763)
);

O2A1O1Ixp33_ASAP7_75t_SL g764 ( 
.A1(n_762),
.A2(n_733),
.B(n_712),
.C(n_709),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_744),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_752),
.Y(n_766)
);

NOR2xp33_ASAP7_75t_L g767 ( 
.A(n_763),
.B(n_722),
.Y(n_767)
);

INVx1_ASAP7_75t_SL g768 ( 
.A(n_760),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_749),
.B(n_737),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_759),
.B(n_737),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_754),
.A2(n_701),
.B1(n_688),
.B2(n_722),
.Y(n_771)
);

OAI21xp5_ASAP7_75t_L g772 ( 
.A1(n_758),
.A2(n_736),
.B(n_741),
.Y(n_772)
);

OAI221xp5_ASAP7_75t_L g773 ( 
.A1(n_746),
.A2(n_740),
.B1(n_739),
.B2(n_731),
.C(n_725),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_744),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_767),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_766),
.B(n_757),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_765),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_767),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_774),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_770),
.Y(n_780)
);

OAI22xp5_ASAP7_75t_L g781 ( 
.A1(n_772),
.A2(n_731),
.B1(n_725),
.B2(n_701),
.Y(n_781)
);

NAND3xp33_ASAP7_75t_L g782 ( 
.A(n_781),
.B(n_764),
.C(n_773),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_775),
.B(n_768),
.Y(n_783)
);

OA22x2_ASAP7_75t_L g784 ( 
.A1(n_778),
.A2(n_771),
.B1(n_769),
.B2(n_754),
.Y(n_784)
);

AOI222xp33_ASAP7_75t_L g785 ( 
.A1(n_781),
.A2(n_761),
.B1(n_747),
.B2(n_756),
.C1(n_753),
.C2(n_734),
.Y(n_785)
);

OAI221xp5_ASAP7_75t_L g786 ( 
.A1(n_776),
.A2(n_757),
.B1(n_754),
.B2(n_750),
.C(n_743),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_780),
.A2(n_755),
.B1(n_757),
.B2(n_701),
.Y(n_787)
);

NAND4xp25_ASAP7_75t_L g788 ( 
.A(n_782),
.B(n_777),
.C(n_779),
.D(n_734),
.Y(n_788)
);

NAND4xp25_ASAP7_75t_L g789 ( 
.A(n_785),
.B(n_691),
.C(n_750),
.D(n_755),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_784),
.B(n_745),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_783),
.B(n_751),
.C(n_698),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_787),
.B(n_786),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_792),
.A2(n_751),
.B(n_755),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_788),
.B(n_748),
.Y(n_794)
);

NOR4xp75_ASAP7_75t_L g795 ( 
.A(n_790),
.B(n_700),
.C(n_645),
.D(n_745),
.Y(n_795)
);

NAND4xp75_ASAP7_75t_L g796 ( 
.A(n_793),
.B(n_794),
.C(n_795),
.D(n_789),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_794),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_793),
.B(n_791),
.Y(n_798)
);

OAI21xp5_ASAP7_75t_L g799 ( 
.A1(n_798),
.A2(n_742),
.B(n_655),
.Y(n_799)
);

XNOR2xp5_ASAP7_75t_L g800 ( 
.A(n_797),
.B(n_796),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_798),
.B(n_742),
.Y(n_801)
);

XOR2xp5_ASAP7_75t_L g802 ( 
.A(n_796),
.B(n_691),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_797),
.B(n_748),
.Y(n_803)
);

BUFx2_ASAP7_75t_L g804 ( 
.A(n_802),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_803),
.Y(n_805)
);

OAI22x1_ASAP7_75t_L g806 ( 
.A1(n_800),
.A2(n_759),
.B1(n_720),
.B2(n_669),
.Y(n_806)
);

OAI22xp5_ASAP7_75t_L g807 ( 
.A1(n_799),
.A2(n_688),
.B1(n_627),
.B2(n_715),
.Y(n_807)
);

NAND5xp2_ASAP7_75t_L g808 ( 
.A(n_801),
.B(n_655),
.C(n_667),
.D(n_668),
.E(n_580),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_R g809 ( 
.A(n_804),
.B(n_661),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_805),
.B(n_714),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_806),
.B(n_714),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_808),
.Y(n_812)
);

INVxp67_ASAP7_75t_L g813 ( 
.A(n_812),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_SL g814 ( 
.A1(n_810),
.A2(n_807),
.B1(n_645),
.B2(n_580),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_811),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_809),
.Y(n_816)
);

AO21x2_ASAP7_75t_L g817 ( 
.A1(n_809),
.A2(n_563),
.B(n_621),
.Y(n_817)
);

OAI21xp5_ASAP7_75t_L g818 ( 
.A1(n_813),
.A2(n_664),
.B(n_618),
.Y(n_818)
);

AOI21x1_ASAP7_75t_L g819 ( 
.A1(n_816),
.A2(n_621),
.B(n_620),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_815),
.B(n_715),
.Y(n_820)
);

OR2x2_ASAP7_75t_L g821 ( 
.A(n_817),
.B(n_716),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_820),
.A2(n_814),
.B1(n_697),
.B2(n_680),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_821),
.A2(n_563),
.B(n_564),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_819),
.Y(n_824)
);

XNOR2x1_ASAP7_75t_L g825 ( 
.A(n_824),
.B(n_818),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_L g826 ( 
.A1(n_825),
.A2(n_822),
.B1(n_823),
.B2(n_661),
.Y(n_826)
);

AOI221xp5_ASAP7_75t_L g827 ( 
.A1(n_826),
.A2(n_661),
.B1(n_620),
.B2(n_618),
.C(n_611),
.Y(n_827)
);


endmodule