module fake_jpeg_30428_n_447 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_447);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_447;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g19 ( 
.A(n_18),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_18),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

CKINVDCx5p33_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_47),
.Y(n_95)
);

BUFx12_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_25),
.B(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_49),
.B(n_52),
.Y(n_122)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_50),
.Y(n_137)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_53),
.B(n_58),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_21),
.Y(n_55)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_57),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_25),
.B(n_17),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_59),
.B(n_61),
.Y(n_136)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_22),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_70),
.Y(n_97)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_28),
.Y(n_68)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_71),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_32),
.Y(n_72)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_73),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_76),
.Y(n_102)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_26),
.B(n_8),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_79),
.B(n_92),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_36),
.Y(n_81)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_36),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_85),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_40),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_39),
.Y(n_140)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

BUFx12f_ASAP7_75t_L g128 ( 
.A(n_88),
.Y(n_128)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_89),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_33),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_90),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_91),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_26),
.B(n_7),
.Y(n_92)
);

OAI21xp33_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_41),
.B(n_23),
.Y(n_103)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_103),
.A2(n_30),
.B(n_23),
.C(n_48),
.Y(n_163)
);

CKINVDCx11_ASAP7_75t_R g114 ( 
.A(n_48),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_114),
.Y(n_165)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_84),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_120),
.B(n_126),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_81),
.B(n_29),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_121),
.B(n_27),
.Y(n_172)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_69),
.A2(n_20),
.B1(n_46),
.B2(n_19),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_135),
.A2(n_20),
.B1(n_61),
.B2(n_42),
.Y(n_153)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_139),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_39),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_112),
.Y(n_146)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_146),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_151),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_148),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_67),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_149),
.B(n_158),
.Y(n_200)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_141),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_150),
.Y(n_198)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_31),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_97),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_152),
.B(n_154),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_172),
.B1(n_27),
.B2(n_46),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_97),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_95),
.Y(n_155)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_155),
.Y(n_194)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_118),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_118),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_117),
.B(n_64),
.C(n_73),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_66),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_159),
.B(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_111),
.Y(n_160)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_108),
.Y(n_161)
);

CKINVDCx12_ASAP7_75t_R g162 ( 
.A(n_93),
.Y(n_162)
);

BUFx24_ASAP7_75t_L g193 ( 
.A(n_162),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_163),
.A2(n_178),
.B1(n_103),
.B2(n_140),
.Y(n_195)
);

INVx8_ASAP7_75t_L g164 ( 
.A(n_98),
.Y(n_164)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_138),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_124),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_167),
.Y(n_204)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_168),
.B(n_169),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g169 ( 
.A(n_127),
.Y(n_169)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_102),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_171),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_115),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.Y(n_185)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_101),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_31),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_175),
.B(n_177),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_105),
.B(n_63),
.Y(n_176)
);

AND2x2_ASAP7_75t_SL g205 ( 
.A(n_176),
.B(n_109),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_132),
.B(n_29),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g178 ( 
.A(n_133),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_176),
.A2(n_121),
.B1(n_116),
.B2(n_94),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_180),
.A2(n_190),
.B1(n_203),
.B2(n_113),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_159),
.B(n_132),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_192),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_91),
.B1(n_85),
.B2(n_83),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_122),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_197),
.Y(n_216)
);

OA22x2_ASAP7_75t_L g203 ( 
.A1(n_163),
.A2(n_99),
.B1(n_131),
.B2(n_134),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_187),
.B(n_151),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_208),
.B(n_222),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_209),
.Y(n_236)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_212),
.Y(n_254)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_213),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_192),
.B(n_149),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_214),
.B(n_215),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_200),
.B(n_149),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_158),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_217),
.B(n_229),
.C(n_205),
.Y(n_242)
);

OR2x6_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_176),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_218),
.A2(n_201),
.B(n_203),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_150),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_220),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_189),
.B(n_145),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_155),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_221),
.B(n_226),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_183),
.B(n_144),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_223),
.Y(n_247)
);

OAI32xp33_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_160),
.A3(n_146),
.B1(n_143),
.B2(n_166),
.Y(n_224)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_224),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_225),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_186),
.B(n_143),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_227),
.A2(n_82),
.B1(n_99),
.B2(n_131),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g228 ( 
.A(n_194),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_195),
.C(n_205),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_173),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_165),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_231),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_230),
.A2(n_218),
.B(n_229),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_257),
.Y(n_264)
);

OR2x2_ASAP7_75t_SL g265 ( 
.A(n_233),
.B(n_207),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_218),
.A2(n_180),
.B1(n_203),
.B2(n_190),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_238),
.A2(n_213),
.B1(n_217),
.B2(n_214),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_242),
.B(n_207),
.C(n_220),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_218),
.A2(n_198),
.B1(n_204),
.B2(n_191),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_246),
.A2(n_250),
.B1(n_255),
.B2(n_256),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_198),
.B(n_199),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_249),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_216),
.A2(n_227),
.B1(n_211),
.B2(n_218),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_204),
.B1(n_191),
.B2(n_206),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_219),
.A2(n_215),
.B(n_216),
.Y(n_253)
);

INVx13_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g255 ( 
.A1(n_224),
.A2(n_164),
.B1(n_129),
.B2(n_123),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_209),
.A2(n_129),
.B1(n_113),
.B2(n_156),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_202),
.B(n_206),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_254),
.Y(n_258)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_258),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_237),
.B(n_222),
.Y(n_259)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_259),
.Y(n_289)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_261),
.A2(n_238),
.B1(n_240),
.B2(n_196),
.Y(n_301)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_265),
.A2(n_196),
.B(n_178),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_266),
.Y(n_309)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_236),
.Y(n_268)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_268),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_274),
.C(n_276),
.Y(n_290)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_241),
.Y(n_270)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_270),
.Y(n_315)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_243),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_271),
.B(n_277),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_237),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_278),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_242),
.B(n_221),
.C(n_226),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_287),
.B1(n_249),
.B2(n_248),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_231),
.C(n_188),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

NOR3xp33_ASAP7_75t_L g278 ( 
.A(n_243),
.B(n_212),
.C(n_210),
.Y(n_278)
);

MAJx2_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_193),
.C(n_188),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_232),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_245),
.B(n_212),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_280),
.B(n_283),
.Y(n_291)
);

BUFx6f_ASAP7_75t_SL g281 ( 
.A(n_256),
.Y(n_281)
);

INVxp33_ASAP7_75t_L g295 ( 
.A(n_281),
.Y(n_295)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_246),
.B(n_251),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_282),
.B(n_72),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_210),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_284),
.B(n_234),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_239),
.B(n_223),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_285),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_SL g286 ( 
.A(n_240),
.B(n_252),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g293 ( 
.A(n_286),
.B(n_244),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_248),
.A2(n_235),
.B1(n_255),
.B2(n_250),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_288),
.A2(n_314),
.B1(n_316),
.B2(n_171),
.Y(n_337)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_281),
.A2(n_244),
.B1(n_253),
.B2(n_246),
.Y(n_294)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_294),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_296),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_297),
.B(n_305),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_274),
.B(n_233),
.C(n_257),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_276),
.C(n_264),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_301),
.B(n_303),
.Y(n_328)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_284),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_304),
.A2(n_313),
.B(n_194),
.Y(n_334)
);

MAJx2_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_193),
.C(n_107),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_168),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_307),
.B(n_279),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_258),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_312),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_282),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_287),
.A2(n_182),
.B1(n_184),
.B2(n_157),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_263),
.A2(n_184),
.B1(n_182),
.B2(n_46),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g317 ( 
.A(n_311),
.Y(n_317)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_317),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_318),
.B(n_323),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_301),
.A2(n_272),
.B1(n_312),
.B2(n_262),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_319),
.A2(n_303),
.B1(n_292),
.B2(n_295),
.Y(n_356)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_264),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_296),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_325),
.B(n_338),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_268),
.Y(n_326)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_326),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_327),
.B(n_90),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_290),
.B(n_265),
.C(n_270),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_329),
.B(n_330),
.C(n_339),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_290),
.B(n_267),
.C(n_272),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_291),
.B(n_271),
.Y(n_331)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_300),
.A2(n_267),
.B(n_161),
.Y(n_332)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_332),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_334),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_179),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_336),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_337),
.A2(n_306),
.B1(n_310),
.B2(n_309),
.Y(n_352)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_293),
.B(n_7),
.C(n_14),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_299),
.B(n_305),
.C(n_307),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_181),
.C(n_167),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_341),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_288),
.B(n_181),
.C(n_104),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_321),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_345),
.B(n_349),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_314),
.B1(n_313),
.B2(n_315),
.Y(n_346)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_346),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_333),
.A2(n_328),
.B1(n_335),
.B2(n_327),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_355),
.Y(n_365)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_334),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_330),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_169),
.Y(n_376)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_340),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_359),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_322),
.Y(n_357)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_357),
.Y(n_378)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_319),
.A2(n_295),
.B1(n_298),
.B2(n_174),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_362),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_341),
.A2(n_42),
.B1(n_56),
.B2(n_54),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_323),
.B(n_318),
.Y(n_366)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_366),
.Y(n_385)
);

BUFx12_ASAP7_75t_L g368 ( 
.A(n_350),
.Y(n_368)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_368),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_351),
.B(n_339),
.C(n_324),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_371),
.B(n_382),
.C(n_364),
.Y(n_392)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_354),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_372),
.B(n_375),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_361),
.A2(n_324),
.B(n_30),
.Y(n_373)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_373),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_358),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g398 ( 
.A(n_376),
.B(n_169),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_350),
.B(n_9),
.Y(n_377)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_377),
.Y(n_390)
);

INVx3_ASAP7_75t_L g380 ( 
.A(n_360),
.Y(n_380)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_380),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_355),
.B(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_381),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_142),
.C(n_106),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_347),
.Y(n_383)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_383),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g384 ( 
.A(n_343),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_384),
.A2(n_348),
.B1(n_342),
.B2(n_359),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_388),
.B(n_398),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_375),
.A2(n_369),
.B1(n_370),
.B2(n_367),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_391),
.A2(n_377),
.B1(n_368),
.B2(n_98),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_392),
.B(n_367),
.C(n_382),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_371),
.B(n_353),
.C(n_364),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_393),
.A2(n_397),
.B(n_380),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_381),
.B(n_342),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_396),
.B(n_368),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_379),
.A2(n_110),
.B(n_130),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_400),
.B(n_401),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_395),
.A2(n_378),
.B1(n_366),
.B2(n_374),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_402),
.B(n_412),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_399),
.A2(n_365),
.B(n_373),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_403),
.A2(n_410),
.B(n_411),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_393),
.B(n_365),
.C(n_374),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_404),
.B(n_407),
.C(n_408),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_405),
.Y(n_423)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_398),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_392),
.B(n_385),
.C(n_396),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_42),
.C(n_51),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_387),
.A2(n_12),
.B(n_16),
.Y(n_410)
);

AOI21x1_ASAP7_75t_L g411 ( 
.A1(n_389),
.A2(n_11),
.B(n_13),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_50),
.C(n_137),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_405),
.A2(n_386),
.B(n_394),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_414),
.B(n_418),
.Y(n_426)
);

XOR2x2_ASAP7_75t_L g417 ( 
.A(n_403),
.B(n_390),
.Y(n_417)
);

INVxp33_ASAP7_75t_L g424 ( 
.A(n_417),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_409),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_419),
.B(n_421),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_410),
.B(n_88),
.C(n_128),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_88),
.C(n_128),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_422),
.B(n_416),
.Y(n_428)
);

AOI322xp5_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_41),
.A3(n_33),
.B1(n_6),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_427),
.B(n_429),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_428),
.B(n_430),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_415),
.B(n_41),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_420),
.B(n_5),
.C(n_12),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_418),
.B(n_5),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_431),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_422),
.B(n_3),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_432),
.A2(n_3),
.B(n_9),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g434 ( 
.A1(n_426),
.A2(n_417),
.B(n_413),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_438),
.Y(n_439)
);

NOR3xp33_ASAP7_75t_L g436 ( 
.A(n_424),
.B(n_425),
.C(n_421),
.Y(n_436)
);

AOI322xp5_ASAP7_75t_L g440 ( 
.A1(n_436),
.A2(n_424),
.A3(n_433),
.B1(n_437),
.B2(n_435),
.C1(n_432),
.C2(n_33),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g442 ( 
.A(n_440),
.B(n_0),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_435),
.B(n_33),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_441),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_442),
.Y(n_444)
);

NOR4xp25_ASAP7_75t_L g445 ( 
.A(n_444),
.B(n_439),
.C(n_443),
.D(n_2),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_445),
.A2(n_0),
.B1(n_1),
.B2(n_90),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_446),
.B(n_0),
.Y(n_447)
);


endmodule