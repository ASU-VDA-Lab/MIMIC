module fake_jpeg_30720_n_219 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_15),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_44),
.Y(n_75)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_16),
.B(n_15),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_47),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_23),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_16),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_34),
.Y(n_69)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_18),
.B(n_0),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_51),
.B(n_20),
.Y(n_67)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_57),
.Y(n_87)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_59),
.Y(n_84)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_67),
.Y(n_96)
);

NOR2x1_ASAP7_75t_L g64 ( 
.A(n_43),
.B(n_37),
.Y(n_64)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_64),
.B(n_78),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_28),
.B1(n_23),
.B2(n_37),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_68),
.B1(n_73),
.B2(n_80),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_58),
.A2(n_23),
.B1(n_35),
.B2(n_27),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_69),
.B(n_70),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_52),
.B(n_19),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_54),
.B(n_19),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_71),
.B(n_72),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_34),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_59),
.B1(n_56),
.B2(n_41),
.Y(n_73)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_41),
.A2(n_20),
.B(n_33),
.C(n_32),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_22),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_21),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_36),
.B1(n_30),
.B2(n_27),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_57),
.A2(n_33),
.B1(n_32),
.B2(n_24),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_100),
.Y(n_128)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_88),
.Y(n_92)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_93),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_36),
.B1(n_30),
.B2(n_24),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_117),
.B1(n_87),
.B2(n_82),
.Y(n_121)
);

AND2x6_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_18),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g134 ( 
.A1(n_97),
.A2(n_11),
.B(n_12),
.C(n_4),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_78),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_101),
.Y(n_123)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_106),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_21),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_103),
.B(n_112),
.C(n_113),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_80),
.A2(n_73),
.B(n_90),
.C(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_104),
.B(n_111),
.Y(n_127)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_83),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_105),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_84),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_108),
.B1(n_81),
.B2(n_75),
.Y(n_141)
);

OR2x6_ASAP7_75t_L g108 ( 
.A(n_87),
.B(n_1),
.Y(n_108)
);

CKINVDCx5p33_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_109),
.B(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_60),
.B(n_1),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_110),
.B(n_119),
.Y(n_130)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_3),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_65),
.B(n_3),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_74),
.B(n_9),
.Y(n_114)
);

INVx13_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_95),
.B1(n_96),
.B2(n_108),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_87),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_82),
.B1(n_62),
.B2(n_77),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_120),
.A2(n_121),
.B1(n_133),
.B2(n_138),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_141),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_110),
.B(n_82),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_139),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_62),
.B1(n_86),
.B2(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_137),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_107),
.A2(n_108),
.B(n_118),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_135),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_98),
.B(n_11),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_104),
.B1(n_93),
.B2(n_92),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_108),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_101),
.A2(n_86),
.B1(n_77),
.B2(n_81),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_119),
.B1(n_102),
.B2(n_77),
.Y(n_155)
);

XNOR2x1_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_103),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_142),
.B(n_113),
.C(n_111),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_112),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_128),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_151),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_152),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_153),
.B(n_154),
.Y(n_169)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_130),
.B(n_99),
.C(n_91),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_L g170 ( 
.A(n_156),
.B(n_158),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_112),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_133),
.Y(n_159)
);

OR2x2_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_145),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_126),
.B(n_109),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_160),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_147),
.A2(n_127),
.B(n_135),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_167),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

INVx13_ASAP7_75t_L g181 ( 
.A(n_164),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_131),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_147),
.A2(n_159),
.B(n_161),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_171),
.B(n_177),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_144),
.B(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_172),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_173),
.B(n_175),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_124),
.Y(n_175)
);

A2O1A1O1Ixp25_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_141),
.B(n_97),
.C(n_132),
.D(n_126),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_166),
.B(n_143),
.C(n_146),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_178),
.B(n_189),
.C(n_170),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_121),
.B1(n_145),
.B2(n_141),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_179),
.A2(n_180),
.B1(n_182),
.B2(n_188),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_174),
.A2(n_164),
.B1(n_163),
.B2(n_173),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_174),
.A2(n_157),
.B1(n_123),
.B2(n_156),
.Y(n_182)
);

AO221x1_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_151),
.B1(n_125),
.B2(n_136),
.C(n_105),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_125),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_172),
.B1(n_175),
.B2(n_171),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_123),
.C(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_185),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_190),
.B(n_191),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_180),
.A2(n_162),
.B(n_167),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_192),
.A2(n_197),
.B(n_184),
.C(n_168),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_194),
.B(n_184),
.Y(n_202)
);

NOR3xp33_ASAP7_75t_SL g195 ( 
.A(n_186),
.B(n_177),
.C(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_195),
.B(n_196),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_187),
.B(n_169),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_182),
.B(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_170),
.C(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_202),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_192),
.A2(n_179),
.B1(n_188),
.B2(n_185),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_203),
.B(n_204),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_194),
.B(n_168),
.Y(n_205)
);

FAx1_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_198),
.CI(n_193),
.CON(n_207),
.SN(n_207)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_181),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_207),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_203),
.A2(n_195),
.B(n_181),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_209),
.A2(n_199),
.B(n_200),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_212),
.B(n_214),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_209),
.A2(n_202),
.B(n_205),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_213),
.Y(n_215)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_6),
.A3(n_75),
.B1(n_85),
.B2(n_115),
.C1(n_201),
.C2(n_206),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_216),
.B(n_211),
.C(n_208),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_217),
.B(n_218),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_215),
.B(n_207),
.Y(n_218)
);


endmodule