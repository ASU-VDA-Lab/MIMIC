module fake_jpeg_2310_n_423 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_423);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_423;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx4f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_SL g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_2),
.Y(n_44)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_47),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_26),
.B(n_16),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_78),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

BUFx8_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_50),
.A2(n_44),
.B1(n_23),
.B2(n_33),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_26),
.B(n_15),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_52),
.B(n_81),
.Y(n_101)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_53),
.Y(n_115)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g105 ( 
.A(n_54),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_55),
.Y(n_125)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_63),
.Y(n_139)
);

INVx2_ASAP7_75t_SL g64 ( 
.A(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_64),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_69),
.Y(n_120)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_34),
.Y(n_70)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_72),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_31),
.Y(n_75)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_77),
.Y(n_106)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_20),
.Y(n_78)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_79),
.B(n_80),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_17),
.B(n_19),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_21),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_82),
.B(n_83),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_16),
.Y(n_83)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_84),
.B(n_86),
.Y(n_129)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_85),
.Y(n_117)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_31),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_90),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_39),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_88),
.Y(n_134)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_39),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_89),
.B(n_91),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_99),
.B(n_131),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_66),
.A2(n_21),
.B1(n_37),
.B2(n_40),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_51),
.A2(n_40),
.B1(n_42),
.B2(n_31),
.Y(n_114)
);

AO22x1_ASAP7_75t_SL g170 ( 
.A1(n_114),
.A2(n_122),
.B1(n_128),
.B2(n_69),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_60),
.A2(n_35),
.B1(n_21),
.B2(n_40),
.Y(n_122)
);

HAxp5_ASAP7_75t_SL g124 ( 
.A(n_45),
.B(n_24),
.CON(n_124),
.SN(n_124)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_124),
.A2(n_24),
.B(n_20),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_40),
.C(n_37),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_127),
.B(n_24),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_65),
.A2(n_56),
.B1(n_85),
.B2(n_35),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_37),
.B1(n_23),
.B2(n_44),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_32),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_136),
.B(n_137),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_32),
.Y(n_137)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_141),
.Y(n_194)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_104),
.B(n_47),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_146),
.B(n_151),
.Y(n_186)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_105),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_147),
.Y(n_196)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_148),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_25),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_154),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_98),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_158),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_126),
.B(n_25),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_25),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_169),
.Y(n_189)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_120),
.Y(n_156)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_123),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_157),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

A2O1A1Ixp33_ASAP7_75t_SL g212 ( 
.A1(n_159),
.A2(n_162),
.B(n_182),
.C(n_139),
.Y(n_212)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

A2O1A1Ixp33_ASAP7_75t_L g161 ( 
.A1(n_101),
.A2(n_33),
.B(n_64),
.C(n_28),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_161),
.B(n_163),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_127),
.A2(n_124),
.B(n_129),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_108),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_164),
.B(n_165),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_133),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_97),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_132),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_171),
.Y(n_195)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_97),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_117),
.B(n_41),
.Y(n_169)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_98),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_123),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_172),
.A2(n_173),
.B1(n_175),
.B2(n_181),
.Y(n_208)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_125),
.B(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_174),
.B(n_177),
.Y(n_197)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

AOI21xp33_ASAP7_75t_L g176 ( 
.A1(n_98),
.A2(n_41),
.B(n_20),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_SL g188 ( 
.A(n_176),
.B(n_41),
.C(n_30),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_102),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_111),
.B(n_91),
.Y(n_178)
);

AND2x2_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_111),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_100),
.B(n_62),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_179),
.B(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_102),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_140),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_139),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

OA22x2_ASAP7_75t_L g192 ( 
.A1(n_183),
.A2(n_130),
.B1(n_140),
.B2(n_107),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_187),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_188),
.B(n_198),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_152),
.A2(n_112),
.B1(n_131),
.B2(n_134),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_210),
.B1(n_163),
.B2(n_161),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_192),
.Y(n_220)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_142),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_198)
);

OAI32xp33_ASAP7_75t_L g205 ( 
.A1(n_152),
.A2(n_118),
.A3(n_119),
.B1(n_103),
.B2(n_135),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_205),
.B(n_212),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_152),
.A2(n_106),
.B1(n_76),
.B2(n_88),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_207),
.A2(n_142),
.B1(n_181),
.B2(n_154),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_162),
.A2(n_95),
.B1(n_109),
.B2(n_92),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_231),
.B1(n_233),
.B2(n_207),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_226),
.Y(n_250)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_216),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_210),
.A2(n_169),
.B1(n_170),
.B2(n_155),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_223),
.B1(n_189),
.B2(n_184),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_227),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_199),
.A2(n_153),
.B(n_149),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_212),
.B(n_188),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_170),
.B1(n_150),
.B2(n_143),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_209),
.B(n_172),
.Y(n_224)
);

INVxp33_ASAP7_75t_L g244 ( 
.A(n_224),
.Y(n_244)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_225),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_203),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_202),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_228),
.B(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_167),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_189),
.A2(n_95),
.B1(n_92),
.B2(n_109),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_186),
.A2(n_171),
.B1(n_157),
.B2(n_178),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_232),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_77),
.B1(n_67),
.B2(n_90),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_234),
.Y(n_248)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_223),
.B1(n_222),
.B2(n_229),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_236),
.A2(n_246),
.B1(n_251),
.B2(n_256),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_237),
.A2(n_239),
.B1(n_220),
.B2(n_198),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_238),
.A2(n_194),
.B(n_201),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_217),
.A2(n_195),
.B1(n_212),
.B2(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_230),
.B(n_206),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_237),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_229),
.A2(n_197),
.B1(n_212),
.B2(n_206),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_187),
.C(n_212),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_178),
.Y(n_272)
);

BUFx5_ASAP7_75t_L g249 ( 
.A(n_216),
.Y(n_249)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_249),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_222),
.A2(n_205),
.B1(n_198),
.B2(n_211),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_215),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_228),
.B(n_187),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_254),
.B(n_227),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_213),
.A2(n_198),
.B1(n_211),
.B2(n_187),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_258),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_238),
.A2(n_215),
.B(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_259),
.A2(n_270),
.B(n_273),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_220),
.B1(n_231),
.B2(n_226),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_260),
.A2(n_274),
.B1(n_243),
.B2(n_242),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g296 ( 
.A(n_262),
.B(n_272),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_L g263 ( 
.A1(n_253),
.A2(n_224),
.B(n_232),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_263),
.B(n_266),
.Y(n_298)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

OAI21xp33_ASAP7_75t_L g266 ( 
.A1(n_253),
.A2(n_233),
.B(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_247),
.Y(n_267)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_267),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_271),
.B1(n_192),
.B2(n_241),
.Y(n_287)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_208),
.B(n_190),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_239),
.A2(n_246),
.B1(n_255),
.B2(n_236),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_245),
.A2(n_255),
.B1(n_250),
.B2(n_254),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_256),
.A2(n_218),
.B1(n_192),
.B2(n_194),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_275),
.A2(n_255),
.B(n_240),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_244),
.B(n_193),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_251),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_141),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_278),
.B(n_243),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_248),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_279),
.Y(n_290)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_280),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_282),
.B(n_286),
.Y(n_309)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_284),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_278),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_273),
.A2(n_242),
.B(n_249),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_288),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_261),
.A2(n_241),
.B1(n_218),
.B2(n_192),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_173),
.C(n_166),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_289),
.B(n_272),
.C(n_262),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_147),
.B(n_145),
.Y(n_291)
);

AOI221xp5_ASAP7_75t_L g307 ( 
.A1(n_291),
.A2(n_302),
.B1(n_290),
.B2(n_280),
.C(n_282),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_271),
.A2(n_193),
.B1(n_201),
.B2(n_200),
.Y(n_293)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_293),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_261),
.A2(n_200),
.B1(n_185),
.B2(n_160),
.Y(n_295)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_295),
.Y(n_316)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_257),
.A2(n_144),
.B1(n_148),
.B2(n_156),
.Y(n_299)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

NOR2x1_ASAP7_75t_L g302 ( 
.A(n_264),
.B(n_183),
.Y(n_302)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_302),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_292),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_303),
.B(n_304),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_317),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_311),
.B1(n_288),
.B2(n_293),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_300),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_296),
.C(n_289),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_314),
.C(n_318),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_285),
.B(n_275),
.C(n_257),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_294),
.B(n_258),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_281),
.B(n_279),
.C(n_268),
.Y(n_318)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_294),
.Y(n_321)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_321),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_SL g322 ( 
.A(n_281),
.B(n_260),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g330 ( 
.A(n_322),
.B(n_291),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_297),
.B(n_270),
.C(n_274),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_283),
.B(n_175),
.C(n_265),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_283),
.B(n_265),
.C(n_168),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_298),
.B(n_182),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_326),
.B(n_299),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_309),
.A2(n_286),
.B(n_302),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g352 ( 
.A1(n_327),
.A2(n_341),
.B(n_315),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_330),
.B(n_333),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_318),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_331),
.B(n_336),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_308),
.A2(n_287),
.B1(n_284),
.B2(n_290),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_332),
.A2(n_314),
.B1(n_325),
.B2(n_312),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_334),
.A2(n_340),
.B1(n_343),
.B2(n_304),
.Y(n_355)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_335),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_317),
.B(n_295),
.Y(n_336)
);

AO21x1_ASAP7_75t_L g337 ( 
.A1(n_320),
.A2(n_277),
.B(n_301),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g363 ( 
.A(n_337),
.Y(n_363)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_319),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_339),
.Y(n_359)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_322),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_310),
.A2(n_301),
.B1(n_35),
.B2(n_139),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_313),
.A2(n_28),
.B(n_30),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_323),
.A2(n_28),
.B1(n_30),
.B2(n_79),
.Y(n_343)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_326),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_344),
.B(n_12),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g346 ( 
.A(n_316),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_346),
.B(n_336),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_324),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_347),
.A2(n_80),
.B1(n_61),
.B2(n_54),
.Y(n_362)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_351),
.Y(n_366)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_354),
.Y(n_369)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_355),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_332),
.A2(n_303),
.B1(n_306),
.B2(n_89),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_360),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_342),
.B(n_125),
.C(n_55),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_357),
.B(n_364),
.C(n_348),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_358),
.B(n_362),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_342),
.B(n_73),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_347),
.A2(n_73),
.B1(n_86),
.B2(n_75),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_361),
.A2(n_362),
.B(n_353),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_348),
.B(n_72),
.C(n_18),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_328),
.B(n_13),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_13),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_359),
.A2(n_327),
.B(n_337),
.Y(n_367)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_367),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_368),
.B(n_376),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_349),
.B(n_345),
.C(n_328),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_370),
.B(n_379),
.Y(n_385)
);

AOI211xp5_ASAP7_75t_L g372 ( 
.A1(n_363),
.A2(n_330),
.B(n_329),
.C(n_345),
.Y(n_372)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_372),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_351),
.A2(n_333),
.B(n_341),
.Y(n_373)
);

XNOR2x1_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_374),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_378),
.B(n_12),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_360),
.B(n_18),
.C(n_13),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_364),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g394 ( 
.A(n_380),
.B(n_381),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_350),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_368),
.B(n_350),
.Y(n_384)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_384),
.B(n_377),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_366),
.B(n_365),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_386),
.B(n_388),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_357),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g389 ( 
.A(n_369),
.B(n_12),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_389),
.B(n_391),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_390),
.B(n_379),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_0),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_387),
.B(n_369),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_396),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_385),
.B(n_375),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_383),
.A2(n_372),
.B(n_373),
.Y(n_397)
);

AO21x1_ASAP7_75t_L g407 ( 
.A1(n_397),
.A2(n_400),
.B(n_11),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_376),
.C(n_374),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g405 ( 
.A(n_399),
.B(n_401),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_384),
.B(n_380),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_398),
.B(n_381),
.Y(n_402)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_402),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_400),
.A2(n_390),
.B1(n_361),
.B2(n_2),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_404),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_407),
.B(n_409),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_394),
.A2(n_0),
.B(n_1),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_SL g412 ( 
.A1(n_408),
.A2(n_11),
.B(n_3),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_1),
.C(n_3),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_406),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_411)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_412),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_405),
.A2(n_1),
.B(n_6),
.Y(n_415)
);

AOI321xp33_ASAP7_75t_L g416 ( 
.A1(n_415),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C(n_11),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_416),
.B(n_417),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_410),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_418),
.B(n_402),
.C(n_414),
.Y(n_420)
);

O2A1O1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_420),
.A2(n_413),
.B(n_8),
.C(n_10),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_419),
.Y(n_422)
);

NAND2x1_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_6),
.Y(n_423)
);


endmodule