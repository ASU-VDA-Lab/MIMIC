module real_aes_17007_n_3 (n_0, n_2, n_1, n_3);
input n_0;
input n_2;
input n_1;
output n_3;
wire n_13;
wire n_4;
wire n_5;
wire n_15;
wire n_7;
wire n_8;
wire n_6;
wire n_9;
wire n_12;
wire n_14;
wire n_10;
wire n_11;
INVx2_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
AOI22xp33_ASAP7_75t_L g3 ( .A1(n_1), .A2(n_4), .B1(n_11), .B2(n_14), .Y(n_3) );
INVx1_ASAP7_75t_L g15 ( .A(n_2), .Y(n_15) );
BUFx2_ASAP7_75t_L g4 ( .A(n_5), .Y(n_4) );
INVx1_ASAP7_75t_L g13 ( .A(n_5), .Y(n_13) );
INVx2_ASAP7_75t_L g5 ( .A(n_6), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_7), .Y(n_6) );
BUFx2_ASAP7_75t_L g7 ( .A(n_8), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_9), .Y(n_8) );
INVx2_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
BUFx3_ASAP7_75t_L g11 ( .A(n_12), .Y(n_11) );
BUFx8_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
INVx1_ASAP7_75t_L g14 ( .A(n_15), .Y(n_14) );
endmodule