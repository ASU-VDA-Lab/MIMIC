module fake_jpeg_11436_n_578 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_578);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_387;
wire n_270;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_332;
wire n_92;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_14),
.Y(n_29)
);

CKINVDCx14_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_SL g37 ( 
.A(n_11),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_7),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_9),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_7),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_74),
.Y(n_127)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_59),
.Y(n_135)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

CKINVDCx12_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx16f_ASAP7_75t_L g182 ( 
.A(n_61),
.Y(n_182)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_27),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_63),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_64),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_65),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_66),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

INVx5_ASAP7_75t_L g178 ( 
.A(n_68),
.Y(n_178)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_27),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_70),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_71),
.Y(n_189)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_31),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_72),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_18),
.B(n_9),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_73),
.B(n_114),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_37),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_75),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_38),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_85),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_77),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_78),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_79),
.Y(n_194)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_31),
.Y(n_81)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_81),
.Y(n_133)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_82),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_18),
.B(n_10),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_83),
.B(n_102),
.Y(n_163)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_38),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx8_ASAP7_75t_L g157 ( 
.A(n_86),
.Y(n_157)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_48),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_87),
.Y(n_161)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_43),
.Y(n_88)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g89 ( 
.A(n_48),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_89),
.B(n_36),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_90),
.B(n_91),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_50),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_20),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_94),
.Y(n_167)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_95),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_96),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_50),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_103),
.Y(n_134)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_28),
.B(n_16),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_34),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_104),
.Y(n_148)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_32),
.Y(n_107)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_31),
.Y(n_108)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_108),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_109),
.Y(n_150)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_45),
.Y(n_111)
);

INVx11_ASAP7_75t_L g145 ( 
.A(n_111),
.Y(n_145)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_55),
.Y(n_112)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_113),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_28),
.B(n_8),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_46),
.Y(n_115)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_32),
.Y(n_116)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_116),
.Y(n_184)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_32),
.Y(n_117)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx16f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

BUFx12_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_55),
.Y(n_119)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_21),
.Y(n_120)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_121),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_106),
.A2(n_46),
.B1(n_25),
.B2(n_47),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_124),
.A2(n_154),
.B1(n_30),
.B2(n_98),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_104),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_130),
.B(n_144),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_115),
.A2(n_25),
.B1(n_47),
.B2(n_46),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_136),
.A2(n_139),
.B1(n_152),
.B2(n_96),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_109),
.A2(n_25),
.B1(n_47),
.B2(n_54),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_118),
.B(n_40),
.Y(n_144)
);

INVx11_ASAP7_75t_L g151 ( 
.A(n_89),
.Y(n_151)
);

INVx11_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_68),
.A2(n_36),
.B1(n_54),
.B2(n_55),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_92),
.B(n_40),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_153),
.B(n_164),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_154),
.B(n_95),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_49),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_72),
.B(n_29),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_168),
.B(n_175),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_81),
.B(n_39),
.Y(n_169)
);

NOR2x1_ASAP7_75t_L g220 ( 
.A(n_169),
.B(n_183),
.Y(n_220)
);

INVx11_ASAP7_75t_L g171 ( 
.A(n_82),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_171),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_108),
.B(n_29),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_119),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_176),
.B(n_67),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_84),
.B(n_39),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_121),
.B(n_49),
.Y(n_190)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_190),
.B(n_66),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_64),
.A2(n_36),
.B(n_53),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_87),
.C(n_33),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_198),
.B(n_233),
.Y(n_277)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_187),
.Y(n_199)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_199),
.Y(n_321)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_125),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_201),
.Y(n_281)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_202),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_L g204 ( 
.A1(n_163),
.A2(n_21),
.B(n_53),
.C(n_42),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_204),
.B(n_214),
.Y(n_314)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_141),
.A2(n_36),
.B1(n_26),
.B2(n_23),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_205),
.Y(n_282)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_207),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g280 ( 
.A(n_208),
.Y(n_280)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx4_ASAP7_75t_L g306 ( 
.A(n_209),
.Y(n_306)
);

CKINVDCx9p33_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

INVx4_ASAP7_75t_SL g295 ( 
.A(n_210),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_133),
.Y(n_211)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_211),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_141),
.A2(n_23),
.B1(n_26),
.B2(n_41),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_212),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_167),
.A2(n_41),
.B1(n_42),
.B2(n_94),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_213),
.A2(n_251),
.B1(n_252),
.B2(n_256),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_134),
.B(n_196),
.Y(n_214)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_215),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_142),
.B(n_52),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_216),
.B(n_217),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_160),
.B(n_52),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g218 ( 
.A(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_218),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_219),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_222),
.A2(n_265),
.B1(n_266),
.B2(n_194),
.Y(n_311)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_224),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_177),
.B(n_51),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_225),
.B(n_226),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_131),
.B(n_51),
.Y(n_226)
);

CKINVDCx12_ASAP7_75t_R g227 ( 
.A(n_182),
.Y(n_227)
);

INVx4_ASAP7_75t_SL g307 ( 
.A(n_227),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

INVx8_ASAP7_75t_L g267 ( 
.A(n_228),
.Y(n_267)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_229),
.Y(n_289)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_230),
.Y(n_302)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_148),
.Y(n_231)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_231),
.Y(n_320)
);

OAI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_152),
.A2(n_173),
.B1(n_167),
.B2(n_186),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_232),
.A2(n_178),
.B1(n_143),
.B2(n_126),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_137),
.B(n_55),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_146),
.B(n_0),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_234),
.B(n_249),
.Y(n_308)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_184),
.A2(n_70),
.B1(n_79),
.B2(n_78),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_236),
.A2(n_239),
.B1(n_260),
.B2(n_210),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_145),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_238),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_62),
.B1(n_65),
.B2(n_97),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_128),
.B(n_35),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_159),
.B(n_35),
.Y(n_241)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_195),
.Y(n_242)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_242),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g243 ( 
.A(n_145),
.Y(n_243)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_243),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_244),
.A2(n_198),
.B(n_234),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_155),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_245),
.B(n_247),
.Y(n_290)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_195),
.Y(n_246)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_246),
.Y(n_310)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_123),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g248 ( 
.A(n_155),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_248),
.B(n_250),
.Y(n_298)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_126),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_135),
.B(n_33),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_161),
.A2(n_111),
.B1(n_101),
.B2(n_75),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_156),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_147),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_253),
.B(n_254),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_165),
.B(n_30),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_181),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_255),
.B(n_257),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_156),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_185),
.B(n_13),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_122),
.B(n_129),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_258),
.B(n_264),
.Y(n_316)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_147),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_261),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_123),
.Y(n_261)
);

CKINVDCx12_ASAP7_75t_R g262 ( 
.A(n_138),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_263),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_161),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_170),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_188),
.A2(n_86),
.B1(n_77),
.B2(n_71),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g268 ( 
.A(n_244),
.B(n_179),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_268),
.B(n_198),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_296),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_283),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_241),
.B(n_162),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_286),
.B(n_305),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_157),
.B1(n_180),
.B2(n_173),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_292),
.A2(n_299),
.B1(n_221),
.B2(n_203),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_266),
.A2(n_172),
.B1(n_132),
.B2(n_194),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g334 ( 
.A1(n_293),
.A2(n_301),
.B1(n_312),
.B2(n_315),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_223),
.A2(n_178),
.B1(n_143),
.B2(n_188),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_221),
.B(n_203),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_220),
.A2(n_174),
.B(n_0),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_236),
.A2(n_180),
.B1(n_157),
.B2(n_191),
.Y(n_299)
);

OAI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_222),
.A2(n_172),
.B1(n_192),
.B2(n_191),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_220),
.B(n_234),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_311),
.B(n_243),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_200),
.A2(n_192),
.B1(n_189),
.B2(n_170),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_240),
.A2(n_189),
.B1(n_3),
.B2(n_4),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_204),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_318),
.B(n_2),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_319),
.B(n_268),
.C(n_277),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_324),
.B(n_310),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_325),
.B(n_363),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_280),
.B(n_206),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_326),
.B(n_341),
.Y(n_373)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_274),
.Y(n_327)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_328),
.A2(n_347),
.B(n_348),
.Y(n_367)
);

INVx13_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g384 ( 
.A(n_329),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_314),
.B(n_233),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_SL g386 ( 
.A(n_330),
.B(n_279),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_290),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_331),
.B(n_346),
.Y(n_382)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_273),
.Y(n_332)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_332),
.Y(n_370)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_333),
.B(n_335),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_233),
.C(n_258),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_274),
.Y(n_336)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_336),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_277),
.B(n_258),
.C(n_211),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_337),
.B(n_359),
.Y(n_371)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_273),
.Y(n_338)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_338),
.Y(n_394)
);

INVx13_ASAP7_75t_L g339 ( 
.A(n_307),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_339),
.Y(n_383)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_275),
.Y(n_340)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_276),
.B(n_211),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_342),
.A2(n_293),
.B1(n_316),
.B2(n_310),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_286),
.B(n_218),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_343),
.B(n_345),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_272),
.B(n_218),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_313),
.Y(n_346)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_282),
.A2(n_261),
.B(n_199),
.Y(n_348)
);

CKINVDCx6p67_ASAP7_75t_R g349 ( 
.A(n_307),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_349),
.B(n_350),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_317),
.Y(n_350)
);

INVx13_ASAP7_75t_L g351 ( 
.A(n_300),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g376 ( 
.A(n_351),
.B(n_353),
.Y(n_376)
);

AOI32xp33_ASAP7_75t_L g352 ( 
.A1(n_305),
.A2(n_237),
.A3(n_215),
.B1(n_259),
.B2(n_253),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g378 ( 
.A1(n_352),
.A2(n_296),
.B(n_285),
.Y(n_378)
);

BUFx12f_ASAP7_75t_L g353 ( 
.A(n_300),
.Y(n_353)
);

INVx13_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_354),
.B(n_356),
.Y(n_381)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_275),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_355),
.B(n_357),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_276),
.B(n_219),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_272),
.B(n_229),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g358 ( 
.A1(n_314),
.A2(n_231),
.B(n_219),
.C(n_249),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_294),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_277),
.B(n_224),
.C(n_207),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_271),
.B(n_247),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_360),
.B(n_361),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_308),
.B(n_230),
.Y(n_361)
);

CKINVDCx10_ASAP7_75t_R g362 ( 
.A(n_295),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_362),
.B(n_297),
.Y(n_398)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_316),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_334),
.A2(n_269),
.B1(n_283),
.B2(n_282),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_365),
.A2(n_369),
.B1(n_374),
.B2(n_388),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_334),
.A2(n_278),
.B1(n_285),
.B2(n_309),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_344),
.A2(n_352),
.B1(n_345),
.B2(n_357),
.Y(n_374)
);

OAI21xp33_ASAP7_75t_SL g423 ( 
.A1(n_377),
.A2(n_325),
.B(n_349),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_378),
.B(n_379),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_323),
.A2(n_304),
.B(n_298),
.Y(n_379)
);

XNOR2x1_ASAP7_75t_SL g380 ( 
.A(n_333),
.B(n_308),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_335),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_324),
.B(n_308),
.Y(n_385)
);

XNOR2x1_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_392),
.Y(n_413)
);

CKINVDCx14_ASAP7_75t_R g411 ( 
.A(n_386),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_387),
.A2(n_355),
.B1(n_336),
.B2(n_327),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_344),
.A2(n_201),
.B1(n_256),
.B2(n_252),
.Y(n_388)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_323),
.A2(n_316),
.B(n_318),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_390),
.B(n_328),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_L g395 ( 
.A(n_322),
.B(n_295),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_395),
.B(n_397),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_343),
.B(n_291),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_398),
.B(n_349),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_322),
.B(n_291),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_337),
.C(n_359),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_410),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_389),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_401),
.B(n_409),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_377),
.A2(n_323),
.B1(n_363),
.B2(n_347),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_402),
.B(n_417),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_SL g403 ( 
.A(n_386),
.B(n_347),
.C(n_330),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_403),
.B(n_416),
.Y(n_449)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_404),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_374),
.A2(n_346),
.B1(n_342),
.B2(n_331),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_406),
.A2(n_425),
.B1(n_387),
.B2(n_393),
.Y(n_433)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_407),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_408),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_350),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_410),
.B(n_412),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_368),
.B(n_361),
.C(n_348),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g441 ( 
.A(n_415),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_382),
.B(n_340),
.Y(n_416)
);

AND2x6_ASAP7_75t_L g417 ( 
.A(n_380),
.B(n_358),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_366),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_418),
.B(n_420),
.Y(n_442)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_384),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_419),
.Y(n_444)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_396),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_396),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_421),
.Y(n_462)
);

MAJx2_ASAP7_75t_L g422 ( 
.A(n_368),
.B(n_349),
.C(n_362),
.Y(n_422)
);

MAJx2_ASAP7_75t_L g455 ( 
.A(n_422),
.B(n_385),
.C(n_399),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_423),
.A2(n_367),
.B(n_390),
.Y(n_440)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_397),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_426),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_369),
.A2(n_281),
.B1(n_267),
.B2(n_332),
.Y(n_425)
);

AND2x6_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_378),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_391),
.B(n_288),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_427),
.B(n_428),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_381),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_372),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_395),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_371),
.B(n_288),
.C(n_270),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_431),
.B(n_432),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_371),
.B(n_270),
.C(n_284),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_433),
.A2(n_447),
.B1(n_448),
.B2(n_457),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_435),
.B(n_413),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_429),
.B(n_372),
.Y(n_438)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_438),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_SL g481 ( 
.A1(n_440),
.A2(n_445),
.B(n_452),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_414),
.A2(n_367),
.B(n_429),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_405),
.A2(n_364),
.B1(n_375),
.B2(n_365),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_405),
.A2(n_406),
.B1(n_424),
.B2(n_430),
.Y(n_448)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

NOR2x1_ASAP7_75t_L g452 ( 
.A(n_402),
.B(n_364),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_400),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_431),
.B(n_375),
.Y(n_456)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_456),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_425),
.A2(n_393),
.B1(n_392),
.B2(n_388),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_411),
.A2(n_383),
.B1(n_384),
.B2(n_394),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_458),
.A2(n_419),
.B1(n_297),
.B2(n_267),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_404),
.B(n_394),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_459),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_420),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_460),
.B(n_320),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g461 ( 
.A1(n_414),
.A2(n_383),
.B(n_376),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_461),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_463),
.B(n_465),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_451),
.B(n_432),
.C(n_412),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_466),
.B(n_474),
.C(n_476),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_SL g467 ( 
.A(n_436),
.B(n_414),
.C(n_426),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g510 ( 
.A1(n_467),
.A2(n_471),
.B(n_483),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_449),
.B(n_353),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_468),
.B(n_469),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_449),
.B(n_353),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_SL g471 ( 
.A(n_443),
.B(n_403),
.C(n_417),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_439),
.A2(n_422),
.B1(n_413),
.B2(n_370),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_472),
.A2(n_475),
.B1(n_478),
.B2(n_479),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g474 ( 
.A(n_451),
.B(n_370),
.C(n_321),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_446),
.B(n_435),
.C(n_456),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g478 ( 
.A1(n_441),
.A2(n_353),
.B1(n_321),
.B2(n_303),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_448),
.A2(n_281),
.B1(n_338),
.B2(n_264),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_437),
.A2(n_354),
.B1(n_228),
.B2(n_329),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_480),
.A2(n_444),
.B1(n_462),
.B2(n_454),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_482),
.B(n_437),
.Y(n_503)
);

AOI22x1_ASAP7_75t_L g483 ( 
.A1(n_450),
.A2(n_354),
.B1(n_329),
.B2(n_339),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_434),
.B(n_306),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_484),
.B(n_486),
.Y(n_493)
);

CKINVDCx16_ASAP7_75t_R g486 ( 
.A(n_458),
.Y(n_486)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_488),
.Y(n_497)
);

FAx1_ASAP7_75t_SL g489 ( 
.A(n_467),
.B(n_436),
.CI(n_443),
.CON(n_489),
.SN(n_489)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_489),
.B(n_500),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_463),
.B(n_446),
.Y(n_490)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_490),
.B(n_502),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g492 ( 
.A(n_475),
.Y(n_492)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_476),
.B(n_461),
.C(n_455),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_496),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_445),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_495),
.B(n_499),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_487),
.B(n_453),
.Y(n_496)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_477),
.Y(n_498)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_498),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_472),
.B(n_440),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_474),
.B(n_433),
.C(n_457),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_501),
.A2(n_481),
.B1(n_483),
.B2(n_303),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_465),
.B(n_447),
.C(n_459),
.Y(n_502)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_503),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_473),
.B(n_460),
.C(n_442),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_507),
.A2(n_351),
.B1(n_320),
.B2(n_289),
.Y(n_522)
);

A2O1A1Ixp33_ASAP7_75t_L g508 ( 
.A1(n_485),
.A2(n_452),
.B(n_438),
.C(n_442),
.Y(n_508)
);

OAI321xp33_ASAP7_75t_L g513 ( 
.A1(n_508),
.A2(n_481),
.A3(n_470),
.B1(n_483),
.B2(n_479),
.C(n_482),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_470),
.B(n_452),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_509),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_506),
.A2(n_464),
.B1(n_473),
.B2(n_454),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g533 ( 
.A(n_512),
.B(n_516),
.Y(n_533)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_513),
.Y(n_530)
);

INVxp33_ASAP7_75t_L g514 ( 
.A(n_493),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_525),
.Y(n_532)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_515),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_492),
.A2(n_246),
.B1(n_306),
.B2(n_242),
.Y(n_516)
);

BUFx12_ASAP7_75t_L g520 ( 
.A(n_489),
.Y(n_520)
);

CKINVDCx16_ASAP7_75t_R g539 ( 
.A(n_520),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_522),
.B(n_497),
.Y(n_540)
);

BUFx24_ASAP7_75t_SL g525 ( 
.A(n_489),
.Y(n_525)
);

AOI22x1_ASAP7_75t_L g526 ( 
.A1(n_508),
.A2(n_289),
.B1(n_287),
.B2(n_302),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_526),
.B(n_507),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_528),
.B(n_519),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_518),
.B(n_491),
.C(n_490),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_531),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_491),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_523),
.B(n_500),
.C(n_495),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_535),
.B(n_536),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_523),
.B(n_494),
.C(n_510),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_517),
.B(n_502),
.C(n_509),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_537),
.A2(n_541),
.B(n_527),
.Y(n_542)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_524),
.B(n_504),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g545 ( 
.A(n_538),
.B(n_519),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_540),
.A2(n_514),
.B1(n_521),
.B2(n_520),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_511),
.B(n_505),
.C(n_499),
.Y(n_541)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_548),
.Y(n_553)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_544),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_545),
.B(n_549),
.Y(n_555)
);

BUFx24_ASAP7_75t_SL g546 ( 
.A(n_530),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g559 ( 
.A(n_546),
.B(n_552),
.Y(n_559)
);

XNOR2x1_ASAP7_75t_SL g548 ( 
.A(n_541),
.B(n_505),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_534),
.B(n_520),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_550),
.B(n_551),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_529),
.B(n_526),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g552 ( 
.A(n_535),
.B(n_287),
.C(n_302),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_544),
.A2(n_539),
.B1(n_536),
.B2(n_537),
.Y(n_554)
);

OR2x2_ASAP7_75t_L g567 ( 
.A(n_554),
.B(n_561),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_543),
.B(n_532),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_560),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_533),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_SL g561 ( 
.A(n_549),
.B(n_303),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_557),
.A2(n_238),
.B1(n_209),
.B2(n_263),
.Y(n_562)
);

AO21x1_ASAP7_75t_L g570 ( 
.A1(n_562),
.A2(n_559),
.B(n_8),
.Y(n_570)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_553),
.A2(n_303),
.B(n_243),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_563),
.A2(n_566),
.B(n_556),
.Y(n_568)
);

XNOR2x1_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_237),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g571 ( 
.A(n_565),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_2),
.C(n_5),
.Y(n_566)
);

AOI21xp33_ASAP7_75t_L g573 ( 
.A1(n_568),
.A2(n_569),
.B(n_570),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_564),
.B(n_555),
.Y(n_569)
);

AOI322xp5_ASAP7_75t_L g572 ( 
.A1(n_571),
.A2(n_564),
.A3(n_567),
.B1(n_11),
.B2(n_12),
.C1(n_13),
.C2(n_7),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g574 ( 
.A(n_572),
.B(n_8),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g575 ( 
.A(n_574),
.B(n_573),
.C(n_13),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_575),
.A2(n_11),
.B1(n_14),
.B2(n_15),
.Y(n_576)
);

OAI21xp33_ASAP7_75t_L g577 ( 
.A1(n_576),
.A2(n_15),
.B(n_16),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_15),
.B(n_16),
.Y(n_578)
);


endmodule