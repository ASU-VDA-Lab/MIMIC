module fake_jpeg_23795_n_64 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_64);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_64;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_3),
.Y(n_8)
);

CKINVDCx20_ASAP7_75t_R g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_1),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g20 ( 
.A1(n_8),
.A2(n_0),
.B1(n_7),
.B2(n_5),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_20),
.B(n_21),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g21 ( 
.A(n_8),
.B(n_4),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_11),
.B1(n_18),
.B2(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_21),
.B(n_14),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_17),
.B(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g35 ( 
.A(n_27),
.B(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_26),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_28),
.B(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_24),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_34),
.Y(n_41)
);

XNOR2x2_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_13),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_32),
.B1(n_35),
.B2(n_16),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_16),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_24),
.A2(n_5),
.B(n_6),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_22),
.A2(n_15),
.B(n_9),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_23),
.B(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_36),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_42),
.B(n_12),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_44),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_31),
.C(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_47),
.B(n_50),
.C(n_41),
.Y(n_51)
);

FAx1_ASAP7_75t_SL g49 ( 
.A(n_42),
.B(n_32),
.CI(n_12),
.CON(n_49),
.SN(n_49)
);

XNOR2x1_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_45),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_54),
.C(n_46),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_48),
.A2(n_45),
.B1(n_38),
.B2(n_39),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_52),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_53),
.B(n_47),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_56),
.A2(n_49),
.B1(n_12),
.B2(n_7),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_54),
.C(n_46),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_59),
.C(n_49),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_55),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_SL g63 ( 
.A1(n_62),
.A2(n_61),
.B(n_6),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_63),
.B(n_12),
.Y(n_64)
);


endmodule