module fake_jpeg_23583_n_332 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_332);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_332;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_SL g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_41),
.B(n_43),
.Y(n_69)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_20),
.B(n_8),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_46),
.Y(n_67)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_48),
.B(n_49),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_27),
.B(n_0),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_51),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_52),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_19),
.B1(n_35),
.B2(n_32),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_56),
.B1(n_61),
.B2(n_72),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_19),
.B1(n_35),
.B2(n_32),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_29),
.Y(n_60)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_39),
.A2(n_35),
.B1(n_32),
.B2(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx11_ASAP7_75t_L g98 ( 
.A(n_62),
.Y(n_98)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_64),
.Y(n_115)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_66),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_27),
.B1(n_37),
.B2(n_24),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_45),
.A2(n_37),
.B1(n_24),
.B2(n_20),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_78),
.B1(n_81),
.B2(n_84),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_42),
.A2(n_37),
.B1(n_24),
.B2(n_38),
.Y(n_78)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_79),
.Y(n_119)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_80),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_45),
.A2(n_20),
.B1(n_22),
.B2(n_17),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_82),
.Y(n_104)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_83),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_38),
.B1(n_17),
.B2(n_23),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_49),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_93),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

BUFx2_ASAP7_75t_SL g136 ( 
.A(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_76),
.B(n_49),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_54),
.A2(n_21),
.B1(n_26),
.B2(n_38),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_96),
.A2(n_101),
.B1(n_112),
.B2(n_9),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_81),
.B(n_48),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_97),
.B(n_99),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_53),
.B(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_53),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_22),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_21),
.B1(n_17),
.B2(n_23),
.Y(n_101)
);

AOI21xp33_ASAP7_75t_SL g102 ( 
.A1(n_83),
.A2(n_25),
.B(n_50),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g150 ( 
.A1(n_102),
.A2(n_113),
.B(n_118),
.C(n_7),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_61),
.A2(n_51),
.B1(n_23),
.B2(n_26),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_103),
.A2(n_26),
.B1(n_31),
.B2(n_28),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_57),
.B(n_50),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_109),
.C(n_56),
.Y(n_139)
);

AND2x4_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_25),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_108),
.A2(n_70),
.B(n_33),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_43),
.C(n_36),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_52),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_114),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_73),
.A2(n_22),
.B1(n_36),
.B2(n_34),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_69),
.A2(n_43),
.B(n_34),
.C(n_31),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_55),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_67),
.B(n_66),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_116),
.B(n_117),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_33),
.Y(n_117)
);

OR2x2_ASAP7_75t_SL g118 ( 
.A(n_64),
.B(n_11),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_52),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_121),
.B(n_79),
.Y(n_130)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_124),
.B(n_127),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_125),
.B(n_88),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_126),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g127 ( 
.A(n_86),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_128),
.A2(n_148),
.B1(n_156),
.B2(n_118),
.Y(n_170)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_115),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_134),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_130),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_28),
.B(n_33),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_131),
.A2(n_138),
.B(n_106),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_33),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_145),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g137 ( 
.A(n_108),
.B(n_15),
.Y(n_137)
);

A2O1A1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_137),
.A2(n_149),
.B(n_128),
.C(n_138),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_105),
.A2(n_33),
.B(n_1),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_121),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_114),
.A2(n_82),
.B1(n_80),
.B2(n_75),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_140),
.A2(n_87),
.B1(n_119),
.B2(n_94),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_108),
.A2(n_68),
.B1(n_77),
.B2(n_75),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_141),
.Y(n_175)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_143),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g143 ( 
.A(n_109),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_144),
.B(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_99),
.B(n_97),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_97),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_89),
.B(n_65),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_147),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_87),
.A2(n_77),
.B1(n_68),
.B2(n_62),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_149),
.A2(n_150),
.B(n_113),
.Y(n_161)
);

AO21x2_ASAP7_75t_L g151 ( 
.A1(n_85),
.A2(n_70),
.B(n_1),
.Y(n_151)
);

OAI22x1_ASAP7_75t_L g181 ( 
.A1(n_151),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_0),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_153),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_91),
.B(n_0),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_104),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_186),
.B(n_190),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g193 ( 
.A1(n_162),
.A2(n_170),
.B1(n_181),
.B2(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_132),
.B(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_167),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_120),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_151),
.A2(n_90),
.B1(n_106),
.B2(n_104),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_168),
.A2(n_140),
.B1(n_151),
.B2(n_142),
.Y(n_192)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_145),
.B(n_91),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_171),
.B(n_173),
.Y(n_212)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_126),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_176),
.Y(n_219)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_178),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_151),
.A2(n_94),
.B1(n_98),
.B2(n_90),
.Y(n_179)
);

CKINVDCx14_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_182),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_123),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_183),
.B(n_107),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_124),
.C(n_144),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_185),
.B(n_10),
.Y(n_220)
);

OAI31xp33_ASAP7_75t_L g206 ( 
.A1(n_187),
.A2(n_152),
.A3(n_129),
.B(n_95),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_95),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_122),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_133),
.B(n_2),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_191),
.B(n_150),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_192),
.A2(n_193),
.B1(n_200),
.B2(n_207),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_188),
.B(n_133),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_194),
.A2(n_202),
.B(n_206),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_195),
.B(n_177),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_197),
.A2(n_221),
.B(n_222),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_122),
.Y(n_199)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_175),
.A2(n_155),
.B1(n_139),
.B2(n_135),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_158),
.B(n_131),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_164),
.B(n_153),
.Y(n_204)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_172),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_205),
.B(n_210),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_181),
.A2(n_162),
.B1(n_183),
.B2(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_209),
.Y(n_242)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_180),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_211),
.B(n_218),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_88),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_213),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g216 ( 
.A(n_173),
.B(n_10),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_165),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_220),
.B(n_185),
.C(n_171),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_158),
.B(n_111),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_217),
.A2(n_175),
.B(n_163),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_223),
.A2(n_245),
.B1(n_215),
.B2(n_203),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_224),
.B(n_237),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_219),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_226),
.B(n_233),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_173),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_243),
.Y(n_249)
);

AOI31xp33_ASAP7_75t_SL g231 ( 
.A1(n_216),
.A2(n_161),
.A3(n_187),
.B(n_190),
.Y(n_231)
);

NAND3xp33_ASAP7_75t_L g252 ( 
.A(n_231),
.B(n_196),
.C(n_222),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_235),
.B(n_241),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_192),
.A2(n_168),
.B1(n_166),
.B2(n_174),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_238),
.A2(n_239),
.B1(n_244),
.B2(n_221),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_197),
.A2(n_166),
.B1(n_174),
.B2(n_176),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_219),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_208),
.A2(n_184),
.B(n_159),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_199),
.A2(n_169),
.B1(n_178),
.B2(n_111),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_218),
.A2(n_189),
.B1(n_2),
.B2(n_4),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_203),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_189),
.C(n_2),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_204),
.C(n_202),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_200),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_251),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_231),
.B(n_208),
.Y(n_251)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_243),
.C(n_237),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_253),
.A2(n_254),
.B1(n_267),
.B2(n_229),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_232),
.A2(n_206),
.B1(n_211),
.B2(n_196),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_220),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_260),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_256),
.B(n_257),
.C(n_258),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_194),
.C(n_202),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_227),
.B(n_194),
.C(n_205),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_240),
.B(n_210),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_244),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_225),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_236),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_239),
.B(n_198),
.Y(n_263)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_263),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_227),
.A2(n_201),
.B1(n_198),
.B2(n_214),
.Y(n_265)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_265),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_238),
.A2(n_201),
.B1(n_214),
.B2(n_5),
.Y(n_267)
);

AO21x1_ASAP7_75t_L g298 ( 
.A1(n_270),
.A2(n_3),
.B(n_4),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_271),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_266),
.B(n_230),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_272),
.B(n_279),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_273),
.A2(n_285),
.B1(n_242),
.B2(n_264),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_247),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_275),
.B(n_284),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g277 ( 
.A1(n_263),
.A2(n_236),
.B(n_223),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_282),
.B(n_230),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_233),
.Y(n_279)
);

XNOR2x1_ASAP7_75t_L g281 ( 
.A(n_260),
.B(n_234),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_281),
.B(n_251),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_229),
.B(n_225),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_256),
.B(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_283),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_234),
.Y(n_284)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_281),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_297),
.Y(n_302)
);

NAND2xp67_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_252),
.Y(n_287)
);

FAx1_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_298),
.CI(n_270),
.CON(n_304),
.SN(n_304)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_289),
.B(n_295),
.C(n_296),
.Y(n_301)
);

OAI221xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_280),
.B1(n_274),
.B2(n_269),
.C(n_284),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_276),
.B(n_249),
.C(n_255),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_249),
.Y(n_296)
);

INVx13_ASAP7_75t_L g299 ( 
.A(n_268),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_282),
.Y(n_300)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_295),
.B(n_276),
.C(n_269),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_303),
.B(n_307),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_298),
.Y(n_310)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_287),
.A2(n_274),
.B(n_6),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_309),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_5),
.C(n_12),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_291),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_308),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_14),
.C(n_15),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_310),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_317),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_302),
.A2(n_299),
.B1(n_289),
.B2(n_288),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_306),
.A2(n_296),
.B1(n_288),
.B2(n_16),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_SL g318 ( 
.A(n_315),
.B(n_301),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_318),
.A2(n_316),
.B(n_313),
.Y(n_323)
);

OR2x2_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_14),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_321),
.A2(n_311),
.B(n_312),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_323),
.B(n_324),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_322),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_325),
.B(n_317),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_320),
.C(n_310),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g329 ( 
.A(n_328),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_329),
.A2(n_326),
.B(n_319),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_15),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_331),
.B(n_16),
.Y(n_332)
);


endmodule