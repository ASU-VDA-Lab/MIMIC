module fake_ariane_1437_n_2442 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_225, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_226, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_224, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_229, n_70, n_222, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_227, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_232, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_228, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_231, n_192, n_28, n_80, n_146, n_230, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_223, n_35, n_54, n_25, n_2442);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_225;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_226;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_224;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_229;
input n_70;
input n_222;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_227;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_232;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_228;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_231;
input n_192;
input n_28;
input n_80;
input n_146;
input n_230;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_223;
input n_35;
input n_54;
input n_25;

output n_2442;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1507;
wire n_1486;
wire n_1938;
wire n_589;
wire n_1174;
wire n_2346;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2334;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_2407;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_717;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_2436;
wire n_2376;
wire n_2367;
wire n_1706;
wire n_2207;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_2374;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_2380;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_279;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_2288;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_2323;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_2317;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2342;
wire n_2200;
wire n_259;
wire n_953;
wire n_1364;
wire n_2390;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_2322;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_2370;
wire n_495;
wire n_267;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2359;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_2301;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_2433;
wire n_352;
wire n_899;
wire n_1703;
wire n_2332;
wire n_2391;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_2427;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_1924;
wire n_438;
wire n_1654;
wire n_1560;
wire n_2341;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_2382;
wire n_237;
wire n_2043;
wire n_780;
wire n_2349;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2326;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_2245;
wire n_249;
wire n_1108;
wire n_851;
wire n_444;
wire n_355;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_2426;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_2398;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_2415;
wire n_436;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_274;
wire n_1083;
wire n_337;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_2439;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2365;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_2333;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_2435;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_2293;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_2400;
wire n_632;
wire n_477;
wire n_650;
wire n_2388;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1908;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_2302;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_2294;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_2363;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_2328;
wire n_347;
wire n_2434;
wire n_1042;
wire n_1234;
wire n_2311;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_2287;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_2438;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_2335;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2404;
wire n_2168;
wire n_552;
wire n_348;
wire n_2312;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_720;
wire n_926;
wire n_1943;
wire n_2296;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2146;
wire n_1868;
wire n_1501;
wire n_2241;
wire n_2373;
wire n_1173;
wire n_2350;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_2327;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_2437;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_2399;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_600;
wire n_481;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_677;
wire n_604;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_874;
wire n_2286;
wire n_2023;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_2418;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_2338;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_321;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_2379;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_2300;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_2284;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_2366;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_2292;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_2306;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_2424;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2414;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2337;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_1804;
wire n_2106;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_2348;
wire n_1281;
wire n_516;
wire n_2364;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_2307;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_2295;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_2412;
wire n_374;
wire n_1352;
wire n_2405;
wire n_1824;
wire n_643;
wire n_1492;
wire n_2383;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_2416;
wire n_819;
wire n_2386;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_2353;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_2325;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_2298;
wire n_1149;
wire n_1505;
wire n_2408;
wire n_2320;
wire n_979;
wire n_2329;
wire n_1642;
wire n_2417;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_2354;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_2368;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_2352;
wire n_1256;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_354;
wire n_725;
wire n_2377;
wire n_1577;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2410;
wire n_2314;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2203;
wire n_2133;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_2001;
wire n_1047;
wire n_1472;
wire n_2413;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_2285;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_2403;
wire n_1367;
wire n_2044;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_2310;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_1511;
wire n_2177;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_2343;
wire n_775;
wire n_667;
wire n_2419;
wire n_1049;
wire n_2330;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_2411;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_2309;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_2431;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_2401;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_2331;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_810;
wire n_1290;
wire n_1959;
wire n_617;
wire n_2396;
wire n_543;
wire n_1362;
wire n_1559;
wire n_2121;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_2371;
wire n_1978;
wire n_571;
wire n_414;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_2313;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_2303;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2441;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_540;
wire n_692;
wire n_2054;
wire n_1857;
wire n_2315;
wire n_984;
wire n_1687;
wire n_2073;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1910;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_2093;
wire n_2340;
wire n_2018;
wire n_1772;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_2305;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_2428;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_2425;
wire n_2394;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_2356;
wire n_1601;
wire n_1057;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_2385;
wire n_2387;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_2291;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_2402;
wire n_318;
wire n_1458;
wire n_679;
wire n_244;
wire n_1630;
wire n_663;
wire n_1720;
wire n_2409;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_2344;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_2392;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_2321;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_2000;
wire n_1268;
wire n_385;
wire n_2395;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2440;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1323;
wire n_1235;
wire n_2375;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_2420;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_2358;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_2355;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_2324;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_2397;
wire n_369;
wire n_240;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_2351;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_2347;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_2362;
wire n_1615;
wire n_1236;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_2372;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_2422;
wire n_1334;
wire n_654;
wire n_2290;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2429;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_2339;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_838;
wire n_383;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_2360;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_2432;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_2430;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_2297;
wire n_371;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_2381;
wire n_1967;
wire n_2384;
wire n_2179;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2205;
wire n_2183;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2357;
wire n_2029;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_2421;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_2318;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_2361;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_2316;
wire n_1010;
wire n_882;
wire n_2304;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_548;
wire n_289;
wire n_2336;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2319;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_2345;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_180),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_178),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_166),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_218),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_0),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_106),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_151),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_35),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_162),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_205),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_216),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_195),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_20),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_160),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_48),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_62),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_124),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_214),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_35),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_110),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_99),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_185),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_93),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_44),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_58),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_188),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_78),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_155),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_219),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_112),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_9),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_147),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_172),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_140),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_119),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_93),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_108),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_31),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_176),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_42),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_189),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_34),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_69),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_114),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_152),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_157),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_196),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_92),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_105),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_38),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_22),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_204),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_26),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_22),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_133),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_1),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

BUFx8_ASAP7_75t_SL g298 ( 
.A(n_44),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_19),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_83),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_202),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_25),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_229),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_210),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_182),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_215),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_14),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_49),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_130),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_111),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_39),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_103),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_137),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_23),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_144),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_63),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_34),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_127),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_26),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_154),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_65),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_37),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_6),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_161),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_164),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_65),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_31),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_19),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_90),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_163),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_121),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_63),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_199),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_168),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_7),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_132),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_120),
.Y(n_338)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_58),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_194),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_95),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_86),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_191),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_126),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_125),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_105),
.Y(n_346)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_21),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_33),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_217),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_30),
.Y(n_350)
);

CKINVDCx14_ASAP7_75t_R g351 ( 
.A(n_156),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_1),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_208),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_16),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_141),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_29),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_21),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_181),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_36),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_66),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_97),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_77),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_139),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_17),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_118),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_223),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_222),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_82),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_23),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_116),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_173),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_39),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_76),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_30),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_11),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_54),
.Y(n_376)
);

CKINVDCx14_ASAP7_75t_R g377 ( 
.A(n_212),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_170),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_82),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_103),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_158),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_165),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_4),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_198),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_60),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_177),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_37),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_104),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_24),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_122),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_56),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_206),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_150),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_49),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_184),
.Y(n_395)
);

CKINVDCx16_ASAP7_75t_R g396 ( 
.A(n_42),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_131),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_129),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_128),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_200),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_2),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_7),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_203),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_134),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_99),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_43),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_95),
.Y(n_407)
);

BUFx6f_ASAP7_75t_L g408 ( 
.A(n_29),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_87),
.Y(n_409)
);

BUFx5_ASAP7_75t_L g410 ( 
.A(n_169),
.Y(n_410)
);

BUFx10_ASAP7_75t_L g411 ( 
.A(n_104),
.Y(n_411)
);

BUFx10_ASAP7_75t_L g412 ( 
.A(n_32),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_16),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_53),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_153),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_66),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_80),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_142),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_90),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_98),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_56),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_232),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_230),
.Y(n_423)
);

CKINVDCx14_ASAP7_75t_R g424 ( 
.A(n_107),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_60),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_53),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_113),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_201),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_9),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_70),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_149),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_179),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_186),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_227),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_45),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g437 ( 
.A(n_74),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_59),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_81),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_89),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_41),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_192),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_64),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_61),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_38),
.Y(n_445)
);

INVx2_ASAP7_75t_SL g446 ( 
.A(n_96),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_94),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_15),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_97),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_51),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_84),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_67),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_6),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_3),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_71),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_91),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_145),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_413),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_0),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_298),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_413),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_233),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_255),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

CKINVDCx14_ASAP7_75t_R g466 ( 
.A(n_351),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_413),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_336),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_353),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_433),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_239),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_253),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_413),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_413),
.Y(n_474)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_275),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_413),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_314),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_413),
.Y(n_478)
);

INVxp67_ASAP7_75t_SL g479 ( 
.A(n_439),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_316),
.Y(n_480)
);

NOR2xp67_ASAP7_75t_L g481 ( 
.A(n_234),
.B(n_339),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_437),
.Y(n_482)
);

NOR2xp67_ASAP7_75t_L g483 ( 
.A(n_234),
.B(n_2),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_437),
.Y(n_484)
);

INVxp33_ASAP7_75t_SL g485 ( 
.A(n_254),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_259),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_257),
.B(n_3),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_437),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_242),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_437),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_437),
.Y(n_493)
);

INVxp67_ASAP7_75t_SL g494 ( 
.A(n_449),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_263),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_437),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_437),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_449),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_341),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_241),
.Y(n_501)
);

INVxp33_ASAP7_75t_SL g502 ( 
.A(n_266),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_402),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_241),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_270),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_409),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_441),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_243),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_271),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_276),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_245),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_443),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_278),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_280),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_282),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_377),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_245),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_246),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_246),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_424),
.Y(n_520)
);

INVxp33_ASAP7_75t_SL g521 ( 
.A(n_283),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_247),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g523 ( 
.A(n_408),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_247),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_339),
.B(n_4),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_258),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_258),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_288),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_260),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_260),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_268),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_268),
.B(n_272),
.Y(n_532)
);

CKINVDCx14_ASAP7_75t_R g533 ( 
.A(n_287),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_408),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_287),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_272),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_294),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_274),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_408),
.Y(n_539)
);

CKINVDCx20_ASAP7_75t_R g540 ( 
.A(n_287),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_287),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_296),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_274),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_300),
.Y(n_544)
);

INVxp67_ASAP7_75t_L g545 ( 
.A(n_242),
.Y(n_545)
);

BUFx2_ASAP7_75t_L g546 ( 
.A(n_446),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_251),
.Y(n_547)
);

BUFx3_ASAP7_75t_L g548 ( 
.A(n_284),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_277),
.Y(n_549)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_284),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_277),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_286),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_243),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_286),
.Y(n_554)
);

BUFx6f_ASAP7_75t_SL g555 ( 
.A(n_422),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_307),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_295),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_295),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_251),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_301),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_308),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_301),
.B(n_5),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_305),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_311),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_305),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_306),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_312),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_306),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_243),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_330),
.B(n_5),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_330),
.Y(n_571)
);

CKINVDCx16_ASAP7_75t_R g572 ( 
.A(n_411),
.Y(n_572)
);

INVxp33_ASAP7_75t_SL g573 ( 
.A(n_319),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_411),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_321),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_338),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_338),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_343),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_343),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_408),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_344),
.Y(n_581)
);

NOR2xp67_ASAP7_75t_L g582 ( 
.A(n_501),
.B(n_422),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_463),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_468),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_458),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_458),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_461),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_534),
.Y(n_588)
);

BUFx6f_ASAP7_75t_L g589 ( 
.A(n_534),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_461),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_469),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_470),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_464),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_462),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_460),
.Y(n_595)
);

AND2x4_ASAP7_75t_SL g596 ( 
.A(n_550),
.B(n_411),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_462),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_539),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_503),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_477),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_465),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_539),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_499),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_580),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_475),
.B(n_248),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_465),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g607 ( 
.A(n_480),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_467),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_467),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_473),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_473),
.Y(n_611)
);

NAND2xp33_ASAP7_75t_SL g612 ( 
.A(n_459),
.B(n_535),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_474),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_471),
.Y(n_614)
);

INVx3_ASAP7_75t_L g615 ( 
.A(n_580),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_474),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_551),
.B(n_579),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_476),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_551),
.B(n_579),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_500),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_501),
.B(n_504),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_478),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_482),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_506),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_482),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_472),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_484),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_484),
.Y(n_630)
);

BUFx8_ASAP7_75t_L g631 ( 
.A(n_555),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_548),
.B(n_344),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_488),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_486),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_523),
.B(n_345),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_488),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_507),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_489),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_489),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_555),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_495),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_492),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_492),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_493),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_505),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_509),
.Y(n_646)
);

BUFx6f_ASAP7_75t_L g647 ( 
.A(n_493),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_510),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_496),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_513),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_514),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_496),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_497),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_497),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_498),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_515),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_528),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_512),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_537),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_548),
.B(n_446),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_498),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_516),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_504),
.B(n_453),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_511),
.Y(n_664)
);

CKINVDCx16_ASAP7_75t_R g665 ( 
.A(n_508),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_511),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_542),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_517),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_491),
.Y(n_669)
);

CKINVDCx20_ASAP7_75t_R g670 ( 
.A(n_520),
.Y(n_670)
);

NAND2xp33_ASAP7_75t_R g671 ( 
.A(n_544),
.B(n_323),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_517),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_518),
.B(n_519),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_518),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_519),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_522),
.B(n_257),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_556),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_522),
.Y(n_678)
);

BUFx3_ASAP7_75t_L g679 ( 
.A(n_672),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_674),
.Y(n_680)
);

INVx2_ASAP7_75t_SL g681 ( 
.A(n_617),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_617),
.B(n_533),
.Y(n_682)
);

AND2x4_ASAP7_75t_L g683 ( 
.A(n_617),
.B(n_479),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_605),
.B(n_485),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_618),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_596),
.B(n_459),
.Y(n_686)
);

INVx1_ASAP7_75t_SL g687 ( 
.A(n_599),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_673),
.B(n_524),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_618),
.Y(n_689)
);

INVxp67_ASAP7_75t_SL g690 ( 
.A(n_674),
.Y(n_690)
);

BUFx3_ASAP7_75t_L g691 ( 
.A(n_672),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_SL g692 ( 
.A1(n_596),
.A2(n_541),
.B1(n_540),
.B2(n_553),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_619),
.B(n_466),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_674),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_674),
.Y(n_695)
);

BUFx6f_ASAP7_75t_L g696 ( 
.A(n_647),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_623),
.B(n_494),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_618),
.Y(n_698)
);

INVx2_ASAP7_75t_SL g699 ( 
.A(n_619),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_603),
.B(n_502),
.Y(n_700)
);

BUFx6f_ASAP7_75t_L g701 ( 
.A(n_647),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_619),
.B(n_524),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_663),
.B(n_491),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_674),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_674),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_664),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_622),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_622),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_663),
.B(n_490),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_673),
.B(n_526),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_614),
.B(n_561),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_622),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_603),
.B(n_521),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_595),
.Y(n_714)
);

AO22x2_ASAP7_75t_L g715 ( 
.A1(n_663),
.A2(n_487),
.B1(n_532),
.B2(n_570),
.Y(n_715)
);

OR2x2_ASAP7_75t_L g716 ( 
.A(n_669),
.B(n_572),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_625),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_625),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_L g719 ( 
.A(n_673),
.B(n_527),
.Y(n_719)
);

BUFx6f_ASAP7_75t_L g720 ( 
.A(n_647),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_672),
.B(n_573),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_625),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_627),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_623),
.B(n_527),
.Y(n_724)
);

NOR2x1p5_ASAP7_75t_L g725 ( 
.A(n_628),
.B(n_564),
.Y(n_725)
);

BUFx3_ASAP7_75t_L g726 ( 
.A(n_585),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_624),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_627),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_627),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_624),
.Y(n_730)
);

INVx3_ASAP7_75t_L g731 ( 
.A(n_624),
.Y(n_731)
);

BUFx3_ASAP7_75t_L g732 ( 
.A(n_585),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_586),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_664),
.Y(n_734)
);

AND2x6_ASAP7_75t_L g735 ( 
.A(n_623),
.B(n_345),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_642),
.Y(n_736)
);

BUFx10_ASAP7_75t_L g737 ( 
.A(n_634),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_642),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_642),
.Y(n_739)
);

BUFx3_ASAP7_75t_L g740 ( 
.A(n_586),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_644),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_635),
.B(n_567),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_641),
.B(n_575),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_645),
.B(n_483),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_644),
.Y(n_745)
);

AND2x2_ASAP7_75t_SL g746 ( 
.A(n_596),
.B(n_487),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_663),
.B(n_545),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_676),
.B(n_546),
.Y(n_748)
);

AND2x6_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_358),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_675),
.B(n_678),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_644),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_600),
.Y(n_752)
);

INVx3_ASAP7_75t_L g753 ( 
.A(n_624),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_666),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_583),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_666),
.Y(n_756)
);

OR2x2_ASAP7_75t_L g757 ( 
.A(n_669),
.B(n_546),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_666),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_646),
.B(n_525),
.Y(n_759)
);

AND2x2_ASAP7_75t_SL g760 ( 
.A(n_677),
.B(n_562),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_647),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_668),
.Y(n_762)
);

BUFx3_ASAP7_75t_L g763 ( 
.A(n_587),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_668),
.Y(n_764)
);

INVxp33_ASAP7_75t_L g765 ( 
.A(n_677),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_660),
.B(n_547),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

AND2x6_ASAP7_75t_L g768 ( 
.A(n_678),
.B(n_358),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_668),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_660),
.A2(n_529),
.B1(n_531),
.B2(n_530),
.Y(n_770)
);

INVx2_ASAP7_75t_SL g771 ( 
.A(n_631),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_587),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_676),
.B(n_529),
.Y(n_773)
);

BUFx4f_ASAP7_75t_L g774 ( 
.A(n_647),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_635),
.B(n_555),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_640),
.B(n_530),
.Y(n_776)
);

CKINVDCx16_ASAP7_75t_R g777 ( 
.A(n_665),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_654),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_640),
.B(n_633),
.Y(n_779)
);

INVx4_ASAP7_75t_L g780 ( 
.A(n_654),
.Y(n_780)
);

CKINVDCx8_ASAP7_75t_R g781 ( 
.A(n_665),
.Y(n_781)
);

AND2x4_ASAP7_75t_L g782 ( 
.A(n_660),
.B(n_559),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

NAND2x1p5_ASAP7_75t_L g784 ( 
.A(n_676),
.B(n_531),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_590),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_654),
.B(n_410),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_594),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_640),
.B(n_536),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_648),
.B(n_536),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_650),
.B(n_538),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_654),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_654),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_654),
.Y(n_793)
);

AND2x6_ASAP7_75t_L g794 ( 
.A(n_594),
.B(n_363),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_640),
.B(n_538),
.Y(n_795)
);

NAND3x1_ASAP7_75t_L g796 ( 
.A(n_632),
.B(n_264),
.C(n_262),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_651),
.B(n_543),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_633),
.B(n_543),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_597),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_597),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_655),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_656),
.B(n_549),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_655),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_657),
.B(n_549),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_584),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_633),
.Y(n_806)
);

AND3x4_ASAP7_75t_L g807 ( 
.A(n_660),
.B(n_481),
.C(n_379),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_601),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_633),
.B(n_552),
.Y(n_809)
);

INVx2_ASAP7_75t_SL g810 ( 
.A(n_631),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_659),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_601),
.B(n_552),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_667),
.B(n_554),
.Y(n_813)
);

INVx5_ASAP7_75t_L g814 ( 
.A(n_655),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_631),
.B(n_554),
.Y(n_815)
);

INVx3_ASAP7_75t_L g816 ( 
.A(n_655),
.Y(n_816)
);

BUFx6f_ASAP7_75t_L g817 ( 
.A(n_655),
.Y(n_817)
);

AND2x6_ASAP7_75t_L g818 ( 
.A(n_606),
.B(n_363),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_655),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_606),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_671),
.A2(n_335),
.B1(n_346),
.B2(n_289),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_608),
.B(n_557),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_L g823 ( 
.A(n_608),
.B(n_557),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_671),
.A2(n_374),
.B1(n_327),
.B2(n_328),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_661),
.Y(n_825)
);

BUFx3_ASAP7_75t_L g826 ( 
.A(n_609),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_661),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_661),
.Y(n_828)
);

INVxp33_ASAP7_75t_L g829 ( 
.A(n_632),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_591),
.Y(n_830)
);

INVx6_ASAP7_75t_L g831 ( 
.A(n_631),
.Y(n_831)
);

OR2x6_ASAP7_75t_L g832 ( 
.A(n_582),
.B(n_453),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_592),
.B(n_558),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_609),
.B(n_558),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_582),
.A2(n_563),
.B1(n_565),
.B2(n_560),
.Y(n_835)
);

INVx6_ASAP7_75t_L g836 ( 
.A(n_661),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_610),
.B(n_560),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_610),
.B(n_563),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_612),
.B(n_565),
.Y(n_839)
);

A2O1A1Ixp33_ASAP7_75t_L g840 ( 
.A1(n_742),
.A2(n_568),
.B(n_571),
.C(n_566),
.Y(n_840)
);

NOR2x2_ASAP7_75t_L g841 ( 
.A(n_760),
.B(n_322),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_790),
.B(n_611),
.Y(n_842)
);

AOI21xp5_ASAP7_75t_L g843 ( 
.A1(n_779),
.A2(n_613),
.B(n_611),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_726),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_685),
.Y(n_845)
);

NOR2x1p5_ASAP7_75t_L g846 ( 
.A(n_714),
.B(n_593),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_726),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_732),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_688),
.B(n_802),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_732),
.Y(n_850)
);

BUFx6f_ASAP7_75t_L g851 ( 
.A(n_696),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_714),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_733),
.Y(n_853)
);

AOI22xp5_ASAP7_75t_L g854 ( 
.A1(n_760),
.A2(n_616),
.B1(n_620),
.B2(n_613),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_784),
.B(n_616),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_733),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_784),
.B(n_620),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_784),
.B(n_629),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_740),
.Y(n_859)
);

AND2x6_ASAP7_75t_SL g860 ( 
.A(n_700),
.B(n_713),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_690),
.A2(n_630),
.B(n_629),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_685),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_687),
.Y(n_863)
);

INVx3_ASAP7_75t_L g864 ( 
.A(n_740),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_829),
.B(n_630),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_775),
.B(n_636),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_773),
.B(n_636),
.Y(n_867)
);

NAND2xp33_ASAP7_75t_L g868 ( 
.A(n_688),
.B(n_638),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_773),
.B(n_638),
.Y(n_869)
);

INVx3_ASAP7_75t_L g870 ( 
.A(n_763),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_765),
.B(n_703),
.Y(n_871)
);

BUFx12f_ASAP7_75t_L g872 ( 
.A(n_737),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_689),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_721),
.B(n_639),
.Y(n_874)
);

INVx4_ASAP7_75t_L g875 ( 
.A(n_831),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_763),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_703),
.B(n_569),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_688),
.B(n_639),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_783),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_735),
.A2(n_568),
.B1(n_571),
.B2(n_566),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_689),
.Y(n_881)
);

BUFx6f_ASAP7_75t_SL g882 ( 
.A(n_737),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_822),
.B(n_643),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_789),
.B(n_643),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_797),
.B(n_649),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_804),
.B(n_649),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_783),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_823),
.B(n_652),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_735),
.A2(n_653),
.B1(n_652),
.B2(n_359),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_837),
.B(n_653),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_831),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_813),
.B(n_661),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_698),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_681),
.B(n_661),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_838),
.B(n_724),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_710),
.B(n_576),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_831),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_698),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_735),
.A2(n_715),
.B1(n_684),
.B2(n_807),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_703),
.B(n_574),
.Y(n_900)
);

NAND2x1p5_ASAP7_75t_L g901 ( 
.A(n_679),
.B(n_577),
.Y(n_901)
);

AOI22xp33_ASAP7_75t_L g902 ( 
.A1(n_735),
.A2(n_578),
.B1(n_581),
.B2(n_577),
.Y(n_902)
);

AND2x6_ASAP7_75t_SL g903 ( 
.A(n_755),
.B(n_262),
.Y(n_903)
);

AND2x2_ASAP7_75t_SL g904 ( 
.A(n_686),
.B(n_248),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_716),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_776),
.A2(n_581),
.B(n_578),
.Y(n_906)
);

AND2x6_ASAP7_75t_L g907 ( 
.A(n_709),
.B(n_367),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_826),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_719),
.B(n_615),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_681),
.B(n_615),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_826),
.Y(n_911)
);

AOI22xp33_ASAP7_75t_L g912 ( 
.A1(n_735),
.A2(n_347),
.B1(n_379),
.B2(n_322),
.Y(n_912)
);

AO221x1_ASAP7_75t_L g913 ( 
.A1(n_715),
.A2(n_408),
.B1(n_421),
.B2(n_290),
.C(n_291),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_772),
.Y(n_914)
);

INVx2_ASAP7_75t_SL g915 ( 
.A(n_716),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_699),
.B(n_615),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_SL g917 ( 
.A(n_755),
.B(n_662),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_699),
.B(n_615),
.Y(n_918)
);

NAND2xp33_ASAP7_75t_L g919 ( 
.A(n_735),
.B(n_410),
.Y(n_919)
);

INVxp67_ASAP7_75t_L g920 ( 
.A(n_811),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_683),
.B(n_235),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_683),
.B(n_273),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_683),
.B(n_444),
.Y(n_923)
);

INVx8_ASAP7_75t_L g924 ( 
.A(n_794),
.Y(n_924)
);

AO22x1_ASAP7_75t_L g925 ( 
.A1(n_807),
.A2(n_329),
.B1(n_342),
.B2(n_326),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_SL g926 ( 
.A(n_727),
.B(n_367),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_SL g927 ( 
.A1(n_686),
.A2(n_621),
.B1(n_626),
.B2(n_607),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_702),
.A2(n_290),
.B(n_291),
.C(n_264),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_723),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_715),
.A2(n_444),
.B1(n_412),
.B2(n_421),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_727),
.B(n_393),
.Y(n_931)
);

INVx2_ASAP7_75t_SL g932 ( 
.A(n_757),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_SL g933 ( 
.A(n_727),
.B(n_393),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_715),
.A2(n_412),
.B1(n_421),
.B2(n_399),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_723),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_697),
.B(n_293),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_811),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_679),
.B(n_397),
.Y(n_938)
);

AOI22xp33_ASAP7_75t_L g939 ( 
.A1(n_749),
.A2(n_768),
.B1(n_818),
.B2(n_794),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_728),
.Y(n_940)
);

NOR2x1p5_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_348),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_709),
.B(n_747),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_730),
.B(n_399),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_682),
.B(n_350),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_730),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_693),
.B(n_352),
.Y(n_946)
);

AND2x2_ASAP7_75t_L g947 ( 
.A(n_709),
.B(n_670),
.Y(n_947)
);

AOI22xp33_ASAP7_75t_L g948 ( 
.A1(n_749),
.A2(n_412),
.B1(n_421),
.B2(n_429),
.Y(n_948)
);

HB1xp67_ASAP7_75t_L g949 ( 
.A(n_752),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_747),
.B(n_429),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_747),
.B(n_442),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_772),
.Y(n_952)
);

INVx3_ASAP7_75t_L g953 ( 
.A(n_730),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_748),
.B(n_658),
.Y(n_954)
);

NAND2x1p5_ASAP7_75t_L g955 ( 
.A(n_691),
.B(n_442),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_706),
.B(n_293),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_731),
.B(n_310),
.Y(n_957)
);

AOI21x1_ASAP7_75t_L g958 ( 
.A1(n_785),
.A2(n_598),
.B(n_588),
.Y(n_958)
);

NAND2xp33_ASAP7_75t_L g959 ( 
.A(n_794),
.B(n_818),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_785),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_787),
.A2(n_800),
.B1(n_808),
.B2(n_799),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_734),
.B(n_297),
.Y(n_962)
);

BUFx6f_ASAP7_75t_L g963 ( 
.A(n_696),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_833),
.B(n_839),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_770),
.B(n_766),
.Y(n_965)
);

OR2x6_ASAP7_75t_L g966 ( 
.A(n_771),
.B(n_637),
.Y(n_966)
);

AOI22xp5_ASAP7_75t_L g967 ( 
.A1(n_766),
.A2(n_238),
.B1(n_244),
.B2(n_236),
.Y(n_967)
);

INVx4_ASAP7_75t_L g968 ( 
.A(n_831),
.Y(n_968)
);

INVx2_ASAP7_75t_SL g969 ( 
.A(n_757),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_766),
.B(n_297),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_815),
.B(n_354),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_696),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_748),
.B(n_299),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_782),
.A2(n_746),
.B1(n_768),
.B2(n_749),
.Y(n_974)
);

BUFx8_ASAP7_75t_L g975 ( 
.A(n_771),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_782),
.B(n_299),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_782),
.B(n_731),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_731),
.B(n_302),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_753),
.B(n_310),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_691),
.B(n_357),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_810),
.B(n_302),
.Y(n_981)
);

NOR2xp33_ASAP7_75t_L g982 ( 
.A(n_753),
.B(n_806),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_728),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_787),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_746),
.B(n_317),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_753),
.B(n_360),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_749),
.A2(n_250),
.B1(n_252),
.B2(n_249),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_805),
.Y(n_988)
);

OAI22xp33_ASAP7_75t_L g989 ( 
.A1(n_824),
.A2(n_821),
.B1(n_832),
.B2(n_810),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_799),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_806),
.B(n_317),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_736),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_806),
.B(n_332),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_750),
.B(n_332),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_749),
.A2(n_421),
.B1(n_602),
.B2(n_598),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_800),
.B(n_356),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_788),
.B(n_362),
.Y(n_997)
);

BUFx8_ASAP7_75t_L g998 ( 
.A(n_749),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_768),
.A2(n_588),
.B1(n_602),
.B2(n_598),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_808),
.B(n_356),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_696),
.B(n_340),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_820),
.A2(n_426),
.B1(n_394),
.B2(n_456),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_SL g1003 ( 
.A(n_696),
.B(n_340),
.Y(n_1003)
);

AND2x4_ASAP7_75t_L g1004 ( 
.A(n_832),
.B(n_361),
.Y(n_1004)
);

AOI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_768),
.A2(n_265),
.B1(n_457),
.B2(n_261),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_820),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_754),
.Y(n_1007)
);

AOI22xp33_ASAP7_75t_L g1008 ( 
.A1(n_768),
.A2(n_588),
.B1(n_602),
.B2(n_380),
.Y(n_1008)
);

AND2x2_ASAP7_75t_SL g1009 ( 
.A(n_777),
.B(n_361),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_737),
.Y(n_1010)
);

INVx2_ASAP7_75t_SL g1011 ( 
.A(n_725),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_865),
.B(n_835),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_SL g1013 ( 
.A(n_852),
.B(n_743),
.C(n_711),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_949),
.Y(n_1014)
);

INVx3_ASAP7_75t_L g1015 ( 
.A(n_851),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_865),
.B(n_812),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_985),
.B(n_830),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_842),
.B(n_834),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_914),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_952),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_852),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_960),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_845),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_874),
.B(n_798),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_872),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_845),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_872),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_984),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_R g1029 ( 
.A(n_917),
.B(n_781),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_997),
.A2(n_809),
.B(n_369),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_851),
.Y(n_1031)
);

BUFx2_ASAP7_75t_L g1032 ( 
.A(n_954),
.Y(n_1032)
);

AND2x2_ASAP7_75t_SL g1033 ( 
.A(n_904),
.B(n_754),
.Y(n_1033)
);

INVxp67_ASAP7_75t_SL g1034 ( 
.A(n_868),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_990),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_882),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_897),
.B(n_832),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_1006),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_862),
.Y(n_1039)
);

OR2x6_ASAP7_75t_L g1040 ( 
.A(n_924),
.B(n_832),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_1007),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_924),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_920),
.B(n_781),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_871),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_895),
.B(n_768),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_897),
.B(n_744),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_884),
.B(n_794),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_851),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_910),
.Y(n_1049)
);

BUFx6f_ASAP7_75t_L g1050 ( 
.A(n_851),
.Y(n_1050)
);

BUFx2_ASAP7_75t_L g1051 ( 
.A(n_947),
.Y(n_1051)
);

INVx3_ASAP7_75t_SL g1052 ( 
.A(n_966),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_975),
.Y(n_1053)
);

NAND2x1p5_ASAP7_75t_L g1054 ( 
.A(n_875),
.B(n_780),
.Y(n_1054)
);

OA22x2_ASAP7_75t_L g1055 ( 
.A1(n_899),
.A2(n_796),
.B1(n_759),
.B2(n_758),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_884),
.A2(n_795),
.B(n_708),
.C(n_712),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_916),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_961),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_862),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_885),
.B(n_794),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_885),
.B(n_794),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_886),
.B(n_818),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_963),
.Y(n_1063)
);

BUFx2_ASAP7_75t_L g1064 ( 
.A(n_905),
.Y(n_1064)
);

BUFx3_ASAP7_75t_L g1065 ( 
.A(n_975),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_873),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_873),
.Y(n_1067)
);

NOR3xp33_ASAP7_75t_SL g1068 ( 
.A(n_1002),
.B(n_372),
.C(n_368),
.Y(n_1068)
);

AOI22x1_ASAP7_75t_L g1069 ( 
.A1(n_843),
.A2(n_758),
.B1(n_762),
.B2(n_756),
.Y(n_1069)
);

HB1xp67_ASAP7_75t_L g1070 ( 
.A(n_932),
.Y(n_1070)
);

INVx1_ASAP7_75t_SL g1071 ( 
.A(n_863),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_924),
.Y(n_1072)
);

NAND2xp33_ASAP7_75t_SL g1073 ( 
.A(n_849),
.B(n_780),
.Y(n_1073)
);

AND2x4_ASAP7_75t_L g1074 ( 
.A(n_875),
.B(n_891),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_886),
.B(n_818),
.Y(n_1075)
);

BUFx3_ASAP7_75t_L g1076 ( 
.A(n_975),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_963),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_969),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_882),
.Y(n_1079)
);

AOI22xp33_ASAP7_75t_L g1080 ( 
.A1(n_904),
.A2(n_818),
.B1(n_692),
.B2(n_762),
.Y(n_1080)
);

OR2x2_ASAP7_75t_SL g1081 ( 
.A(n_942),
.B(n_796),
.Y(n_1081)
);

INVx3_ASAP7_75t_SL g1082 ( 
.A(n_966),
.Y(n_1082)
);

OR2x6_ASAP7_75t_L g1083 ( 
.A(n_924),
.B(n_756),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_901),
.Y(n_1084)
);

NOR3xp33_ASAP7_75t_L g1085 ( 
.A(n_937),
.B(n_376),
.C(n_364),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_918),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_936),
.B(n_764),
.Y(n_1087)
);

NOR2xp33_ASAP7_75t_R g1088 ( 
.A(n_1010),
.B(n_695),
.Y(n_1088)
);

NOR3xp33_ASAP7_75t_SL g1089 ( 
.A(n_927),
.B(n_375),
.C(n_373),
.Y(n_1089)
);

HB1xp67_ASAP7_75t_L g1090 ( 
.A(n_915),
.Y(n_1090)
);

BUFx6f_ASAP7_75t_L g1091 ( 
.A(n_963),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_974),
.B(n_701),
.Y(n_1092)
);

INVx1_ASAP7_75t_SL g1093 ( 
.A(n_988),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_963),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_881),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_977),
.B(n_707),
.Y(n_1096)
);

BUFx6f_ASAP7_75t_L g1097 ( 
.A(n_972),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_881),
.Y(n_1098)
);

NOR2xp33_ASAP7_75t_L g1099 ( 
.A(n_860),
.B(n_780),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_972),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_936),
.B(n_764),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_965),
.A2(n_769),
.B1(n_741),
.B2(n_751),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_966),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_867),
.Y(n_1105)
);

BUFx6f_ASAP7_75t_L g1106 ( 
.A(n_972),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_944),
.B(n_708),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_1009),
.Y(n_1108)
);

NOR3xp33_ASAP7_75t_SL g1109 ( 
.A(n_946),
.B(n_385),
.C(n_383),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_936),
.B(n_769),
.Y(n_1110)
);

INVx1_ASAP7_75t_SL g1111 ( 
.A(n_877),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_846),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_L g1113 ( 
.A(n_989),
.B(n_792),
.Y(n_1113)
);

INVx3_ASAP7_75t_L g1114 ( 
.A(n_945),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_944),
.B(n_712),
.Y(n_1115)
);

INVx3_ASAP7_75t_L g1116 ( 
.A(n_945),
.Y(n_1116)
);

NOR3xp33_ASAP7_75t_SL g1117 ( 
.A(n_986),
.B(n_391),
.C(n_388),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_893),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_869),
.B(n_717),
.Y(n_1119)
);

BUFx4f_ASAP7_75t_L g1120 ( 
.A(n_907),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_981),
.B(n_718),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_849),
.B(n_864),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_973),
.B(n_718),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_1009),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_900),
.Y(n_1125)
);

INVx5_ASAP7_75t_L g1126 ( 
.A(n_875),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_981),
.B(n_722),
.Y(n_1127)
);

AOI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_907),
.A2(n_836),
.B1(n_695),
.B2(n_819),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_893),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_996),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_981),
.B(n_722),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_898),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_945),
.Y(n_1133)
);

AND2x6_ASAP7_75t_L g1134 ( 
.A(n_998),
.B(n_729),
.Y(n_1134)
);

INVx3_ASAP7_75t_L g1135 ( 
.A(n_953),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_923),
.B(n_729),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_921),
.B(n_738),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_922),
.B(n_738),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_907),
.B(n_739),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_903),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_907),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_891),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_998),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1000),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_891),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_844),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_907),
.B(n_980),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_847),
.Y(n_1148)
);

AND2x4_ASAP7_75t_L g1149 ( 
.A(n_968),
.B(n_695),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_980),
.B(n_739),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_848),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_SL g1152 ( 
.A(n_864),
.B(n_701),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_898),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_929),
.Y(n_1154)
);

INVx2_ASAP7_75t_SL g1155 ( 
.A(n_901),
.Y(n_1155)
);

AO22x1_ASAP7_75t_L g1156 ( 
.A1(n_998),
.A2(n_376),
.B1(n_380),
.B2(n_364),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_968),
.Y(n_1157)
);

AND2x2_ASAP7_75t_L g1158 ( 
.A(n_1004),
.B(n_745),
.Y(n_1158)
);

AND2x2_ASAP7_75t_L g1159 ( 
.A(n_1004),
.B(n_970),
.Y(n_1159)
);

INVx6_ASAP7_75t_L g1160 ( 
.A(n_968),
.Y(n_1160)
);

BUFx3_ASAP7_75t_L g1161 ( 
.A(n_864),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_929),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_938),
.Y(n_1163)
);

O2A1O1Ixp5_ASAP7_75t_L g1164 ( 
.A1(n_866),
.A2(n_774),
.B(n_792),
.C(n_825),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_953),
.Y(n_1165)
);

INVx5_ASAP7_75t_L g1166 ( 
.A(n_870),
.Y(n_1166)
);

NOR2xp33_ASAP7_75t_R g1167 ( 
.A(n_1011),
.B(n_816),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_SL g1168 ( 
.A(n_986),
.B(n_405),
.C(n_401),
.Y(n_1168)
);

BUFx3_ASAP7_75t_L g1169 ( 
.A(n_870),
.Y(n_1169)
);

INVx3_ASAP7_75t_SL g1170 ( 
.A(n_841),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_L g1171 ( 
.A(n_964),
.B(n_792),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_896),
.B(n_745),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_841),
.Y(n_1173)
);

AND2x4_ASAP7_75t_L g1174 ( 
.A(n_870),
.B(n_825),
.Y(n_1174)
);

INVx4_ASAP7_75t_L g1175 ( 
.A(n_908),
.Y(n_1175)
);

O2A1O1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_840),
.A2(n_387),
.B(n_389),
.C(n_455),
.Y(n_1176)
);

OR2x4_ASAP7_75t_L g1177 ( 
.A(n_964),
.B(n_387),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_SL g1178 ( 
.A(n_967),
.B(n_414),
.C(n_406),
.Y(n_1178)
);

AND2x2_ASAP7_75t_L g1179 ( 
.A(n_1004),
.B(n_736),
.Y(n_1179)
);

NOR3xp33_ASAP7_75t_SL g1180 ( 
.A(n_956),
.B(n_419),
.C(n_417),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_908),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_953),
.Y(n_1182)
);

AND2x4_ASAP7_75t_L g1183 ( 
.A(n_908),
.B(n_825),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_935),
.Y(n_1184)
);

NOR3xp33_ASAP7_75t_SL g1185 ( 
.A(n_962),
.B(n_430),
.C(n_425),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_925),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_935),
.Y(n_1187)
);

OR2x2_ASAP7_75t_L g1188 ( 
.A(n_976),
.B(n_741),
.Y(n_1188)
);

NOR3xp33_ASAP7_75t_SL g1189 ( 
.A(n_994),
.B(n_436),
.C(n_431),
.Y(n_1189)
);

OR2x6_ASAP7_75t_L g1190 ( 
.A(n_938),
.B(n_751),
.Y(n_1190)
);

INVx3_ASAP7_75t_L g1191 ( 
.A(n_940),
.Y(n_1191)
);

HB1xp67_ASAP7_75t_L g1192 ( 
.A(n_955),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_939),
.B(n_701),
.Y(n_1193)
);

OR2x6_ASAP7_75t_L g1194 ( 
.A(n_955),
.B(n_761),
.Y(n_1194)
);

INVx2_ASAP7_75t_L g1195 ( 
.A(n_940),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_SL g1196 ( 
.A(n_889),
.B(n_701),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_983),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_983),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_971),
.A2(n_836),
.B1(n_816),
.B2(n_827),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_992),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_883),
.B(n_819),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_850),
.Y(n_1202)
);

OR2x6_ASAP7_75t_SL g1203 ( 
.A(n_950),
.B(n_447),
.Y(n_1203)
);

AOI21xp33_ASAP7_75t_L g1204 ( 
.A1(n_1055),
.A2(n_971),
.B(n_919),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1016),
.A2(n_840),
.B(n_890),
.C(n_888),
.Y(n_1205)
);

NAND2x1p5_ASAP7_75t_L g1206 ( 
.A(n_1120),
.B(n_853),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1105),
.B(n_951),
.Y(n_1207)
);

OAI21x1_ASAP7_75t_L g1208 ( 
.A1(n_1069),
.A2(n_958),
.B(n_1001),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1120),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1018),
.B(n_854),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1143),
.B(n_1037),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1159),
.B(n_856),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_SL g1213 ( 
.A1(n_1058),
.A2(n_857),
.B(n_855),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1022),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1069),
.A2(n_1003),
.B(n_1001),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1164),
.A2(n_1003),
.B(n_861),
.Y(n_1216)
);

OAI21xp33_ASAP7_75t_L g1217 ( 
.A1(n_1030),
.A2(n_902),
.B(n_880),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1034),
.A2(n_959),
.B(n_878),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1058),
.A2(n_979),
.B(n_957),
.Y(n_1219)
);

INVx4_ASAP7_75t_L g1220 ( 
.A(n_1042),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1159),
.B(n_859),
.Y(n_1221)
);

NOR2x1_ASAP7_75t_SL g1222 ( 
.A(n_1083),
.B(n_858),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1130),
.B(n_876),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1045),
.A2(n_919),
.B(n_894),
.Y(n_1224)
);

OAI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1122),
.A2(n_979),
.B(n_957),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1147),
.B(n_1047),
.Y(n_1226)
);

AND2x2_ASAP7_75t_L g1227 ( 
.A(n_1017),
.B(n_941),
.Y(n_1227)
);

BUFx12f_ASAP7_75t_L g1228 ( 
.A(n_1027),
.Y(n_1228)
);

NAND2x1p5_ASAP7_75t_L g1229 ( 
.A(n_1120),
.B(n_879),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1092),
.A2(n_992),
.B(n_991),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1028),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1144),
.B(n_887),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1056),
.A2(n_894),
.A3(n_892),
.B(n_911),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1023),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1055),
.A2(n_993),
.B(n_978),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_SL g1236 ( 
.A(n_1060),
.B(n_892),
.Y(n_1236)
);

AO31x2_ASAP7_75t_L g1237 ( 
.A1(n_1107),
.A2(n_705),
.A3(n_680),
.B(n_694),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1038),
.Y(n_1238)
);

NOR2xp67_ASAP7_75t_L g1239 ( 
.A(n_1021),
.B(n_906),
.Y(n_1239)
);

NOR2xp67_ASAP7_75t_SL g1240 ( 
.A(n_1021),
.B(n_926),
.Y(n_1240)
);

NOR2x1_ASAP7_75t_SL g1241 ( 
.A(n_1083),
.B(n_926),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1171),
.A2(n_982),
.B(n_909),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_1029),
.Y(n_1243)
);

A2O1A1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1113),
.A2(n_928),
.B(n_982),
.C(n_912),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1017),
.B(n_930),
.Y(n_1245)
);

BUFx12f_ASAP7_75t_L g1246 ( 
.A(n_1027),
.Y(n_1246)
);

OAI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1115),
.A2(n_933),
.B(n_931),
.Y(n_1247)
);

INVx1_ASAP7_75t_SL g1248 ( 
.A(n_1014),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1033),
.B(n_934),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1055),
.A2(n_767),
.B(n_761),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1176),
.A2(n_778),
.B(n_767),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1024),
.A2(n_774),
.B(n_931),
.Y(n_1252)
);

AOI221x1_ASAP7_75t_L g1253 ( 
.A1(n_1073),
.A2(n_680),
.B1(n_704),
.B2(n_705),
.C(n_694),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_1036),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_1150),
.A2(n_1191),
.B(n_1154),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1191),
.A2(n_791),
.B(n_778),
.Y(n_1256)
);

AO21x1_ASAP7_75t_L g1257 ( 
.A1(n_1073),
.A2(n_943),
.B(n_933),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1191),
.A2(n_793),
.B(n_791),
.Y(n_1258)
);

OA22x2_ASAP7_75t_L g1259 ( 
.A1(n_1108),
.A2(n_913),
.B1(n_1005),
.B2(n_987),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1023),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1033),
.B(n_1008),
.Y(n_1261)
);

AOI21x1_ASAP7_75t_L g1262 ( 
.A1(n_1152),
.A2(n_704),
.B(n_793),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1087),
.B(n_948),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1026),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1025),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1067),
.A2(n_828),
.B(n_827),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1087),
.B(n_819),
.Y(n_1267)
);

AO21x1_ASAP7_75t_L g1268 ( 
.A1(n_1061),
.A2(n_786),
.B(n_828),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1102),
.B(n_827),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1102),
.B(n_701),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1119),
.A2(n_801),
.B(n_720),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1110),
.B(n_720),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1067),
.A2(n_999),
.B(n_995),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1110),
.B(n_720),
.Y(n_1274)
);

OAI22xp5_ASAP7_75t_L g1275 ( 
.A1(n_1019),
.A2(n_836),
.B1(n_454),
.B2(n_420),
.Y(n_1275)
);

BUFx2_ASAP7_75t_L g1276 ( 
.A(n_1125),
.Y(n_1276)
);

AO31x2_ASAP7_75t_L g1277 ( 
.A1(n_1062),
.A2(n_455),
.A3(n_438),
.B(n_440),
.Y(n_1277)
);

AND2x4_ASAP7_75t_L g1278 ( 
.A(n_1143),
.B(n_814),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1019),
.A2(n_1035),
.B1(n_1020),
.B2(n_1075),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1123),
.B(n_720),
.Y(n_1280)
);

CKINVDCx6p67_ASAP7_75t_R g1281 ( 
.A(n_1025),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_1154),
.A2(n_407),
.B(n_389),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1026),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1039),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_SL g1285 ( 
.A(n_1181),
.B(n_720),
.Y(n_1285)
);

OAI21x1_ASAP7_75t_L g1286 ( 
.A1(n_1197),
.A2(n_416),
.B(n_407),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_SL g1287 ( 
.A1(n_1175),
.A2(n_420),
.B(n_416),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1123),
.B(n_801),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1020),
.A2(n_836),
.B1(n_440),
.B2(n_454),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1039),
.Y(n_1290)
);

BUFx4f_ASAP7_75t_SL g1291 ( 
.A(n_1093),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1172),
.A2(n_803),
.B(n_801),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1012),
.B(n_801),
.Y(n_1293)
);

NAND2x1_ASAP7_75t_L g1294 ( 
.A(n_1042),
.B(n_801),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_SL g1295 ( 
.A(n_1036),
.B(n_448),
.Y(n_1295)
);

CKINVDCx5p33_ASAP7_75t_R g1296 ( 
.A(n_1079),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1035),
.A2(n_445),
.B1(n_438),
.B2(n_450),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1201),
.A2(n_817),
.B(n_803),
.Y(n_1298)
);

INVx2_ASAP7_75t_L g1299 ( 
.A(n_1059),
.Y(n_1299)
);

AO31x2_ASAP7_75t_L g1300 ( 
.A1(n_1059),
.A2(n_445),
.A3(n_786),
.B(n_604),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1096),
.A2(n_814),
.B(n_452),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1197),
.A2(n_817),
.B(n_803),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1200),
.A2(n_817),
.B(n_803),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1200),
.A2(n_817),
.B(n_803),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1066),
.A2(n_817),
.B(n_814),
.Y(n_1305)
);

AOI21xp33_ASAP7_75t_L g1306 ( 
.A1(n_1111),
.A2(n_1127),
.B(n_1121),
.Y(n_1306)
);

AO31x2_ASAP7_75t_L g1307 ( 
.A1(n_1066),
.A2(n_604),
.A3(n_589),
.B(n_814),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1158),
.B(n_451),
.Y(n_1308)
);

AO31x2_ASAP7_75t_L g1309 ( 
.A1(n_1095),
.A2(n_604),
.A3(n_589),
.B(n_814),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1158),
.B(n_8),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1126),
.A2(n_267),
.B(n_256),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1126),
.A2(n_279),
.B(n_269),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1095),
.A2(n_410),
.B(n_589),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_SL g1314 ( 
.A(n_1181),
.B(n_589),
.Y(n_1314)
);

AOI211x1_ASAP7_75t_L g1315 ( 
.A1(n_1041),
.A2(n_8),
.B(n_10),
.C(n_11),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1126),
.A2(n_285),
.B(n_281),
.Y(n_1316)
);

CKINVDCx5p33_ASAP7_75t_R g1317 ( 
.A(n_1079),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1049),
.A2(n_1086),
.B(n_1057),
.Y(n_1318)
);

BUFx3_ASAP7_75t_L g1319 ( 
.A(n_1053),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1098),
.A2(n_410),
.B(n_589),
.Y(n_1320)
);

AOI21xp5_ASAP7_75t_L g1321 ( 
.A1(n_1126),
.A2(n_1183),
.B(n_1174),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1098),
.A2(n_303),
.B(n_292),
.Y(n_1322)
);

OAI21x1_ASAP7_75t_L g1323 ( 
.A1(n_1118),
.A2(n_410),
.B(n_604),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1118),
.A2(n_1132),
.A3(n_1153),
.B(n_1129),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1146),
.Y(n_1325)
);

INVx2_ASAP7_75t_L g1326 ( 
.A(n_1129),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_SL g1327 ( 
.A(n_1181),
.B(n_589),
.Y(n_1327)
);

AOI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1174),
.A2(n_378),
.B(n_435),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1071),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1108),
.B(n_604),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1148),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1199),
.A2(n_381),
.B(n_434),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1141),
.A2(n_1175),
.B1(n_1131),
.B2(n_1072),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1174),
.A2(n_1183),
.B(n_1175),
.Y(n_1334)
);

OAI21x1_ASAP7_75t_L g1335 ( 
.A1(n_1132),
.A2(n_1162),
.B(n_1153),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1183),
.A2(n_370),
.B(n_432),
.Y(n_1336)
);

NAND2x1p5_ASAP7_75t_L g1337 ( 
.A(n_1042),
.B(n_604),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1162),
.Y(n_1338)
);

A2O1A1Ixp33_ASAP7_75t_L g1339 ( 
.A1(n_1109),
.A2(n_237),
.B(n_240),
.C(n_423),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1141),
.A2(n_428),
.B1(n_427),
.B2(n_304),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1151),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1166),
.A2(n_309),
.B(n_418),
.Y(n_1342)
);

AOI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1166),
.A2(n_315),
.B(n_415),
.Y(n_1343)
);

AO31x2_ASAP7_75t_L g1344 ( 
.A1(n_1184),
.A2(n_410),
.A3(n_423),
.B(n_371),
.Y(n_1344)
);

NAND2xp5_ASAP7_75t_L g1345 ( 
.A(n_1044),
.B(n_10),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1184),
.A2(n_410),
.B(n_423),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1072),
.B(n_237),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1139),
.A2(n_404),
.B(n_403),
.Y(n_1348)
);

OR2x6_ASAP7_75t_L g1349 ( 
.A(n_1040),
.B(n_237),
.Y(n_1349)
);

AND2x6_ASAP7_75t_L g1350 ( 
.A(n_1074),
.B(n_237),
.Y(n_1350)
);

INVx4_ASAP7_75t_L g1351 ( 
.A(n_1072),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1187),
.A2(n_410),
.B(n_423),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1124),
.B(n_12),
.Y(n_1353)
);

NOR2x1_ASAP7_75t_SL g1354 ( 
.A(n_1083),
.B(n_237),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1187),
.A2(n_410),
.B(n_423),
.Y(n_1355)
);

NOR2xp33_ASAP7_75t_L g1356 ( 
.A(n_1032),
.B(n_12),
.Y(n_1356)
);

AOI21x1_ASAP7_75t_L g1357 ( 
.A1(n_1193),
.A2(n_240),
.B(n_313),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1195),
.A2(n_400),
.B(n_398),
.Y(n_1358)
);

OAI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1136),
.A2(n_395),
.B(n_392),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1124),
.B(n_13),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1195),
.A2(n_240),
.B(n_313),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_1186),
.Y(n_1362)
);

AOI21xp33_ASAP7_75t_SL g1363 ( 
.A1(n_1043),
.A2(n_13),
.B(n_14),
.Y(n_1363)
);

NAND2x1_ASAP7_75t_L g1364 ( 
.A(n_1160),
.B(n_240),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1044),
.B(n_15),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1198),
.A2(n_240),
.B(n_313),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1166),
.A2(n_390),
.B(n_386),
.Y(n_1367)
);

AOI21xp5_ASAP7_75t_L g1368 ( 
.A1(n_1166),
.A2(n_384),
.B(n_382),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1198),
.A2(n_371),
.B(n_313),
.Y(n_1369)
);

OAI21x1_ASAP7_75t_L g1370 ( 
.A1(n_1015),
.A2(n_371),
.B(n_313),
.Y(n_1370)
);

OAI21x1_ASAP7_75t_L g1371 ( 
.A1(n_1015),
.A2(n_371),
.B(n_221),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1361),
.A2(n_1031),
.B(n_1015),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1204),
.A2(n_1032),
.B1(n_1051),
.B2(n_1125),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1220),
.Y(n_1374)
);

AOI21xp33_ASAP7_75t_L g1375 ( 
.A1(n_1205),
.A2(n_1080),
.B(n_1137),
.Y(n_1375)
);

OA21x2_ASAP7_75t_L g1376 ( 
.A1(n_1255),
.A2(n_1103),
.B(n_1138),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1210),
.B(n_1064),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1249),
.B(n_1179),
.Y(n_1378)
);

AO21x2_ASAP7_75t_L g1379 ( 
.A1(n_1255),
.A2(n_1196),
.B(n_1136),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1211),
.B(n_1040),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1248),
.B(n_1064),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1207),
.B(n_1051),
.Y(n_1382)
);

OAI21x1_ASAP7_75t_L g1383 ( 
.A1(n_1361),
.A2(n_1063),
.B(n_1031),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_L g1384 ( 
.A1(n_1366),
.A2(n_1063),
.B(n_1031),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1291),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1242),
.A2(n_1099),
.B(n_1178),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_L g1387 ( 
.A1(n_1366),
.A2(n_1094),
.B(n_1063),
.Y(n_1387)
);

NAND2x1p5_ASAP7_75t_L g1388 ( 
.A(n_1209),
.B(n_1166),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1268),
.A2(n_1202),
.A3(n_1163),
.B(n_1177),
.Y(n_1389)
);

BUFx10_ASAP7_75t_L g1390 ( 
.A(n_1254),
.Y(n_1390)
);

OAI21x1_ASAP7_75t_L g1391 ( 
.A1(n_1369),
.A2(n_1100),
.B(n_1094),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1214),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1231),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1369),
.A2(n_1100),
.B(n_1094),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1211),
.B(n_1040),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1249),
.A2(n_1186),
.B1(n_1140),
.B2(n_1104),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1346),
.A2(n_1128),
.B(n_1117),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1346),
.A2(n_1100),
.B(n_1114),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1238),
.Y(n_1399)
);

OR2x2_ASAP7_75t_L g1400 ( 
.A(n_1245),
.B(n_1081),
.Y(n_1400)
);

AND2x2_ASAP7_75t_L g1401 ( 
.A(n_1261),
.B(n_1179),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1329),
.B(n_1070),
.Y(n_1402)
);

BUFx8_ASAP7_75t_L g1403 ( 
.A(n_1228),
.Y(n_1403)
);

OR2x2_ASAP7_75t_L g1404 ( 
.A(n_1233),
.B(n_1081),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1352),
.A2(n_1116),
.B(n_1114),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1211),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1265),
.Y(n_1407)
);

OA21x2_ASAP7_75t_L g1408 ( 
.A1(n_1352),
.A2(n_1168),
.B(n_1188),
.Y(n_1408)
);

BUFx10_ASAP7_75t_L g1409 ( 
.A(n_1254),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1355),
.A2(n_1116),
.B(n_1114),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1355),
.A2(n_1133),
.B(n_1116),
.Y(n_1411)
);

AND2x4_ASAP7_75t_SL g1412 ( 
.A(n_1281),
.B(n_1040),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1325),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1233),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1208),
.A2(n_1135),
.B(n_1133),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1324),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1331),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1208),
.A2(n_1135),
.B(n_1133),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1341),
.Y(n_1419)
);

BUFx4_ASAP7_75t_R g1420 ( 
.A(n_1241),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1223),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1356),
.B(n_1078),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1324),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1233),
.B(n_1163),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1313),
.A2(n_1165),
.B(n_1135),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1232),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1313),
.A2(n_1182),
.B(n_1165),
.Y(n_1427)
);

AOI21x1_ASAP7_75t_L g1428 ( 
.A1(n_1226),
.A2(n_1190),
.B(n_1194),
.Y(n_1428)
);

INVx2_ASAP7_75t_L g1429 ( 
.A(n_1324),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1320),
.A2(n_1182),
.B(n_1165),
.Y(n_1430)
);

BUFx12f_ASAP7_75t_L g1431 ( 
.A(n_1228),
.Y(n_1431)
);

OAI221xp5_ASAP7_75t_L g1432 ( 
.A1(n_1356),
.A2(n_1085),
.B1(n_1013),
.B2(n_1068),
.C(n_1089),
.Y(n_1432)
);

OAI21x1_ASAP7_75t_L g1433 ( 
.A1(n_1320),
.A2(n_1323),
.B(n_1216),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1209),
.B(n_1037),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1323),
.A2(n_1182),
.B(n_1054),
.Y(n_1435)
);

A2O1A1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1244),
.A2(n_1188),
.B(n_1155),
.C(n_1084),
.Y(n_1436)
);

BUFx3_ASAP7_75t_L g1437 ( 
.A(n_1265),
.Y(n_1437)
);

AO32x2_ASAP7_75t_L g1438 ( 
.A1(n_1279),
.A2(n_1084),
.A3(n_1155),
.B1(n_1177),
.B2(n_1156),
.Y(n_1438)
);

INVx2_ASAP7_75t_L g1439 ( 
.A(n_1324),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1234),
.Y(n_1440)
);

BUFx8_ASAP7_75t_L g1441 ( 
.A(n_1246),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1227),
.A2(n_1173),
.B1(n_1104),
.B2(n_1170),
.Y(n_1442)
);

BUFx2_ASAP7_75t_L g1443 ( 
.A(n_1233),
.Y(n_1443)
);

AO31x2_ASAP7_75t_L g1444 ( 
.A1(n_1257),
.A2(n_1177),
.A3(n_1190),
.B(n_1156),
.Y(n_1444)
);

INVx3_ASAP7_75t_SL g1445 ( 
.A(n_1296),
.Y(n_1445)
);

BUFx12f_ASAP7_75t_L g1446 ( 
.A(n_1246),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1216),
.A2(n_1054),
.B(n_1192),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1215),
.A2(n_1054),
.B(n_1050),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1319),
.B(n_1278),
.Y(n_1449)
);

INVx3_ASAP7_75t_L g1450 ( 
.A(n_1220),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1349),
.B(n_1190),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1215),
.A2(n_1101),
.B(n_1106),
.Y(n_1452)
);

OAI221xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1217),
.A2(n_1203),
.B1(n_1090),
.B2(n_1053),
.C(n_1065),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1220),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1307),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1276),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1234),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1243),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_L g1459 ( 
.A1(n_1261),
.A2(n_1170),
.B1(n_1037),
.B2(n_1052),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1240),
.A2(n_1112),
.B1(n_1140),
.B2(n_1046),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1281),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1360),
.B(n_1190),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1335),
.Y(n_1463)
);

NAND3xp33_ASAP7_75t_L g1464 ( 
.A(n_1363),
.B(n_1189),
.C(n_1180),
.Y(n_1464)
);

OA21x2_ASAP7_75t_L g1465 ( 
.A1(n_1253),
.A2(n_1185),
.B(n_1149),
.Y(n_1465)
);

INVx3_ASAP7_75t_L g1466 ( 
.A(n_1351),
.Y(n_1466)
);

NAND3xp33_ASAP7_75t_L g1467 ( 
.A(n_1359),
.B(n_1046),
.C(n_1194),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1307),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1319),
.B(n_1065),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1260),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1260),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1370),
.A2(n_1149),
.B(n_1046),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1264),
.Y(n_1473)
);

AND2x4_ASAP7_75t_L g1474 ( 
.A(n_1278),
.B(n_1076),
.Y(n_1474)
);

CKINVDCx11_ASAP7_75t_R g1475 ( 
.A(n_1296),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1360),
.B(n_1194),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1264),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1370),
.A2(n_1106),
.B(n_1091),
.Y(n_1478)
);

INVxp67_ASAP7_75t_L g1479 ( 
.A(n_1353),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1224),
.A2(n_1149),
.B(n_1194),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1335),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1351),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1362),
.Y(n_1483)
);

INVx1_ASAP7_75t_SL g1484 ( 
.A(n_1362),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1278),
.B(n_1076),
.Y(n_1485)
);

OAI21x1_ASAP7_75t_L g1486 ( 
.A1(n_1302),
.A2(n_1101),
.B(n_1091),
.Y(n_1486)
);

NAND2x1p5_ASAP7_75t_L g1487 ( 
.A(n_1351),
.B(n_1074),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1283),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1302),
.A2(n_1101),
.B(n_1091),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1318),
.B(n_1052),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_1317),
.Y(n_1491)
);

INVx3_ASAP7_75t_L g1492 ( 
.A(n_1206),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1235),
.A2(n_1304),
.B(n_1303),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1330),
.B(n_1161),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1243),
.B(n_1082),
.Y(n_1495)
);

OAI21x1_ASAP7_75t_L g1496 ( 
.A1(n_1303),
.A2(n_1304),
.B(n_1266),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1222),
.B(n_1161),
.Y(n_1497)
);

AOI21xp5_ASAP7_75t_L g1498 ( 
.A1(n_1218),
.A2(n_1077),
.B(n_1050),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1283),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1206),
.Y(n_1500)
);

INVx4_ASAP7_75t_L g1501 ( 
.A(n_1350),
.Y(n_1501)
);

OAI21xp5_ASAP7_75t_L g1502 ( 
.A1(n_1244),
.A2(n_1169),
.B(n_1074),
.Y(n_1502)
);

OAI21x1_ASAP7_75t_L g1503 ( 
.A1(n_1266),
.A2(n_1106),
.B(n_1091),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1285),
.B(n_1048),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1256),
.A2(n_1106),
.B(n_1091),
.Y(n_1505)
);

CKINVDCx5p33_ASAP7_75t_R g1506 ( 
.A(n_1317),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1284),
.Y(n_1507)
);

OAI22xp5_ASAP7_75t_L g1508 ( 
.A1(n_1239),
.A2(n_1203),
.B1(n_1169),
.B2(n_1112),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1284),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1290),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1212),
.B(n_1181),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1221),
.B(n_1082),
.Y(n_1512)
);

AND2x4_ASAP7_75t_L g1513 ( 
.A(n_1349),
.B(n_1048),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1310),
.A2(n_1181),
.B1(n_1160),
.B2(n_1048),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1256),
.A2(n_1101),
.B(n_1077),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1345),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1290),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1365),
.Y(n_1518)
);

BUFx2_ASAP7_75t_SL g1519 ( 
.A(n_1350),
.Y(n_1519)
);

OAI21x1_ASAP7_75t_L g1520 ( 
.A1(n_1258),
.A2(n_1097),
.B(n_1077),
.Y(n_1520)
);

BUFx3_ASAP7_75t_L g1521 ( 
.A(n_1229),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1308),
.Y(n_1522)
);

OAI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1263),
.A2(n_1160),
.B1(n_1142),
.B2(n_1157),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1235),
.A2(n_366),
.B(n_320),
.Y(n_1524)
);

OAI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1258),
.A2(n_1097),
.B(n_1077),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_1307),
.Y(n_1526)
);

INVxp33_ASAP7_75t_L g1527 ( 
.A(n_1295),
.Y(n_1527)
);

CKINVDCx6p67_ASAP7_75t_R g1528 ( 
.A(n_1349),
.Y(n_1528)
);

A2O1A1Ixp33_ASAP7_75t_L g1529 ( 
.A1(n_1247),
.A2(n_1142),
.B(n_1157),
.C(n_1145),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_L g1530 ( 
.A(n_1285),
.B(n_1048),
.Y(n_1530)
);

OAI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1305),
.A2(n_1097),
.B(n_1077),
.Y(n_1531)
);

AOI21xp33_ASAP7_75t_SL g1532 ( 
.A1(n_1297),
.A2(n_17),
.B(n_18),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1229),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1299),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1280),
.A2(n_1160),
.B1(n_1048),
.B2(n_1097),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1337),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1299),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1306),
.A2(n_1134),
.B1(n_1167),
.B2(n_1088),
.Y(n_1538)
);

XOR2xp5_ASAP7_75t_L g1539 ( 
.A(n_1259),
.B(n_1050),
.Y(n_1539)
);

AO21x2_ASAP7_75t_L g1540 ( 
.A1(n_1213),
.A2(n_1134),
.B(n_1097),
.Y(n_1540)
);

OA21x2_ASAP7_75t_L g1541 ( 
.A1(n_1219),
.A2(n_349),
.B(n_324),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1267),
.Y(n_1542)
);

NAND2x1p5_ASAP7_75t_L g1543 ( 
.A(n_1334),
.B(n_1050),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1226),
.A2(n_1134),
.B(n_1145),
.Y(n_1544)
);

BUFx8_ASAP7_75t_L g1545 ( 
.A(n_1350),
.Y(n_1545)
);

INVx4_ASAP7_75t_L g1546 ( 
.A(n_1350),
.Y(n_1546)
);

NOR2xp33_ASAP7_75t_L g1547 ( 
.A(n_1340),
.B(n_318),
.Y(n_1547)
);

AOI21xp5_ASAP7_75t_L g1548 ( 
.A1(n_1252),
.A2(n_1157),
.B(n_1145),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1288),
.A2(n_1157),
.B1(n_1145),
.B2(n_1142),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1259),
.A2(n_1134),
.B1(n_1145),
.B2(n_1142),
.Y(n_1550)
);

AOI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1333),
.A2(n_1134),
.B1(n_1157),
.B2(n_1142),
.Y(n_1551)
);

OAI21x1_ASAP7_75t_L g1552 ( 
.A1(n_1305),
.A2(n_1134),
.B(n_371),
.Y(n_1552)
);

NAND2x1p5_ASAP7_75t_L g1553 ( 
.A(n_1321),
.B(n_109),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1275),
.A2(n_365),
.B1(n_355),
.B2(n_337),
.C(n_334),
.Y(n_1554)
);

NOR2x1_ASAP7_75t_SL g1555 ( 
.A(n_1349),
.B(n_20),
.Y(n_1555)
);

AOI21xp5_ASAP7_75t_L g1556 ( 
.A1(n_1271),
.A2(n_333),
.B(n_331),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_1475),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1518),
.A2(n_1339),
.B1(n_1301),
.B2(n_1269),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1377),
.B(n_1326),
.Y(n_1559)
);

AO31x2_ASAP7_75t_L g1560 ( 
.A1(n_1414),
.A2(n_1339),
.A3(n_1293),
.B(n_1292),
.Y(n_1560)
);

OR2x2_ASAP7_75t_L g1561 ( 
.A(n_1400),
.B(n_1277),
.Y(n_1561)
);

INVx2_ASAP7_75t_L g1562 ( 
.A(n_1537),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1392),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_SL g1564 ( 
.A1(n_1386),
.A2(n_1287),
.B(n_1354),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1518),
.A2(n_1432),
.B1(n_1522),
.B2(n_1422),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1522),
.A2(n_1272),
.B1(n_1270),
.B2(n_1274),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1475),
.Y(n_1567)
);

NAND3xp33_ASAP7_75t_SL g1568 ( 
.A(n_1532),
.B(n_1332),
.C(n_1328),
.Y(n_1568)
);

AOI21xp33_ASAP7_75t_L g1569 ( 
.A1(n_1547),
.A2(n_1348),
.B(n_1322),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1537),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1393),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1479),
.B(n_24),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1381),
.Y(n_1573)
);

OAI22xp5_ASAP7_75t_L g1574 ( 
.A1(n_1453),
.A2(n_1373),
.B1(n_1460),
.B2(n_1516),
.Y(n_1574)
);

INVx4_ASAP7_75t_L g1575 ( 
.A(n_1461),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1502),
.B(n_1236),
.Y(n_1576)
);

AO21x2_ASAP7_75t_L g1577 ( 
.A1(n_1529),
.A2(n_1357),
.B(n_1262),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1375),
.A2(n_1371),
.B(n_1286),
.C(n_1282),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1399),
.Y(n_1579)
);

BUFx6f_ASAP7_75t_L g1580 ( 
.A(n_1380),
.Y(n_1580)
);

BUFx3_ASAP7_75t_L g1581 ( 
.A(n_1407),
.Y(n_1581)
);

AOI21xp5_ASAP7_75t_L g1582 ( 
.A1(n_1498),
.A2(n_1298),
.B(n_1327),
.Y(n_1582)
);

AND2x2_ASAP7_75t_L g1583 ( 
.A(n_1401),
.B(n_25),
.Y(n_1583)
);

OR2x6_ASAP7_75t_L g1584 ( 
.A(n_1451),
.B(n_1250),
.Y(n_1584)
);

AOI22xp33_ASAP7_75t_L g1585 ( 
.A1(n_1401),
.A2(n_1322),
.B1(n_1358),
.B2(n_1289),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1413),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1380),
.B(n_1326),
.Y(n_1587)
);

BUFx8_ASAP7_75t_SL g1588 ( 
.A(n_1431),
.Y(n_1588)
);

OAI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1400),
.A2(n_1347),
.B1(n_1364),
.B2(n_1315),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1378),
.B(n_1382),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1417),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1419),
.Y(n_1592)
);

NAND2xp33_ASAP7_75t_SL g1593 ( 
.A(n_1374),
.B(n_1294),
.Y(n_1593)
);

NAND2xp33_ASAP7_75t_R g1594 ( 
.A(n_1451),
.B(n_1322),
.Y(n_1594)
);

O2A1O1Ixp33_ASAP7_75t_SL g1595 ( 
.A1(n_1436),
.A2(n_1314),
.B(n_1327),
.C(n_1336),
.Y(n_1595)
);

INVxp67_ASAP7_75t_SL g1596 ( 
.A(n_1463),
.Y(n_1596)
);

INVxp67_ASAP7_75t_SL g1597 ( 
.A(n_1463),
.Y(n_1597)
);

OAI22xp5_ASAP7_75t_L g1598 ( 
.A1(n_1542),
.A2(n_1347),
.B1(n_1314),
.B2(n_1337),
.Y(n_1598)
);

NAND2x1p5_ASAP7_75t_L g1599 ( 
.A(n_1501),
.B(n_1338),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1467),
.A2(n_1368),
.B1(n_1367),
.B2(n_1342),
.Y(n_1600)
);

CKINVDCx16_ASAP7_75t_R g1601 ( 
.A(n_1431),
.Y(n_1601)
);

OAI22xp33_ASAP7_75t_L g1602 ( 
.A1(n_1404),
.A2(n_1451),
.B1(n_1512),
.B2(n_1490),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1378),
.A2(n_1358),
.B1(n_1338),
.B2(n_1273),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1456),
.A2(n_1343),
.B1(n_1358),
.B2(n_1316),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1421),
.B(n_1277),
.Y(n_1605)
);

AOI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1462),
.A2(n_1350),
.B1(n_1312),
.B2(n_1311),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1440),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1426),
.B(n_1277),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1449),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1416),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1476),
.B(n_27),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1476),
.B(n_27),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1462),
.B(n_1396),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1539),
.A2(n_1273),
.B1(n_1350),
.B2(n_1282),
.Y(n_1614)
);

INVx3_ASAP7_75t_L g1615 ( 
.A(n_1449),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1380),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1457),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1539),
.A2(n_1404),
.B1(n_1550),
.B2(n_1459),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1478),
.A2(n_1230),
.B(n_1251),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1483),
.B(n_28),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1484),
.B(n_28),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1449),
.B(n_32),
.Y(n_1622)
);

OAI211xp5_ASAP7_75t_L g1623 ( 
.A1(n_1464),
.A2(n_1286),
.B(n_325),
.C(n_1225),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1407),
.Y(n_1624)
);

BUFx3_ASAP7_75t_L g1625 ( 
.A(n_1437),
.Y(n_1625)
);

NOR3xp33_ASAP7_75t_SL g1626 ( 
.A(n_1491),
.B(n_33),
.C(n_36),
.Y(n_1626)
);

AND2x4_ASAP7_75t_L g1627 ( 
.A(n_1395),
.B(n_1250),
.Y(n_1627)
);

BUFx2_ASAP7_75t_L g1628 ( 
.A(n_1437),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1433),
.A2(n_1251),
.B(n_1225),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1513),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1470),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1385),
.Y(n_1632)
);

HB1xp67_ASAP7_75t_L g1633 ( 
.A(n_1455),
.Y(n_1633)
);

INVxp67_ASAP7_75t_L g1634 ( 
.A(n_1511),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1469),
.B(n_40),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1402),
.B(n_1277),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1458),
.B(n_1237),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1471),
.Y(n_1638)
);

BUFx2_ASAP7_75t_L g1639 ( 
.A(n_1469),
.Y(n_1639)
);

AND2x4_ASAP7_75t_L g1640 ( 
.A(n_1395),
.B(n_1307),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1473),
.Y(n_1641)
);

OR2x6_ASAP7_75t_L g1642 ( 
.A(n_1519),
.B(n_1273),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1477),
.Y(n_1643)
);

CKINVDCx14_ASAP7_75t_R g1644 ( 
.A(n_1461),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1436),
.A2(n_1237),
.B1(n_41),
.B2(n_43),
.C(n_45),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1488),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1499),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_SL g1648 ( 
.A(n_1527),
.B(n_40),
.C(n_46),
.Y(n_1648)
);

AND2x4_ASAP7_75t_L g1649 ( 
.A(n_1395),
.B(n_1412),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1403),
.Y(n_1650)
);

AOI21xp5_ASAP7_75t_L g1651 ( 
.A1(n_1480),
.A2(n_1237),
.B(n_1309),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1414),
.A2(n_1300),
.B1(n_1344),
.B2(n_50),
.Y(n_1652)
);

OAI22xp5_ASAP7_75t_L g1653 ( 
.A1(n_1527),
.A2(n_46),
.B1(n_47),
.B2(n_50),
.Y(n_1653)
);

OAI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1508),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1424),
.B(n_1511),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1443),
.A2(n_1344),
.A3(n_1300),
.B(n_1309),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1507),
.Y(n_1657)
);

CKINVDCx20_ASAP7_75t_R g1658 ( 
.A(n_1403),
.Y(n_1658)
);

AOI211xp5_ASAP7_75t_L g1659 ( 
.A1(n_1554),
.A2(n_1458),
.B(n_1495),
.C(n_1442),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1509),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1510),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1538),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_1662)
);

BUFx6f_ASAP7_75t_L g1663 ( 
.A(n_1406),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1412),
.B(n_1309),
.Y(n_1664)
);

AOI22xp33_ASAP7_75t_L g1665 ( 
.A1(n_1443),
.A2(n_1300),
.B1(n_1344),
.B2(n_59),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1517),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1474),
.B(n_1485),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1469),
.B(n_55),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1556),
.A2(n_57),
.B1(n_61),
.B2(n_62),
.C(n_64),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1474),
.B(n_1344),
.Y(n_1670)
);

AOI22xp33_ASAP7_75t_SL g1671 ( 
.A1(n_1545),
.A2(n_1300),
.B1(n_67),
.B2(n_68),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1434),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_L g1673 ( 
.A1(n_1552),
.A2(n_231),
.B(n_228),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_L g1674 ( 
.A1(n_1529),
.A2(n_71),
.B(n_72),
.Y(n_1674)
);

INVx5_ASAP7_75t_L g1675 ( 
.A(n_1501),
.Y(n_1675)
);

AOI22xp33_ASAP7_75t_L g1676 ( 
.A1(n_1424),
.A2(n_72),
.B1(n_73),
.B2(n_74),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_L g1677 ( 
.A1(n_1545),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_SL g1678 ( 
.A(n_1523),
.B(n_75),
.Y(n_1678)
);

AO32x2_ASAP7_75t_L g1679 ( 
.A1(n_1514),
.A2(n_78),
.A3(n_79),
.B1(n_80),
.B2(n_81),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1534),
.Y(n_1680)
);

OAI22xp5_ASAP7_75t_L g1681 ( 
.A1(n_1528),
.A2(n_79),
.B1(n_83),
.B2(n_84),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1494),
.B(n_85),
.Y(n_1682)
);

OAI221xp5_ASAP7_75t_L g1683 ( 
.A1(n_1465),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.C(n_88),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1445),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1513),
.Y(n_1685)
);

OAI22xp33_ASAP7_75t_L g1686 ( 
.A1(n_1528),
.A2(n_88),
.B1(n_89),
.B2(n_91),
.Y(n_1686)
);

CKINVDCx20_ASAP7_75t_R g1687 ( 
.A(n_1403),
.Y(n_1687)
);

OAI22xp5_ASAP7_75t_L g1688 ( 
.A1(n_1487),
.A2(n_92),
.B1(n_94),
.B2(n_96),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1423),
.Y(n_1689)
);

O2A1O1Ixp33_ASAP7_75t_SL g1690 ( 
.A1(n_1450),
.A2(n_98),
.B(n_100),
.C(n_101),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1423),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1474),
.B(n_100),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1485),
.B(n_101),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1494),
.A2(n_102),
.B1(n_115),
.B2(n_117),
.C(n_123),
.Y(n_1694)
);

BUFx3_ASAP7_75t_L g1695 ( 
.A(n_1485),
.Y(n_1695)
);

NOR2x1_ASAP7_75t_SL g1696 ( 
.A(n_1374),
.B(n_102),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_L g1697 ( 
.A1(n_1465),
.A2(n_226),
.B1(n_136),
.B2(n_143),
.C(n_146),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1429),
.Y(n_1698)
);

AOI22xp33_ASAP7_75t_L g1699 ( 
.A1(n_1545),
.A2(n_225),
.B1(n_148),
.B2(n_159),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1513),
.Y(n_1700)
);

INVx1_ASAP7_75t_SL g1701 ( 
.A(n_1445),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1487),
.A2(n_135),
.B1(n_183),
.B2(n_187),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1548),
.A2(n_224),
.B(n_197),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1390),
.B(n_193),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1390),
.B(n_207),
.Y(n_1705)
);

AOI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1434),
.A2(n_209),
.B1(n_213),
.B2(n_220),
.Y(n_1706)
);

NAND2xp33_ASAP7_75t_R g1707 ( 
.A(n_1472),
.B(n_1465),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1434),
.A2(n_1406),
.B1(n_1546),
.B2(n_1501),
.Y(n_1708)
);

BUFx2_ASAP7_75t_L g1709 ( 
.A(n_1497),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1497),
.B(n_1521),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1406),
.B(n_1444),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1429),
.Y(n_1712)
);

BUFx2_ASAP7_75t_L g1713 ( 
.A(n_1497),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1446),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1390),
.B(n_1409),
.Y(n_1715)
);

BUFx2_ASAP7_75t_L g1716 ( 
.A(n_1406),
.Y(n_1716)
);

BUFx3_ASAP7_75t_L g1717 ( 
.A(n_1409),
.Y(n_1717)
);

INVx6_ASAP7_75t_L g1718 ( 
.A(n_1409),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1546),
.A2(n_1551),
.B1(n_1446),
.B2(n_1374),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1439),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1444),
.B(n_1491),
.Y(n_1721)
);

AND2x4_ASAP7_75t_L g1722 ( 
.A(n_1521),
.B(n_1492),
.Y(n_1722)
);

INVx3_ASAP7_75t_L g1723 ( 
.A(n_1492),
.Y(n_1723)
);

AOI22xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1555),
.A2(n_1546),
.B1(n_1438),
.B2(n_1524),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_SL g1725 ( 
.A1(n_1438),
.A2(n_1524),
.B1(n_1541),
.B2(n_1553),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1444),
.B(n_1506),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1506),
.B(n_1444),
.Y(n_1727)
);

OR2x6_ASAP7_75t_L g1728 ( 
.A(n_1428),
.B(n_1553),
.Y(n_1728)
);

OR2x6_ASAP7_75t_L g1729 ( 
.A(n_1553),
.B(n_1492),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1444),
.B(n_1389),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1441),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1500),
.B(n_1533),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1439),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1441),
.Y(n_1734)
);

AOI22xp33_ASAP7_75t_L g1735 ( 
.A1(n_1524),
.A2(n_1379),
.B1(n_1541),
.B2(n_1376),
.Y(n_1735)
);

INVx3_ASAP7_75t_SL g1736 ( 
.A(n_1441),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_L g1737 ( 
.A(n_1420),
.B(n_1533),
.Y(n_1737)
);

INVx3_ASAP7_75t_L g1738 ( 
.A(n_1500),
.Y(n_1738)
);

OR2x2_ASAP7_75t_L g1739 ( 
.A(n_1389),
.B(n_1504),
.Y(n_1739)
);

INVx2_ASAP7_75t_L g1740 ( 
.A(n_1481),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_L g1741 ( 
.A1(n_1379),
.A2(n_1541),
.B1(n_1376),
.B2(n_1468),
.Y(n_1741)
);

BUFx2_ASAP7_75t_L g1742 ( 
.A(n_1504),
.Y(n_1742)
);

INVx2_ASAP7_75t_SL g1743 ( 
.A(n_1500),
.Y(n_1743)
);

INVx3_ASAP7_75t_L g1744 ( 
.A(n_1533),
.Y(n_1744)
);

AOI22xp33_ASAP7_75t_L g1745 ( 
.A1(n_1376),
.A2(n_1455),
.B1(n_1526),
.B2(n_1468),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1450),
.B(n_1482),
.Y(n_1746)
);

INVx6_ASAP7_75t_L g1747 ( 
.A(n_1420),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1481),
.Y(n_1748)
);

AND2x6_ASAP7_75t_L g1749 ( 
.A(n_1536),
.B(n_1450),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1389),
.B(n_1454),
.Y(n_1750)
);

NOR2x1p5_ASAP7_75t_L g1751 ( 
.A(n_1454),
.B(n_1466),
.Y(n_1751)
);

INVx1_ASAP7_75t_SL g1752 ( 
.A(n_1504),
.Y(n_1752)
);

CKINVDCx5p33_ASAP7_75t_R g1753 ( 
.A(n_1454),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1389),
.B(n_1482),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1563),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1590),
.B(n_1389),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1634),
.B(n_1526),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1634),
.B(n_1655),
.Y(n_1758)
);

CKINVDCx5p33_ASAP7_75t_R g1759 ( 
.A(n_1588),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1677),
.A2(n_1482),
.B1(n_1466),
.B2(n_1530),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1727),
.B(n_1438),
.Y(n_1761)
);

AOI22xp33_ASAP7_75t_L g1762 ( 
.A1(n_1618),
.A2(n_1574),
.B1(n_1686),
.B2(n_1676),
.Y(n_1762)
);

AOI22xp33_ASAP7_75t_L g1763 ( 
.A1(n_1618),
.A2(n_1408),
.B1(n_1544),
.B2(n_1397),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_SL g1764 ( 
.A1(n_1686),
.A2(n_1535),
.B1(n_1549),
.B2(n_1466),
.C(n_1438),
.Y(n_1764)
);

BUFx4f_ASAP7_75t_SL g1765 ( 
.A(n_1650),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1676),
.A2(n_1408),
.B1(n_1544),
.B2(n_1397),
.Y(n_1766)
);

OAI221xp5_ASAP7_75t_L g1767 ( 
.A1(n_1565),
.A2(n_1408),
.B1(n_1397),
.B2(n_1530),
.C(n_1543),
.Y(n_1767)
);

OAI21x1_ASAP7_75t_L g1768 ( 
.A1(n_1619),
.A2(n_1496),
.B(n_1552),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1683),
.A2(n_1747),
.B1(n_1558),
.B2(n_1613),
.Y(n_1769)
);

BUFx2_ASAP7_75t_L g1770 ( 
.A(n_1750),
.Y(n_1770)
);

AOI221xp5_ASAP7_75t_L g1771 ( 
.A1(n_1648),
.A2(n_1438),
.B1(n_1544),
.B2(n_1540),
.C(n_1536),
.Y(n_1771)
);

OAI322xp33_ASAP7_75t_L g1772 ( 
.A1(n_1672),
.A2(n_1530),
.A3(n_1543),
.B1(n_1388),
.B2(n_1536),
.C1(n_1540),
.C2(n_1493),
.Y(n_1772)
);

OAI22xp33_ASAP7_75t_L g1773 ( 
.A1(n_1681),
.A2(n_1543),
.B1(n_1388),
.B2(n_1472),
.Y(n_1773)
);

INVx1_ASAP7_75t_SL g1774 ( 
.A(n_1684),
.Y(n_1774)
);

AOI22xp5_ASAP7_75t_SL g1775 ( 
.A1(n_1658),
.A2(n_1687),
.B1(n_1644),
.B2(n_1731),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1571),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1701),
.Y(n_1777)
);

AO221x2_ASAP7_75t_L g1778 ( 
.A1(n_1653),
.A2(n_1540),
.B1(n_1418),
.B2(n_1415),
.C(n_1472),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1614),
.A2(n_1447),
.B1(n_1493),
.B2(n_1398),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1677),
.B(n_1626),
.C(n_1669),
.Y(n_1780)
);

AOI221xp5_ASAP7_75t_L g1781 ( 
.A1(n_1645),
.A2(n_1493),
.B1(n_1447),
.B2(n_1398),
.C(n_1411),
.Y(n_1781)
);

AND2x4_ASAP7_75t_L g1782 ( 
.A(n_1640),
.B(n_1452),
.Y(n_1782)
);

HB1xp67_ASAP7_75t_L g1783 ( 
.A(n_1624),
.Y(n_1783)
);

OAI22xp5_ASAP7_75t_L g1784 ( 
.A1(n_1626),
.A2(n_1418),
.B1(n_1415),
.B2(n_1452),
.Y(n_1784)
);

CKINVDCx14_ASAP7_75t_R g1785 ( 
.A(n_1644),
.Y(n_1785)
);

OAI22xp5_ASAP7_75t_L g1786 ( 
.A1(n_1566),
.A2(n_1435),
.B1(n_1448),
.B2(n_1430),
.Y(n_1786)
);

OAI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1747),
.A2(n_1435),
.B1(n_1448),
.B2(n_1531),
.Y(n_1787)
);

OAI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1682),
.A2(n_1425),
.B1(n_1427),
.B2(n_1430),
.Y(n_1788)
);

AOI22xp33_ASAP7_75t_SL g1789 ( 
.A1(n_1747),
.A2(n_1486),
.B1(n_1489),
.B2(n_1384),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_SL g1790 ( 
.A1(n_1736),
.A2(n_1601),
.B1(n_1575),
.B2(n_1731),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1573),
.B(n_1486),
.Y(n_1791)
);

AOI22xp33_ASAP7_75t_L g1792 ( 
.A1(n_1614),
.A2(n_1411),
.B1(n_1410),
.B2(n_1405),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1721),
.B(n_1410),
.Y(n_1793)
);

OAI22xp33_ASAP7_75t_L g1794 ( 
.A1(n_1654),
.A2(n_1405),
.B1(n_1425),
.B2(n_1427),
.Y(n_1794)
);

BUFx6f_ASAP7_75t_L g1795 ( 
.A(n_1675),
.Y(n_1795)
);

OAI211xp5_ASAP7_75t_SL g1796 ( 
.A1(n_1726),
.A2(n_1503),
.B(n_1520),
.C(n_1515),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1682),
.A2(n_1525),
.B1(n_1520),
.B2(n_1515),
.Y(n_1797)
);

OAI211xp5_ASAP7_75t_L g1798 ( 
.A1(n_1690),
.A2(n_1525),
.B(n_1505),
.C(n_1384),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1579),
.B(n_1505),
.Y(n_1799)
);

AOI22xp33_ASAP7_75t_L g1800 ( 
.A1(n_1561),
.A2(n_1372),
.B1(n_1383),
.B2(n_1387),
.Y(n_1800)
);

AOI22xp33_ASAP7_75t_L g1801 ( 
.A1(n_1568),
.A2(n_1569),
.B1(n_1602),
.B2(n_1671),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1586),
.Y(n_1802)
);

OAI221xp5_ASAP7_75t_L g1803 ( 
.A1(n_1659),
.A2(n_1372),
.B1(n_1383),
.B2(n_1387),
.C(n_1391),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1605),
.Y(n_1804)
);

OAI21x1_ASAP7_75t_L g1805 ( 
.A1(n_1582),
.A2(n_1391),
.B(n_1394),
.Y(n_1805)
);

OAI22xp33_ASAP7_75t_L g1806 ( 
.A1(n_1662),
.A2(n_1394),
.B1(n_1678),
.B2(n_1706),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1740),
.Y(n_1807)
);

INVx6_ASAP7_75t_L g1808 ( 
.A(n_1580),
.Y(n_1808)
);

AOI322xp5_ASAP7_75t_L g1809 ( 
.A1(n_1602),
.A2(n_1671),
.A3(n_1678),
.B1(n_1583),
.B2(n_1725),
.C1(n_1585),
.C2(n_1636),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1587),
.A2(n_1640),
.B1(n_1711),
.B2(n_1725),
.Y(n_1810)
);

CKINVDCx5p33_ASAP7_75t_R g1811 ( 
.A(n_1588),
.Y(n_1811)
);

AOI21x1_ASAP7_75t_L g1812 ( 
.A1(n_1651),
.A2(n_1629),
.B(n_1604),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1633),
.B(n_1730),
.Y(n_1813)
);

AOI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1587),
.A2(n_1585),
.B1(n_1608),
.B2(n_1627),
.Y(n_1814)
);

AOI21x1_ASAP7_75t_L g1815 ( 
.A1(n_1629),
.A2(n_1564),
.B(n_1674),
.Y(n_1815)
);

AOI22xp33_ASAP7_75t_SL g1816 ( 
.A1(n_1697),
.A2(n_1623),
.B1(n_1696),
.B2(n_1612),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1592),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1627),
.A2(n_1724),
.B1(n_1631),
.B2(n_1617),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1633),
.B(n_1754),
.Y(n_1819)
);

AOI22xp33_ASAP7_75t_L g1820 ( 
.A1(n_1724),
.A2(n_1603),
.B1(n_1694),
.B2(n_1611),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1591),
.Y(n_1821)
);

OA21x2_ASAP7_75t_L g1822 ( 
.A1(n_1578),
.A2(n_1735),
.B(n_1741),
.Y(n_1822)
);

OR2x2_ASAP7_75t_SL g1823 ( 
.A(n_1637),
.B(n_1718),
.Y(n_1823)
);

OA21x2_ASAP7_75t_L g1824 ( 
.A1(n_1578),
.A2(n_1735),
.B(n_1741),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1603),
.A2(n_1642),
.B1(n_1670),
.B2(n_1699),
.Y(n_1825)
);

AOI21xp5_ASAP7_75t_L g1826 ( 
.A1(n_1595),
.A2(n_1593),
.B(n_1576),
.Y(n_1826)
);

AOI222xp33_ASAP7_75t_L g1827 ( 
.A1(n_1688),
.A2(n_1572),
.B1(n_1699),
.B2(n_1576),
.C1(n_1620),
.C2(n_1621),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_L g1828 ( 
.A1(n_1642),
.A2(n_1584),
.B1(n_1641),
.B2(n_1643),
.Y(n_1828)
);

INVx4_ASAP7_75t_SL g1829 ( 
.A(n_1749),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1559),
.B(n_1628),
.Y(n_1830)
);

AOI22xp33_ASAP7_75t_L g1831 ( 
.A1(n_1642),
.A2(n_1584),
.B1(n_1680),
.B2(n_1657),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1740),
.Y(n_1832)
);

AOI21xp5_ASAP7_75t_L g1833 ( 
.A1(n_1595),
.A2(n_1593),
.B(n_1719),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1607),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1719),
.A2(n_1729),
.B(n_1728),
.Y(n_1835)
);

AOI22xp33_ASAP7_75t_L g1836 ( 
.A1(n_1584),
.A2(n_1660),
.B1(n_1638),
.B2(n_1646),
.Y(n_1836)
);

AOI22xp33_ASAP7_75t_L g1837 ( 
.A1(n_1647),
.A2(n_1661),
.B1(n_1666),
.B2(n_1664),
.Y(n_1837)
);

OAI222xp33_ASAP7_75t_L g1838 ( 
.A1(n_1652),
.A2(n_1665),
.B1(n_1589),
.B2(n_1693),
.C1(n_1692),
.C2(n_1728),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_L g1839 ( 
.A1(n_1632),
.A2(n_1753),
.B1(n_1718),
.B2(n_1736),
.Y(n_1839)
);

OAI22xp33_ASAP7_75t_L g1840 ( 
.A1(n_1606),
.A2(n_1575),
.B1(n_1639),
.B2(n_1667),
.Y(n_1840)
);

BUFx4f_ASAP7_75t_SL g1841 ( 
.A(n_1734),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1718),
.A2(n_1589),
.B1(n_1717),
.B2(n_1751),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1664),
.A2(n_1710),
.B1(n_1713),
.B2(n_1709),
.Y(n_1843)
);

INVx4_ASAP7_75t_L g1844 ( 
.A(n_1749),
.Y(n_1844)
);

AOI221xp5_ASAP7_75t_L g1845 ( 
.A1(n_1690),
.A2(n_1652),
.B1(n_1665),
.B2(n_1702),
.C(n_1600),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1635),
.A2(n_1668),
.B1(n_1745),
.B2(n_1705),
.C(n_1704),
.Y(n_1846)
);

AOI22xp33_ASAP7_75t_L g1847 ( 
.A1(n_1710),
.A2(n_1722),
.B1(n_1700),
.B2(n_1685),
.Y(n_1847)
);

AOI21xp5_ASAP7_75t_L g1848 ( 
.A1(n_1729),
.A2(n_1728),
.B(n_1598),
.Y(n_1848)
);

OAI221xp5_ASAP7_75t_L g1849 ( 
.A1(n_1594),
.A2(n_1707),
.B1(n_1622),
.B2(n_1752),
.C(n_1703),
.Y(n_1849)
);

OAI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1594),
.A2(n_1707),
.B1(n_1743),
.B2(n_1717),
.C(n_1625),
.Y(n_1850)
);

OAI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1708),
.A2(n_1737),
.B1(n_1714),
.B2(n_1581),
.Y(n_1851)
);

OAI22xp5_ASAP7_75t_L g1852 ( 
.A1(n_1708),
.A2(n_1737),
.B1(n_1625),
.B2(n_1581),
.Y(n_1852)
);

INVx1_ASAP7_75t_SL g1853 ( 
.A(n_1715),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1679),
.B(n_1742),
.Y(n_1854)
);

OAI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1557),
.A2(n_1567),
.B1(n_1746),
.B2(n_1609),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1722),
.A2(n_1700),
.B1(n_1630),
.B2(n_1685),
.Y(n_1856)
);

AND2x4_ASAP7_75t_L g1857 ( 
.A(n_1630),
.B(n_1675),
.Y(n_1857)
);

AOI22xp33_ASAP7_75t_L g1858 ( 
.A1(n_1562),
.A2(n_1570),
.B1(n_1580),
.B2(n_1616),
.Y(n_1858)
);

AOI211xp5_ASAP7_75t_L g1859 ( 
.A1(n_1679),
.A2(n_1663),
.B(n_1732),
.C(n_1716),
.Y(n_1859)
);

AOI22xp33_ASAP7_75t_L g1860 ( 
.A1(n_1570),
.A2(n_1580),
.B1(n_1616),
.B2(n_1649),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1580),
.A2(n_1616),
.B1(n_1649),
.B2(n_1663),
.Y(n_1861)
);

BUFx6f_ASAP7_75t_L g1862 ( 
.A(n_1675),
.Y(n_1862)
);

NAND2xp5_ASAP7_75t_L g1863 ( 
.A(n_1609),
.B(n_1615),
.Y(n_1863)
);

AOI22xp33_ASAP7_75t_SL g1864 ( 
.A1(n_1679),
.A2(n_1675),
.B1(n_1616),
.B2(n_1695),
.Y(n_1864)
);

AOI221xp5_ASAP7_75t_L g1865 ( 
.A1(n_1745),
.A2(n_1679),
.B1(n_1596),
.B2(n_1597),
.C(n_1748),
.Y(n_1865)
);

BUFx3_ASAP7_75t_L g1866 ( 
.A(n_1695),
.Y(n_1866)
);

AOI222xp33_ASAP7_75t_L g1867 ( 
.A1(n_1732),
.A2(n_1689),
.B1(n_1691),
.B2(n_1733),
.C1(n_1720),
.C2(n_1712),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1615),
.B(n_1656),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1596),
.B(n_1597),
.Y(n_1869)
);

AOI22xp5_ASAP7_75t_L g1870 ( 
.A1(n_1663),
.A2(n_1729),
.B1(n_1749),
.B2(n_1744),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1698),
.Y(n_1871)
);

OAI221xp5_ASAP7_75t_L g1872 ( 
.A1(n_1723),
.A2(n_1738),
.B1(n_1744),
.B2(n_1663),
.C(n_1599),
.Y(n_1872)
);

BUFx2_ASAP7_75t_L g1873 ( 
.A(n_1749),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1610),
.A2(n_1738),
.B1(n_1723),
.B2(n_1749),
.Y(n_1874)
);

AOI22xp33_ASAP7_75t_L g1875 ( 
.A1(n_1599),
.A2(n_1577),
.B1(n_1746),
.B2(n_1629),
.Y(n_1875)
);

INVx3_ASAP7_75t_L g1876 ( 
.A(n_1560),
.Y(n_1876)
);

AOI22xp33_ASAP7_75t_L g1877 ( 
.A1(n_1577),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1560),
.B(n_1673),
.Y(n_1878)
);

AOI22xp33_ASAP7_75t_L g1879 ( 
.A1(n_1560),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1879)
);

INVx1_ASAP7_75t_SL g1880 ( 
.A(n_1684),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1634),
.B(n_1655),
.Y(n_1881)
);

OAI211xp5_ASAP7_75t_SL g1882 ( 
.A1(n_1626),
.A2(n_1109),
.B(n_988),
.C(n_1013),
.Y(n_1882)
);

OA21x2_ASAP7_75t_L g1883 ( 
.A1(n_1578),
.A2(n_1735),
.B(n_1619),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1677),
.A2(n_1518),
.B1(n_760),
.B2(n_899),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_L g1885 ( 
.A(n_1677),
.B(n_1676),
.C(n_1626),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1563),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1887)
);

AOI221xp5_ASAP7_75t_L g1888 ( 
.A1(n_1686),
.A2(n_925),
.B1(n_1676),
.B2(n_1683),
.C(n_1297),
.Y(n_1888)
);

OA21x2_ASAP7_75t_L g1889 ( 
.A1(n_1578),
.A2(n_1735),
.B(n_1619),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1655),
.B(n_1633),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1581),
.Y(n_1891)
);

AOI22xp33_ASAP7_75t_SL g1892 ( 
.A1(n_1574),
.A2(n_1055),
.B1(n_464),
.B2(n_596),
.Y(n_1892)
);

AOI22xp33_ASAP7_75t_SL g1893 ( 
.A1(n_1574),
.A2(n_1055),
.B1(n_464),
.B2(n_596),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1578),
.A2(n_1034),
.B(n_1595),
.Y(n_1894)
);

AOI22xp33_ASAP7_75t_L g1895 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1895)
);

AOI21xp5_ASAP7_75t_L g1896 ( 
.A1(n_1578),
.A2(n_1034),
.B(n_1595),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1563),
.Y(n_1897)
);

BUFx2_ASAP7_75t_L g1898 ( 
.A(n_1750),
.Y(n_1898)
);

AOI22xp33_ASAP7_75t_L g1899 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1899)
);

A2O1A1Ixp33_ASAP7_75t_L g1900 ( 
.A1(n_1645),
.A2(n_1204),
.B(n_899),
.C(n_1386),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1558),
.A2(n_760),
.B(n_1386),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1574),
.A2(n_927),
.B1(n_1522),
.B2(n_760),
.Y(n_1902)
);

AOI22xp33_ASAP7_75t_SL g1903 ( 
.A1(n_1574),
.A2(n_1055),
.B1(n_464),
.B2(n_596),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1563),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1906)
);

AOI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1634),
.B(n_1655),
.Y(n_1908)
);

BUFx12f_ASAP7_75t_L g1909 ( 
.A(n_1650),
.Y(n_1909)
);

OA21x2_ASAP7_75t_L g1910 ( 
.A1(n_1578),
.A2(n_1735),
.B(n_1619),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1563),
.Y(n_1911)
);

AOI22xp33_ASAP7_75t_SL g1912 ( 
.A1(n_1574),
.A2(n_1055),
.B1(n_464),
.B2(n_596),
.Y(n_1912)
);

NOR2xp67_ASAP7_75t_L g1913 ( 
.A(n_1575),
.B(n_1458),
.Y(n_1913)
);

OAI21xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1677),
.A2(n_1676),
.B(n_1751),
.Y(n_1914)
);

AOI22xp33_ASAP7_75t_L g1915 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1915)
);

AOI22xp33_ASAP7_75t_L g1916 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1916)
);

AOI221xp5_ASAP7_75t_L g1917 ( 
.A1(n_1686),
.A2(n_925),
.B1(n_1676),
.B2(n_1683),
.C(n_1297),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1918)
);

AOI221xp5_ASAP7_75t_L g1919 ( 
.A1(n_1686),
.A2(n_925),
.B1(n_1676),
.B2(n_1683),
.C(n_1297),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1634),
.B(n_1655),
.Y(n_1920)
);

OAI22xp33_ASAP7_75t_L g1921 ( 
.A1(n_1686),
.A2(n_899),
.B1(n_1672),
.B2(n_1055),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1922)
);

AOI22xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1574),
.A2(n_1055),
.B1(n_464),
.B2(n_596),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1590),
.B(n_1573),
.Y(n_1924)
);

HB1xp67_ASAP7_75t_L g1925 ( 
.A(n_1634),
.Y(n_1925)
);

AOI21xp33_ASAP7_75t_L g1926 ( 
.A1(n_1594),
.A2(n_1574),
.B(n_1569),
.Y(n_1926)
);

INVx3_ASAP7_75t_L g1927 ( 
.A(n_1739),
.Y(n_1927)
);

AOI22xp33_ASAP7_75t_L g1928 ( 
.A1(n_1618),
.A2(n_1055),
.B1(n_1124),
.B2(n_1108),
.Y(n_1928)
);

AO21x2_ASAP7_75t_L g1929 ( 
.A1(n_1926),
.A2(n_1812),
.B(n_1878),
.Y(n_1929)
);

AND2x2_ASAP7_75t_L g1930 ( 
.A(n_1799),
.B(n_1793),
.Y(n_1930)
);

BUFx3_ASAP7_75t_L g1931 ( 
.A(n_1823),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1807),
.Y(n_1932)
);

INVx2_ASAP7_75t_L g1933 ( 
.A(n_1807),
.Y(n_1933)
);

AND2x2_ASAP7_75t_L g1934 ( 
.A(n_1799),
.B(n_1793),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1832),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1770),
.B(n_1898),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1834),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1819),
.B(n_1761),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1819),
.B(n_1761),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1755),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1776),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1802),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1817),
.Y(n_1944)
);

HB1xp67_ASAP7_75t_L g1945 ( 
.A(n_1813),
.Y(n_1945)
);

INVx4_ASAP7_75t_L g1946 ( 
.A(n_1844),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1886),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1948)
);

OR2x2_ASAP7_75t_L g1949 ( 
.A(n_1890),
.B(n_1813),
.Y(n_1949)
);

HB1xp67_ASAP7_75t_L g1950 ( 
.A(n_1925),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1897),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1905),
.Y(n_1952)
);

BUFx2_ASAP7_75t_L g1953 ( 
.A(n_1823),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1812),
.Y(n_1954)
);

HB1xp67_ASAP7_75t_L g1955 ( 
.A(n_1890),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1770),
.B(n_1898),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1911),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_L g1958 ( 
.A(n_1804),
.B(n_1756),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1871),
.Y(n_1959)
);

BUFx3_ASAP7_75t_L g1960 ( 
.A(n_1873),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1804),
.Y(n_1961)
);

BUFx2_ASAP7_75t_L g1962 ( 
.A(n_1783),
.Y(n_1962)
);

BUFx3_ASAP7_75t_L g1963 ( 
.A(n_1873),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1821),
.Y(n_1964)
);

INVx2_ASAP7_75t_SL g1965 ( 
.A(n_1891),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1782),
.B(n_1881),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1881),
.B(n_1908),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1830),
.B(n_1908),
.Y(n_1968)
);

BUFx2_ASAP7_75t_L g1969 ( 
.A(n_1891),
.Y(n_1969)
);

AND2x2_ASAP7_75t_L g1970 ( 
.A(n_1920),
.B(n_1757),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1791),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1920),
.B(n_1854),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1854),
.B(n_1757),
.Y(n_1973)
);

NAND2xp5_ASAP7_75t_L g1974 ( 
.A(n_1859),
.B(n_1764),
.Y(n_1974)
);

NOR2xp33_ASAP7_75t_L g1975 ( 
.A(n_1774),
.B(n_1777),
.Y(n_1975)
);

AND2x2_ASAP7_75t_L g1976 ( 
.A(n_1883),
.B(n_1889),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1869),
.B(n_1865),
.Y(n_1977)
);

BUFx2_ASAP7_75t_L g1978 ( 
.A(n_1866),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1880),
.B(n_1841),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1869),
.Y(n_1980)
);

INVx3_ASAP7_75t_L g1981 ( 
.A(n_1883),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1771),
.B(n_1887),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1868),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1868),
.Y(n_1984)
);

INVx3_ASAP7_75t_L g1985 ( 
.A(n_1883),
.Y(n_1985)
);

OR2x2_ASAP7_75t_L g1986 ( 
.A(n_1927),
.B(n_1922),
.Y(n_1986)
);

INVxp67_ASAP7_75t_L g1987 ( 
.A(n_1803),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1889),
.B(n_1910),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1889),
.B(n_1910),
.Y(n_1989)
);

AND2x4_ASAP7_75t_L g1990 ( 
.A(n_1829),
.B(n_1844),
.Y(n_1990)
);

AND2x4_ASAP7_75t_L g1991 ( 
.A(n_1829),
.B(n_1857),
.Y(n_1991)
);

AND2x2_ASAP7_75t_L g1992 ( 
.A(n_1910),
.B(n_1876),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_L g1993 ( 
.A(n_1924),
.B(n_1840),
.Y(n_1993)
);

AOI21xp5_ASAP7_75t_L g1994 ( 
.A1(n_1894),
.A2(n_1896),
.B(n_1833),
.Y(n_1994)
);

OR2x2_ASAP7_75t_L g1995 ( 
.A(n_1822),
.B(n_1824),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1876),
.B(n_1822),
.Y(n_1996)
);

AND2x2_ASAP7_75t_L g1997 ( 
.A(n_1876),
.B(n_1822),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1867),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1826),
.B(n_1797),
.Y(n_1999)
);

INVx1_ASAP7_75t_L g2000 ( 
.A(n_1863),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1778),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1778),
.Y(n_2002)
);

INVx4_ASAP7_75t_L g2003 ( 
.A(n_1795),
.Y(n_2003)
);

AND2x4_ASAP7_75t_L g2004 ( 
.A(n_1857),
.B(n_1835),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1836),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1853),
.B(n_1810),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1788),
.B(n_1864),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1824),
.B(n_1800),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1824),
.B(n_1779),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1778),
.B(n_1792),
.Y(n_2010)
);

INVxp67_ASAP7_75t_L g2011 ( 
.A(n_1767),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1837),
.Y(n_2012)
);

NAND2x1p5_ASAP7_75t_L g2013 ( 
.A(n_1795),
.B(n_1862),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1957),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1957),
.Y(n_2015)
);

NAND4xp25_ASAP7_75t_SL g2016 ( 
.A(n_2010),
.B(n_1885),
.C(n_1780),
.D(n_1902),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1938),
.B(n_1875),
.Y(n_2017)
);

BUFx3_ASAP7_75t_L g2018 ( 
.A(n_1978),
.Y(n_2018)
);

AOI22xp33_ASAP7_75t_L g2019 ( 
.A1(n_1998),
.A2(n_1762),
.B1(n_1921),
.B2(n_1892),
.Y(n_2019)
);

AOI22xp5_ASAP7_75t_L g2020 ( 
.A1(n_2011),
.A2(n_1914),
.B1(n_1884),
.B2(n_1901),
.Y(n_2020)
);

CKINVDCx20_ASAP7_75t_R g2021 ( 
.A(n_1979),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1938),
.B(n_1789),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_SL g2023 ( 
.A(n_2002),
.B(n_1842),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1932),
.Y(n_2024)
);

AND2x2_ASAP7_75t_SL g2025 ( 
.A(n_1953),
.B(n_1801),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1938),
.B(n_1828),
.Y(n_2026)
);

AO21x1_ASAP7_75t_SL g2027 ( 
.A1(n_2007),
.A2(n_1838),
.B(n_1818),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1955),
.Y(n_2028)
);

BUFx2_ASAP7_75t_L g2029 ( 
.A(n_1969),
.Y(n_2029)
);

NAND3xp33_ASAP7_75t_L g2030 ( 
.A(n_1987),
.B(n_1809),
.C(n_1845),
.Y(n_2030)
);

AOI21xp5_ASAP7_75t_L g2031 ( 
.A1(n_1994),
.A2(n_1900),
.B(n_1806),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1955),
.B(n_1852),
.Y(n_2032)
);

INVxp67_ASAP7_75t_L g2033 ( 
.A(n_1962),
.Y(n_2033)
);

INVxp67_ASAP7_75t_SL g2034 ( 
.A(n_1936),
.Y(n_2034)
);

OAI21x1_ASAP7_75t_L g2035 ( 
.A1(n_1954),
.A2(n_1815),
.B(n_1805),
.Y(n_2035)
);

AOI22xp33_ASAP7_75t_L g2036 ( 
.A1(n_1998),
.A2(n_1912),
.B1(n_1923),
.B2(n_1893),
.Y(n_2036)
);

OAI31xp33_ASAP7_75t_L g2037 ( 
.A1(n_2011),
.A2(n_1849),
.A3(n_1900),
.B(n_1882),
.Y(n_2037)
);

OAI31xp33_ASAP7_75t_L g2038 ( 
.A1(n_1974),
.A2(n_1850),
.A3(n_1773),
.B(n_1904),
.Y(n_2038)
);

NAND2xp33_ASAP7_75t_R g2039 ( 
.A(n_1953),
.B(n_1759),
.Y(n_2039)
);

INVx2_ASAP7_75t_SL g2040 ( 
.A(n_1950),
.Y(n_2040)
);

AO21x1_ASAP7_75t_SL g2041 ( 
.A1(n_2007),
.A2(n_1763),
.B(n_1766),
.Y(n_2041)
);

AOI33xp33_ASAP7_75t_L g2042 ( 
.A1(n_2002),
.A2(n_1903),
.A3(n_1769),
.B1(n_1888),
.B2(n_1917),
.B3(n_1919),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_1932),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1939),
.B(n_1831),
.Y(n_2044)
);

NAND3xp33_ASAP7_75t_L g2045 ( 
.A(n_1987),
.B(n_1827),
.C(n_1846),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1932),
.Y(n_2046)
);

HB1xp67_ASAP7_75t_L g2047 ( 
.A(n_1945),
.Y(n_2047)
);

NAND3xp33_ASAP7_75t_L g2048 ( 
.A(n_2001),
.B(n_1820),
.C(n_1816),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1950),
.B(n_1839),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1961),
.Y(n_2050)
);

INVx4_ASAP7_75t_L g2051 ( 
.A(n_1946),
.Y(n_2051)
);

AOI22xp33_ASAP7_75t_SL g2052 ( 
.A1(n_2010),
.A2(n_1851),
.B1(n_1848),
.B2(n_1785),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1933),
.Y(n_2053)
);

AOI222xp33_ASAP7_75t_L g2054 ( 
.A1(n_1982),
.A2(n_1928),
.B1(n_1918),
.B2(n_1895),
.C1(n_1916),
.C2(n_1915),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2001),
.A2(n_1899),
.B1(n_1906),
.B2(n_1907),
.Y(n_2055)
);

OAI211xp5_ASAP7_75t_L g2056 ( 
.A1(n_2002),
.A2(n_1785),
.B(n_1913),
.C(n_1815),
.Y(n_2056)
);

OAI22xp5_ASAP7_75t_L g2057 ( 
.A1(n_1974),
.A2(n_2010),
.B1(n_1999),
.B2(n_1993),
.Y(n_2057)
);

INVx2_ASAP7_75t_L g2058 ( 
.A(n_1933),
.Y(n_2058)
);

AND2x6_ASAP7_75t_SL g2059 ( 
.A(n_1975),
.B(n_1759),
.Y(n_2059)
);

AO21x2_ASAP7_75t_L g2060 ( 
.A1(n_1976),
.A2(n_1787),
.B(n_1798),
.Y(n_2060)
);

BUFx6f_ASAP7_75t_L g2061 ( 
.A(n_2013),
.Y(n_2061)
);

AOI221xp5_ASAP7_75t_L g2062 ( 
.A1(n_1982),
.A2(n_1772),
.B1(n_1877),
.B2(n_1879),
.C(n_1825),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_1993),
.A2(n_1870),
.B1(n_1760),
.B2(n_1862),
.Y(n_2063)
);

AOI22xp33_ASAP7_75t_SL g2064 ( 
.A1(n_2009),
.A2(n_1775),
.B1(n_1808),
.B2(n_1855),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_1961),
.Y(n_2065)
);

NOR2xp33_ASAP7_75t_R g2066 ( 
.A(n_1946),
.B(n_1811),
.Y(n_2066)
);

OAI211xp5_ASAP7_75t_L g2067 ( 
.A1(n_1999),
.A2(n_1811),
.B(n_1874),
.C(n_1781),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1939),
.B(n_1786),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_1939),
.B(n_1814),
.Y(n_2069)
);

OAI22xp5_ASAP7_75t_L g2070 ( 
.A1(n_1994),
.A2(n_1847),
.B1(n_1856),
.B2(n_1790),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_1949),
.B(n_1843),
.Y(n_2071)
);

AND2x4_ASAP7_75t_L g2072 ( 
.A(n_1931),
.B(n_1795),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_1935),
.Y(n_2073)
);

AOI22xp33_ASAP7_75t_SL g2074 ( 
.A1(n_2009),
.A2(n_1808),
.B1(n_1862),
.B2(n_1784),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_1945),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_1937),
.Y(n_2076)
);

OAI22xp5_ASAP7_75t_L g2077 ( 
.A1(n_1968),
.A2(n_1872),
.B1(n_1861),
.B2(n_1862),
.Y(n_2077)
);

INVx4_ASAP7_75t_L g2078 ( 
.A(n_1946),
.Y(n_2078)
);

INVx2_ASAP7_75t_L g2079 ( 
.A(n_1935),
.Y(n_2079)
);

NAND3xp33_ASAP7_75t_L g2080 ( 
.A(n_1977),
.B(n_1796),
.C(n_1858),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2000),
.B(n_1794),
.Y(n_2081)
);

AOI221xp5_ASAP7_75t_L g2082 ( 
.A1(n_1977),
.A2(n_1860),
.B1(n_1909),
.B2(n_1765),
.C(n_1808),
.Y(n_2082)
);

AOI33xp33_ASAP7_75t_L g2083 ( 
.A1(n_1976),
.A2(n_1768),
.A3(n_1909),
.B1(n_1988),
.B2(n_1989),
.B3(n_2008),
.Y(n_2083)
);

OAI33xp33_ASAP7_75t_L g2084 ( 
.A1(n_1958),
.A2(n_1768),
.A3(n_1956),
.B1(n_1936),
.B2(n_2000),
.B3(n_2005),
.Y(n_2084)
);

OAI211xp5_ASAP7_75t_L g2085 ( 
.A1(n_1976),
.A2(n_1989),
.B(n_1988),
.C(n_2008),
.Y(n_2085)
);

AND2x4_ASAP7_75t_L g2086 ( 
.A(n_1931),
.B(n_2004),
.Y(n_2086)
);

NAND2xp33_ASAP7_75t_SL g2087 ( 
.A(n_1946),
.B(n_1962),
.Y(n_2087)
);

AOI21xp33_ASAP7_75t_L g2088 ( 
.A1(n_1995),
.A2(n_2005),
.B(n_2009),
.Y(n_2088)
);

AOI22xp33_ASAP7_75t_L g2089 ( 
.A1(n_2012),
.A2(n_2008),
.B1(n_2006),
.B2(n_1995),
.Y(n_2089)
);

AOI22xp33_ASAP7_75t_L g2090 ( 
.A1(n_2012),
.A2(n_2006),
.B1(n_1995),
.B2(n_1931),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1937),
.Y(n_2091)
);

AOI222xp33_ASAP7_75t_SL g2092 ( 
.A1(n_1940),
.A2(n_1943),
.B1(n_1951),
.B2(n_1952),
.C1(n_1947),
.C2(n_1941),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_1940),
.Y(n_2093)
);

NAND3xp33_ASAP7_75t_L g2094 ( 
.A(n_1988),
.B(n_1989),
.C(n_1971),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_1956),
.B(n_1967),
.Y(n_2095)
);

NOR2xp33_ASAP7_75t_L g2096 ( 
.A(n_1968),
.B(n_1965),
.Y(n_2096)
);

NAND2xp5_ASAP7_75t_L g2097 ( 
.A(n_1967),
.B(n_1949),
.Y(n_2097)
);

OAI221xp5_ASAP7_75t_L g2098 ( 
.A1(n_1971),
.A2(n_1985),
.B1(n_1981),
.B2(n_1958),
.C(n_1964),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1941),
.Y(n_2099)
);

HB1xp67_ASAP7_75t_L g2100 ( 
.A(n_2047),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_2034),
.B(n_1980),
.Y(n_2101)
);

INVx1_ASAP7_75t_SL g2102 ( 
.A(n_2029),
.Y(n_2102)
);

AND2x4_ASAP7_75t_L g2103 ( 
.A(n_2086),
.B(n_1991),
.Y(n_2103)
);

AND2x4_ASAP7_75t_L g2104 ( 
.A(n_2086),
.B(n_2072),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2014),
.Y(n_2105)
);

AND2x4_ASAP7_75t_L g2106 ( 
.A(n_2086),
.B(n_1991),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_L g2107 ( 
.A(n_2015),
.B(n_1980),
.Y(n_2107)
);

AND2x2_ASAP7_75t_L g2108 ( 
.A(n_2022),
.B(n_1967),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2022),
.B(n_1930),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_L g2110 ( 
.A(n_2083),
.B(n_2040),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2050),
.Y(n_2111)
);

INVx1_ASAP7_75t_L g2112 ( 
.A(n_2065),
.Y(n_2112)
);

AND2x2_ASAP7_75t_L g2113 ( 
.A(n_2068),
.B(n_1930),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2068),
.B(n_1930),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2028),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_2075),
.Y(n_2116)
);

INVx2_ASAP7_75t_L g2117 ( 
.A(n_2024),
.Y(n_2117)
);

AND2x2_ASAP7_75t_L g2118 ( 
.A(n_2083),
.B(n_1934),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2040),
.B(n_2057),
.Y(n_2119)
);

AND2x2_ASAP7_75t_L g2120 ( 
.A(n_2017),
.B(n_1934),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_2076),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_L g2122 ( 
.A(n_2094),
.B(n_1934),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2096),
.B(n_1943),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_2021),
.Y(n_2124)
);

OR2x2_ASAP7_75t_L g2125 ( 
.A(n_2097),
.B(n_1973),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_2091),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2093),
.Y(n_2127)
);

HB1xp67_ASAP7_75t_L g2128 ( 
.A(n_2033),
.Y(n_2128)
);

NAND2xp5_ASAP7_75t_SL g2129 ( 
.A(n_2064),
.B(n_2004),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_2024),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_2096),
.B(n_1944),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2099),
.Y(n_2132)
);

INVx1_ASAP7_75t_L g2133 ( 
.A(n_2043),
.Y(n_2133)
);

AND2x2_ASAP7_75t_L g2134 ( 
.A(n_2017),
.B(n_1942),
.Y(n_2134)
);

BUFx6f_ASAP7_75t_L g2135 ( 
.A(n_2061),
.Y(n_2135)
);

AND2x2_ASAP7_75t_L g2136 ( 
.A(n_2018),
.B(n_1942),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2032),
.B(n_1944),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2046),
.Y(n_2138)
);

HB1xp67_ASAP7_75t_L g2139 ( 
.A(n_2098),
.Y(n_2139)
);

AND2x2_ASAP7_75t_L g2140 ( 
.A(n_2018),
.B(n_1942),
.Y(n_2140)
);

OR2x6_ASAP7_75t_L g2141 ( 
.A(n_2031),
.B(n_1990),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2095),
.B(n_1973),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2081),
.B(n_1947),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2046),
.Y(n_2144)
);

INVx2_ASAP7_75t_L g2145 ( 
.A(n_2053),
.Y(n_2145)
);

INVx1_ASAP7_75t_L g2146 ( 
.A(n_2053),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2058),
.Y(n_2147)
);

AND2x2_ASAP7_75t_L g2148 ( 
.A(n_2085),
.B(n_1948),
.Y(n_2148)
);

INVx2_ASAP7_75t_SL g2149 ( 
.A(n_2061),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2026),
.B(n_1948),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_SL g2151 ( 
.A(n_2066),
.B(n_2004),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2026),
.B(n_1948),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_2069),
.B(n_1951),
.Y(n_2153)
);

AND2x2_ASAP7_75t_L g2154 ( 
.A(n_2044),
.B(n_1966),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_2069),
.B(n_1952),
.Y(n_2155)
);

NAND2x1p5_ASAP7_75t_L g2156 ( 
.A(n_2051),
.B(n_1990),
.Y(n_2156)
);

INVx1_ASAP7_75t_L g2157 ( 
.A(n_2073),
.Y(n_2157)
);

NAND2xp5_ASAP7_75t_L g2158 ( 
.A(n_2044),
.B(n_1970),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_2021),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2049),
.B(n_1966),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2079),
.Y(n_2161)
);

HB1xp67_ASAP7_75t_L g2162 ( 
.A(n_2071),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_2080),
.B(n_1970),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2079),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2060),
.B(n_1970),
.Y(n_2165)
);

HB1xp67_ASAP7_75t_L g2166 ( 
.A(n_2060),
.Y(n_2166)
);

AND2x2_ASAP7_75t_L g2167 ( 
.A(n_2074),
.B(n_1966),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2061),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_2117),
.Y(n_2169)
);

HB1xp67_ASAP7_75t_L g2170 ( 
.A(n_2100),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2117),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2163),
.B(n_1972),
.Y(n_2172)
);

INVx1_ASAP7_75t_L g2173 ( 
.A(n_2111),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2111),
.Y(n_2174)
);

AND2x2_ASAP7_75t_L g2175 ( 
.A(n_2148),
.B(n_2118),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2121),
.Y(n_2176)
);

INVx2_ASAP7_75t_L g2177 ( 
.A(n_2117),
.Y(n_2177)
);

INVxp67_ASAP7_75t_SL g2178 ( 
.A(n_2166),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2143),
.B(n_2020),
.Y(n_2179)
);

INVx1_ASAP7_75t_L g2180 ( 
.A(n_2112),
.Y(n_2180)
);

INVx2_ASAP7_75t_SL g2181 ( 
.A(n_2124),
.Y(n_2181)
);

INVx2_ASAP7_75t_L g2182 ( 
.A(n_2130),
.Y(n_2182)
);

INVx3_ASAP7_75t_R g2183 ( 
.A(n_2103),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_2141),
.B(n_2051),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_2124),
.B(n_2059),
.Y(n_2185)
);

HB1xp67_ASAP7_75t_L g2186 ( 
.A(n_2128),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2112),
.Y(n_2187)
);

AOI22xp5_ASAP7_75t_L g2188 ( 
.A1(n_2139),
.A2(n_2016),
.B1(n_2025),
.B2(n_2030),
.Y(n_2188)
);

AND2x2_ASAP7_75t_L g2189 ( 
.A(n_2148),
.B(n_1978),
.Y(n_2189)
);

AND2x2_ASAP7_75t_L g2190 ( 
.A(n_2118),
.B(n_1960),
.Y(n_2190)
);

OAI322xp33_ASAP7_75t_L g2191 ( 
.A1(n_2163),
.A2(n_2045),
.A3(n_2048),
.B1(n_2023),
.B2(n_2025),
.C1(n_1972),
.C2(n_2055),
.Y(n_2191)
);

NOR2x1p5_ASAP7_75t_L g2192 ( 
.A(n_2124),
.B(n_1960),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_2130),
.Y(n_2193)
);

NAND2x1p5_ASAP7_75t_L g2194 ( 
.A(n_2151),
.B(n_2078),
.Y(n_2194)
);

AND2x2_ASAP7_75t_L g2195 ( 
.A(n_2109),
.B(n_1960),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_2130),
.Y(n_2196)
);

OR2x2_ASAP7_75t_L g2197 ( 
.A(n_2158),
.B(n_1986),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2121),
.Y(n_2198)
);

INVx1_ASAP7_75t_L g2199 ( 
.A(n_2126),
.Y(n_2199)
);

NAND3xp33_ASAP7_75t_L g2200 ( 
.A(n_2110),
.B(n_2037),
.C(n_2038),
.Y(n_2200)
);

NAND2x1_ASAP7_75t_SL g2201 ( 
.A(n_2104),
.B(n_2072),
.Y(n_2201)
);

AND2x2_ASAP7_75t_L g2202 ( 
.A(n_2109),
.B(n_1963),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2143),
.B(n_1959),
.Y(n_2203)
);

OAI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2141),
.A2(n_2052),
.B1(n_2023),
.B2(n_2067),
.Y(n_2204)
);

OR2x2_ASAP7_75t_L g2205 ( 
.A(n_2158),
.B(n_1986),
.Y(n_2205)
);

OR2x2_ASAP7_75t_L g2206 ( 
.A(n_2101),
.B(n_1983),
.Y(n_2206)
);

INVx1_ASAP7_75t_L g2207 ( 
.A(n_2126),
.Y(n_2207)
);

NAND2xp5_ASAP7_75t_L g2208 ( 
.A(n_2137),
.B(n_1959),
.Y(n_2208)
);

NAND2xp5_ASAP7_75t_L g2209 ( 
.A(n_2137),
.B(n_1969),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2120),
.B(n_1963),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2127),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2127),
.Y(n_2212)
);

INVx1_ASAP7_75t_SL g2213 ( 
.A(n_2159),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2132),
.Y(n_2214)
);

INVx1_ASAP7_75t_L g2215 ( 
.A(n_2132),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2105),
.Y(n_2216)
);

AND2x4_ASAP7_75t_L g2217 ( 
.A(n_2141),
.B(n_2078),
.Y(n_2217)
);

NAND2xp5_ASAP7_75t_L g2218 ( 
.A(n_2123),
.B(n_1983),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2123),
.B(n_1984),
.Y(n_2219)
);

INVxp67_ASAP7_75t_SL g2220 ( 
.A(n_2119),
.Y(n_2220)
);

OR2x2_ASAP7_75t_L g2221 ( 
.A(n_2101),
.B(n_1984),
.Y(n_2221)
);

AND2x4_ASAP7_75t_L g2222 ( 
.A(n_2141),
.B(n_2078),
.Y(n_2222)
);

AND2x4_ASAP7_75t_L g2223 ( 
.A(n_2141),
.B(n_1991),
.Y(n_2223)
);

BUFx2_ASAP7_75t_L g2224 ( 
.A(n_2103),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_2169),
.Y(n_2225)
);

AOI21xp33_ASAP7_75t_SL g2226 ( 
.A1(n_2185),
.A2(n_2039),
.B(n_2119),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2220),
.B(n_2113),
.Y(n_2227)
);

OR2x2_ASAP7_75t_L g2228 ( 
.A(n_2172),
.B(n_2153),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2179),
.B(n_2113),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_2173),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2186),
.B(n_2114),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2170),
.B(n_2114),
.Y(n_2232)
);

INVx1_ASAP7_75t_L g2233 ( 
.A(n_2173),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2174),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2174),
.Y(n_2235)
);

NOR3xp33_ASAP7_75t_L g2236 ( 
.A(n_2200),
.B(n_2084),
.C(n_2056),
.Y(n_2236)
);

AND2x2_ASAP7_75t_L g2237 ( 
.A(n_2224),
.B(n_2108),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2180),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_2180),
.Y(n_2239)
);

CKINVDCx16_ASAP7_75t_R g2240 ( 
.A(n_2188),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2187),
.Y(n_2241)
);

OR2x6_ASAP7_75t_L g2242 ( 
.A(n_2181),
.B(n_1990),
.Y(n_2242)
);

INVxp67_ASAP7_75t_L g2243 ( 
.A(n_2181),
.Y(n_2243)
);

INVx3_ASAP7_75t_L g2244 ( 
.A(n_2223),
.Y(n_2244)
);

AND2x2_ASAP7_75t_L g2245 ( 
.A(n_2224),
.B(n_2108),
.Y(n_2245)
);

INVx1_ASAP7_75t_SL g2246 ( 
.A(n_2213),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_SL g2247 ( 
.A(n_2223),
.B(n_2104),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_2172),
.B(n_2153),
.Y(n_2248)
);

AOI22xp33_ASAP7_75t_L g2249 ( 
.A1(n_2204),
.A2(n_2041),
.B1(n_2027),
.B2(n_2062),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_2203),
.B(n_2160),
.Y(n_2250)
);

BUFx2_ASAP7_75t_L g2251 ( 
.A(n_2201),
.Y(n_2251)
);

NAND2xp33_ASAP7_75t_SL g2252 ( 
.A(n_2192),
.B(n_2066),
.Y(n_2252)
);

O2A1O1Ixp33_ASAP7_75t_L g2253 ( 
.A1(n_2191),
.A2(n_2110),
.B(n_2165),
.C(n_2129),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_2175),
.B(n_2160),
.Y(n_2254)
);

INVx2_ASAP7_75t_SL g2255 ( 
.A(n_2201),
.Y(n_2255)
);

OR2x2_ASAP7_75t_L g2256 ( 
.A(n_2197),
.B(n_2155),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2175),
.B(n_2120),
.Y(n_2257)
);

AND2x2_ASAP7_75t_L g2258 ( 
.A(n_2189),
.B(n_2103),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_SL g2259 ( 
.A(n_2223),
.B(n_2104),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_R g2260 ( 
.A(n_2184),
.B(n_2039),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2169),
.Y(n_2261)
);

AND2x2_ASAP7_75t_L g2262 ( 
.A(n_2189),
.B(n_2103),
.Y(n_2262)
);

OR2x2_ASAP7_75t_L g2263 ( 
.A(n_2197),
.B(n_2155),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_2171),
.Y(n_2264)
);

BUFx2_ASAP7_75t_L g2265 ( 
.A(n_2194),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2187),
.Y(n_2266)
);

INVx2_ASAP7_75t_L g2267 ( 
.A(n_2171),
.Y(n_2267)
);

AND2x4_ASAP7_75t_L g2268 ( 
.A(n_2184),
.B(n_2106),
.Y(n_2268)
);

INVx1_ASAP7_75t_L g2269 ( 
.A(n_2198),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_2198),
.Y(n_2270)
);

OR2x2_ASAP7_75t_L g2271 ( 
.A(n_2205),
.B(n_2165),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2190),
.A2(n_2162),
.B1(n_2089),
.B2(n_2070),
.Y(n_2272)
);

AND2x2_ASAP7_75t_L g2273 ( 
.A(n_2190),
.B(n_2106),
.Y(n_2273)
);

NAND2xp5_ASAP7_75t_SL g2274 ( 
.A(n_2184),
.B(n_2104),
.Y(n_2274)
);

NAND2xp5_ASAP7_75t_L g2275 ( 
.A(n_2208),
.B(n_2131),
.Y(n_2275)
);

NOR4xp25_ASAP7_75t_SL g2276 ( 
.A(n_2178),
.B(n_2087),
.C(n_2115),
.D(n_2116),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2209),
.B(n_2131),
.Y(n_2277)
);

AO22x1_ASAP7_75t_L g2278 ( 
.A1(n_2217),
.A2(n_2159),
.B1(n_2222),
.B2(n_2167),
.Y(n_2278)
);

HB1xp67_ASAP7_75t_L g2279 ( 
.A(n_2176),
.Y(n_2279)
);

AND2x2_ASAP7_75t_L g2280 ( 
.A(n_2217),
.B(n_2106),
.Y(n_2280)
);

NAND2xp33_ASAP7_75t_L g2281 ( 
.A(n_2260),
.B(n_2236),
.Y(n_2281)
);

NAND3xp33_ASAP7_75t_L g2282 ( 
.A(n_2253),
.B(n_2042),
.C(n_2092),
.Y(n_2282)
);

NAND2xp5_ASAP7_75t_L g2283 ( 
.A(n_2246),
.B(n_2211),
.Y(n_2283)
);

OAI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2249),
.A2(n_2122),
.B1(n_2194),
.B2(n_2205),
.Y(n_2284)
);

AOI22xp5_ASAP7_75t_L g2285 ( 
.A1(n_2240),
.A2(n_2090),
.B1(n_2019),
.B2(n_2082),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2279),
.Y(n_2286)
);

NAND2xp5_ASAP7_75t_L g2287 ( 
.A(n_2229),
.B(n_2212),
.Y(n_2287)
);

NAND2xp5_ASAP7_75t_L g2288 ( 
.A(n_2243),
.B(n_2216),
.Y(n_2288)
);

AOI22xp33_ASAP7_75t_L g2289 ( 
.A1(n_2272),
.A2(n_2036),
.B1(n_2054),
.B2(n_1929),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2230),
.Y(n_2290)
);

AOI221xp5_ASAP7_75t_L g2291 ( 
.A1(n_2226),
.A2(n_2088),
.B1(n_2122),
.B2(n_2216),
.C(n_2218),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2230),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2233),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_2227),
.B(n_2199),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_2251),
.Y(n_2295)
);

OAI22xp5_ASAP7_75t_L g2296 ( 
.A1(n_2276),
.A2(n_2194),
.B1(n_2167),
.B2(n_2222),
.Y(n_2296)
);

OAI22xp33_ASAP7_75t_L g2297 ( 
.A1(n_2251),
.A2(n_2063),
.B1(n_1985),
.B2(n_1981),
.Y(n_2297)
);

NOR2xp67_ASAP7_75t_L g2298 ( 
.A(n_2255),
.B(n_2217),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_L g2299 ( 
.A(n_2255),
.B(n_2183),
.Y(n_2299)
);

CKINVDCx14_ASAP7_75t_R g2300 ( 
.A(n_2252),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2233),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2257),
.B(n_2199),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2235),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2235),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_2266),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2266),
.Y(n_2306)
);

INVx1_ASAP7_75t_SL g2307 ( 
.A(n_2252),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2265),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_2269),
.Y(n_2309)
);

OAI221xp5_ASAP7_75t_L g2310 ( 
.A1(n_2271),
.A2(n_2221),
.B1(n_2206),
.B2(n_2177),
.C(n_2193),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2269),
.Y(n_2311)
);

NOR2xp33_ASAP7_75t_L g2312 ( 
.A(n_2254),
.B(n_2183),
.Y(n_2312)
);

OR2x2_ASAP7_75t_L g2313 ( 
.A(n_2228),
.B(n_2206),
.Y(n_2313)
);

AOI22xp33_ASAP7_75t_L g2314 ( 
.A1(n_2225),
.A2(n_1929),
.B1(n_1981),
.B2(n_1985),
.Y(n_2314)
);

O2A1O1Ixp5_ASAP7_75t_SL g2315 ( 
.A1(n_2244),
.A2(n_2207),
.B(n_2214),
.C(n_2215),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2234),
.Y(n_2316)
);

INVx2_ASAP7_75t_SL g2317 ( 
.A(n_2268),
.Y(n_2317)
);

OAI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2265),
.A2(n_2042),
.B(n_2222),
.Y(n_2318)
);

AOI21xp5_ASAP7_75t_L g2319 ( 
.A1(n_2278),
.A2(n_2107),
.B(n_2215),
.Y(n_2319)
);

NAND3xp33_ASAP7_75t_L g2320 ( 
.A(n_2278),
.B(n_2214),
.C(n_2207),
.Y(n_2320)
);

NAND2xp33_ASAP7_75t_SL g2321 ( 
.A(n_2237),
.B(n_2195),
.Y(n_2321)
);

INVx1_ASAP7_75t_L g2322 ( 
.A(n_2238),
.Y(n_2322)
);

INVx1_ASAP7_75t_L g2323 ( 
.A(n_2290),
.Y(n_2323)
);

AOI22xp5_ASAP7_75t_L g2324 ( 
.A1(n_2289),
.A2(n_2282),
.B1(n_2281),
.B2(n_2285),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2292),
.Y(n_2325)
);

OR2x2_ASAP7_75t_L g2326 ( 
.A(n_2313),
.B(n_2287),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2293),
.Y(n_2327)
);

O2A1O1Ixp33_ASAP7_75t_SL g2328 ( 
.A1(n_2307),
.A2(n_2274),
.B(n_2247),
.C(n_2259),
.Y(n_2328)
);

INVx1_ASAP7_75t_L g2329 ( 
.A(n_2301),
.Y(n_2329)
);

O2A1O1Ixp33_ASAP7_75t_L g2330 ( 
.A1(n_2318),
.A2(n_2241),
.B(n_2270),
.C(n_2239),
.Y(n_2330)
);

OAI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2289),
.A2(n_2242),
.B1(n_2231),
.B2(n_2244),
.Y(n_2331)
);

AOI221xp5_ASAP7_75t_L g2332 ( 
.A1(n_2291),
.A2(n_2275),
.B1(n_2277),
.B2(n_2261),
.C(n_2225),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2303),
.Y(n_2333)
);

NOR3xp33_ASAP7_75t_L g2334 ( 
.A(n_2295),
.B(n_2244),
.C(n_2271),
.Y(n_2334)
);

NAND2xp5_ASAP7_75t_L g2335 ( 
.A(n_2286),
.B(n_2257),
.Y(n_2335)
);

NAND4xp25_ASAP7_75t_L g2336 ( 
.A(n_2308),
.B(n_2245),
.C(n_2237),
.D(n_2232),
.Y(n_2336)
);

HB1xp67_ASAP7_75t_L g2337 ( 
.A(n_2283),
.Y(n_2337)
);

AOI32xp33_ASAP7_75t_L g2338 ( 
.A1(n_2297),
.A2(n_2245),
.A3(n_2228),
.B1(n_2248),
.B2(n_2258),
.Y(n_2338)
);

AOI221xp5_ASAP7_75t_L g2339 ( 
.A1(n_2314),
.A2(n_2297),
.B1(n_2284),
.B2(n_2310),
.C(n_2320),
.Y(n_2339)
);

OA21x2_ASAP7_75t_L g2340 ( 
.A1(n_2319),
.A2(n_2264),
.B(n_2261),
.Y(n_2340)
);

OAI211xp5_ASAP7_75t_SL g2341 ( 
.A1(n_2300),
.A2(n_2102),
.B(n_2250),
.C(n_2248),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2316),
.B(n_2322),
.Y(n_2342)
);

AOI22xp5_ASAP7_75t_L g2343 ( 
.A1(n_2312),
.A2(n_2267),
.B1(n_2264),
.B2(n_2242),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2288),
.B(n_2256),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2304),
.Y(n_2345)
);

OAI221xp5_ASAP7_75t_L g2346 ( 
.A1(n_2314),
.A2(n_2299),
.B1(n_2296),
.B2(n_2312),
.C(n_2298),
.Y(n_2346)
);

NAND2xp5_ASAP7_75t_L g2347 ( 
.A(n_2302),
.B(n_2256),
.Y(n_2347)
);

INVx1_ASAP7_75t_L g2348 ( 
.A(n_2305),
.Y(n_2348)
);

OAI22xp33_ASAP7_75t_L g2349 ( 
.A1(n_2299),
.A2(n_2242),
.B1(n_2263),
.B2(n_1981),
.Y(n_2349)
);

INVx1_ASAP7_75t_L g2350 ( 
.A(n_2306),
.Y(n_2350)
);

INVxp67_ASAP7_75t_L g2351 ( 
.A(n_2317),
.Y(n_2351)
);

AOI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_2321),
.A2(n_2267),
.B1(n_2242),
.B2(n_2077),
.Y(n_2352)
);

AOI22xp5_ASAP7_75t_L g2353 ( 
.A1(n_2300),
.A2(n_1929),
.B1(n_2193),
.B2(n_2182),
.Y(n_2353)
);

INVx1_ASAP7_75t_SL g2354 ( 
.A(n_2337),
.Y(n_2354)
);

NOR2x1_ASAP7_75t_L g2355 ( 
.A(n_2341),
.B(n_2309),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2351),
.B(n_2280),
.Y(n_2356)
);

INVx1_ASAP7_75t_SL g2357 ( 
.A(n_2326),
.Y(n_2357)
);

NAND2xp5_ASAP7_75t_SL g2358 ( 
.A(n_2338),
.B(n_2268),
.Y(n_2358)
);

NAND2xp5_ASAP7_75t_L g2359 ( 
.A(n_2324),
.B(n_2294),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2334),
.B(n_2315),
.Y(n_2360)
);

NAND2xp33_ASAP7_75t_SL g2361 ( 
.A(n_2342),
.B(n_2311),
.Y(n_2361)
);

INVx2_ASAP7_75t_L g2362 ( 
.A(n_2340),
.Y(n_2362)
);

INVxp67_ASAP7_75t_L g2363 ( 
.A(n_2346),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2344),
.B(n_2263),
.Y(n_2364)
);

NAND2xp33_ASAP7_75t_L g2365 ( 
.A(n_2335),
.B(n_2273),
.Y(n_2365)
);

AND2x2_ASAP7_75t_L g2366 ( 
.A(n_2347),
.B(n_2280),
.Y(n_2366)
);

NAND2xp5_ASAP7_75t_L g2367 ( 
.A(n_2330),
.B(n_2258),
.Y(n_2367)
);

NAND3xp33_ASAP7_75t_L g2368 ( 
.A(n_2339),
.B(n_2268),
.C(n_2262),
.Y(n_2368)
);

NAND2xp5_ASAP7_75t_L g2369 ( 
.A(n_2336),
.B(n_2262),
.Y(n_2369)
);

NOR2xp33_ASAP7_75t_L g2370 ( 
.A(n_2336),
.B(n_2328),
.Y(n_2370)
);

NAND2xp5_ASAP7_75t_L g2371 ( 
.A(n_2323),
.B(n_2273),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_2325),
.B(n_2327),
.Y(n_2372)
);

INVx2_ASAP7_75t_SL g2373 ( 
.A(n_2340),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2329),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2333),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2345),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2348),
.Y(n_2377)
);

AOI31xp33_ASAP7_75t_L g2378 ( 
.A1(n_2370),
.A2(n_2354),
.A3(n_2357),
.B(n_2363),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_2366),
.B(n_2350),
.Y(n_2379)
);

NOR3xp33_ASAP7_75t_L g2380 ( 
.A(n_2360),
.B(n_2331),
.C(n_2332),
.Y(n_2380)
);

AOI21xp5_ASAP7_75t_L g2381 ( 
.A1(n_2361),
.A2(n_2343),
.B(n_2353),
.Y(n_2381)
);

OAI211xp5_ASAP7_75t_L g2382 ( 
.A1(n_2355),
.A2(n_2352),
.B(n_2102),
.C(n_2087),
.Y(n_2382)
);

OAI21xp5_ASAP7_75t_L g2383 ( 
.A1(n_2373),
.A2(n_2349),
.B(n_2195),
.Y(n_2383)
);

OAI221xp5_ASAP7_75t_L g2384 ( 
.A1(n_2373),
.A2(n_2196),
.B1(n_2177),
.B2(n_2182),
.C(n_1985),
.Y(n_2384)
);

AOI22xp5_ASAP7_75t_L g2385 ( 
.A1(n_2362),
.A2(n_1929),
.B1(n_2196),
.B2(n_2135),
.Y(n_2385)
);

NOR2xp33_ASAP7_75t_SL g2386 ( 
.A(n_2356),
.B(n_2156),
.Y(n_2386)
);

NAND2xp5_ASAP7_75t_L g2387 ( 
.A(n_2366),
.B(n_2134),
.Y(n_2387)
);

NOR3xp33_ASAP7_75t_L g2388 ( 
.A(n_2359),
.B(n_2168),
.C(n_2219),
.Y(n_2388)
);

INVxp67_ASAP7_75t_L g2389 ( 
.A(n_2362),
.Y(n_2389)
);

O2A1O1Ixp33_ASAP7_75t_L g2390 ( 
.A1(n_2377),
.A2(n_2221),
.B(n_1954),
.C(n_2107),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_2356),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2361),
.A2(n_1992),
.B1(n_1954),
.B2(n_2115),
.C(n_2116),
.Y(n_2392)
);

NOR4xp25_ASAP7_75t_L g2393 ( 
.A(n_2378),
.B(n_2376),
.C(n_2375),
.D(n_2377),
.Y(n_2393)
);

NOR2xp33_ASAP7_75t_L g2394 ( 
.A(n_2391),
.B(n_2364),
.Y(n_2394)
);

OAI21xp5_ASAP7_75t_L g2395 ( 
.A1(n_2381),
.A2(n_2382),
.B(n_2380),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2379),
.Y(n_2396)
);

AOI22xp5_ASAP7_75t_L g2397 ( 
.A1(n_2389),
.A2(n_2358),
.B1(n_2367),
.B2(n_2368),
.Y(n_2397)
);

AOI221xp5_ASAP7_75t_L g2398 ( 
.A1(n_2389),
.A2(n_2376),
.B1(n_2375),
.B2(n_2374),
.C(n_2372),
.Y(n_2398)
);

NAND2xp5_ASAP7_75t_SL g2399 ( 
.A(n_2386),
.B(n_2369),
.Y(n_2399)
);

AOI211xp5_ASAP7_75t_L g2400 ( 
.A1(n_2383),
.A2(n_2365),
.B(n_2371),
.C(n_2202),
.Y(n_2400)
);

INVxp67_ASAP7_75t_L g2401 ( 
.A(n_2387),
.Y(n_2401)
);

OAI211xp5_ASAP7_75t_SL g2402 ( 
.A1(n_2392),
.A2(n_2365),
.B(n_2105),
.C(n_1954),
.Y(n_2402)
);

AOI222xp33_ASAP7_75t_L g2403 ( 
.A1(n_2384),
.A2(n_1996),
.B1(n_1997),
.B2(n_1992),
.C1(n_1964),
.C2(n_2147),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2388),
.B(n_2202),
.Y(n_2404)
);

NAND4xp25_ASAP7_75t_SL g2405 ( 
.A(n_2390),
.B(n_2210),
.C(n_2140),
.D(n_2136),
.Y(n_2405)
);

NOR2x1_ASAP7_75t_L g2406 ( 
.A(n_2396),
.B(n_2210),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2393),
.B(n_2385),
.Y(n_2407)
);

HB1xp67_ASAP7_75t_SL g2408 ( 
.A(n_2394),
.Y(n_2408)
);

NOR4xp25_ASAP7_75t_L g2409 ( 
.A(n_2395),
.B(n_2134),
.C(n_2152),
.D(n_2150),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2404),
.B(n_2150),
.Y(n_2410)
);

HB1xp67_ASAP7_75t_L g2411 ( 
.A(n_2401),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2398),
.Y(n_2412)
);

INVx3_ASAP7_75t_L g2413 ( 
.A(n_2397),
.Y(n_2413)
);

NAND2xp5_ASAP7_75t_SL g2414 ( 
.A(n_2413),
.B(n_2407),
.Y(n_2414)
);

AND2x4_ASAP7_75t_L g2415 ( 
.A(n_2406),
.B(n_2399),
.Y(n_2415)
);

NOR2x1_ASAP7_75t_L g2416 ( 
.A(n_2413),
.B(n_2412),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2413),
.B(n_2400),
.Y(n_2417)
);

NOR2xp33_ASAP7_75t_L g2418 ( 
.A(n_2408),
.B(n_2405),
.Y(n_2418)
);

AO21x1_ASAP7_75t_L g2419 ( 
.A1(n_2407),
.A2(n_2402),
.B(n_2403),
.Y(n_2419)
);

AND2x2_ASAP7_75t_L g2420 ( 
.A(n_2411),
.B(n_2136),
.Y(n_2420)
);

AOI22xp33_ASAP7_75t_L g2421 ( 
.A1(n_2410),
.A2(n_2135),
.B1(n_2168),
.B2(n_1996),
.Y(n_2421)
);

NAND3xp33_ASAP7_75t_SL g2422 ( 
.A(n_2414),
.B(n_2409),
.C(n_2410),
.Y(n_2422)
);

NAND3xp33_ASAP7_75t_SL g2423 ( 
.A(n_2417),
.B(n_2152),
.C(n_2154),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_2415),
.B(n_2106),
.Y(n_2424)
);

NAND4xp25_ASAP7_75t_L g2425 ( 
.A(n_2418),
.B(n_2140),
.C(n_1963),
.D(n_2003),
.Y(n_2425)
);

OAI221xp5_ASAP7_75t_L g2426 ( 
.A1(n_2416),
.A2(n_2156),
.B1(n_2135),
.B2(n_2149),
.C(n_2154),
.Y(n_2426)
);

NAND3xp33_ASAP7_75t_SL g2427 ( 
.A(n_2419),
.B(n_2156),
.C(n_2142),
.Y(n_2427)
);

NAND3xp33_ASAP7_75t_SL g2428 ( 
.A(n_2426),
.B(n_2420),
.C(n_2421),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2424),
.B(n_2135),
.Y(n_2429)
);

BUFx2_ASAP7_75t_L g2430 ( 
.A(n_2425),
.Y(n_2430)
);

NAND2xp5_ASAP7_75t_L g2431 ( 
.A(n_2427),
.B(n_2135),
.Y(n_2431)
);

HB1xp67_ASAP7_75t_L g2432 ( 
.A(n_2431),
.Y(n_2432)
);

OAI22xp5_ASAP7_75t_L g2433 ( 
.A1(n_2432),
.A2(n_2429),
.B1(n_2430),
.B2(n_2422),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2433),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2433),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2434),
.B(n_2423),
.Y(n_2436)
);

AOI21xp33_ASAP7_75t_SL g2437 ( 
.A1(n_2435),
.A2(n_2428),
.B(n_2142),
.Y(n_2437)
);

AOI22xp33_ASAP7_75t_L g2438 ( 
.A1(n_2436),
.A2(n_2135),
.B1(n_2149),
.B2(n_2138),
.Y(n_2438)
);

AOI222xp33_ASAP7_75t_L g2439 ( 
.A1(n_2437),
.A2(n_2164),
.B1(n_2133),
.B2(n_2144),
.C1(n_2146),
.C2(n_2157),
.Y(n_2439)
);

AOI22xp33_ASAP7_75t_L g2440 ( 
.A1(n_2438),
.A2(n_2138),
.B1(n_2161),
.B2(n_2145),
.Y(n_2440)
);

OAI221xp5_ASAP7_75t_L g2441 ( 
.A1(n_2440),
.A2(n_2439),
.B1(n_2149),
.B2(n_2125),
.C(n_2013),
.Y(n_2441)
);

AOI211xp5_ASAP7_75t_L g2442 ( 
.A1(n_2441),
.A2(n_2125),
.B(n_1990),
.C(n_2035),
.Y(n_2442)
);


endmodule