module fake_jpeg_10520_n_208 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_208);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_208;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx12_ASAP7_75t_R g33 ( 
.A(n_16),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_42),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_34),
.A2(n_32),
.B1(n_28),
.B2(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_16),
.B(n_1),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_38),
.Y(n_47)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_2),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_39),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_27),
.Y(n_41)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_32),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

AND2x2_ASAP7_75t_SL g49 ( 
.A(n_43),
.B(n_17),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_17),
.C(n_32),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_26),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_52),
.B(n_34),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_35),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_55),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_56),
.A2(n_37),
.B1(n_36),
.B2(n_19),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_59),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_61),
.A2(n_21),
.B1(n_28),
.B2(n_20),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_33),
.B(n_22),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_64),
.B(n_25),
.Y(n_65)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_47),
.A2(n_21),
.B(n_26),
.C(n_31),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_68),
.Y(n_95)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_67),
.B(n_77),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_23),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_72),
.B(n_82),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_48),
.A2(n_19),
.B1(n_24),
.B2(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_73),
.B(n_83),
.Y(n_98)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AND2x4_ASAP7_75t_L g78 ( 
.A(n_49),
.B(n_42),
.Y(n_78)
);

MAJx2_ASAP7_75t_L g97 ( 
.A(n_78),
.B(n_57),
.C(n_64),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_66),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_47),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_48),
.A2(n_50),
.B1(n_56),
.B2(n_53),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_50),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_91),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_87),
.B(n_89),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_79),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_78),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_45),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_55),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_101),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g94 ( 
.A1(n_78),
.A2(n_53),
.A3(n_42),
.B1(n_57),
.B2(n_63),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_94),
.A2(n_97),
.B(n_44),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_77),
.B1(n_74),
.B2(n_76),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_99),
.B(n_102),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_81),
.B(n_22),
.Y(n_100)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_100),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_68),
.B(n_46),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_29),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_103),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_75),
.B(n_57),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_30),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_73),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_105),
.B(n_30),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_89),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_107),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_102),
.A2(n_65),
.B1(n_60),
.B2(n_80),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_108),
.A2(n_114),
.B1(n_120),
.B2(n_104),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_67),
.B(n_60),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_111),
.A2(n_112),
.B(n_118),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_20),
.B(n_28),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_117),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_95),
.A2(n_76),
.B1(n_74),
.B2(n_71),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_70),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_71),
.B1(n_24),
.B2(n_29),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_18),
.C(n_25),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_121),
.B(n_88),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_124),
.B(n_125),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_98),
.A2(n_18),
.B1(n_25),
.B2(n_23),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_98),
.B1(n_101),
.B2(n_93),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_127),
.B(n_131),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_109),
.B(n_86),
.Y(n_129)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_124),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_135),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_133),
.A2(n_140),
.B(n_144),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_109),
.B(n_95),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_137),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_85),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_93),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_139),
.Y(n_158)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_125),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_116),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_114),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_123),
.B(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_122),
.C(n_117),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_145),
.B(n_149),
.C(n_152),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_141),
.A2(n_118),
.B(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_130),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_128),
.A2(n_107),
.B1(n_122),
.B2(n_119),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_148),
.A2(n_120),
.B1(n_115),
.B2(n_30),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_119),
.C(n_111),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_127),
.B(n_128),
.C(n_137),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_129),
.B(n_97),
.C(n_99),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_154),
.B(n_155),
.C(n_160),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_141),
.B(n_135),
.C(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_115),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_157),
.B(n_132),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_133),
.B(n_96),
.Y(n_160)
);

AO221x1_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_87),
.B1(n_90),
.B2(n_138),
.C(n_139),
.Y(n_161)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_161),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_162),
.B(n_167),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_163),
.B(n_150),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_136),
.B(n_142),
.C(n_94),
.D(n_131),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_173),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_153),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_159),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_147),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_152),
.A2(n_130),
.B(n_112),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_169),
.A2(n_155),
.B1(n_154),
.B2(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_156),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_170),
.B(n_15),
.Y(n_183)
);

AOI221xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_15),
.B1(n_13),
.B2(n_23),
.C(n_30),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_145),
.B(n_121),
.C(n_126),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_172),
.B(n_149),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_166),
.C(n_164),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_176),
.B(n_183),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_169),
.B(n_172),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_165),
.Y(n_185)
);

AOI31xp67_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_173),
.A3(n_4),
.B(n_6),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_168),
.A2(n_25),
.B1(n_4),
.B2(n_5),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_182),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_187)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_184),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_185),
.B(n_189),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_186),
.B(n_188),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_187),
.A2(n_190),
.B1(n_182),
.B2(n_177),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_180),
.B(n_165),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_181),
.A2(n_166),
.B1(n_6),
.B2(n_7),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_175),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_191),
.B(n_174),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_196),
.A2(n_3),
.B(n_8),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_185),
.C(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_200),
.C(n_201),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_192),
.B(n_187),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g202 ( 
.A1(n_199),
.A2(n_195),
.B1(n_197),
.B2(n_193),
.Y(n_202)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_202),
.A2(n_9),
.A3(n_11),
.B1(n_12),
.B2(n_193),
.C1(n_186),
.C2(n_184),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_9),
.B(n_10),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_11),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_205),
.B(n_206),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_207),
.B(n_203),
.Y(n_208)
);


endmodule