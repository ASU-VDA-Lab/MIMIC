module fake_jpeg_1763_n_150 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_150);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_150;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_21),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_34),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_33),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_51),
.B1(n_40),
.B2(n_43),
.Y(n_64)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_44),
.B(n_32),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_56),
.A2(n_57),
.B1(n_58),
.B2(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_41),
.B(n_1),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_63),
.B(n_64),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_54),
.A2(n_47),
.B1(n_43),
.B2(n_40),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_66),
.A2(n_56),
.B1(n_51),
.B2(n_45),
.Y(n_80)
);

INVx5_ASAP7_75t_SL g68 ( 
.A(n_59),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_47),
.Y(n_74)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_69),
.Y(n_72)
);

CKINVDCx6p67_ASAP7_75t_R g70 ( 
.A(n_56),
.Y(n_70)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_58),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_57),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_77),
.B(n_79),
.Y(n_91)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_68),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_48),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_61),
.B1(n_66),
.B2(n_45),
.Y(n_90)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_60),
.Y(n_82)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_82),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_67),
.B(n_50),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_36),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_62),
.C(n_50),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_84),
.B(n_27),
.C(n_26),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_60),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_86),
.B(n_90),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_81),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_61),
.B1(n_38),
.B2(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_93),
.A2(n_60),
.B1(n_4),
.B2(n_6),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_96),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g96 ( 
.A(n_73),
.B(n_1),
.CI(n_2),
.CON(n_96),
.SN(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_42),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_97),
.B(n_7),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_85),
.A2(n_72),
.B(n_82),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_98),
.A2(n_103),
.B(n_8),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_84),
.B(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_101),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_37),
.Y(n_101)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_86),
.CON(n_103),
.SN(n_103)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_105),
.B(n_10),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_31),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_110),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_3),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_87),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_109),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_88),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_112),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_111),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_114),
.A2(n_118),
.B1(n_123),
.B2(n_125),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_116),
.B(n_119),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_124),
.Y(n_129)
);

INVx1_ASAP7_75t_SL g119 ( 
.A(n_99),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_120),
.B(n_127),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_102),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_100),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_102),
.A2(n_16),
.B(n_25),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_107),
.C(n_106),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_131),
.C(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_103),
.C(n_104),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_123),
.A2(n_105),
.B1(n_104),
.B2(n_109),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_133),
.A2(n_118),
.B1(n_119),
.B2(n_114),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_28),
.C(n_24),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_124),
.B(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_139),
.B(n_140),
.C(n_135),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_129),
.A2(n_130),
.B(n_128),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_141),
.B(n_136),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_144),
.B(n_145),
.C(n_142),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_143),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_146),
.A2(n_145),
.B(n_18),
.Y(n_147)
);

NOR2xp67_ASAP7_75t_SL g148 ( 
.A(n_147),
.B(n_14),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_14),
.B(n_15),
.Y(n_149)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_149),
.B(n_15),
.Y(n_150)
);


endmodule