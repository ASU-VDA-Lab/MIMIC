module fake_jpeg_30554_n_70 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_70);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_70;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_66;

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_1),
.B(n_21),
.Y(n_24)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_17),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_27),
.A2(n_29),
.B1(n_25),
.B2(n_30),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_31),
.B(n_29),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_26),
.B(n_27),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_30),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_28),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

NAND3xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_2),
.C(n_3),
.Y(n_42)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_0),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_4),
.C(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_37),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_39),
.A2(n_42),
.B1(n_31),
.B2(n_34),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_25),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_46),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_43),
.B(n_45),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_3),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_48),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_42),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_49),
.B(n_8),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_50),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_14),
.B(n_15),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_55),
.A2(n_59),
.B1(n_54),
.B2(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_16),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_10),
.C(n_12),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_57),
.B(n_58),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_23),
.B1(n_18),
.B2(n_19),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_61),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_65),
.B(n_57),
.C(n_59),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_66),
.B(n_63),
.C(n_62),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_67),
.B1(n_60),
.B2(n_55),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_69),
.A2(n_51),
.B(n_20),
.Y(n_70)
);


endmodule