module fake_jpeg_19287_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_7),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_SL g10 ( 
.A(n_7),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

BUFx12_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_0),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_1),
.B(n_5),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_0),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_10),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_10),
.B(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_19),
.B(n_20),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_1),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_21),
.Y(n_25)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_27),
.B(n_20),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_32),
.Y(n_37)
);

A2O1A1O1Ixp25_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_26),
.B(n_23),
.C(n_19),
.D(n_12),
.Y(n_30)
);

NOR2xp67_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_35),
.B1(n_31),
.B2(n_33),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_2),
.B(n_3),
.Y(n_35)
);

XNOR2x1_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_12),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.C(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_14),
.B1(n_11),
.B2(n_9),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_22),
.B1(n_16),
.B2(n_12),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_40),
.A2(n_12),
.B1(n_8),
.B2(n_15),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_16),
.C(n_9),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_42),
.B(n_43),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_11),
.B(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_44),
.B(n_38),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_37),
.C(n_41),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_37),
.C(n_43),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_48),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g52 ( 
.A(n_50),
.B(n_40),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_46),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.C(n_9),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_2),
.B(n_3),
.Y(n_54)
);

O2A1O1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_54),
.A2(n_11),
.B(n_14),
.C(n_29),
.Y(n_55)
);


endmodule