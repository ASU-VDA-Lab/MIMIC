module fake_netlist_6_4711_n_1151 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_212, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_218, n_70, n_120, n_214, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1151);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_212;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_214;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1151;

wire n_992;
wire n_591;
wire n_435;
wire n_1115;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_1030;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_1008;
wire n_1027;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_1079;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_1033;
wire n_316;
wire n_419;
wire n_304;
wire n_700;
wire n_694;
wire n_1103;
wire n_933;
wire n_740;
wire n_1038;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_1061;
wire n_384;
wire n_297;
wire n_627;
wire n_595;
wire n_524;
wire n_342;
wire n_820;
wire n_1044;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_1072;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_1065;
wire n_815;
wire n_350;
wire n_1100;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_1128;
wire n_382;
wire n_673;
wire n_1020;
wire n_1009;
wire n_1042;
wire n_1071;
wire n_628;
wire n_1067;
wire n_883;
wire n_557;
wire n_823;
wire n_1132;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_1074;
wire n_898;
wire n_1032;
wire n_845;
wire n_255;
wire n_807;
wire n_1036;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_1138;
wire n_893;
wire n_925;
wire n_485;
wire n_1099;
wire n_1026;
wire n_443;
wire n_1101;
wire n_246;
wire n_892;
wire n_768;
wire n_1097;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_1130;
wire n_1127;
wire n_238;
wire n_1095;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_1120;
wire n_369;
wire n_894;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_1024;
wire n_669;
wire n_447;
wire n_872;
wire n_1139;
wire n_300;
wire n_222;
wire n_718;
wire n_248;
wire n_517;
wire n_1018;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_1105;
wire n_621;
wire n_305;
wire n_1037;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_1078;
wire n_504;
wire n_1140;
wire n_314;
wire n_923;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_1015;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1057;
wire n_1147;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_1005;
wire n_991;
wire n_957;
wire n_235;
wire n_1143;
wire n_536;
wire n_895;
wire n_1126;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_1108;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_1119;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_1116;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_989;
wire n_843;
wire n_797;
wire n_666;
wire n_1016;
wire n_371;
wire n_795;
wire n_770;
wire n_940;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_538;
wire n_1035;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_953;
wire n_448;
wire n_886;
wire n_1017;
wire n_844;
wire n_1004;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_1022;
wire n_1083;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_1112;
wire n_454;
wire n_638;
wire n_234;
wire n_910;
wire n_901;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_1117;
wire n_1087;
wire n_752;
wire n_908;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_1049;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_1043;
wire n_1011;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_1088;
wire n_708;
wire n_919;
wire n_1081;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_1084;
wire n_1104;
wire n_907;
wire n_854;
wire n_1058;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_1122;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_1109;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_1148;
wire n_293;
wire n_1054;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_1070;
wire n_1085;
wire n_232;
wire n_650;
wire n_998;
wire n_1046;
wire n_717;
wire n_1145;
wire n_330;
wire n_771;
wire n_1121;
wire n_470;
wire n_475;
wire n_924;
wire n_1102;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_551;
wire n_258;
wire n_699;
wire n_456;
wire n_1149;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1073;
wire n_1000;
wire n_279;
wire n_686;
wire n_1041;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_594;
wire n_565;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_1062;
wire n_619;
wire n_885;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_1090;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_1142;
wire n_503;
wire n_716;
wire n_623;
wire n_1048;
wire n_1123;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_934;
wire n_482;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_1137;
wire n_433;
wire n_500;
wire n_942;
wire n_792;
wire n_880;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_1144;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_1068;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_1075;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_959;
wire n_879;
wire n_237;
wire n_584;
wire n_1110;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_707;
wire n_322;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_1133;
wire n_635;
wire n_787;
wire n_311;
wire n_1064;
wire n_403;
wire n_1080;
wire n_723;
wire n_253;
wire n_634;
wire n_1051;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_1141;
wire n_1146;
wire n_386;
wire n_249;
wire n_764;
wire n_1039;
wire n_556;
wire n_1034;
wire n_1086;
wire n_1066;
wire n_692;
wire n_733;
wire n_754;
wire n_1136;
wire n_941;
wire n_975;
wire n_1031;
wire n_487;
wire n_550;
wire n_241;
wire n_1125;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_1107;
wire n_560;
wire n_1014;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_1092;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_1060;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_1111;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_1053;
wire n_530;
wire n_277;
wire n_520;
wire n_1029;
wire n_418;
wire n_1093;
wire n_618;
wire n_1055;
wire n_790;
wire n_1106;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_518;
wire n_299;
wire n_679;
wire n_1069;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_1047;
wire n_1010;
wire n_355;
wire n_426;
wire n_317;
wire n_1040;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_1131;
wire n_1052;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_1006;
wire n_373;
wire n_1012;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_1089;
wire n_1135;
wire n_401;
wire n_324;
wire n_743;
wire n_816;
wire n_766;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_1019;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_1096;
wire n_1063;
wire n_729;
wire n_1091;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_438;
wire n_267;
wire n_1124;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_1059;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_1077;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_1082;
wire n_259;
wire n_1113;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_457;
wire n_391;
wire n_1098;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_1050;
wire n_379;
wire n_778;
wire n_1025;
wire n_1134;
wire n_332;
wire n_891;
wire n_336;
wire n_1150;
wire n_398;
wire n_410;
wire n_1129;
wire n_566;
wire n_554;
wire n_602;
wire n_1013;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_664;
wire n_949;
wire n_678;
wire n_1007;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g219 ( 
.A(n_207),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_194),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_16),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_31),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_29),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_73),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_69),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_47),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_103),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_82),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_67),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_38),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_61),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_63),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_129),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_18),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_6),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_20),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_198),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_27),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g244 ( 
.A(n_14),
.Y(n_244)
);

BUFx10_ASAP7_75t_L g245 ( 
.A(n_164),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_109),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_125),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_28),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_209),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_159),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_65),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_169),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_153),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_218),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_130),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_4),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_160),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_88),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_77),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_131),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_208),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_202),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_182),
.Y(n_264)
);

INVx2_ASAP7_75t_SL g265 ( 
.A(n_119),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_200),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_186),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_81),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_13),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_143),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_148),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_18),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_8),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_2),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_157),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_94),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_14),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_16),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_9),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_80),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_46),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_28),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_135),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_215),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_189),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_146),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_6),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_102),
.Y(n_290)
);

INVx2_ASAP7_75t_SL g291 ( 
.A(n_176),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_118),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_154),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_244),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_284),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_240),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_279),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_220),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_280),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_268),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_245),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_219),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_268),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g305 ( 
.A(n_222),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_221),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_234),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_283),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_259),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_223),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

INVxp33_ASAP7_75t_SL g313 ( 
.A(n_236),
.Y(n_313)
);

OR2x2_ASAP7_75t_L g314 ( 
.A(n_289),
.B(n_237),
.Y(n_314)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_239),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_283),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_269),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_226),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_271),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_272),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

INVx4_ASAP7_75t_R g322 ( 
.A(n_291),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_224),
.Y(n_323)
);

BUFx3_ASAP7_75t_L g324 ( 
.A(n_245),
.Y(n_324)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_250),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_226),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_266),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_225),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_226),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_291),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_292),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_229),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_238),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_229),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_229),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_229),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_227),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_248),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_257),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_228),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_245),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_304),
.Y(n_345)
);

OA21x2_ASAP7_75t_L g346 ( 
.A1(n_318),
.A2(n_329),
.B(n_327),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_333),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

INVx6_ASAP7_75t_L g349 ( 
.A(n_326),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g350 ( 
.A(n_326),
.Y(n_350)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_314),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_301),
.Y(n_352)
);

OA21x2_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_336),
.B(n_334),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_343),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_326),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_330),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_330),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_330),
.Y(n_359)
);

AND2x4_ASAP7_75t_L g360 ( 
.A(n_331),
.B(n_265),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_304),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_337),
.Y(n_363)
);

NOR2x1_ASAP7_75t_L g364 ( 
.A(n_302),
.B(n_260),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_338),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_295),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_295),
.Y(n_367)
);

AND2x4_ASAP7_75t_L g368 ( 
.A(n_306),
.B(n_247),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_310),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_312),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_344),
.B(n_270),
.Y(n_373)
);

BUFx2_ASAP7_75t_L g374 ( 
.A(n_305),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_305),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_320),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_230),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_311),
.B(n_293),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_297),
.Y(n_382)
);

INVx5_ASAP7_75t_L g383 ( 
.A(n_302),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_298),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

BUFx3_ASAP7_75t_L g386 ( 
.A(n_344),
.Y(n_386)
);

BUFx3_ASAP7_75t_L g387 ( 
.A(n_344),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_296),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_324),
.Y(n_390)
);

INVx6_ASAP7_75t_L g391 ( 
.A(n_344),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_296),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_308),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_344),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_341),
.B(n_30),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_332),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_324),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_323),
.Y(n_400)
);

INVx2_ASAP7_75t_SL g401 ( 
.A(n_328),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_340),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_357),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_354),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_388),
.B(n_335),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_354),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_393),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_393),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_400),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_370),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_371),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_400),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_315),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_352),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_R g415 ( 
.A(n_399),
.B(n_316),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_401),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_345),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_R g418 ( 
.A(n_399),
.B(n_231),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_372),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_401),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_345),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_362),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_R g423 ( 
.A(n_351),
.B(n_232),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_382),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_362),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_382),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_355),
.Y(n_428)
);

INVx3_ASAP7_75t_L g429 ( 
.A(n_348),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_389),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_374),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_402),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_402),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_388),
.B(n_313),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_379),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_388),
.B(n_233),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_384),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_355),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_381),
.Y(n_439)
);

INVx3_ASAP7_75t_L g440 ( 
.A(n_348),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_374),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_390),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_398),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_384),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_398),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_398),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_398),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_348),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_376),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_369),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_398),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_388),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_355),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_R g454 ( 
.A(n_392),
.B(n_235),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_358),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_388),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_389),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_397),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_369),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_397),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_383),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_377),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_377),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_358),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_377),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_373),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_383),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_383),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g469 ( 
.A(n_364),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_383),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_353),
.Y(n_471)
);

AND2x6_ASAP7_75t_L g472 ( 
.A(n_394),
.B(n_32),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_377),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_383),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_359),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_368),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_435),
.B(n_386),
.Y(n_478)
);

AOI22xp33_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_396),
.B1(n_386),
.B2(n_395),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_439),
.B(n_387),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_471),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_413),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_432),
.B(n_315),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_457),
.Y(n_484)
);

INVx5_ASAP7_75t_L g485 ( 
.A(n_472),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_368),
.Y(n_486)
);

OAI21xp33_ASAP7_75t_SL g487 ( 
.A1(n_471),
.A2(n_394),
.B(n_325),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_430),
.Y(n_488)
);

OR2x6_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_360),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_433),
.B(n_368),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_459),
.B(n_385),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_452),
.B(n_387),
.Y(n_492)
);

AND2x4_ASAP7_75t_L g493 ( 
.A(n_424),
.B(n_385),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_SL g494 ( 
.A(n_416),
.B(n_396),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_458),
.B(n_395),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_325),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_426),
.Y(n_497)
);

AND2x6_ASAP7_75t_L g498 ( 
.A(n_434),
.B(n_360),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_294),
.Y(n_499)
);

INVx6_ASAP7_75t_L g500 ( 
.A(n_427),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_444),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_420),
.B(n_391),
.Y(n_503)
);

AND2x2_ASAP7_75t_SL g504 ( 
.A(n_405),
.B(n_360),
.Y(n_504)
);

INVx1_ASAP7_75t_SL g505 ( 
.A(n_431),
.Y(n_505)
);

BUFx6f_ASAP7_75t_L g506 ( 
.A(n_472),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_423),
.B(n_375),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_456),
.B(n_443),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_403),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_410),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_455),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_472),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_396),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_419),
.B(n_396),
.Y(n_514)
);

BUFx10_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_464),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_406),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_445),
.B(n_375),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_475),
.Y(n_519)
);

AOI22xp33_ASAP7_75t_L g520 ( 
.A1(n_472),
.A2(n_396),
.B1(n_346),
.B2(n_391),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_428),
.Y(n_521)
);

INVx6_ASAP7_75t_L g522 ( 
.A(n_427),
.Y(n_522)
);

INVx2_ASAP7_75t_SL g523 ( 
.A(n_442),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_438),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_453),
.Y(n_525)
);

AND2x2_ASAP7_75t_SL g526 ( 
.A(n_415),
.B(n_378),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_476),
.B(n_391),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_462),
.Y(n_528)
);

INVx4_ASAP7_75t_L g529 ( 
.A(n_446),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_466),
.B(n_391),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_429),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_447),
.B(n_378),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_463),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_451),
.B(n_380),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_465),
.B(n_473),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_436),
.B(n_273),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_472),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_429),
.Y(n_538)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_441),
.Y(n_539)
);

INVx3_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_477),
.B(n_396),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_440),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_436),
.B(n_274),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_448),
.B(n_346),
.Y(n_544)
);

BUFx6f_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

AND2x6_ASAP7_75t_L g546 ( 
.A(n_448),
.B(n_380),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_423),
.B(n_241),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_409),
.B(n_347),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_427),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_418),
.B(n_242),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_454),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_412),
.B(n_347),
.Y(n_552)
);

NAND2x1p5_ASAP7_75t_L g553 ( 
.A(n_418),
.B(n_346),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_474),
.B(n_346),
.Y(n_554)
);

INVx1_ASAP7_75t_SL g555 ( 
.A(n_417),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_407),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_422),
.B(n_275),
.Y(n_557)
);

AND2x6_ASAP7_75t_L g558 ( 
.A(n_415),
.B(n_359),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_449),
.B(n_366),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_461),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_504),
.A2(n_414),
.B1(n_468),
.B2(n_467),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_523),
.B(n_421),
.Y(n_563)
);

AND2x4_ASAP7_75t_L g564 ( 
.A(n_518),
.B(n_425),
.Y(n_564)
);

AO22x2_ASAP7_75t_L g565 ( 
.A1(n_555),
.A2(n_408),
.B1(n_1),
.B2(n_2),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_481),
.Y(n_566)
);

NAND2x1p5_ASAP7_75t_L g567 ( 
.A(n_529),
.B(n_366),
.Y(n_567)
);

AO22x2_ASAP7_75t_L g568 ( 
.A1(n_505),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g569 ( 
.A(n_483),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_484),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_518),
.B(n_470),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_499),
.B(n_281),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_503),
.B(n_353),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_532),
.B(n_534),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_491),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_497),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_536),
.A2(n_353),
.B1(n_365),
.B2(n_363),
.Y(n_579)
);

INVxp67_ASAP7_75t_L g580 ( 
.A(n_496),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_538),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_532),
.B(n_367),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_534),
.B(n_367),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_545),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_498),
.A2(n_277),
.B1(n_249),
.B2(n_251),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_478),
.B(n_246),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_498),
.A2(n_285),
.B1(n_253),
.B2(n_254),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_480),
.B(n_252),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_507),
.B(n_353),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_527),
.B(n_363),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_493),
.Y(n_591)
);

OAI221xp5_ASAP7_75t_L g592 ( 
.A1(n_543),
.A2(n_482),
.B1(n_501),
.B2(n_502),
.C(n_510),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_542),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_493),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g595 ( 
.A(n_556),
.Y(n_595)
);

INVxp67_ASAP7_75t_L g596 ( 
.A(n_560),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_535),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_511),
.Y(n_599)
);

INVxp67_ASAP7_75t_L g600 ( 
.A(n_548),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_526),
.B(n_365),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_517),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_516),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_486),
.B(n_33),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_519),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_551),
.B(n_255),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_521),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_533),
.Y(n_609)
);

AO22x2_ASAP7_75t_L g610 ( 
.A1(n_557),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_531),
.Y(n_611)
);

AO22x2_ASAP7_75t_L g612 ( 
.A1(n_488),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_486),
.B(n_34),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_524),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_545),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_525),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_540),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_549),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_552),
.B(n_256),
.Y(n_619)
);

NOR2x1_ASAP7_75t_L g620 ( 
.A(n_529),
.B(n_361),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_544),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_508),
.B(n_258),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_559),
.B(n_261),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_492),
.B(n_263),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_SL g625 ( 
.A(n_530),
.B(n_267),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_500),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_546),
.Y(n_627)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_539),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_546),
.Y(n_629)
);

AND2x2_ASAP7_75t_L g630 ( 
.A(n_552),
.B(n_276),
.Y(n_630)
);

O2A1O1Ixp33_ASAP7_75t_L g631 ( 
.A1(n_573),
.A2(n_490),
.B(n_495),
.C(n_547),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_577),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_564),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_584),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_575),
.A2(n_600),
.B1(n_569),
.B2(n_607),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_579),
.A2(n_520),
.B(n_479),
.Y(n_636)
);

AOI21xp5_ASAP7_75t_L g637 ( 
.A1(n_574),
.A2(n_494),
.B(n_485),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_575),
.B(n_515),
.Y(n_638)
);

NOR2xp67_ASAP7_75t_L g639 ( 
.A(n_592),
.B(n_487),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_580),
.A2(n_550),
.B(n_489),
.C(n_561),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_597),
.B(n_621),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_598),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g643 ( 
.A(n_596),
.B(n_515),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_564),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_597),
.B(n_498),
.Y(n_645)
);

NOR3xp33_ASAP7_75t_L g646 ( 
.A(n_628),
.B(n_541),
.C(n_554),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_601),
.B(n_558),
.Y(n_647)
);

AOI21x1_ASAP7_75t_L g648 ( 
.A1(n_589),
.A2(n_489),
.B(n_553),
.Y(n_648)
);

OAI321xp33_ASAP7_75t_L g649 ( 
.A1(n_623),
.A2(n_537),
.A3(n_512),
.B1(n_506),
.B2(n_558),
.C(n_11),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_566),
.A2(n_514),
.B(n_513),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_622),
.B(n_558),
.Y(n_651)
);

OAI21xp5_ASAP7_75t_L g652 ( 
.A1(n_566),
.A2(n_514),
.B(n_513),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_606),
.Y(n_653)
);

AOI22xp5_ASAP7_75t_L g654 ( 
.A1(n_604),
.A2(n_514),
.B1(n_513),
.B2(n_537),
.Y(n_654)
);

AOI21xp5_ASAP7_75t_L g655 ( 
.A1(n_590),
.A2(n_485),
.B(n_545),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_602),
.B(n_506),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_624),
.A2(n_485),
.B(n_506),
.Y(n_657)
);

AOI21xp5_ASAP7_75t_L g658 ( 
.A1(n_570),
.A2(n_537),
.B(n_512),
.Y(n_658)
);

AND2x2_ASAP7_75t_SL g659 ( 
.A(n_604),
.B(n_613),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_609),
.A2(n_512),
.B1(n_500),
.B2(n_522),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_593),
.Y(n_661)
);

OAI22x1_ASAP7_75t_L g662 ( 
.A1(n_562),
.A2(n_282),
.B1(n_286),
.B2(n_287),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_582),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_582),
.B(n_288),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_583),
.B(n_546),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_627),
.A2(n_522),
.B(n_36),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_583),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_591),
.A2(n_290),
.B1(n_349),
.B2(n_350),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_584),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g670 ( 
.A1(n_611),
.A2(n_349),
.B(n_37),
.Y(n_670)
);

INVx11_ASAP7_75t_L g671 ( 
.A(n_595),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_627),
.A2(n_39),
.B(n_35),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_619),
.B(n_5),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_571),
.B(n_40),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_603),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_SL g676 ( 
.A1(n_629),
.A2(n_113),
.B(n_217),
.C(n_216),
.Y(n_676)
);

NOR2x1_ASAP7_75t_L g677 ( 
.A(n_563),
.B(n_348),
.Y(n_677)
);

AOI21xp5_ASAP7_75t_L g678 ( 
.A1(n_586),
.A2(n_356),
.B(n_350),
.Y(n_678)
);

O2A1O1Ixp5_ASAP7_75t_L g679 ( 
.A1(n_588),
.A2(n_625),
.B(n_629),
.C(n_618),
.Y(n_679)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_611),
.A2(n_349),
.B(n_42),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_605),
.A2(n_349),
.B(n_43),
.Y(n_681)
);

AOI21xp33_ASAP7_75t_L g682 ( 
.A1(n_594),
.A2(n_7),
.B(n_9),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_613),
.B(n_350),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_614),
.A2(n_44),
.B(n_41),
.Y(n_684)
);

NAND2xp33_ASAP7_75t_L g685 ( 
.A(n_584),
.B(n_350),
.Y(n_685)
);

A2O1A1Ixp33_ASAP7_75t_L g686 ( 
.A1(n_576),
.A2(n_361),
.B(n_356),
.C(n_350),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_578),
.B(n_10),
.Y(n_687)
);

AOI21xp5_ASAP7_75t_L g688 ( 
.A1(n_572),
.A2(n_615),
.B(n_581),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_615),
.Y(n_689)
);

AND2x6_ASAP7_75t_L g690 ( 
.A(n_620),
.B(n_356),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_616),
.Y(n_691)
);

INVx5_ASAP7_75t_L g692 ( 
.A(n_615),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_671),
.Y(n_693)
);

INVx5_ASAP7_75t_L g694 ( 
.A(n_634),
.Y(n_694)
);

NAND2x1_ASAP7_75t_SL g695 ( 
.A(n_656),
.B(n_630),
.Y(n_695)
);

AOI222xp33_ASAP7_75t_L g696 ( 
.A1(n_673),
.A2(n_565),
.B1(n_568),
.B2(n_610),
.C1(n_612),
.C2(n_641),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_692),
.B(n_581),
.Y(n_697)
);

AOI21xp5_ASAP7_75t_L g698 ( 
.A1(n_636),
.A2(n_637),
.B(n_651),
.Y(n_698)
);

O2A1O1Ixp5_ASAP7_75t_L g699 ( 
.A1(n_681),
.A2(n_617),
.B(n_626),
.C(n_608),
.Y(n_699)
);

INVx2_ASAP7_75t_SL g700 ( 
.A(n_633),
.Y(n_700)
);

O2A1O1Ixp5_ASAP7_75t_L g701 ( 
.A1(n_670),
.A2(n_599),
.B(n_585),
.C(n_587),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_663),
.B(n_563),
.Y(n_702)
);

O2A1O1Ixp33_ASAP7_75t_L g703 ( 
.A1(n_631),
.A2(n_567),
.B(n_610),
.C(n_565),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_R g704 ( 
.A(n_659),
.B(n_45),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_634),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_661),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_634),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_646),
.B(n_612),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_657),
.A2(n_361),
.B(n_356),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_642),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_635),
.B(n_10),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_647),
.B(n_568),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_653),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_643),
.B(n_356),
.Y(n_715)
);

AOI21xp5_ASAP7_75t_L g716 ( 
.A1(n_645),
.A2(n_361),
.B(n_49),
.Y(n_716)
);

BUFx3_ASAP7_75t_L g717 ( 
.A(n_644),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_654),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_R g719 ( 
.A(n_692),
.B(n_48),
.Y(n_719)
);

INVxp67_ASAP7_75t_SL g720 ( 
.A(n_675),
.Y(n_720)
);

AOI21xp5_ASAP7_75t_L g721 ( 
.A1(n_655),
.A2(n_361),
.B(n_51),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_667),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_640),
.A2(n_12),
.B(n_15),
.C(n_17),
.Y(n_723)
);

INVx2_ASAP7_75t_SL g724 ( 
.A(n_638),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_691),
.Y(n_725)
);

A2O1A1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_684),
.A2(n_15),
.B(n_17),
.C(n_19),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_687),
.Y(n_727)
);

AOI21xp5_ASAP7_75t_L g728 ( 
.A1(n_650),
.A2(n_652),
.B(n_639),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_664),
.B(n_19),
.Y(n_729)
);

AOI21xp5_ASAP7_75t_L g730 ( 
.A1(n_639),
.A2(n_121),
.B(n_213),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_669),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_683),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_665),
.B(n_21),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_669),
.Y(n_734)
);

BUFx2_ASAP7_75t_L g735 ( 
.A(n_689),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_662),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_689),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_649),
.B(n_23),
.Y(n_738)
);

O2A1O1Ixp5_ASAP7_75t_L g739 ( 
.A1(n_680),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_739)
);

BUFx2_ASAP7_75t_SL g740 ( 
.A(n_692),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_660),
.Y(n_741)
);

OAI21x1_ASAP7_75t_L g742 ( 
.A1(n_666),
.A2(n_124),
.B(n_212),
.Y(n_742)
);

O2A1O1Ixp5_ASAP7_75t_SL g743 ( 
.A1(n_682),
.A2(n_25),
.B(n_26),
.C(n_27),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_677),
.B(n_50),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_672),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_648),
.Y(n_746)
);

O2A1O1Ixp33_ASAP7_75t_L g747 ( 
.A1(n_679),
.A2(n_676),
.B(n_686),
.C(n_688),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_685),
.A2(n_52),
.B(n_53),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_658),
.B(n_214),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_668),
.B(n_54),
.Y(n_750)
);

OAI21x1_ASAP7_75t_L g751 ( 
.A1(n_678),
.A2(n_55),
.B(n_56),
.Y(n_751)
);

AOI21xp5_ASAP7_75t_L g752 ( 
.A1(n_674),
.A2(n_57),
.B(n_58),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_690),
.A2(n_59),
.B1(n_60),
.B2(n_62),
.Y(n_753)
);

BUFx3_ASAP7_75t_L g754 ( 
.A(n_717),
.Y(n_754)
);

INVx3_ASAP7_75t_L g755 ( 
.A(n_697),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_710),
.Y(n_756)
);

INVx5_ASAP7_75t_L g757 ( 
.A(n_694),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_714),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_694),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_694),
.Y(n_760)
);

INVx1_ASAP7_75t_SL g761 ( 
.A(n_702),
.Y(n_761)
);

BUFx3_ASAP7_75t_L g762 ( 
.A(n_693),
.Y(n_762)
);

NAND2x1p5_ASAP7_75t_L g763 ( 
.A(n_724),
.B(n_690),
.Y(n_763)
);

INVx1_ASAP7_75t_SL g764 ( 
.A(n_735),
.Y(n_764)
);

INVx3_ASAP7_75t_SL g765 ( 
.A(n_700),
.Y(n_765)
);

INVx1_ASAP7_75t_SL g766 ( 
.A(n_695),
.Y(n_766)
);

INVx4_ASAP7_75t_L g767 ( 
.A(n_705),
.Y(n_767)
);

BUFx6f_ASAP7_75t_L g768 ( 
.A(n_705),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_712),
.B(n_64),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_725),
.Y(n_770)
);

INVx1_ASAP7_75t_SL g771 ( 
.A(n_740),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_713),
.B(n_66),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_711),
.Y(n_773)
);

BUFx3_ASAP7_75t_L g774 ( 
.A(n_707),
.Y(n_774)
);

BUFx12f_ASAP7_75t_L g775 ( 
.A(n_697),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_707),
.Y(n_776)
);

BUFx3_ASAP7_75t_L g777 ( 
.A(n_734),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_706),
.Y(n_778)
);

BUFx6f_ASAP7_75t_L g779 ( 
.A(n_737),
.Y(n_779)
);

AND2x4_ASAP7_75t_L g780 ( 
.A(n_722),
.B(n_690),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_720),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_727),
.B(n_690),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_731),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_719),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

BUFx5_ASAP7_75t_L g786 ( 
.A(n_745),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_708),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_708),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_699),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_728),
.B(n_70),
.Y(n_790)
);

INVx5_ASAP7_75t_L g791 ( 
.A(n_746),
.Y(n_791)
);

INVx1_ASAP7_75t_SL g792 ( 
.A(n_704),
.Y(n_792)
);

BUFx2_ASAP7_75t_L g793 ( 
.A(n_741),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_733),
.Y(n_794)
);

INVxp67_ASAP7_75t_SL g795 ( 
.A(n_747),
.Y(n_795)
);

INVx4_ASAP7_75t_L g796 ( 
.A(n_746),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_729),
.Y(n_797)
);

NAND2x1p5_ASAP7_75t_L g798 ( 
.A(n_715),
.B(n_71),
.Y(n_798)
);

AND2x4_ASAP7_75t_L g799 ( 
.A(n_723),
.B(n_72),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_703),
.B(n_211),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_746),
.Y(n_801)
);

INVx5_ASAP7_75t_L g802 ( 
.A(n_753),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_698),
.B(n_74),
.Y(n_803)
);

INVxp67_ASAP7_75t_SL g804 ( 
.A(n_742),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_751),
.Y(n_805)
);

BUFx2_ASAP7_75t_SL g806 ( 
.A(n_753),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_744),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_718),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_739),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_749),
.Y(n_810)
);

NAND2x1p5_ASAP7_75t_L g811 ( 
.A(n_730),
.B(n_75),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_701),
.Y(n_812)
);

INVx5_ASAP7_75t_L g813 ( 
.A(n_718),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_732),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_736),
.B(n_76),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_721),
.B(n_78),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_732),
.Y(n_817)
);

BUFx6f_ASAP7_75t_SL g818 ( 
.A(n_743),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_738),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_696),
.B(n_79),
.Y(n_820)
);

INVx5_ASAP7_75t_L g821 ( 
.A(n_726),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_750),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_696),
.Y(n_823)
);

NAND2x1p5_ASAP7_75t_L g824 ( 
.A(n_757),
.B(n_752),
.Y(n_824)
);

OAI21x1_ASAP7_75t_L g825 ( 
.A1(n_803),
.A2(n_709),
.B(n_716),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_773),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_781),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_787),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_785),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_793),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_819),
.B(n_752),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_822),
.A2(n_748),
.B(n_84),
.Y(n_832)
);

OAI21x1_ASAP7_75t_L g833 ( 
.A1(n_803),
.A2(n_83),
.B(n_85),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_788),
.B(n_86),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_817),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_835)
);

A2O1A1Ixp33_ASAP7_75t_L g836 ( 
.A1(n_821),
.A2(n_91),
.B(n_92),
.C(n_93),
.Y(n_836)
);

AOI22x1_ASAP7_75t_L g837 ( 
.A1(n_817),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_761),
.B(n_98),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_754),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_768),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_757),
.Y(n_841)
);

INVx1_ASAP7_75t_SL g842 ( 
.A(n_764),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_SL g843 ( 
.A1(n_800),
.A2(n_99),
.B(n_100),
.C(n_101),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_761),
.B(n_104),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_788),
.B(n_105),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_794),
.B(n_106),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_788),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_756),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_758),
.Y(n_849)
);

OAI21x1_ASAP7_75t_L g850 ( 
.A1(n_812),
.A2(n_107),
.B(n_108),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_810),
.B(n_110),
.Y(n_851)
);

OAI21x1_ASAP7_75t_L g852 ( 
.A1(n_789),
.A2(n_790),
.B(n_804),
.Y(n_852)
);

AO31x2_ASAP7_75t_L g853 ( 
.A1(n_809),
.A2(n_111),
.A3(n_112),
.B(n_114),
.Y(n_853)
);

OAI21xp5_ASAP7_75t_L g854 ( 
.A1(n_790),
.A2(n_115),
.B(n_116),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_770),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_804),
.A2(n_117),
.B(n_120),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_778),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_823),
.B(n_122),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_SL g859 ( 
.A(n_802),
.B(n_126),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_783),
.Y(n_860)
);

OA21x2_ASAP7_75t_L g861 ( 
.A1(n_795),
.A2(n_127),
.B(n_128),
.Y(n_861)
);

CKINVDCx6p67_ASAP7_75t_R g862 ( 
.A(n_765),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_768),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_797),
.A2(n_132),
.B1(n_133),
.B2(n_134),
.Y(n_864)
);

O2A1O1Ixp33_ASAP7_75t_SL g865 ( 
.A1(n_800),
.A2(n_136),
.B(n_137),
.C(n_138),
.Y(n_865)
);

OAI21x1_ASAP7_75t_L g866 ( 
.A1(n_811),
.A2(n_139),
.B(n_140),
.Y(n_866)
);

INVx3_ASAP7_75t_L g867 ( 
.A(n_768),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_811),
.A2(n_144),
.B(n_145),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_797),
.A2(n_147),
.B1(n_149),
.B2(n_150),
.Y(n_869)
);

BUFx3_ASAP7_75t_L g870 ( 
.A(n_754),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_813),
.A2(n_821),
.B1(n_802),
.B2(n_807),
.Y(n_871)
);

OA21x2_ASAP7_75t_L g872 ( 
.A1(n_795),
.A2(n_151),
.B(n_152),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_783),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_777),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_777),
.Y(n_875)
);

OAI21xp5_ASAP7_75t_L g876 ( 
.A1(n_799),
.A2(n_155),
.B(n_156),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_806),
.B(n_158),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_820),
.B(n_161),
.Y(n_878)
);

OAI21x1_ASAP7_75t_L g879 ( 
.A1(n_816),
.A2(n_162),
.B(n_163),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_779),
.Y(n_880)
);

OAI21x1_ASAP7_75t_L g881 ( 
.A1(n_816),
.A2(n_165),
.B(n_166),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_779),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_801),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_767),
.Y(n_884)
);

INVx2_ASAP7_75t_SL g885 ( 
.A(n_762),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_807),
.B(n_167),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_807),
.B(n_168),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_SL g888 ( 
.A1(n_813),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_801),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_825),
.A2(n_763),
.B(n_782),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_826),
.B(n_813),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_830),
.B(n_813),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_828),
.Y(n_893)
);

OAI21x1_ASAP7_75t_L g894 ( 
.A1(n_852),
.A2(n_763),
.B(n_782),
.Y(n_894)
);

AOI21x1_ASAP7_75t_L g895 ( 
.A1(n_831),
.A2(n_799),
.B(n_772),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_870),
.Y(n_896)
);

AOI22xp33_ASAP7_75t_SL g897 ( 
.A1(n_859),
.A2(n_821),
.B1(n_802),
.B2(n_808),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_847),
.Y(n_898)
);

AOI22xp33_ASAP7_75t_SL g899 ( 
.A1(n_859),
.A2(n_769),
.B1(n_815),
.B2(n_814),
.Y(n_899)
);

BUFx2_ASAP7_75t_L g900 ( 
.A(n_827),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_829),
.B(n_786),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_862),
.Y(n_902)
);

INVx2_ASAP7_75t_SL g903 ( 
.A(n_841),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_849),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_841),
.Y(n_905)
);

INVxp67_ASAP7_75t_SL g906 ( 
.A(n_873),
.Y(n_906)
);

AOI22xp33_ASAP7_75t_L g907 ( 
.A1(n_876),
.A2(n_766),
.B1(n_818),
.B2(n_792),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_841),
.Y(n_908)
);

CKINVDCx11_ASAP7_75t_R g909 ( 
.A(n_842),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_855),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_857),
.Y(n_911)
);

INVx1_ASAP7_75t_SL g912 ( 
.A(n_842),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_848),
.B(n_766),
.Y(n_913)
);

INVx1_ASAP7_75t_SL g914 ( 
.A(n_875),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_860),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_831),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_853),
.Y(n_917)
);

OA21x2_ASAP7_75t_L g918 ( 
.A1(n_832),
.A2(n_818),
.B(n_780),
.Y(n_918)
);

BUFx3_ASAP7_75t_L g919 ( 
.A(n_883),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_889),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_874),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_853),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_853),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_839),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_861),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_861),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_872),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_872),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_824),
.Y(n_929)
);

OAI22xp33_ASAP7_75t_L g930 ( 
.A1(n_876),
.A2(n_792),
.B1(n_784),
.B2(n_771),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_824),
.Y(n_931)
);

AO21x2_ASAP7_75t_L g932 ( 
.A1(n_832),
.A2(n_780),
.B(n_786),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_833),
.Y(n_933)
);

AO21x1_ASAP7_75t_SL g934 ( 
.A1(n_854),
.A2(n_786),
.B(n_791),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_850),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_856),
.A2(n_798),
.B(n_755),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_911),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_912),
.B(n_914),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_912),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_909),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_902),
.Y(n_941)
);

BUFx2_ASAP7_75t_L g942 ( 
.A(n_896),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_896),
.Y(n_943)
);

OAI22xp5_ASAP7_75t_L g944 ( 
.A1(n_899),
.A2(n_877),
.B1(n_888),
.B2(n_836),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_904),
.Y(n_945)
);

AOI22xp33_ASAP7_75t_L g946 ( 
.A1(n_907),
.A2(n_864),
.B1(n_869),
.B2(n_878),
.Y(n_946)
);

CKINVDCx20_ASAP7_75t_R g947 ( 
.A(n_896),
.Y(n_947)
);

HB1xp67_ASAP7_75t_L g948 ( 
.A(n_900),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_R g949 ( 
.A(n_918),
.B(n_877),
.Y(n_949)
);

NAND2xp33_ASAP7_75t_R g950 ( 
.A(n_918),
.B(n_877),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_921),
.B(n_885),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_904),
.Y(n_952)
);

INVx2_ASAP7_75t_SL g953 ( 
.A(n_924),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_897),
.A2(n_835),
.B1(n_837),
.B2(n_871),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_921),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_921),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_918),
.B(n_881),
.Y(n_957)
);

BUFx8_ASAP7_75t_SL g958 ( 
.A(n_919),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_892),
.B(n_880),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_910),
.Y(n_960)
);

BUFx3_ASAP7_75t_L g961 ( 
.A(n_919),
.Y(n_961)
);

HB1xp67_ASAP7_75t_L g962 ( 
.A(n_900),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_919),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_892),
.B(n_882),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_924),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_895),
.B(n_765),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_939),
.B(n_914),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_945),
.Y(n_968)
);

OR2x2_ASAP7_75t_SL g969 ( 
.A(n_938),
.B(n_918),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_942),
.B(n_916),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_958),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_952),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_948),
.B(n_916),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_937),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_937),
.Y(n_975)
);

AND2x2_ASAP7_75t_L g976 ( 
.A(n_962),
.B(n_916),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_961),
.B(n_929),
.Y(n_977)
);

INVx1_ASAP7_75t_SL g978 ( 
.A(n_940),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_960),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_961),
.Y(n_980)
);

INVx4_ASAP7_75t_R g981 ( 
.A(n_953),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_959),
.Y(n_982)
);

OR2x2_ASAP7_75t_L g983 ( 
.A(n_957),
.B(n_925),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_964),
.Y(n_984)
);

AND2x2_ASAP7_75t_L g985 ( 
.A(n_957),
.B(n_929),
.Y(n_985)
);

OR2x2_ASAP7_75t_L g986 ( 
.A(n_957),
.B(n_925),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_955),
.Y(n_987)
);

OR2x2_ASAP7_75t_L g988 ( 
.A(n_957),
.B(n_926),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_983),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_987),
.B(n_965),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_967),
.B(n_951),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_979),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_969),
.A2(n_946),
.B1(n_944),
.B2(n_947),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_974),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_979),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_968),
.Y(n_996)
);

AOI22xp5_ASAP7_75t_L g997 ( 
.A1(n_971),
.A2(n_949),
.B1(n_950),
.B2(n_954),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_974),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_R g999 ( 
.A(n_980),
.B(n_966),
.Y(n_999)
);

OAI21x1_ASAP7_75t_L g1000 ( 
.A1(n_983),
.A2(n_928),
.B(n_927),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_970),
.B(n_955),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_982),
.B(n_956),
.Y(n_1002)
);

NOR2x1_ASAP7_75t_SL g1003 ( 
.A(n_971),
.B(n_934),
.Y(n_1003)
);

NAND4xp25_ASAP7_75t_L g1004 ( 
.A(n_986),
.B(n_846),
.C(n_913),
.D(n_858),
.Y(n_1004)
);

INVx2_ASAP7_75t_L g1005 ( 
.A(n_986),
.Y(n_1005)
);

BUFx2_ASAP7_75t_L g1006 ( 
.A(n_971),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_1006),
.Y(n_1007)
);

OAI211xp5_ASAP7_75t_L g1008 ( 
.A1(n_997),
.A2(n_971),
.B(n_854),
.C(n_895),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_1002),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_993),
.B(n_978),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_989),
.Y(n_1011)
);

OR2x2_ASAP7_75t_L g1012 ( 
.A(n_1005),
.B(n_984),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_1003),
.B(n_985),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_1001),
.B(n_985),
.Y(n_1014)
);

INVx2_ASAP7_75t_L g1015 ( 
.A(n_995),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_996),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_995),
.B(n_972),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_1000),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_1013),
.B(n_980),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_1016),
.Y(n_1020)
);

NAND2x1p5_ASAP7_75t_L g1021 ( 
.A(n_1007),
.B(n_757),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_977),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_1015),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_1017),
.Y(n_1024)
);

NAND2x1p5_ASAP7_75t_L g1025 ( 
.A(n_1009),
.B(n_757),
.Y(n_1025)
);

INVxp67_ASAP7_75t_L g1026 ( 
.A(n_1010),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_1017),
.Y(n_1027)
);

OAI22xp5_ASAP7_75t_L g1028 ( 
.A1(n_1026),
.A2(n_1010),
.B1(n_1008),
.B2(n_947),
.Y(n_1028)
);

AOI32xp33_ASAP7_75t_L g1029 ( 
.A1(n_1019),
.A2(n_1011),
.A3(n_930),
.B1(n_1008),
.B2(n_1018),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_1025),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_1025),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_1022),
.B(n_1012),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_1026),
.B(n_992),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_1033),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_1032),
.B(n_1023),
.Y(n_1035)
);

INVx4_ASAP7_75t_L g1036 ( 
.A(n_1030),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_1028),
.B(n_1020),
.Y(n_1037)
);

INVx4_ASAP7_75t_L g1038 ( 
.A(n_1031),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_1029),
.B(n_1024),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_1032),
.B(n_1027),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_1033),
.B(n_1021),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1033),
.B(n_1021),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_1033),
.Y(n_1043)
);

OR2x2_ASAP7_75t_L g1044 ( 
.A(n_1035),
.B(n_991),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_1036),
.B(n_990),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_1038),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_1037),
.B(n_941),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_1040),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_1040),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_1039),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_1034),
.B(n_990),
.Y(n_1051)
);

BUFx3_ASAP7_75t_L g1052 ( 
.A(n_1049),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_1050),
.A2(n_1043),
.B1(n_1041),
.B2(n_999),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_1047),
.A2(n_1045),
.B(n_1051),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_1048),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1046),
.B(n_1042),
.Y(n_1056)
);

OR2x2_ASAP7_75t_L g1057 ( 
.A(n_1044),
.B(n_1018),
.Y(n_1057)
);

OAI22xp5_ASAP7_75t_L g1058 ( 
.A1(n_1050),
.A2(n_941),
.B1(n_943),
.B2(n_988),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_1052),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_1055),
.B(n_994),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_1056),
.Y(n_1061)
);

AND2x4_ASAP7_75t_L g1062 ( 
.A(n_1053),
.B(n_977),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1054),
.B(n_994),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_SL g1064 ( 
.A(n_1059),
.B(n_1058),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1061),
.B(n_1057),
.Y(n_1065)
);

OAI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1062),
.A2(n_887),
.B(n_886),
.Y(n_1066)
);

INVx1_ASAP7_75t_SL g1067 ( 
.A(n_1063),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_1060),
.Y(n_1068)
);

NAND2x1_ASAP7_75t_SL g1069 ( 
.A(n_1060),
.B(n_999),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_1068),
.B(n_998),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_1065),
.Y(n_1071)
);

AOI222xp33_ASAP7_75t_L g1072 ( 
.A1(n_1064),
.A2(n_771),
.B1(n_844),
.B2(n_886),
.C1(n_887),
.C2(n_851),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_1067),
.B(n_998),
.Y(n_1073)
);

AOI221xp5_ASAP7_75t_L g1074 ( 
.A1(n_1066),
.A2(n_865),
.B1(n_843),
.B2(n_764),
.C(n_1004),
.Y(n_1074)
);

AND2x2_ASAP7_75t_L g1075 ( 
.A(n_1069),
.B(n_982),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_1071),
.Y(n_1076)
);

OAI211xp5_ASAP7_75t_L g1077 ( 
.A1(n_1073),
.A2(n_851),
.B(n_858),
.C(n_760),
.Y(n_1077)
);

NAND4xp75_ASAP7_75t_L g1078 ( 
.A(n_1070),
.B(n_838),
.C(n_845),
.D(n_834),
.Y(n_1078)
);

AOI221xp5_ASAP7_75t_L g1079 ( 
.A1(n_1075),
.A2(n_844),
.B1(n_988),
.B2(n_845),
.C(n_834),
.Y(n_1079)
);

INVxp67_ASAP7_75t_SL g1080 ( 
.A(n_1072),
.Y(n_1080)
);

OR2x2_ASAP7_75t_L g1081 ( 
.A(n_1074),
.B(n_970),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_1071),
.A2(n_933),
.B(n_879),
.Y(n_1082)
);

NOR4xp75_ASAP7_75t_L g1083 ( 
.A(n_1073),
.B(n_981),
.C(n_863),
.D(n_840),
.Y(n_1083)
);

AOI211xp5_ASAP7_75t_L g1084 ( 
.A1(n_1076),
.A2(n_759),
.B(n_760),
.C(n_866),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_1080),
.B(n_958),
.Y(n_1085)
);

AND4x1_ASAP7_75t_L g1086 ( 
.A(n_1079),
.B(n_759),
.C(n_931),
.D(n_775),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_1081),
.B(n_774),
.Y(n_1087)
);

OAI321xp33_ASAP7_75t_L g1088 ( 
.A1(n_1077),
.A2(n_759),
.A3(n_798),
.B1(n_903),
.B2(n_905),
.C(n_931),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_1082),
.A2(n_776),
.B(n_868),
.C(n_908),
.Y(n_1089)
);

AOI211xp5_ASAP7_75t_L g1090 ( 
.A1(n_1083),
.A2(n_908),
.B(n_903),
.C(n_905),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1078),
.B(n_975),
.Y(n_1091)
);

AOI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_1085),
.A2(n_933),
.B(n_175),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_1086),
.Y(n_1093)
);

AOI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_1087),
.A2(n_963),
.B1(n_863),
.B2(n_867),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_1091),
.B(n_963),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_1088),
.B(n_840),
.Y(n_1096)
);

AOI32xp33_ASAP7_75t_L g1097 ( 
.A1(n_1090),
.A2(n_908),
.A3(n_976),
.B1(n_973),
.B2(n_867),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_1084),
.A2(n_920),
.B1(n_898),
.B2(n_933),
.Y(n_1098)
);

AND2x2_ASAP7_75t_L g1099 ( 
.A(n_1089),
.B(n_976),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1085),
.Y(n_1100)
);

NAND3xp33_ASAP7_75t_L g1101 ( 
.A(n_1085),
.B(n_767),
.C(n_779),
.Y(n_1101)
);

OAI211xp5_ASAP7_75t_SL g1102 ( 
.A1(n_1100),
.A2(n_174),
.B(n_177),
.C(n_178),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1095),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_1099),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1101),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_1093),
.B(n_973),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_1094),
.B(n_920),
.Y(n_1107)
);

OAI211xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1092),
.A2(n_179),
.B(n_180),
.C(n_181),
.Y(n_1108)
);

NOR2x1_ASAP7_75t_L g1109 ( 
.A(n_1096),
.B(n_884),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_1097),
.B(n_920),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1098),
.B(n_898),
.Y(n_1111)
);

INVx2_ASAP7_75t_SL g1112 ( 
.A(n_1095),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1095),
.Y(n_1113)
);

NAND4xp75_ASAP7_75t_L g1114 ( 
.A(n_1100),
.B(n_185),
.C(n_187),
.D(n_188),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_1106),
.B(n_975),
.Y(n_1115)
);

BUFx2_ASAP7_75t_L g1116 ( 
.A(n_1109),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_1112),
.Y(n_1117)
);

BUFx2_ASAP7_75t_L g1118 ( 
.A(n_1104),
.Y(n_1118)
);

CKINVDCx14_ASAP7_75t_R g1119 ( 
.A(n_1103),
.Y(n_1119)
);

OAI22x1_ASAP7_75t_SL g1120 ( 
.A1(n_1113),
.A2(n_884),
.B1(n_192),
.B2(n_193),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_1114),
.Y(n_1121)
);

INVx1_ASAP7_75t_SL g1122 ( 
.A(n_1105),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_SL g1123 ( 
.A(n_1107),
.Y(n_1123)
);

AO22x2_ASAP7_75t_L g1124 ( 
.A1(n_1122),
.A2(n_1110),
.B1(n_1111),
.B2(n_1108),
.Y(n_1124)
);

AO22x2_ASAP7_75t_L g1125 ( 
.A1(n_1119),
.A2(n_1102),
.B1(n_926),
.B2(n_928),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1118),
.A2(n_755),
.B(n_891),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1117),
.A2(n_890),
.B(n_915),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1123),
.A2(n_1121),
.B1(n_1116),
.B2(n_1115),
.Y(n_1128)
);

OAI21xp33_ASAP7_75t_SL g1129 ( 
.A1(n_1120),
.A2(n_936),
.B(n_906),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1117),
.B(n_915),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1124),
.Y(n_1131)
);

AOI222xp33_ASAP7_75t_L g1132 ( 
.A1(n_1129),
.A2(n_1128),
.B1(n_1125),
.B2(n_1130),
.C1(n_1126),
.C2(n_1127),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1128),
.A2(n_936),
.B(n_894),
.Y(n_1133)
);

INVxp67_ASAP7_75t_SL g1134 ( 
.A(n_1131),
.Y(n_1134)
);

OAI22x1_ASAP7_75t_L g1135 ( 
.A1(n_1134),
.A2(n_1132),
.B1(n_1133),
.B2(n_791),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_1135),
.B(n_934),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1136),
.B(n_191),
.Y(n_1137)
);

OAI22xp33_ASAP7_75t_L g1138 ( 
.A1(n_1136),
.A2(n_791),
.B1(n_796),
.B2(n_801),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1136),
.Y(n_1139)
);

AOI222xp33_ASAP7_75t_SL g1140 ( 
.A1(n_1139),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.C1(n_199),
.C2(n_201),
.Y(n_1140)
);

AOI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1137),
.A2(n_932),
.B1(n_891),
.B2(n_928),
.Y(n_1141)
);

XOR2x1_ASAP7_75t_L g1142 ( 
.A(n_1138),
.B(n_203),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1139),
.A2(n_922),
.B1(n_935),
.B2(n_917),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_SL g1144 ( 
.A1(n_1142),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_1144)
);

AOI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1140),
.A2(n_932),
.B1(n_927),
.B2(n_791),
.Y(n_1145)
);

AOI31xp33_ASAP7_75t_L g1146 ( 
.A1(n_1143),
.A2(n_210),
.A3(n_935),
.B(n_922),
.Y(n_1146)
);

AOI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1141),
.A2(n_932),
.B1(n_935),
.B2(n_901),
.Y(n_1147)
);

AO21x2_ASAP7_75t_L g1148 ( 
.A1(n_1146),
.A2(n_1144),
.B(n_1145),
.Y(n_1148)
);

AOI221xp5_ASAP7_75t_L g1149 ( 
.A1(n_1147),
.A2(n_910),
.B1(n_893),
.B2(n_923),
.C(n_917),
.Y(n_1149)
);

AOI221xp5_ASAP7_75t_L g1150 ( 
.A1(n_1148),
.A2(n_893),
.B1(n_923),
.B2(n_917),
.C(n_911),
.Y(n_1150)
);

AOI211xp5_ASAP7_75t_L g1151 ( 
.A1(n_1150),
.A2(n_1149),
.B(n_805),
.C(n_923),
.Y(n_1151)
);


endmodule