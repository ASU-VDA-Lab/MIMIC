module fake_jpeg_30269_n_480 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_480);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_480;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

OR2x2_ASAP7_75t_L g17 ( 
.A(n_3),
.B(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_49),
.Y(n_129)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_51),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_17),
.B(n_8),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_59),
.B(n_61),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_22),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_60),
.B(n_65),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_17),
.B(n_8),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_62),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_43),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_66),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_17),
.B(n_8),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_67),
.B(n_70),
.Y(n_113)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_69),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_7),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_71),
.Y(n_146)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_73),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_75),
.Y(n_105)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_7),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_77),
.B(n_81),
.Y(n_143)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_33),
.Y(n_80)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_19),
.B(n_7),
.Y(n_81)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_82),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_33),
.Y(n_83)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_21),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_87),
.B(n_47),
.Y(n_109)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_88),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_20),
.B(n_9),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_89),
.B(n_23),
.Y(n_150)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_90),
.Y(n_153)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_41),
.Y(n_92)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_92),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_21),
.Y(n_94)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_95),
.Y(n_148)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_96),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_46),
.Y(n_97)
);

BUFx8_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_21),
.Y(n_99)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_99),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_49),
.A2(n_47),
.B1(n_20),
.B2(n_40),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_101),
.A2(n_32),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

AO22x1_ASAP7_75t_SL g107 ( 
.A1(n_54),
.A2(n_98),
.B1(n_51),
.B2(n_95),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_107),
.B(n_109),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_62),
.B1(n_92),
.B2(n_57),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_111),
.A2(n_152),
.B1(n_80),
.B2(n_86),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_115),
.B(n_37),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_52),
.B(n_29),
.C(n_23),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_121),
.B(n_34),
.C(n_26),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g122 ( 
.A(n_58),
.Y(n_122)
);

INVx11_ASAP7_75t_L g180 ( 
.A(n_122),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_93),
.A2(n_39),
.B1(n_46),
.B2(n_35),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_139),
.B1(n_58),
.B2(n_39),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_97),
.A2(n_39),
.B1(n_35),
.B2(n_38),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_150),
.B(n_40),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_63),
.A2(n_35),
.B1(n_39),
.B2(n_22),
.Y(n_152)
);

INVx13_ASAP7_75t_L g154 ( 
.A(n_75),
.Y(n_154)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_154),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_79),
.Y(n_155)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_155),
.Y(n_163)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_105),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g216 ( 
.A(n_158),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_160),
.A2(n_166),
.B1(n_210),
.B2(n_100),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_110),
.Y(n_161)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_162),
.B(n_177),
.Y(n_227)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_165),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_141),
.A2(n_69),
.B1(n_64),
.B2(n_91),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_167),
.A2(n_172),
.B1(n_186),
.B2(n_129),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_132),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_168),
.B(n_197),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_113),
.B(n_29),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g219 ( 
.A(n_169),
.B(n_195),
.Y(n_219)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_170),
.Y(n_236)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_171),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_131),
.A2(n_38),
.B1(n_39),
.B2(n_84),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_103),
.Y(n_173)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_173),
.Y(n_220)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_128),
.A2(n_74),
.B1(n_82),
.B2(n_38),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_174),
.A2(n_207),
.B1(n_142),
.B2(n_148),
.Y(n_224)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_120),
.Y(n_175)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_175),
.Y(n_243)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_106),
.Y(n_176)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_113),
.A2(n_22),
.B(n_44),
.C(n_25),
.Y(n_177)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_127),
.Y(n_178)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_178),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx8_ASAP7_75t_L g217 ( 
.A(n_179),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g181 ( 
.A(n_126),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_190),
.Y(n_212)
);

AO22x2_ASAP7_75t_L g183 ( 
.A1(n_123),
.A2(n_32),
.B1(n_44),
.B2(n_25),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g215 ( 
.A1(n_183),
.A2(n_139),
.B1(n_152),
.B2(n_111),
.Y(n_215)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_133),
.Y(n_184)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

BUFx6f_ASAP7_75t_SL g185 ( 
.A(n_122),
.Y(n_185)
);

BUFx4f_ASAP7_75t_SL g252 ( 
.A(n_185),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_131),
.A2(n_39),
.B1(n_28),
.B2(n_27),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_188),
.Y(n_250)
);

BUFx4f_ASAP7_75t_L g189 ( 
.A(n_155),
.Y(n_189)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_189),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_25),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_191),
.Y(n_237)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_153),
.Y(n_192)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_193),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_199),
.Y(n_245)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_147),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_135),
.Y(n_196)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_196),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_143),
.B(n_37),
.Y(n_197)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_136),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_112),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_200),
.B(n_208),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_108),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_201),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_112),
.B(n_34),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_204),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_L g203 ( 
.A1(n_107),
.A2(n_44),
.B(n_28),
.C(n_27),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_205),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_26),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_116),
.B(n_28),
.C(n_27),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_149),
.A2(n_32),
.B1(n_45),
.B2(n_42),
.Y(n_207)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_134),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_122),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_211),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_117),
.B(n_10),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_215),
.A2(n_158),
.B(n_208),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_207),
.A2(n_140),
.B(n_2),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_223),
.A2(n_45),
.B(n_42),
.Y(n_286)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_224),
.A2(n_191),
.B1(n_178),
.B2(n_176),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_159),
.A2(n_119),
.B1(n_100),
.B2(n_157),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_225),
.A2(n_232),
.B1(n_233),
.B2(n_241),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_189),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_229),
.B(n_249),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_231),
.A2(n_248),
.B1(n_193),
.B2(n_190),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_174),
.A2(n_119),
.B1(n_157),
.B2(n_145),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_166),
.A2(n_142),
.B1(n_145),
.B2(n_144),
.Y(n_233)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_170),
.B1(n_195),
.B2(n_196),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_203),
.A2(n_144),
.B1(n_138),
.B2(n_137),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_L g248 ( 
.A1(n_183),
.A2(n_138),
.B1(n_137),
.B2(n_118),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_201),
.Y(n_249)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_250),
.Y(n_256)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_256),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_215),
.A2(n_160),
.B1(n_183),
.B2(n_167),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_257),
.A2(n_262),
.B1(n_278),
.B2(n_293),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_258),
.Y(n_323)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_259),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g260 ( 
.A(n_246),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_260),
.B(n_279),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_261),
.A2(n_263),
.B1(n_274),
.B2(n_283),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_215),
.A2(n_183),
.B1(n_172),
.B2(n_186),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_245),
.Y(n_264)
);

OR2x2_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_270),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g265 ( 
.A1(n_223),
.A2(n_169),
.B(n_177),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_265),
.A2(n_288),
.B(n_244),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_239),
.B(n_163),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_266),
.B(n_267),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_239),
.B(n_181),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g327 ( 
.A1(n_269),
.A2(n_281),
.B(n_286),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_219),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_212),
.B(n_179),
.C(n_154),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_271),
.B(n_287),
.C(n_236),
.Y(n_294)
);

INVx3_ASAP7_75t_SL g272 ( 
.A(n_217),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_272),
.Y(n_300)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_228),
.Y(n_273)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_273),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_231),
.A2(n_248),
.B1(n_227),
.B2(n_241),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_222),
.B(n_198),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_276),
.B(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_234),
.Y(n_277)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_277),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_225),
.A2(n_224),
.B1(n_232),
.B2(n_255),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_247),
.B(n_219),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_280),
.B(n_282),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_221),
.A2(n_218),
.B(n_212),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_220),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_212),
.A2(n_198),
.B1(n_180),
.B2(n_118),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_254),
.A2(n_180),
.B1(n_2),
.B2(n_3),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_290),
.B1(n_240),
.B2(n_238),
.Y(n_314)
);

AO21x2_ASAP7_75t_L g285 ( 
.A1(n_221),
.A2(n_45),
.B(n_42),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_285),
.A2(n_244),
.B1(n_230),
.B2(n_251),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_214),
.C(n_226),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_243),
.A2(n_45),
.B1(n_2),
.B2(n_4),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_218),
.B(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_291),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_216),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_234),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_238),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_292),
.B(n_242),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_216),
.A2(n_230),
.B1(n_237),
.B2(n_213),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g329 ( 
.A(n_294),
.B(n_287),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_268),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_295),
.Y(n_333)
);

NAND3xp33_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_214),
.C(n_237),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_298),
.B(n_288),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_303),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_266),
.B(n_236),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_302),
.B(n_319),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_282),
.B(n_242),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g304 ( 
.A(n_263),
.B(n_213),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_304),
.A2(n_324),
.B(n_285),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_306),
.A2(n_323),
.B1(n_312),
.B2(n_295),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_314),
.B1(n_321),
.B2(n_275),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g357 ( 
.A(n_312),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_280),
.B(n_251),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_313),
.B(n_11),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_264),
.B(n_240),
.Y(n_315)
);

A2O1A1O1Ixp25_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_322),
.B(n_289),
.C(n_268),
.D(n_273),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_257),
.A2(n_253),
.B1(n_252),
.B2(n_10),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_316),
.A2(n_259),
.B1(n_285),
.B2(n_14),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_SL g319 ( 
.A(n_267),
.B(n_265),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_274),
.A2(n_252),
.B1(n_9),
.B2(n_11),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_276),
.B(n_5),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_286),
.A2(n_252),
.B(n_9),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_271),
.B(n_5),
.C(n_11),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_326),
.C(n_256),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_281),
.B(n_16),
.C(n_12),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_329),
.B(n_335),
.C(n_302),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_330),
.A2(n_341),
.B1(n_342),
.B2(n_349),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_304),
.A2(n_262),
.B1(n_269),
.B2(n_278),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_331),
.A2(n_338),
.B1(n_350),
.B2(n_306),
.Y(n_365)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_297),
.Y(n_334)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_319),
.B(n_308),
.Y(n_335)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_299),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_337),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_304),
.A2(n_275),
.B1(n_286),
.B2(n_261),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_283),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g379 ( 
.A(n_339),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_340),
.A2(n_352),
.B(n_356),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_305),
.A2(n_284),
.B1(n_290),
.B2(n_272),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_277),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g366 ( 
.A(n_343),
.B(n_344),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_299),
.B(n_292),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_308),
.B(n_285),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_345),
.B(n_296),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_346),
.A2(n_300),
.B(n_311),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_318),
.Y(n_347)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_347),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_313),
.B(n_291),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_348),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_305),
.A2(n_272),
.B1(n_285),
.B2(n_279),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_310),
.A2(n_293),
.B1(n_279),
.B2(n_285),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_351),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_301),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g373 ( 
.A1(n_353),
.A2(n_300),
.B1(n_322),
.B2(n_296),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_354),
.Y(n_378)
);

OA22x2_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_12),
.B1(n_14),
.B2(n_15),
.Y(n_355)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_355),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_315),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_294),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_358),
.B(n_359),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_329),
.B(n_327),
.C(n_320),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_363),
.B(n_368),
.C(n_377),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_328),
.B(n_327),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_364),
.B(n_369),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_365),
.A2(n_373),
.B1(n_333),
.B2(n_353),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_337),
.A2(n_309),
.B(n_310),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_367),
.A2(n_376),
.B(n_382),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_357),
.B(n_320),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_303),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_372),
.B(n_345),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_325),
.C(n_317),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_L g382 ( 
.A1(n_339),
.A2(n_326),
.B(n_307),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_346),
.A2(n_321),
.B(n_317),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_383),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_L g384 ( 
.A1(n_339),
.A2(n_307),
.B(n_297),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_384),
.B(n_338),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_385),
.B(n_396),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_374),
.A2(n_331),
.B1(n_330),
.B2(n_350),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_386),
.A2(n_383),
.B1(n_367),
.B2(n_380),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_370),
.B(n_333),
.Y(n_388)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_388),
.Y(n_412)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_366),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_392),
.B(n_394),
.Y(n_410)
);

OA22x2_ASAP7_75t_L g424 ( 
.A1(n_393),
.A2(n_403),
.B1(n_404),
.B2(n_380),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_361),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_356),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_395),
.B(n_399),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_358),
.B(n_359),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_352),
.C(n_332),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_406),
.C(n_372),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_398),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_332),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_361),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_400),
.B(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_360),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_402),
.B(n_379),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_362),
.A2(n_314),
.B1(n_334),
.B2(n_355),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_365),
.A2(n_355),
.B1(n_336),
.B2(n_354),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_318),
.C(n_355),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_14),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_SL g417 ( 
.A(n_407),
.B(n_369),
.Y(n_417)
);

XNOR2x1_ASAP7_75t_L g430 ( 
.A(n_408),
.B(n_422),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_409),
.A2(n_413),
.B1(n_387),
.B2(n_393),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_387),
.A2(n_379),
.B1(n_374),
.B2(n_371),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_389),
.B(n_363),
.C(n_377),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_414),
.B(n_396),
.C(n_389),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_399),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_417),
.B(n_419),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_388),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_390),
.B(n_382),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_425),
.Y(n_427)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_421),
.Y(n_438)
);

XNOR2x1_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_368),
.Y(n_422)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_424),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_395),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_432),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_428),
.B(n_386),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_417),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_410),
.B(n_378),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_414),
.B(n_397),
.C(n_391),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_433),
.B(n_437),
.C(n_439),
.Y(n_446)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_412),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_435),
.B(n_440),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_408),
.B(n_406),
.C(n_405),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_411),
.B(n_405),
.C(n_384),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

NOR3xp33_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_378),
.C(n_413),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_441),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_442),
.B(n_443),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_430),
.B(n_411),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_435),
.B(n_404),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_444),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_434),
.A2(n_403),
.B1(n_423),
.B2(n_424),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_445),
.B(n_450),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_434),
.A2(n_423),
.B1(n_424),
.B2(n_385),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_448),
.B(n_449),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_431),
.B(n_422),
.C(n_407),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_375),
.Y(n_452)
);

CKINVDCx14_ASAP7_75t_R g459 ( 
.A(n_452),
.Y(n_459)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_447),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_454),
.B(n_455),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_446),
.B(n_438),
.Y(n_455)
);

OAI21xp5_ASAP7_75t_SL g458 ( 
.A1(n_444),
.A2(n_429),
.B(n_439),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g463 ( 
.A(n_458),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_446),
.B(n_427),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_461),
.B(n_450),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_L g465 ( 
.A1(n_456),
.A2(n_451),
.B1(n_448),
.B2(n_436),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_465),
.B(n_466),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_457),
.B(n_442),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_460),
.A2(n_437),
.B(n_433),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_467),
.B(n_468),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_464),
.A2(n_463),
.B(n_458),
.Y(n_471)
);

AO21x1_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_472),
.B(n_453),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_463),
.A2(n_462),
.B(n_459),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_469),
.A2(n_453),
.B(n_462),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g476 ( 
.A(n_473),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_474),
.B(n_470),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_475),
.B(n_428),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_477),
.A2(n_476),
.B(n_375),
.Y(n_478)
);

A2O1A1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_478),
.A2(n_430),
.B(n_443),
.C(n_15),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_479),
.B(n_15),
.Y(n_480)
);


endmodule