module fake_jpeg_29086_n_237 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_237);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_237;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_46),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_23),
.Y(n_41)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_35),
.B(n_17),
.Y(n_46)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_28),
.Y(n_48)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_22),
.Y(n_59)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_51),
.Y(n_57)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_22),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_37),
.C(n_31),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_36),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_63),
.B(n_67),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_39),
.B(n_21),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_68),
.B(n_70),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_29),
.B1(n_18),
.B2(n_34),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_81),
.B1(n_49),
.B2(n_42),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_30),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_26),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_20),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_50),
.B(n_30),
.Y(n_73)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp33_ASAP7_75t_SL g74 ( 
.A(n_47),
.B(n_18),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_74),
.A2(n_37),
.B(n_31),
.Y(n_99)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_50),
.B(n_21),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_18),
.B1(n_34),
.B2(n_24),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_66),
.B1(n_71),
.B2(n_62),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_64),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_97),
.Y(n_115)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_72),
.A2(n_50),
.A3(n_33),
.B1(n_32),
.B2(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_89),
.B(n_97),
.Y(n_114)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_90),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_96),
.Y(n_121)
);

A2O1A1Ixp33_ASAP7_75t_SL g94 ( 
.A1(n_74),
.A2(n_48),
.B(n_43),
.C(n_42),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_82),
.B(n_76),
.C(n_66),
.Y(n_123)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_108),
.B(n_65),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_55),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_103),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_80),
.A2(n_43),
.B1(n_48),
.B2(n_44),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_109),
.B1(n_110),
.B2(n_0),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_33),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_64),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_105),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_77),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_77),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_71),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_32),
.B1(n_20),
.B2(n_24),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_80),
.A2(n_27),
.B1(n_19),
.B2(n_25),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_54),
.A2(n_27),
.B1(n_25),
.B2(n_34),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_56),
.Y(n_111)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_54),
.B(n_27),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_25),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_120),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_112),
.A2(n_79),
.B1(n_76),
.B2(n_62),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_118),
.B1(n_128),
.B2(n_132),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_108),
.Y(n_120)
);

AO22x1_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_94),
.B1(n_102),
.B2(n_89),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_85),
.B(n_65),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_124),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_98),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_93),
.B(n_0),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_84),
.B(n_0),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_135),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_94),
.A2(n_1),
.B1(n_4),
.B2(n_6),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_88),
.B1(n_95),
.B2(n_106),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_91),
.B(n_1),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_4),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_103),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_136),
.B(n_92),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_127),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_101),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_142),
.B(n_145),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_98),
.C(n_91),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_143),
.B(n_122),
.C(n_126),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_144),
.B(n_148),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_146),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_149),
.B(n_151),
.Y(n_162)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_125),
.Y(n_152)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_116),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_130),
.Y(n_154)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_129),
.B(n_115),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_155),
.B(n_156),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_129),
.B(n_113),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_134),
.B1(n_117),
.B2(n_110),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_115),
.B(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_159),
.B(n_122),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_137),
.Y(n_160)
);

AO221x1_ASAP7_75t_L g164 ( 
.A1(n_160),
.A2(n_105),
.B1(n_124),
.B2(n_130),
.C(n_137),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_144),
.A2(n_120),
.B1(n_128),
.B2(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_164),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_171),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_172),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_147),
.B(n_131),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_174),
.C(n_145),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_111),
.C(n_90),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_135),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_176),
.B(n_177),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_155),
.B(n_132),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_138),
.B(n_133),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_178),
.B(n_160),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_SL g182 ( 
.A1(n_179),
.A2(n_144),
.B(n_123),
.C(n_139),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_182),
.A2(n_184),
.B(n_196),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_147),
.Y(n_183)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_183),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_179),
.A2(n_158),
.B(n_140),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_185),
.B(n_191),
.C(n_195),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_179),
.A2(n_143),
.B(n_150),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_184),
.B(n_173),
.Y(n_204)
);

AOI322xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_139),
.A3(n_156),
.B1(n_150),
.B2(n_151),
.C1(n_157),
.C2(n_123),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_175),
.B(n_154),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_190),
.B(n_167),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_170),
.B(n_133),
.C(n_83),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_193),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_109),
.C(n_12),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_6),
.B(n_7),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_181),
.A2(n_161),
.B1(n_180),
.B2(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_197),
.A2(n_186),
.B1(n_182),
.B2(n_195),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_207),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_204),
.B(n_205),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_174),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_165),
.C(n_177),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_206),
.B(n_205),
.C(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_192),
.B(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_194),
.B(n_163),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_7),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_215),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_196),
.Y(n_211)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_211),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_213),
.B(n_217),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_199),
.A2(n_182),
.B(n_166),
.Y(n_214)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_214),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_SL g215 ( 
.A1(n_199),
.A2(n_182),
.B(n_166),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_216),
.A2(n_197),
.B1(n_202),
.B2(n_201),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_206),
.B(n_8),
.Y(n_217)
);

BUFx24_ASAP7_75t_SL g219 ( 
.A(n_209),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_221),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_217),
.B(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_10),
.Y(n_229)
);

OAI221xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_204),
.B1(n_223),
.B2(n_218),
.C(n_222),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_225),
.B(n_228),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_222),
.A2(n_212),
.B1(n_215),
.B2(n_198),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_227),
.A2(n_16),
.B1(n_10),
.B2(n_13),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_222),
.B(n_213),
.C(n_212),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_229),
.B(n_14),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_231),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_232),
.A2(n_233),
.B(n_226),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_228),
.A2(n_15),
.B(n_8),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_234),
.B(n_230),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_236),
.B(n_235),
.Y(n_237)
);


endmodule