module fake_jpeg_11078_n_296 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_296);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_296;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_200;
wire n_96;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_8),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx2_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_20),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_44),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_0),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_49),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_20),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_41),
.Y(n_100)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_47),
.Y(n_87)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_18),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_27),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_50),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_51),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_26),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_16),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_54),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_0),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx3_ASAP7_75t_SL g57 ( 
.A(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_58),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_31),
.Y(n_59)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_1),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_61),
.B(n_68),
.Y(n_83)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_62),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g82 ( 
.A(n_64),
.Y(n_82)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_65),
.Y(n_93)
);

INVx3_ASAP7_75t_SL g66 ( 
.A(n_19),
.Y(n_66)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_32),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_48),
.A2(n_25),
.B1(n_27),
.B2(n_39),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_71),
.B1(n_73),
.B2(n_76),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_40),
.B1(n_39),
.B2(n_33),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_33),
.B1(n_40),
.B2(n_22),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_37),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_96),
.B(n_45),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_46),
.A2(n_22),
.B1(n_30),
.B2(n_25),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_30),
.B1(n_56),
.B2(n_57),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_81),
.B(n_95),
.C(n_23),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_42),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_80),
.B(n_34),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_57),
.A2(n_25),
.B1(n_38),
.B2(n_36),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_66),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_95)
);

NAND2xp33_ASAP7_75t_SL g96 ( 
.A(n_67),
.B(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_100),
.B(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_101),
.Y(n_111)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_106),
.B(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_44),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_109),
.B(n_115),
.Y(n_167)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_69),
.Y(n_110)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_112),
.B(n_120),
.Y(n_150)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_72),
.B(n_21),
.Y(n_115)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_117),
.A2(n_104),
.B1(n_97),
.B2(n_105),
.Y(n_141)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_118),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_34),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_125),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_87),
.Y(n_122)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_122),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g124 ( 
.A1(n_74),
.A2(n_1),
.B(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_29),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_126),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_62),
.B1(n_60),
.B2(n_67),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_127),
.A2(n_133),
.B1(n_139),
.B2(n_82),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_91),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_128),
.Y(n_149)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_75),
.Y(n_129)
);

INVx5_ASAP7_75t_SL g156 ( 
.A(n_129),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_105),
.Y(n_130)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_130),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_75),
.B(n_29),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_131),
.B(n_134),
.Y(n_160)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_132),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_84),
.A2(n_66),
.B1(n_50),
.B2(n_63),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_70),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_64),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_2),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_136),
.B(n_140),
.Y(n_147)
);

CKINVDCx9p33_ASAP7_75t_R g137 ( 
.A(n_96),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_137),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_89),
.B(n_3),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_92),
.C(n_85),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_47),
.B1(n_5),
.B2(n_6),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_90),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_141),
.A2(n_151),
.B1(n_162),
.B2(n_127),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_143),
.B(n_148),
.Y(n_192)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_4),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g188 ( 
.A(n_145),
.B(n_124),
.C(n_122),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_138),
.B(n_99),
.C(n_93),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_88),
.B1(n_92),
.B2(n_93),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_107),
.B(n_94),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_94),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_90),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_129),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_117),
.A2(n_88),
.B1(n_92),
.B2(n_103),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_165),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_97),
.B(n_85),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_166),
.A2(n_117),
.B(n_128),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g203 ( 
.A1(n_172),
.A2(n_189),
.B1(n_191),
.B2(n_194),
.Y(n_203)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_155),
.Y(n_173)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_173),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_108),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_174),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_108),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_175),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_176),
.B(n_178),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_177),
.A2(n_165),
.B(n_149),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_126),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_152),
.Y(n_179)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_183),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_130),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_181),
.Y(n_220)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_182),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_147),
.B(n_132),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_148),
.B(n_114),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_160),
.B(n_105),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_186),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_157),
.A2(n_113),
.B1(n_82),
.B2(n_118),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_196),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_166),
.A2(n_116),
.B1(n_110),
.B2(n_9),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_143),
.B(n_5),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_190),
.B(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_157),
.B(n_7),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_141),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_11),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_195),
.B(n_154),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_156),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_170),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_170),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_159),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_205),
.Y(n_230)
);

AND2x2_ASAP7_75t_SL g202 ( 
.A(n_192),
.B(n_184),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_171),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_179),
.B(n_169),
.C(n_146),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_182),
.B(n_190),
.C(n_173),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_208),
.B(n_214),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_213),
.B(n_197),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_145),
.A3(n_169),
.B1(n_144),
.B2(n_168),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_180),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_177),
.A2(n_149),
.B(n_154),
.Y(n_217)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_221),
.B(n_163),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_193),
.A2(n_168),
.B(n_142),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_209),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_223),
.Y(n_251)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_209),
.Y(n_223)
);

NAND4xp25_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_142),
.C(n_176),
.D(n_183),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_224),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_201),
.A2(n_172),
.B1(n_194),
.B2(n_195),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_225),
.A2(n_226),
.B1(n_232),
.B2(n_218),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_216),
.B1(n_201),
.B2(n_219),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_229),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_228),
.B(n_238),
.Y(n_242)
);

AOI21xp33_ASAP7_75t_L g229 ( 
.A1(n_207),
.A2(n_178),
.B(n_198),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_237),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_210),
.B(n_191),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g243 ( 
.A(n_233),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_235),
.A2(n_240),
.B1(n_217),
.B2(n_202),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_158),
.Y(n_236)
);

INVxp33_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx11_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_211),
.B(n_163),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_158),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_239),
.B(n_205),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_241),
.A2(n_244),
.B1(n_247),
.B2(n_249),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_202),
.B1(n_215),
.B2(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_215),
.B1(n_207),
.B2(n_212),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_222),
.A2(n_208),
.B1(n_221),
.B2(n_203),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_252),
.A2(n_240),
.B1(n_227),
.B2(n_228),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_199),
.C(n_214),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_254),
.B(n_237),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_251),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_258),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_249),
.B(n_220),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_263),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_235),
.B(n_231),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_254),
.B(n_230),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_260),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_234),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_262),
.B(n_242),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_232),
.C(n_223),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_265),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_247),
.A2(n_225),
.B1(n_226),
.B2(n_233),
.Y(n_265)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_251),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_266),
.A2(n_253),
.B(n_243),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_241),
.C(n_244),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_273),
.B(n_274),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_242),
.C(n_252),
.Y(n_274)
);

NAND3xp33_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_236),
.C(n_224),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_275),
.A2(n_250),
.B(n_266),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_267),
.A2(n_268),
.B(n_269),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_276),
.A2(n_274),
.B(n_257),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_277),
.B(n_282),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_272),
.B(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_278),
.B(n_280),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_261),
.Y(n_280)
);

NOR2x1_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_264),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_284),
.A2(n_282),
.B(n_278),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_281),
.B(n_265),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_287),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_279),
.B(n_250),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.C(n_286),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_283),
.A2(n_280),
.B(n_258),
.Y(n_289)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_290),
.A2(n_286),
.A3(n_239),
.B1(n_218),
.B2(n_200),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_291),
.Y(n_293)
);

AOI21xp33_ASAP7_75t_L g294 ( 
.A1(n_293),
.A2(n_292),
.B(n_161),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g295 ( 
.A1(n_294),
.A2(n_161),
.A3(n_200),
.B1(n_163),
.B2(n_13),
.C(n_15),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_295),
.B(n_15),
.Y(n_296)
);


endmodule