module fake_netlist_1_6454_n_12 (n_1, n_2, n_0, n_12);
input n_1;
input n_2;
input n_0;
output n_12;
wire n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx3_ASAP7_75t_L g3 ( .A(n_2), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_0), .B(n_1), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
INVx1_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
INVxp67_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
BUFx2_ASAP7_75t_L g8 ( .A(n_5), .Y(n_8) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_7), .B(n_6), .Y(n_9) );
OAI211xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_4), .B(n_8), .C(n_6), .Y(n_10) );
OAI22x1_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_8), .B1(n_1), .B2(n_0), .Y(n_11) );
AO221x1_ASAP7_75t_L g12 ( .A1(n_11), .A2(n_2), .B1(n_3), .B2(n_5), .C(n_8), .Y(n_12) );
endmodule