module real_jpeg_33502_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_682, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_682;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_643;
wire n_656;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_679;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_578;
wire n_328;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_611;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_633;
wire n_497;
wire n_638;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_323;
wire n_176;
wire n_166;
wire n_215;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_594;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_572;
wire n_155;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_642;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_318;
wire n_537;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_534;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_313;
wire n_268;
wire n_42;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_641;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_660;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_625;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g243 ( 
.A(n_0),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_0),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g378 ( 
.A(n_0),
.Y(n_378)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_0),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_1),
.A2(n_312),
.B1(n_313),
.B2(n_315),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_1),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_1),
.A2(n_312),
.B1(n_368),
.B2(n_370),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_1),
.A2(n_312),
.B1(n_510),
.B2(n_514),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_1),
.A2(n_312),
.B1(n_578),
.B2(n_580),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_2),
.Y(n_94)
);

OAI22x1_ASAP7_75t_L g227 ( 
.A1(n_2),
.A2(n_94),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_2),
.A2(n_94),
.B1(n_286),
.B2(n_291),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_2),
.A2(n_94),
.B1(n_385),
.B2(n_389),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_3),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_4),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_4),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_4),
.A2(n_66),
.B1(n_125),
.B2(n_129),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_4),
.A2(n_66),
.B1(n_147),
.B2(n_151),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_4),
.A2(n_66),
.B1(n_249),
.B2(n_252),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g336 ( 
.A1(n_5),
.A2(n_96),
.B1(n_337),
.B2(n_340),
.Y(n_336)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_5),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_5),
.A2(n_340),
.B1(n_419),
.B2(n_421),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g569 ( 
.A1(n_5),
.A2(n_340),
.B1(n_570),
.B2(n_572),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_SL g640 ( 
.A1(n_5),
.A2(n_340),
.B1(n_641),
.B2(n_644),
.Y(n_640)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_6),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_7),
.A2(n_55),
.B1(n_82),
.B2(n_88),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_7),
.A2(n_88),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_7),
.A2(n_88),
.B1(n_255),
.B2(n_259),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_7),
.A2(n_88),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_8),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_8),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_9),
.Y(n_142)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_9),
.Y(n_159)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_10),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_10),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_10),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_11),
.A2(n_360),
.B1(n_363),
.B2(n_366),
.Y(n_359)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_11),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_11),
.A2(n_333),
.B1(n_337),
.B2(n_366),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_11),
.A2(n_366),
.B1(n_550),
.B2(n_553),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_SL g628 ( 
.A1(n_11),
.A2(n_366),
.B1(n_629),
.B2(n_632),
.Y(n_628)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_12),
.Y(n_104)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_12),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_21),
.B(n_679),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g679 ( 
.A(n_13),
.B(n_680),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g262 ( 
.A1(n_14),
.A2(n_263),
.B1(n_267),
.B2(n_268),
.Y(n_262)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_14),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_L g350 ( 
.A1(n_14),
.A2(n_267),
.B1(n_351),
.B2(n_354),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_14),
.A2(n_267),
.B1(n_451),
.B2(n_456),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_SL g533 ( 
.A1(n_14),
.A2(n_267),
.B1(n_304),
.B2(n_534),
.Y(n_533)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_15),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_15),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_15),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_15),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_16),
.A2(n_190),
.B1(n_191),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_16),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_16),
.A2(n_190),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g426 ( 
.A1(n_16),
.A2(n_190),
.B1(n_427),
.B2(n_429),
.Y(n_426)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_17),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_17),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_18),
.A2(n_50),
.B1(n_54),
.B2(n_59),
.Y(n_49)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_18),
.A2(n_59),
.B1(n_167),
.B2(n_170),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_18),
.A2(n_59),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_18),
.A2(n_59),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_19),
.A2(n_332),
.B(n_335),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_19),
.B(n_334),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g439 ( 
.A(n_19),
.Y(n_439)
);

OAI32xp33_ASAP7_75t_L g518 ( 
.A1(n_19),
.A2(n_162),
.A3(n_519),
.B1(n_520),
.B2(n_524),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g557 ( 
.A1(n_19),
.A2(n_439),
.B1(n_558),
.B2(n_559),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_19),
.B(n_138),
.Y(n_575)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_19),
.A2(n_245),
.B1(n_640),
.B2(n_649),
.Y(n_648)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_71),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_69),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.Y(n_23)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_24),
.Y(n_70)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_24),
.B(n_74),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_24),
.B(n_74),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_49),
.B1(n_60),
.B2(n_61),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_25),
.A2(n_60),
.B(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_25),
.A2(n_49),
.B1(n_60),
.B2(n_81),
.Y(n_172)
);

OAI22x1_ASAP7_75t_L g309 ( 
.A1(n_25),
.A2(n_60),
.B1(n_310),
.B2(n_311),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_25),
.A2(n_60),
.B1(n_331),
.B2(n_336),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_25),
.A2(n_60),
.B1(n_311),
.B2(n_447),
.Y(n_471)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_26),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_26),
.A2(n_79),
.B1(n_189),
.B2(n_262),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_38),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_27)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_28),
.Y(n_324)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_29),
.Y(n_412)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_30),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_30),
.Y(n_322)
);

BUFx5_ASAP7_75t_L g423 ( 
.A(n_30),
.Y(n_423)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_31),
.Y(n_403)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_36),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g163 ( 
.A(n_37),
.Y(n_163)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_37),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_37),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_40),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_41),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_41),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_41),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_41),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_48),
.Y(n_53)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_57),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_60),
.B(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_65),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_325),
.B(n_672),
.Y(n_71)
);

NAND3xp33_ASAP7_75t_SL g72 ( 
.A(n_73),
.B(n_176),
.C(n_203),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_73),
.A2(n_673),
.B(n_678),
.Y(n_672)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_172),
.C(n_173),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_75),
.A2(n_76),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_97),
.C(n_134),
.Y(n_76)
);

INVxp67_ASAP7_75t_SL g77 ( 
.A(n_78),
.Y(n_77)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_78),
.B(n_184),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_89),
.B2(n_90),
.Y(n_78)
);

AO22x1_ASAP7_75t_L g187 ( 
.A1(n_79),
.A2(n_90),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

AOI22x1_ASAP7_75t_L g445 ( 
.A1(n_79),
.A2(n_188),
.B1(n_446),
.B2(n_448),
.Y(n_445)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_85),
.Y(n_192)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_98),
.B(n_186),
.C(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_99),
.A2(n_135),
.B1(n_136),
.B2(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_99),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_99),
.A2(n_185),
.B1(n_198),
.B2(n_210),
.Y(n_209)
);

AO21x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_123),
.B(n_124),
.Y(n_99)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_100),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_100),
.A2(n_123),
.B1(n_218),
.B2(n_254),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g284 ( 
.A1(n_100),
.A2(n_123),
.B1(n_254),
.B2(n_285),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_100),
.A2(n_123),
.B1(n_343),
.B2(n_350),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_100),
.A2(n_123),
.B1(n_285),
.B2(n_343),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g507 ( 
.A1(n_100),
.A2(n_123),
.B1(n_350),
.B2(n_508),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_L g567 ( 
.A1(n_100),
.A2(n_123),
.B1(n_549),
.B2(n_568),
.Y(n_567)
);

AO21x2_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_109),
.B(n_114),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_105),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_104),
.Y(n_116)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_107),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g111 ( 
.A(n_108),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_108),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_109),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_111),
.Y(n_346)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_111),
.Y(n_515)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_113),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

OAI22x1_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_117),
.B1(n_120),
.B2(n_122),
.Y(n_114)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_117),
.Y(n_252)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_119),
.Y(n_251)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_119),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_119),
.Y(n_608)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_120),
.Y(n_246)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_120),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g659 ( 
.A(n_120),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_121),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_121),
.Y(n_537)
);

INVx1_ASAP7_75t_SL g214 ( 
.A(n_123),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g646 ( 
.A(n_123),
.B(n_439),
.Y(n_646)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_124),
.Y(n_215)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_127),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_128),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_128),
.Y(n_349)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_133),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_133),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_133),
.Y(n_353)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_133),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_133),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

OA22x2_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_146),
.B1(n_155),
.B2(n_166),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_137),
.A2(n_155),
.B1(n_166),
.B2(n_199),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_137),
.A2(n_155),
.B1(n_359),
.B2(n_367),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g417 ( 
.A1(n_137),
.A2(n_155),
.B1(n_359),
.B2(n_418),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_137),
.A2(n_155),
.B1(n_367),
.B2(n_450),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_137),
.A2(n_155),
.B1(n_319),
.B2(n_450),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_137),
.A2(n_155),
.B1(n_418),
.B2(n_557),
.Y(n_556)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_138),
.A2(n_174),
.B(n_175),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_138),
.A2(n_174),
.B1(n_200),
.B2(n_227),
.Y(n_226)
);

AOI22x1_ASAP7_75t_L g317 ( 
.A1(n_138),
.A2(n_174),
.B1(n_227),
.B2(n_318),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AO21x2_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_156),
.B(n_162),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_142),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_144),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx3_ASAP7_75t_SL g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_149),
.Y(n_362)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_149),
.Y(n_369)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_150),
.Y(n_420)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_151),
.Y(n_519)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

NAND2xp33_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_160),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_163),
.Y(n_171)
);

INVx4_ASAP7_75t_L g558 ( 
.A(n_163),
.Y(n_558)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_169),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_172),
.B(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g673 ( 
.A1(n_177),
.A2(n_674),
.B(n_677),
.Y(n_673)
);

NOR2x1_ASAP7_75t_R g177 ( 
.A(n_178),
.B(n_181),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_178),
.B(n_181),
.Y(n_677)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_186),
.C(n_196),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_183),
.B(n_186),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_190),
.A2(n_344),
.B(n_347),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_190),
.B(n_348),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_196),
.B(n_270),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_198),
.Y(n_210)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_271),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_205),
.A2(n_675),
.B(n_676),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_269),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_206),
.B(n_269),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_211),
.C(n_236),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_208),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_212),
.B(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_212),
.A2(n_213),
.B(n_226),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_226),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_217),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g547 ( 
.A1(n_214),
.A2(n_216),
.B1(n_509),
.B2(n_548),
.Y(n_547)
);

AOI22x1_ASAP7_75t_SL g593 ( 
.A1(n_214),
.A2(n_216),
.B1(n_569),
.B2(n_594),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_218),
.Y(n_217)
);

INVx2_ASAP7_75t_SL g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_224),
.Y(n_602)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_225),
.Y(n_598)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_229),
.Y(n_559)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_239),
.B1(n_260),
.B2(n_682),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_238),
.B(n_278),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_253),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_261),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_239),
.B(n_253),
.Y(n_481)
);

OA21x2_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_244),
.B(n_247),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g626 ( 
.A1(n_240),
.A2(n_383),
.B1(n_627),
.B2(n_635),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx3_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_242),
.A2(n_245),
.B1(n_302),
.B2(n_380),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g639 ( 
.A1(n_242),
.A2(n_245),
.B1(n_628),
.B2(n_640),
.Y(n_639)
);

INVx5_ASAP7_75t_L g656 ( 
.A(n_242),
.Y(n_656)
);

INVx8_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_243),
.B(n_246),
.Y(n_245)
);

INVx8_ASAP7_75t_L g435 ( 
.A(n_243),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_244),
.B(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_245),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_245),
.A2(n_577),
.B1(n_584),
.B2(n_585),
.Y(n_576)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_295),
.B(n_300),
.Y(n_294)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_250),
.Y(n_381)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_251),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_258),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_262),
.Y(n_310)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_264),
.Y(n_334)
);

INVx6_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_272),
.B(n_275),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_279),
.C(n_281),
.Y(n_275)
);

HB1xp67_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_277),
.A2(n_279),
.B1(n_280),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_277),
.Y(n_493)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_282),
.B(n_492),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_308),
.C(n_316),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_283),
.B(n_483),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_294),
.Y(n_283)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_284),
.Y(n_477)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx3_ASAP7_75t_SL g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_293),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_294),
.B(n_477),
.Y(n_476)
);

INVx3_ASAP7_75t_SL g295 ( 
.A(n_296),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_299),
.Y(n_584)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_306),
.Y(n_428)
);

INVx3_ASAP7_75t_L g579 ( 
.A(n_306),
.Y(n_579)
);

BUFx6f_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx6_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_307),
.Y(n_619)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_307),
.Y(n_645)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_308),
.A2(n_309),
.B1(n_317),
.B2(n_484),
.Y(n_483)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_314),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_317),
.Y(n_484)
);

INVxp67_ASAP7_75t_SL g318 ( 
.A(n_319),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_322),
.Y(n_371)
);

INVx4_ASAP7_75t_L g455 ( 
.A(n_322),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_501),
.B(n_666),
.Y(n_325)
);

NAND4xp25_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_464),
.C(n_488),
.D(n_494),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_441),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_328),
.B(n_441),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_372),
.B(n_440),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_329),
.B(n_539),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_341),
.Y(n_329)
);

MAJx2_ASAP7_75t_L g463 ( 
.A(n_330),
.B(n_342),
.C(n_358),
.Y(n_463)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx3_ASAP7_75t_SL g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_335),
.Y(n_413)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_336),
.Y(n_448)
);

INVx11_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

BUFx12f_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_358),
.Y(n_341)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVx2_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx4_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g351 ( 
.A(n_352),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_365),
.Y(n_457)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_370),
.Y(n_397)
);

INVx4_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_415),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_373),
.B(n_415),
.Y(n_440)
);

OA21x2_ASAP7_75t_SL g373 ( 
.A1(n_374),
.A2(n_393),
.B(n_414),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_375),
.A2(n_376),
.B1(n_393),
.B2(n_394),
.Y(n_540)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_395),
.Y(n_414)
);

AO22x1_ASAP7_75t_L g376 ( 
.A1(n_377),
.A2(n_379),
.B1(n_383),
.B2(n_384),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_384),
.B1(n_426),
.B2(n_433),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_383),
.A2(n_426),
.B1(n_529),
.B2(n_533),
.Y(n_528)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_388),
.Y(n_631)
);

BUFx2_ASAP7_75t_L g634 ( 
.A(n_388),
.Y(n_634)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_388),
.Y(n_643)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

BUFx2_ASAP7_75t_SL g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_392),
.Y(n_432)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_396),
.A2(n_398),
.B1(n_404),
.B2(n_413),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_402),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g402 ( 
.A(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_405),
.B(n_409),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

BUFx2_ASAP7_75t_SL g410 ( 
.A(n_411),
.Y(n_410)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

XOR2x2_ASAP7_75t_SL g442 ( 
.A(n_414),
.B(n_443),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_414),
.B(n_445),
.C(n_458),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_415),
.A2(n_416),
.B1(n_540),
.B2(n_541),
.Y(n_539)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_417),
.B(n_424),
.C(n_436),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g505 ( 
.A(n_417),
.B(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_423),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_424),
.A2(n_425),
.B1(n_437),
.B2(n_438),
.Y(n_506)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_434),
.Y(n_433)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_435),
.Y(n_434)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_439),
.B(n_525),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_SL g594 ( 
.A1(n_439),
.A2(n_595),
.B(n_599),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_439),
.B(n_600),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_439),
.B(n_655),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_459),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_442),
.B(n_460),
.C(n_496),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_444),
.A2(n_445),
.B1(n_449),
.B2(n_458),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

XOR2xp5_ASAP7_75t_SL g460 ( 
.A(n_461),
.B(n_462),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_461),
.B(n_462),
.Y(n_469)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_463),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_479),
.Y(n_464)
);

NOR2xp67_ASAP7_75t_SL g667 ( 
.A(n_465),
.B(n_479),
.Y(n_667)
);

AOI22xp33_ASAP7_75t_SL g670 ( 
.A1(n_465),
.A2(n_479),
.B1(n_489),
.B2(n_491),
.Y(n_670)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_475),
.C(n_478),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_500),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_470),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_469),
.B(n_486),
.C(n_487),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_471),
.A2(n_472),
.B1(n_473),
.B2(n_474),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_471),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_472),
.Y(n_474)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_473),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_474),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_476),
.Y(n_500)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_478),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_485),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_481),
.B(n_485),
.C(n_490),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_482),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_489),
.B(n_491),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_497),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g668 ( 
.A(n_495),
.B(n_497),
.C(n_669),
.Y(n_668)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_499),
.Y(n_497)
);

AOI21x1_ASAP7_75t_L g501 ( 
.A1(n_502),
.A2(n_542),
.B(n_665),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_538),
.Y(n_502)
);

NOR2xp67_ASAP7_75t_SL g665 ( 
.A(n_503),
.B(n_538),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_507),
.C(n_516),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g560 ( 
.A1(n_504),
.A2(n_505),
.B1(n_561),
.B2(n_562),
.Y(n_560)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_L g562 ( 
.A1(n_507),
.A2(n_516),
.B1(n_517),
.B2(n_563),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_507),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g508 ( 
.A(n_509),
.Y(n_508)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_517),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_518),
.B(n_527),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_518),
.A2(n_527),
.B1(n_528),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_518),
.Y(n_546)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

HB1xp67_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_523),
.Y(n_554)
);

INVx4_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_532),
.Y(n_531)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_532),
.Y(n_652)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_533),
.Y(n_585)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_540),
.Y(n_541)
);

OAI21x1_ASAP7_75t_L g542 ( 
.A1(n_543),
.A2(n_564),
.B(n_664),
.Y(n_542)
);

NOR2xp67_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_560),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_544),
.B(n_560),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_545),
.B(n_547),
.C(n_555),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_545),
.B(n_587),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_547),
.A2(n_555),
.B1(n_556),
.B2(n_588),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_547),
.Y(n_588)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_SL g550 ( 
.A(n_551),
.Y(n_550)
);

BUFx2_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_562),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g564 ( 
.A1(n_565),
.A2(n_589),
.B(n_663),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_566),
.B(n_586),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_566),
.B(n_586),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_567),
.B(n_574),
.C(n_576),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_567),
.A2(n_574),
.B1(n_575),
.B2(n_623),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_567),
.Y(n_623)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_569),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_571),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_L g621 ( 
.A(n_576),
.B(n_622),
.Y(n_621)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_577),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_582),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_583),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_590),
.A2(n_624),
.B(n_662),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_591),
.B(n_621),
.Y(n_590)
);

OR2x2_ASAP7_75t_L g662 ( 
.A(n_591),
.B(n_621),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_592),
.B(n_603),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_592),
.A2(n_593),
.B1(n_603),
.B2(n_604),
.Y(n_636)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx5_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_599),
.Y(n_614)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_601),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_602),
.Y(n_601)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_604),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_605),
.A2(n_614),
.B1(n_615),
.B2(n_620),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_SL g605 ( 
.A(n_606),
.B(n_609),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

INVx6_ASAP7_75t_L g607 ( 
.A(n_608),
.Y(n_607)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_610),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_611),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_612),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_617),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_618),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_619),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g624 ( 
.A1(n_625),
.A2(n_637),
.B(n_661),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_626),
.B(n_636),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_SL g661 ( 
.A(n_626),
.B(n_636),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_630),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_631),
.Y(n_630)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_633),
.Y(n_632)
);

BUFx2_ASAP7_75t_L g633 ( 
.A(n_634),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_SL g637 ( 
.A1(n_638),
.A2(n_647),
.B(n_660),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_639),
.B(n_646),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_639),
.B(n_646),
.Y(n_660)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_642),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_643),
.Y(n_642)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_645),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_648),
.B(n_653),
.Y(n_647)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_650),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_651),
.Y(n_650)
);

INVx2_ASAP7_75t_SL g651 ( 
.A(n_652),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_SL g653 ( 
.A(n_654),
.B(n_657),
.Y(n_653)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_656),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_658),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_659),
.Y(n_658)
);

O2A1O1Ixp5_ASAP7_75t_L g666 ( 
.A1(n_667),
.A2(n_668),
.B(n_670),
.C(n_671),
.Y(n_666)
);


endmodule