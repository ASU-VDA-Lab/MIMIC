module real_jpeg_6160_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_519;
wire n_205;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_0),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_0),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_0),
.B(n_196),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_0),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_0),
.B(n_229),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_0),
.B(n_270),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_1),
.Y(n_171)
);

INVx8_ASAP7_75t_L g194 ( 
.A(n_1),
.Y(n_194)
);

BUFx5_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g379 ( 
.A(n_1),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_2),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_2),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g178 ( 
.A(n_2),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_2),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_3),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_3),
.B(n_115),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_3),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_3),
.B(n_209),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_3),
.B(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_3),
.B(n_213),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_3),
.B(n_298),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_3),
.B(n_433),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_4),
.B(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_4),
.B(n_176),
.Y(n_175)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_4),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_4),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_4),
.B(n_325),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_4),
.B(n_349),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_4),
.B(n_223),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g549 ( 
.A(n_5),
.Y(n_549)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_6),
.Y(n_64)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_6),
.Y(n_91)
);

BUFx5_ASAP7_75t_L g415 ( 
.A(n_6),
.Y(n_415)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_8),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_8),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_8),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_8),
.B(n_105),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_8),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_8),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_8),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_8),
.B(n_232),
.Y(n_231)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_9),
.Y(n_124)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_9),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_9),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g364 ( 
.A(n_9),
.Y(n_364)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_10),
.Y(n_75)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_11),
.Y(n_191)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_11),
.Y(n_214)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_12),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_13),
.B(n_102),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_13),
.B(n_89),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_13),
.B(n_316),
.Y(n_315)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_13),
.B(n_340),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_13),
.B(n_355),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_13),
.B(n_397),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_13),
.B(n_409),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_14),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_14),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_14),
.B(n_56),
.Y(n_55)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_14),
.B(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_14),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_14),
.B(n_171),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_14),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_15),
.B(n_62),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_15),
.B(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_15),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_15),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_15),
.B(n_334),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_15),
.B(n_364),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g389 ( 
.A(n_15),
.B(n_390),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_15),
.B(n_421),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_16),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_16),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_16),
.B(n_155),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_16),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_16),
.B(n_62),
.Y(n_226)
);

AND2x2_ASAP7_75t_SL g290 ( 
.A(n_16),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_16),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_16),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_17),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_17),
.B(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g243 ( 
.A(n_17),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_17),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_17),
.B(n_295),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_17),
.B(n_325),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_17),
.B(n_382),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_17),
.B(n_423),
.Y(n_422)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_19),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_19),
.B(n_196),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_19),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_19),
.B(n_72),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_19),
.B(n_361),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_19),
.B(n_394),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_19),
.B(n_413),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_24),
.B(n_547),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_22),
.Y(n_548)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

O2A1O1Ixp33_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_44),
.B(n_80),
.C(n_546),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_51),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_27),
.B(n_51),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_42),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_34),
.C(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_29),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_29),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_29),
.A2(n_34),
.B1(n_43),
.B2(n_59),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_30),
.B(n_33),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_32),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_34),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_34),
.B(n_55),
.C(n_61),
.Y(n_77)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_36),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_36),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_37),
.Y(n_180)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_37),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_37),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g78 ( 
.A(n_38),
.B(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_41),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_76),
.C(n_78),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_65),
.C(n_66),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_53),
.B(n_132),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_61),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_55),
.A2(n_60),
.B1(n_71),
.B2(n_125),
.Y(n_129)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_56),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_58),
.Y(n_362)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_58),
.Y(n_399)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_58),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_67),
.C(n_71),
.Y(n_66)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_63),
.B(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_64),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_66),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_67),
.A2(n_68),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_71),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_71),
.A2(n_118),
.B1(n_119),
.B2(n_125),
.Y(n_515)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_73),
.Y(n_145)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_75),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_75),
.Y(n_296)
);

BUFx3_ASAP7_75t_L g358 ( 
.A(n_75),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g391 ( 
.A(n_75),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

AO21x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_136),
.B(n_545),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_133),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_82),
.B(n_133),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_130),
.C(n_131),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g540 ( 
.A1(n_83),
.A2(n_84),
.B1(n_541),
.B2(n_542),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_113),
.C(n_126),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_85),
.A2(n_86),
.B1(n_519),
.B2(n_521),
.Y(n_518)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_98),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_92),
.C(n_98),
.Y(n_130)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_110),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_99),
.B(n_509),
.Y(n_508)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx8_ASAP7_75t_L g247 ( 
.A(n_102),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_103),
.A2(n_104),
.B1(n_110),
.B2(n_111),
.Y(n_509)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_108),
.Y(n_148)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_113),
.A2(n_126),
.B1(n_127),
.B2(n_520),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_113),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_125),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g514 ( 
.A(n_114),
.B(n_515),
.Y(n_514)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_118),
.A2(n_119),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_119),
.B(n_208),
.C(n_212),
.Y(n_516)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_124),
.Y(n_221)
);

BUFx5_ASAP7_75t_L g424 ( 
.A(n_124),
.Y(n_424)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g542 ( 
.A(n_130),
.B(n_131),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_539),
.B(n_544),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_502),
.B(n_536),
.Y(n_137)
);

OAI21x1_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_304),
.B(n_501),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_255),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_140),
.B(n_255),
.Y(n_501)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_205),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_141),
.B(n_206),
.C(n_236),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_173),
.C(n_184),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_142),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_151),
.C(n_160),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_143),
.B(n_487),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_144),
.B(n_147),
.C(n_149),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.Y(n_146)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_148),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g487 ( 
.A1(n_151),
.A2(n_152),
.B1(n_160),
.B2(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_154),
.C(n_156),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_153),
.B(n_156),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_154),
.B(n_477),
.Y(n_476)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx5_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_160),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_161),
.B(n_165),
.C(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_169),
.B1(n_170),
.B2(n_172),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_165),
.Y(n_172)
);

INVx8_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_169),
.B(n_212),
.C(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_169),
.A2(n_170),
.B1(n_212),
.B2(n_215),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_173),
.B(n_184),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_183),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_179),
.B1(n_181),
.B2(n_182),
.Y(n_174)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_175),
.Y(n_181)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_179),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_179),
.B(n_181),
.C(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_179),
.A2(n_182),
.B1(n_245),
.B2(n_248),
.Y(n_244)
);

INVx6_ASAP7_75t_L g395 ( 
.A(n_180),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_182),
.B(n_241),
.C(n_248),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_183),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_195),
.C(n_200),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_185),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_187),
.C(n_192),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_186),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_188),
.B(n_192),
.Y(n_267)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_191),
.Y(n_382)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_194),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_194),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_195),
.B(n_200),
.Y(n_284)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_199),
.Y(n_292)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_204),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_204),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_236),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_216),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_207),
.B(n_217),
.C(n_235),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_211),
.Y(n_207)
);

INVx4_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_212),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_214),
.Y(n_317)
);

BUFx8_ASAP7_75t_L g334 ( 
.A(n_214),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_225),
.B1(n_234),
.B2(n_235),
.Y(n_216)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_217),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.C(n_222),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_218),
.B(n_222),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_221),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_226),
.B(n_228),
.C(n_231),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_231),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_249),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_238),
.B(n_240),
.C(n_249),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_242),
.B(n_251),
.Y(n_250)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

INVx8_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.C(n_253),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_253),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_259),
.C(n_262),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_257),
.B(n_260),
.Y(n_497)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_262),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_282),
.C(n_285),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_264),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_274),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_265),
.A2(n_266),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_268),
.A2(n_269),
.B(n_271),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_268),
.B(n_274),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g445 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.Y(n_445)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_279),
.B(n_445),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_281),
.B(n_375),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g490 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_285),
.Y(n_491)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_297),
.C(n_301),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_287),
.B(n_479),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_293),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_288),
.B(n_457),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g457 ( 
.A1(n_290),
.A2(n_293),
.B1(n_294),
.B2(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_290),
.Y(n_458)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx5_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_297),
.B(n_301),
.Y(n_479)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_300),
.Y(n_340)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_495),
.B(n_500),
.Y(n_304)
);

OAI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_482),
.B(n_494),
.Y(n_305)
);

AOI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_464),
.B(n_481),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_438),
.B(n_463),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_403),
.B(n_437),
.Y(n_308)
);

OAI21x1_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_367),
.B(n_402),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_344),
.B(n_366),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_328),
.B(n_343),
.Y(n_311)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_323),
.B(n_327),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_314),
.B(n_322),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_322),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_324),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_315),
.B(n_318),
.Y(n_329)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_317),
.Y(n_431)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_329),
.B(n_330),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_331),
.A2(n_332),
.B1(n_336),
.B2(n_337),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_331),
.B(n_339),
.C(n_341),
.Y(n_365)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_335),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_333),
.B(n_335),
.Y(n_352)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_341),
.B2(n_342),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_345),
.B(n_365),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_365),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_353),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_352),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_347),
.B(n_352),
.C(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_351),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_351),
.Y(n_372)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_353),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_359),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_354),
.B(n_386),
.C(n_387),
.Y(n_385)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_363),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_360),
.Y(n_386)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_363),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_368),
.B(n_370),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_384),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_371),
.B(n_385),
.C(n_388),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_372),
.B(n_374),
.C(n_377),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_377),
.Y(n_373)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_378),
.A2(n_380),
.B1(n_381),
.B2(n_383),
.Y(n_377)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_378),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_380),
.B(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_392),
.Y(n_388)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_389),
.B(n_396),
.C(n_400),
.Y(n_435)
);

INVx5_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_396),
.B1(n_400),
.B2(n_401),
.Y(n_392)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

INVx5_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g401 ( 
.A(n_396),
.Y(n_401)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_404),
.B(n_436),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_404),
.B(n_436),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_405),
.B(n_418),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_417),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_406),
.B(n_417),
.C(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_416),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_412),
.Y(n_407)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_408),
.Y(n_452)
);

INVx5_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_412),
.Y(n_453)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_416),
.B(n_452),
.C(n_453),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_418),
.Y(n_462)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_419),
.B(n_426),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_419),
.B(n_428),
.C(n_434),
.Y(n_441)
);

BUFx24_ASAP7_75t_SL g550 ( 
.A(n_419),
.Y(n_550)
);

FAx1_ASAP7_75t_SL g419 ( 
.A(n_420),
.B(n_422),
.CI(n_425),
.CON(n_419),
.SN(n_419)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_420),
.B(n_422),
.C(n_425),
.Y(n_449)
);

INVx8_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_428),
.B1(n_434),
.B2(n_435),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_432),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_429),
.B(n_432),
.Y(n_448)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_461),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_439),
.B(n_461),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_440),
.B(n_450),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_442),
.C(n_450),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_444),
.B1(n_446),
.B2(n_447),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_443),
.B(n_473),
.C(n_474),
.Y(n_472)
);

INVx1_ASAP7_75t_SL g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_448),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_449),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_451),
.B(n_454),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_451),
.B(n_455),
.C(n_460),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_455),
.A2(n_456),
.B1(n_459),
.B2(n_460),
.Y(n_454)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_455),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_456),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_480),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_465),
.B(n_480),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_466),
.B(n_471),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_470),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_470),
.C(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_471),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g471 ( 
.A(n_472),
.B(n_475),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_472),
.B(n_476),
.C(n_478),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_478),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g482 ( 
.A(n_483),
.B(n_492),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_483),
.B(n_492),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_485),
.Y(n_483)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_484),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_489),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_486),
.B(n_489),
.C(n_499),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_496),
.B(n_498),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_496),
.B(n_498),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_503),
.B(n_531),
.Y(n_502)
);

OAI21xp33_ASAP7_75t_L g536 ( 
.A1(n_503),
.A2(n_537),
.B(n_538),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.B(n_523),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_504),
.B(n_523),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_L g504 ( 
.A1(n_505),
.A2(n_506),
.B1(n_512),
.B2(n_522),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_505),
.B(n_513),
.C(n_518),
.Y(n_543)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.C(n_510),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_SL g525 ( 
.A(n_507),
.B(n_526),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g526 ( 
.A1(n_508),
.A2(n_510),
.B1(n_511),
.B2(n_527),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_508),
.Y(n_527)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_513),
.B(n_518),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_516),
.C(n_517),
.Y(n_513)
);

XOR2xp5_ASAP7_75t_L g528 ( 
.A(n_514),
.B(n_529),
.Y(n_528)
);

XNOR2xp5_ASAP7_75t_L g529 ( 
.A(n_516),
.B(n_517),
.Y(n_529)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_519),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_528),
.C(n_530),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g533 ( 
.A1(n_524),
.A2(n_525),
.B1(n_528),
.B2(n_534),
.Y(n_533)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_525),
.Y(n_524)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_528),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_530),
.B(n_533),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_532),
.B(n_535),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_532),
.B(n_535),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_540),
.B(n_543),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_540),
.B(n_543),
.Y(n_544)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_542),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_549),
.Y(n_547)
);


endmodule