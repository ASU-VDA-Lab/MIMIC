module fake_jpeg_1146_n_100 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_100);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_SL g12 ( 
.A(n_2),
.B(n_1),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

INVx5_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_2),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_28),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_12),
.B(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_12),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_18),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_4),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OA22x2_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_14),
.B1(n_18),
.B2(n_21),
.Y(n_39)
);

OA21x2_ASAP7_75t_L g59 ( 
.A1(n_39),
.A2(n_41),
.B(n_47),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_13),
.B(n_19),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_45),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_20),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_27),
.A2(n_20),
.B(n_19),
.C(n_17),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_31),
.B(n_11),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_40),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_49),
.A2(n_52),
.B1(n_54),
.B2(n_39),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_40),
.B(n_29),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_46),
.B(n_38),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_51),
.B(n_53),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_41),
.A2(n_29),
.B1(n_14),
.B2(n_15),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_17),
.B1(n_15),
.B2(n_29),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_0),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_60),
.Y(n_66)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_58),
.B(n_47),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_63),
.A2(n_52),
.B1(n_49),
.B2(n_59),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_56),
.B(n_57),
.Y(n_64)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_54),
.Y(n_65)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_65),
.Y(n_78)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_42),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_70),
.B(n_72),
.C(n_60),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_36),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_73),
.B(n_77),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_69),
.A2(n_59),
.B(n_51),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_74),
.A2(n_77),
.B(n_80),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_59),
.C(n_60),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_79),
.B(n_72),
.C(n_70),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_69),
.B(n_62),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_55),
.B1(n_36),
.B2(n_42),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_82),
.B(n_84),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_76),
.C(n_79),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_71),
.C(n_67),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_90),
.B(n_53),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_86),
.A2(n_75),
.B1(n_66),
.B2(n_39),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_92),
.A2(n_94),
.B(n_89),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_35),
.B(n_18),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g97 ( 
.A1(n_95),
.A2(n_35),
.B(n_18),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_91),
.C(n_87),
.Y(n_96)
);

MAJx2_ASAP7_75t_L g98 ( 
.A(n_96),
.B(n_35),
.C(n_5),
.Y(n_98)
);

AOI321xp33_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_98),
.A3(n_5),
.B1(n_8),
.B2(n_9),
.C(n_10),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_0),
.Y(n_100)
);


endmodule