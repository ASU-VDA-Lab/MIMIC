module fake_jpeg_9450_n_63 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_63);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_63;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_27;
wire n_55;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_44;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_4),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_5),
.B(n_7),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_25),
.A2(n_13),
.B1(n_23),
.B2(n_22),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_32),
.A2(n_38),
.B1(n_31),
.B2(n_29),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_30),
.A2(n_11),
.B1(n_19),
.B2(n_18),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_33),
.A2(n_10),
.B1(n_15),
.B2(n_16),
.Y(n_45)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_3),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_26),
.Y(n_35)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_35),
.Y(n_43)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_37),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_27),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_39),
.A2(n_45),
.B1(n_49),
.B2(n_8),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_29),
.B1(n_12),
.B2(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_41),
.A2(n_36),
.B1(n_8),
.B2(n_6),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_9),
.C(n_17),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_44),
.C(n_6),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_0),
.B(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

CKINVDCx14_ASAP7_75t_R g55 ( 
.A(n_48),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_47),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_51),
.Y(n_57)
);

OA21x2_ASAP7_75t_L g51 ( 
.A1(n_39),
.A2(n_41),
.B(n_36),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_53),
.B(n_54),
.C(n_56),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_57),
.C(n_42),
.Y(n_59)
);

AO21x1_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_52),
.B(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_60),
.A2(n_51),
.B1(n_53),
.B2(n_45),
.Y(n_61)
);

OAI321xp33_ASAP7_75t_L g62 ( 
.A1(n_61),
.A2(n_54),
.A3(n_55),
.B1(n_40),
.B2(n_43),
.C(n_24),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_62),
.B(n_40),
.Y(n_63)
);


endmodule