module fake_jpeg_16845_n_145 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_145);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

INVx8_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVxp33_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_8),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_0),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g44 ( 
.A(n_28),
.B(n_30),
.Y(n_44)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_13),
.B(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_25),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_15),
.B1(n_20),
.B2(n_13),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_45),
.B1(n_32),
.B2(n_14),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_29),
.A2(n_27),
.B1(n_18),
.B2(n_14),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g47 ( 
.A(n_36),
.B(n_20),
.Y(n_47)
);

NAND3xp33_ASAP7_75t_L g56 ( 
.A(n_47),
.B(n_36),
.C(n_31),
.Y(n_56)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_31),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_50),
.B(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_16),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_36),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_61),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_45),
.B(n_18),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_55),
.A2(n_40),
.B1(n_46),
.B2(n_25),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_62),
.B(n_64),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_34),
.B1(n_35),
.B2(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_36),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_1),
.B(n_2),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_38),
.A2(n_16),
.B1(n_22),
.B2(n_21),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_42),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_66),
.A2(n_48),
.B1(n_3),
.B2(n_4),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_34),
.B1(n_35),
.B2(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_67),
.A2(n_43),
.B1(n_48),
.B2(n_4),
.Y(n_81)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_57),
.A2(n_46),
.B(n_3),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_68),
.A2(n_75),
.B(n_1),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_69),
.A2(n_65),
.B1(n_48),
.B2(n_5),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_1),
.Y(n_75)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_59),
.B(n_23),
.CI(n_17),
.CON(n_77),
.SN(n_77)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_77),
.B(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_78),
.A2(n_85),
.B1(n_63),
.B2(n_66),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_43),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_80),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_64),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_43),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_87),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_61),
.C(n_62),
.Y(n_87)
);

AOI32xp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_49),
.A3(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_88),
.A2(n_90),
.B(n_100),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_92),
.B(n_98),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_9),
.Y(n_93)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_93),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_94),
.A2(n_84),
.B(n_85),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_10),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_96),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_99),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_70),
.A2(n_65),
.B1(n_6),
.B2(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_75),
.B(n_6),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_6),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_102),
.B(n_106),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_90),
.A2(n_73),
.B(n_68),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g117 ( 
.A1(n_103),
.A2(n_96),
.B(n_75),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_82),
.Y(n_105)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_105),
.Y(n_115)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_99),
.B(n_74),
.C(n_73),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_74),
.Y(n_108)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_89),
.B(n_79),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_112),
.B(n_89),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_110),
.B(n_87),
.C(n_91),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_113),
.B(n_77),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_118),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_102),
.B(n_107),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_111),
.B(n_83),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_119),
.B(n_120),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_79),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_81),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_121),
.A2(n_101),
.B(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_124),
.A2(n_125),
.B(n_117),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_101),
.B(n_98),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_126),
.B(n_77),
.C(n_100),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_113),
.B(n_92),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_118),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_115),
.Y(n_129)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_129),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_130),
.B(n_132),
.C(n_127),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_133),
.Y(n_137)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_133),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_135),
.B(n_136),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_134),
.A2(n_131),
.B1(n_128),
.B2(n_84),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_139),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_137),
.B(n_12),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_138),
.B(n_141),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_137),
.Y(n_145)
);


endmodule