module fake_jpeg_29427_n_98 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_98);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_98;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g10 ( 
.A(n_9),
.Y(n_10)
);

INVx4_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_9),
.B(n_0),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_5),
.B(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_24),
.B(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_0),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_30),
.Y(n_38)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_15),
.B(n_1),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_21),
.A2(n_20),
.B1(n_18),
.B2(n_11),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_22),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_15),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_26),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_19),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_27),
.B(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_23),
.B(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_52),
.B(n_54),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_SL g53 ( 
.A(n_37),
.B(n_10),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_SL g63 ( 
.A(n_53),
.B(n_40),
.C(n_10),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_46),
.A2(n_14),
.B1(n_11),
.B2(n_34),
.Y(n_55)
);

NAND3xp33_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_10),
.C(n_22),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_46),
.A2(n_25),
.B1(n_34),
.B2(n_24),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_56),
.A2(n_49),
.B1(n_35),
.B2(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_58),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_59),
.B(n_49),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_38),
.A2(n_25),
.B1(n_28),
.B2(n_32),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_60),
.A2(n_36),
.B1(n_24),
.B2(n_32),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_37),
.B(n_22),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_22),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_57),
.B1(n_39),
.B2(n_70),
.Y(n_76)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_36),
.B1(n_24),
.B2(n_23),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_39),
.B2(n_36),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_69),
.B(n_72),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_SL g71 ( 
.A(n_58),
.B(n_43),
.C(n_10),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_55),
.B(n_60),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_35),
.Y(n_72)
);

AOI322xp5_ASAP7_75t_SL g73 ( 
.A1(n_71),
.A2(n_52),
.A3(n_51),
.B1(n_53),
.B2(n_61),
.C1(n_56),
.C2(n_16),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_73),
.B(n_80),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_57),
.C(n_54),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_74),
.B(n_70),
.C(n_65),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_78),
.B(n_79),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_83),
.B(n_84),
.C(n_79),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_74),
.B(n_65),
.C(n_68),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_87),
.B(n_89),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_82),
.B(n_77),
.C(n_78),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_77),
.C(n_76),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_90),
.A2(n_86),
.B1(n_77),
.B2(n_24),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_36),
.C(n_10),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_88),
.A2(n_86),
.B(n_64),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_3),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_94),
.B(n_95),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_4),
.A3(n_7),
.B1(n_8),
.B2(n_92),
.C1(n_93),
.C2(n_95),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_7),
.Y(n_98)
);


endmodule