module fake_netlist_6_4470_n_1904 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1904);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1904;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1821;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1851;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_104),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_0),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_5),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_26),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_36),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_53),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_76),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_5),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_165),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_124),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_144),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_140),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_176),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_54),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_90),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_159),
.Y(n_202)
);

BUFx2_ASAP7_75t_R g203 ( 
.A(n_108),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_136),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_138),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_46),
.Y(n_206)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_113),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_131),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_102),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_41),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_158),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_25),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_100),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_42),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_171),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_55),
.Y(n_217)
);

BUFx10_ASAP7_75t_L g218 ( 
.A(n_32),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_147),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_26),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_93),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_59),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_57),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_55),
.Y(n_226)
);

INVxp67_ASAP7_75t_SL g227 ( 
.A(n_44),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_79),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_84),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_33),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_117),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g232 ( 
.A(n_150),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_65),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_51),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_179),
.Y(n_236)
);

BUFx8_ASAP7_75t_SL g237 ( 
.A(n_6),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_58),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_7),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_111),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_20),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_85),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_135),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_101),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_46),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_52),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_128),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_94),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_10),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_11),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_73),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_125),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_175),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_29),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_132),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_87),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_126),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_170),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_96),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_52),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_19),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_71),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_143),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_122),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_134),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_45),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_172),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_61),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_47),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_106),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_25),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_38),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_121),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_164),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_129),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_156),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_80),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_54),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_110),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_181),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_152),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_7),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_47),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_17),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_39),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_127),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_39),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_74),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_9),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_43),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_83),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_36),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_141),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_69),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_154),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_75),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_68),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_35),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_18),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_12),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_133),
.Y(n_303)
);

INVxp67_ASAP7_75t_SL g304 ( 
.A(n_168),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_37),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_49),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_66),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_130),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_28),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_4),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_70),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_162),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_86),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_64),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g316 ( 
.A(n_91),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_116),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_161),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_1),
.Y(n_319)
);

INVx2_ASAP7_75t_SL g320 ( 
.A(n_160),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_142),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_23),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_20),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_115),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_29),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_157),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_169),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_1),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_18),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_105),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_2),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_177),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_109),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_112),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_95),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_120),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_19),
.Y(n_337)
);

INVx2_ASAP7_75t_SL g338 ( 
.A(n_43),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_53),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_28),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_118),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_174),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_49),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_13),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_30),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_67),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_180),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_11),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_166),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_34),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_17),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_50),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_77),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_41),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_42),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_13),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_72),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_57),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_60),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_21),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_44),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_51),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_82),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_4),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_237),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_211),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_194),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_215),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_214),
.B(n_0),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_192),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_197),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_202),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_205),
.Y(n_375)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_204),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g377 ( 
.A(n_215),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_259),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_322),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_275),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_214),
.B(n_2),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_277),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_208),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g384 ( 
.A(n_322),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_245),
.B(n_3),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_284),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_284),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_349),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_232),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_284),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_232),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g393 ( 
.A(n_184),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_224),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_213),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_316),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_231),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_233),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_240),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_243),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_224),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_244),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_248),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_235),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_235),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_325),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_252),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_254),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_245),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_320),
.B(n_6),
.Y(n_410)
);

INVx1_ASAP7_75t_SL g411 ( 
.A(n_225),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_256),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_257),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_261),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_L g417 ( 
.A(n_338),
.B(n_8),
.Y(n_417)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_285),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_265),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_329),
.Y(n_420)
);

HB1xp67_ASAP7_75t_L g421 ( 
.A(n_268),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g422 ( 
.A(n_268),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_267),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_320),
.B(n_8),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_184),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_185),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_272),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_220),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_278),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_220),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_279),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_186),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_281),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_226),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_226),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_282),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_283),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_271),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_288),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_271),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_289),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_290),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_295),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_186),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_308),
.B(n_9),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_234),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_296),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_297),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_289),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_319),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_319),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_308),
.B(n_10),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_345),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_187),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_303),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_432),
.B(n_194),
.Y(n_457)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_421),
.Y(n_458)
);

CKINVDCx6p67_ASAP7_75t_R g459 ( 
.A(n_396),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_365),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_446),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_446),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_446),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_365),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_389),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_424),
.B(n_312),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_386),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_446),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_386),
.B(n_314),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_387),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_196),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_387),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_444),
.B(n_196),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_390),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_390),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_392),
.B(n_315),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_368),
.B(n_444),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_401),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_405),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_405),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_368),
.B(n_207),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_368),
.B(n_317),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_398),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_428),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_394),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_409),
.B(n_207),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_404),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_428),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_430),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_430),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_404),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_417),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_406),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_410),
.B(n_266),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_406),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_445),
.B(n_258),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_412),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_412),
.B(n_258),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_434),
.B(n_318),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_411),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_438),
.Y(n_507)
);

INVx6_ASAP7_75t_L g508 ( 
.A(n_376),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_440),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_440),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_413),
.Y(n_512)
);

AND2x6_ASAP7_75t_L g513 ( 
.A(n_452),
.B(n_234),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_371),
.B(n_209),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_441),
.B(n_326),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_441),
.Y(n_516)
);

HB1xp67_ASAP7_75t_L g517 ( 
.A(n_417),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_413),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_420),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_449),
.Y(n_520)
);

BUFx6f_ASAP7_75t_L g521 ( 
.A(n_420),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_449),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_450),
.Y(n_523)
);

HB1xp67_ASAP7_75t_L g524 ( 
.A(n_377),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_453),
.B(n_327),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_367),
.Y(n_527)
);

INVx3_ASAP7_75t_L g528 ( 
.A(n_453),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_454),
.Y(n_529)
);

BUFx6f_ASAP7_75t_L g530 ( 
.A(n_454),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_399),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_393),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_425),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_381),
.B(n_260),
.Y(n_534)
);

AND2x4_ASAP7_75t_L g535 ( 
.A(n_435),
.B(n_332),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_460),
.Y(n_536)
);

INVx3_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_472),
.Y(n_538)
);

BUFx2_ASAP7_75t_L g539 ( 
.A(n_506),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_500),
.B(n_369),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_514),
.B(n_372),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_455),
.Y(n_542)
);

INVx3_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_460),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g545 ( 
.A(n_506),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_461),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_485),
.B(n_377),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_524),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_500),
.B(n_373),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_472),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_477),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_527),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_534),
.B(n_374),
.Y(n_553)
);

AOI22xp33_ASAP7_75t_L g554 ( 
.A1(n_502),
.A2(n_385),
.B1(n_379),
.B2(n_370),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_534),
.B(n_375),
.Y(n_555)
);

INVxp33_ASAP7_75t_L g556 ( 
.A(n_524),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_464),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_477),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_468),
.B(n_383),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_464),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_485),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_485),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_498),
.Y(n_563)
);

AO22x2_ASAP7_75t_L g564 ( 
.A1(n_502),
.A2(n_384),
.B1(n_338),
.B2(n_358),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_469),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_467),
.B(n_395),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_502),
.A2(n_379),
.B1(n_358),
.B2(n_333),
.Y(n_567)
);

INVx4_ASAP7_75t_SL g568 ( 
.A(n_513),
.Y(n_568)
);

NAND3xp33_ASAP7_75t_L g569 ( 
.A(n_532),
.B(n_400),
.C(n_397),
.Y(n_569)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_468),
.A2(n_407),
.B1(n_448),
.B2(n_447),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_477),
.Y(n_571)
);

INVx4_ASAP7_75t_L g572 ( 
.A(n_474),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_528),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_528),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_498),
.B(n_402),
.Y(n_576)
);

BUFx10_ASAP7_75t_L g577 ( 
.A(n_508),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_467),
.B(n_403),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_486),
.B(n_502),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_528),
.Y(n_580)
);

NOR2xp33_ASAP7_75t_L g581 ( 
.A(n_486),
.B(n_408),
.Y(n_581)
);

INVx6_ASAP7_75t_L g582 ( 
.A(n_508),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_484),
.Y(n_583)
);

OR2x2_ASAP7_75t_L g584 ( 
.A(n_458),
.B(n_422),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_461),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_488),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_488),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_493),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_493),
.Y(n_589)
);

AO21x2_ASAP7_75t_L g590 ( 
.A1(n_471),
.A2(n_191),
.B(n_189),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_508),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_502),
.B(n_415),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_457),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_513),
.Y(n_594)
);

INVx2_ASAP7_75t_SL g595 ( 
.A(n_517),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_474),
.Y(n_596)
);

BUFx2_ASAP7_75t_L g597 ( 
.A(n_458),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_517),
.B(n_422),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_484),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_416),
.Y(n_600)
);

OR2x6_ASAP7_75t_L g601 ( 
.A(n_508),
.B(n_451),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_478),
.B(n_423),
.Y(n_602)
);

BUFx10_ASAP7_75t_L g603 ( 
.A(n_508),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_505),
.B(n_427),
.Y(n_604)
);

INVx4_ASAP7_75t_L g605 ( 
.A(n_474),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_491),
.B(n_431),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_484),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_494),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_478),
.B(n_433),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_532),
.B(n_436),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_513),
.A2(n_333),
.B1(n_332),
.B2(n_189),
.Y(n_611)
);

AND2x6_ASAP7_75t_L g612 ( 
.A(n_457),
.B(n_191),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_505),
.B(n_437),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_484),
.Y(n_614)
);

AOI22xp5_ASAP7_75t_L g615 ( 
.A1(n_491),
.A2(n_429),
.B1(n_419),
.B2(n_442),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_491),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_494),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_528),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_533),
.B(n_439),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_528),
.Y(n_620)
);

INVx4_ASAP7_75t_L g621 ( 
.A(n_474),
.Y(n_621)
);

AND2x6_ASAP7_75t_L g622 ( 
.A(n_457),
.B(n_195),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_484),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_533),
.B(n_443),
.Y(n_624)
);

AOI22xp33_ASAP7_75t_L g625 ( 
.A1(n_513),
.A2(n_264),
.B1(n_198),
.B2(n_357),
.Y(n_625)
);

OR2x6_ASAP7_75t_L g626 ( 
.A(n_508),
.B(n_200),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_484),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_495),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_515),
.B(n_456),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_473),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_495),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_473),
.Y(n_632)
);

BUFx3_ASAP7_75t_L g633 ( 
.A(n_473),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_480),
.B(n_330),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_515),
.B(n_414),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_504),
.B(n_227),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_527),
.Y(n_637)
);

INVxp67_ASAP7_75t_SL g638 ( 
.A(n_480),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_504),
.B(n_195),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_535),
.B(n_366),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_484),
.Y(n_642)
);

INVx4_ASAP7_75t_L g643 ( 
.A(n_474),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_526),
.B(n_334),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_461),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_461),
.Y(n_646)
);

AOI22xp33_ASAP7_75t_L g647 ( 
.A1(n_513),
.A2(n_293),
.B1(n_324),
.B2(n_270),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_489),
.Y(n_648)
);

OR2x6_ASAP7_75t_L g649 ( 
.A(n_535),
.B(n_526),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_489),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_496),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_504),
.B(n_198),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_507),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_487),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_535),
.B(n_391),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_507),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_489),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_509),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_509),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_535),
.B(n_418),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_510),
.Y(n_661)
);

NOR3xp33_ASAP7_75t_L g662 ( 
.A(n_466),
.B(n_348),
.C(n_190),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_489),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_510),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_475),
.B(n_199),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_489),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_511),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_489),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_489),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_511),
.Y(n_670)
);

HB1xp67_ASAP7_75t_L g671 ( 
.A(n_466),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_516),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_516),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_499),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_535),
.B(n_378),
.Y(n_675)
);

BUFx6f_ASAP7_75t_L g676 ( 
.A(n_461),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_466),
.B(n_199),
.Y(n_677)
);

INVxp67_ASAP7_75t_SL g678 ( 
.A(n_465),
.Y(n_678)
);

INVx3_ASAP7_75t_L g679 ( 
.A(n_474),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_513),
.B(n_234),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_520),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_475),
.B(n_269),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_520),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_499),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_499),
.Y(n_685)
);

BUFx10_ASAP7_75t_L g686 ( 
.A(n_487),
.Y(n_686)
);

NAND2xp33_ASAP7_75t_L g687 ( 
.A(n_513),
.B(n_234),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_538),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_638),
.B(n_513),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_579),
.B(n_234),
.Y(n_690)
);

AO221x1_ASAP7_75t_L g691 ( 
.A1(n_564),
.A2(n_353),
.B1(n_276),
.B2(n_293),
.C(n_298),
.Y(n_691)
);

AND2x4_ASAP7_75t_L g692 ( 
.A(n_561),
.B(n_475),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_545),
.B(n_569),
.Y(n_693)
);

O2A1O1Ixp5_ASAP7_75t_L g694 ( 
.A1(n_628),
.A2(n_462),
.B(n_463),
.C(n_479),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_538),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_542),
.B(n_188),
.Y(n_696)
);

O2A1O1Ixp33_ASAP7_75t_L g697 ( 
.A1(n_616),
.A2(n_522),
.B(n_525),
.C(n_529),
.Y(n_697)
);

BUFx6f_ASAP7_75t_SL g698 ( 
.A(n_686),
.Y(n_698)
);

OR2x6_ASAP7_75t_L g699 ( 
.A(n_539),
.B(n_203),
.Y(n_699)
);

AND2x2_ASAP7_75t_SL g700 ( 
.A(n_566),
.B(n_201),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_616),
.B(n_276),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_590),
.A2(n_513),
.B1(n_299),
.B2(n_298),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_581),
.B(n_513),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_604),
.B(n_530),
.Y(n_704)
);

OAI22xp5_ASAP7_75t_SL g705 ( 
.A1(n_552),
.A2(n_380),
.B1(n_382),
.B2(n_388),
.Y(n_705)
);

O2A1O1Ixp33_ASAP7_75t_L g706 ( 
.A1(n_636),
.A2(n_522),
.B(n_529),
.C(n_525),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_561),
.Y(n_707)
);

AO21x2_ASAP7_75t_L g708 ( 
.A1(n_578),
.A2(n_304),
.B(n_216),
.Y(n_708)
);

INVxp67_ASAP7_75t_SL g709 ( 
.A(n_593),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_593),
.Y(n_710)
);

A2O1A1Ixp33_ASAP7_75t_L g711 ( 
.A1(n_553),
.A2(n_613),
.B(n_629),
.C(n_636),
.Y(n_711)
);

O2A1O1Ixp33_ASAP7_75t_L g712 ( 
.A1(n_632),
.A2(n_639),
.B(n_652),
.C(n_562),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_536),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_539),
.B(n_531),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_SL g715 ( 
.A(n_594),
.B(n_276),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_632),
.B(n_530),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_562),
.B(n_530),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_630),
.B(n_530),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_563),
.B(n_193),
.Y(n_719)
);

INVx8_ASAP7_75t_L g720 ( 
.A(n_601),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_630),
.B(n_530),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_536),
.Y(n_722)
);

A2O1A1Ixp33_ASAP7_75t_L g723 ( 
.A1(n_639),
.A2(n_270),
.B(n_307),
.C(n_299),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_633),
.B(n_201),
.Y(n_724)
);

NOR2xp67_ASAP7_75t_L g725 ( 
.A(n_570),
.B(n_615),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_597),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_633),
.B(n_540),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_594),
.B(n_276),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_549),
.B(n_530),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_594),
.B(n_606),
.Y(n_730)
);

AOI22xp5_ASAP7_75t_L g731 ( 
.A1(n_635),
.A2(n_335),
.B1(n_341),
.B2(n_346),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_594),
.B(n_276),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_563),
.B(n_531),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_600),
.B(n_530),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_628),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_SL g736 ( 
.A(n_594),
.B(n_353),
.Y(n_736)
);

NAND2xp33_ASAP7_75t_L g737 ( 
.A(n_612),
.B(n_363),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_595),
.B(n_459),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_602),
.B(n_530),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_631),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_612),
.B(n_353),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_595),
.B(n_459),
.Y(n_742)
);

INVxp67_ASAP7_75t_L g743 ( 
.A(n_597),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_609),
.B(n_490),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_634),
.B(n_490),
.Y(n_745)
);

BUFx6f_ASAP7_75t_L g746 ( 
.A(n_676),
.Y(n_746)
);

NAND3xp33_ASAP7_75t_L g747 ( 
.A(n_660),
.B(n_210),
.C(n_206),
.Y(n_747)
);

NOR3xp33_ASAP7_75t_L g748 ( 
.A(n_655),
.B(n_217),
.C(n_212),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_644),
.B(n_490),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_676),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_649),
.A2(n_264),
.B1(n_357),
.B2(n_347),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_544),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_606),
.B(n_353),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_631),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_592),
.B(n_353),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_654),
.Y(n_756)
);

NOR2xp67_ASAP7_75t_L g757 ( 
.A(n_675),
.B(n_598),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_640),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_640),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_548),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_651),
.B(n_490),
.Y(n_761)
);

NOR2xp67_ASAP7_75t_L g762 ( 
.A(n_598),
.B(n_490),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_574),
.B(n_521),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_550),
.Y(n_764)
);

INVx2_ASAP7_75t_L g765 ( 
.A(n_550),
.Y(n_765)
);

OAI22xp33_ASAP7_75t_L g766 ( 
.A1(n_649),
.A2(n_556),
.B1(n_653),
.B2(n_651),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_574),
.B(n_521),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_649),
.A2(n_555),
.B1(n_541),
.B2(n_612),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_653),
.B(n_492),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_656),
.B(n_492),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_656),
.B(n_492),
.Y(n_771)
);

INVx3_ASAP7_75t_L g772 ( 
.A(n_658),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_658),
.Y(n_773)
);

AND2x6_ASAP7_75t_L g774 ( 
.A(n_575),
.B(n_216),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_575),
.B(n_521),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_659),
.B(n_492),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_659),
.B(n_492),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_548),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_664),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_SL g780 ( 
.A1(n_654),
.A2(n_292),
.B1(n_302),
.B2(n_323),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_590),
.A2(n_253),
.B1(n_347),
.B2(n_342),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_580),
.B(n_521),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_544),
.Y(n_783)
);

AO221x1_ASAP7_75t_L g784 ( 
.A1(n_564),
.A2(n_253),
.B1(n_219),
.B2(n_221),
.C(n_223),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_664),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_580),
.B(n_521),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_649),
.A2(n_342),
.B1(n_221),
.B2(n_223),
.Y(n_787)
);

BUFx2_ASAP7_75t_L g788 ( 
.A(n_671),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_557),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_667),
.B(n_501),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_557),
.Y(n_791)
);

OAI22xp5_ASAP7_75t_L g792 ( 
.A1(n_567),
.A2(n_307),
.B1(n_228),
.B2(n_336),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_590),
.A2(n_321),
.B1(n_219),
.B2(n_336),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_667),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_670),
.B(n_501),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_670),
.Y(n_796)
);

A2O1A1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_652),
.A2(n_228),
.B(n_229),
.C(n_236),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_R g798 ( 
.A(n_552),
.B(n_459),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_681),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_681),
.Y(n_800)
);

INVx2_ASAP7_75t_SL g801 ( 
.A(n_547),
.Y(n_801)
);

INVx2_ASAP7_75t_SL g802 ( 
.A(n_547),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_560),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_683),
.B(n_501),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_560),
.Y(n_805)
);

NOR2xp33_ASAP7_75t_SL g806 ( 
.A(n_584),
.B(n_331),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_683),
.B(n_501),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_551),
.Y(n_808)
);

OR2x6_ASAP7_75t_L g809 ( 
.A(n_677),
.B(n_601),
.Y(n_809)
);

NAND3xp33_ASAP7_75t_L g810 ( 
.A(n_554),
.B(n_251),
.C(n_364),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_586),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_587),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_588),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_589),
.B(n_501),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_551),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_608),
.B(n_617),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_558),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_661),
.B(n_479),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_672),
.B(n_479),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_584),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_673),
.B(n_479),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_565),
.B(n_479),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_618),
.B(n_521),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_558),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_565),
.B(n_499),
.Y(n_825)
);

INVxp67_ASAP7_75t_L g826 ( 
.A(n_610),
.Y(n_826)
);

BUFx6f_ASAP7_75t_L g827 ( 
.A(n_676),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_601),
.B(n_218),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_573),
.B(n_499),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_573),
.B(n_499),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_571),
.Y(n_831)
);

INVxp67_ASAP7_75t_L g832 ( 
.A(n_619),
.Y(n_832)
);

NOR2xp67_ASAP7_75t_L g833 ( 
.A(n_559),
.B(n_481),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_618),
.B(n_499),
.Y(n_834)
);

AOI22xp33_ASAP7_75t_L g835 ( 
.A1(n_612),
.A2(n_249),
.B1(n_324),
.B2(n_321),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_620),
.B(n_512),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_620),
.B(n_521),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_571),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_568),
.B(n_521),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_678),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_665),
.B(n_512),
.Y(n_841)
);

INVxp67_ASAP7_75t_SL g842 ( 
.A(n_679),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_665),
.A2(n_313),
.B(n_229),
.C(n_249),
.Y(n_843)
);

BUFx6f_ASAP7_75t_SL g844 ( 
.A(n_686),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_665),
.B(n_512),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_676),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_601),
.B(n_218),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_582),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_537),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_612),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_612),
.B(n_512),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_568),
.B(n_236),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_622),
.Y(n_853)
);

AND2x6_ASAP7_75t_L g854 ( 
.A(n_583),
.B(n_313),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_L g855 ( 
.A(n_624),
.B(n_222),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_576),
.B(n_230),
.Y(n_856)
);

INVxp67_ASAP7_75t_L g857 ( 
.A(n_677),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_677),
.B(n_218),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_714),
.B(n_677),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_SL g860 ( 
.A(n_756),
.B(n_686),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_704),
.A2(n_596),
.B(n_572),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_696),
.B(n_641),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_711),
.B(n_622),
.Y(n_863)
);

AND2x2_ASAP7_75t_L g864 ( 
.A(n_801),
.B(n_662),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_713),
.Y(n_865)
);

A2O1A1Ixp33_ASAP7_75t_L g866 ( 
.A1(n_711),
.A2(n_682),
.B(n_611),
.C(n_625),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_713),
.Y(n_867)
);

AOI22xp5_ASAP7_75t_L g868 ( 
.A1(n_700),
.A2(n_622),
.B1(n_626),
.B2(n_591),
.Y(n_868)
);

INVx3_ASAP7_75t_L g869 ( 
.A(n_740),
.Y(n_869)
);

INVxp67_ASAP7_75t_L g870 ( 
.A(n_760),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_694),
.A2(n_622),
.B(n_647),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_692),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_700),
.B(n_622),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_727),
.B(n_622),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_734),
.A2(n_596),
.B(n_572),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_740),
.B(n_564),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_722),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_739),
.A2(n_596),
.B(n_572),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_696),
.B(n_637),
.Y(n_879)
);

AOI22xp5_ASAP7_75t_L g880 ( 
.A1(n_768),
.A2(n_626),
.B1(n_591),
.B2(n_582),
.Y(n_880)
);

OAI22xp5_ASAP7_75t_L g881 ( 
.A1(n_781),
.A2(n_564),
.B1(n_626),
.B2(n_362),
.Y(n_881)
);

INVxp67_ASAP7_75t_L g882 ( 
.A(n_788),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_692),
.B(n_577),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_729),
.A2(n_721),
.B(n_718),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_772),
.B(n_537),
.Y(n_885)
);

AO21x1_ASAP7_75t_L g886 ( 
.A1(n_766),
.A2(n_690),
.B(n_755),
.Y(n_886)
);

AND2x4_ASAP7_75t_L g887 ( 
.A(n_710),
.B(n_626),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_745),
.A2(n_621),
.B(n_605),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_772),
.B(n_537),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_781),
.A2(n_309),
.B1(n_355),
.B2(n_354),
.Y(n_890)
);

INVxp67_ASAP7_75t_L g891 ( 
.A(n_733),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_752),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_726),
.B(n_637),
.Y(n_893)
);

AOI21xp5_ASAP7_75t_L g894 ( 
.A1(n_841),
.A2(n_621),
.B(n_605),
.Y(n_894)
);

AOI21xp5_ASAP7_75t_L g895 ( 
.A1(n_845),
.A2(n_621),
.B(n_605),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_783),
.Y(n_896)
);

O2A1O1Ixp33_ASAP7_75t_L g897 ( 
.A1(n_701),
.A2(n_687),
.B(n_680),
.C(n_523),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_709),
.B(n_543),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_735),
.B(n_543),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_783),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_789),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_789),
.Y(n_902)
);

INVx11_ASAP7_75t_L g903 ( 
.A(n_854),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_757),
.B(n_762),
.Y(n_904)
);

HB1xp67_ASAP7_75t_L g905 ( 
.A(n_778),
.Y(n_905)
);

A2O1A1Ixp33_ASAP7_75t_L g906 ( 
.A1(n_712),
.A2(n_687),
.B(n_680),
.C(n_627),
.Y(n_906)
);

OAI22xp5_ASAP7_75t_L g907 ( 
.A1(n_793),
.A2(n_300),
.B1(n_263),
.B2(n_262),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_754),
.B(n_758),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_749),
.A2(n_643),
.B(n_676),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_791),
.Y(n_910)
);

A2O1A1Ixp33_ASAP7_75t_L g911 ( 
.A1(n_706),
.A2(n_623),
.B(n_583),
.C(n_599),
.Y(n_911)
);

NOR3xp33_ASAP7_75t_L g912 ( 
.A(n_705),
.B(n_856),
.C(n_832),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_744),
.A2(n_689),
.B(n_717),
.Y(n_913)
);

BUFx12f_ASAP7_75t_L g914 ( 
.A(n_820),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_791),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_759),
.B(n_543),
.Y(n_916)
);

BUFx2_ASAP7_75t_L g917 ( 
.A(n_743),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_773),
.B(n_546),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_716),
.A2(n_643),
.B(n_627),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_730),
.A2(n_643),
.B(n_642),
.Y(n_920)
);

BUFx6f_ASAP7_75t_L g921 ( 
.A(n_848),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_SL g922 ( 
.A(n_802),
.B(n_826),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_779),
.B(n_546),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_730),
.A2(n_623),
.B(n_642),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_803),
.Y(n_925)
);

BUFx4f_ASAP7_75t_L g926 ( 
.A(n_809),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_741),
.A2(n_599),
.B(n_607),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_803),
.Y(n_928)
);

A2O1A1Ixp33_ASAP7_75t_L g929 ( 
.A1(n_697),
.A2(n_614),
.B(n_607),
.C(n_685),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_785),
.B(n_546),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_738),
.B(n_742),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_703),
.A2(n_614),
.B(n_684),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_707),
.B(n_811),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_851),
.A2(n_685),
.B(n_684),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_842),
.A2(n_650),
.B(n_674),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_690),
.A2(n_650),
.B(n_674),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_794),
.B(n_585),
.Y(n_937)
);

A2O1A1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_855),
.A2(n_669),
.B(n_668),
.C(n_666),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_805),
.Y(n_939)
);

O2A1O1Ixp33_ASAP7_75t_L g940 ( 
.A1(n_701),
.A2(n_523),
.B(n_669),
.C(n_668),
.Y(n_940)
);

O2A1O1Ixp5_ASAP7_75t_L g941 ( 
.A1(n_755),
.A2(n_648),
.B(n_666),
.C(n_663),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_746),
.A2(n_648),
.B(n_663),
.Y(n_942)
);

O2A1O1Ixp33_ASAP7_75t_L g943 ( 
.A1(n_792),
.A2(n_523),
.B(n_657),
.C(n_483),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_805),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_855),
.A2(n_856),
.B(n_719),
.C(n_787),
.Y(n_945)
);

OR2x2_ASAP7_75t_L g946 ( 
.A(n_810),
.B(n_238),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_796),
.B(n_585),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_799),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_812),
.B(n_568),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_766),
.A2(n_591),
.B1(n_582),
.B2(n_657),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_753),
.A2(n_582),
.B1(n_591),
.B2(n_679),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_806),
.B(n_239),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_746),
.A2(n_646),
.B(n_645),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_831),
.Y(n_954)
);

INVx3_ASAP7_75t_L g955 ( 
.A(n_848),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_800),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_840),
.B(n_585),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_719),
.A2(n_679),
.B(n_646),
.C(n_645),
.Y(n_958)
);

NOR2x1_ASAP7_75t_L g959 ( 
.A(n_693),
.B(n_645),
.Y(n_959)
);

OAI21xp5_ASAP7_75t_L g960 ( 
.A1(n_793),
.A2(n_702),
.B(n_761),
.Y(n_960)
);

OAI22xp5_ASAP7_75t_L g961 ( 
.A1(n_835),
.A2(n_344),
.B1(n_242),
.B2(n_247),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_746),
.A2(n_646),
.B(n_465),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_858),
.B(n_218),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_831),
.Y(n_964)
);

O2A1O1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_723),
.A2(n_482),
.B(n_481),
.C(n_483),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_746),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_750),
.A2(n_465),
.B(n_470),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_835),
.A2(n_340),
.B1(n_339),
.B2(n_337),
.Y(n_968)
);

OAI21xp5_ASAP7_75t_L g969 ( 
.A1(n_702),
.A2(n_462),
.B(n_463),
.Y(n_969)
);

AOI21x1_ASAP7_75t_L g970 ( 
.A1(n_763),
.A2(n_463),
.B(n_462),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_747),
.B(n_857),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_769),
.B(n_568),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_699),
.Y(n_973)
);

OAI22xp5_ASAP7_75t_L g974 ( 
.A1(n_751),
.A2(n_306),
.B1(n_305),
.B2(n_301),
.Y(n_974)
);

OAI21xp33_ASAP7_75t_L g975 ( 
.A1(n_731),
.A2(n_294),
.B(n_291),
.Y(n_975)
);

OAI22xp5_ASAP7_75t_L g976 ( 
.A1(n_809),
.A2(n_287),
.B1(n_286),
.B2(n_280),
.Y(n_976)
);

NOR2xp33_ASAP7_75t_L g977 ( 
.A(n_828),
.B(n_241),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_750),
.A2(n_465),
.B(n_470),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_813),
.B(n_577),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_847),
.B(n_250),
.Y(n_980)
);

OAI21xp5_ASAP7_75t_L g981 ( 
.A1(n_770),
.A2(n_776),
.B(n_771),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_809),
.A2(n_274),
.B1(n_273),
.B2(n_255),
.Y(n_982)
);

AO21x1_ASAP7_75t_L g983 ( 
.A1(n_724),
.A2(n_482),
.B(n_497),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_777),
.B(n_790),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_833),
.B(n_577),
.Y(n_985)
);

BUFx6f_ASAP7_75t_L g986 ( 
.A(n_750),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_725),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_750),
.A2(n_465),
.B(n_470),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_753),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_795),
.B(n_512),
.Y(n_990)
);

AND2x6_ASAP7_75t_L g991 ( 
.A(n_850),
.B(n_470),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_827),
.A2(n_470),
.B(n_603),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_688),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_816),
.B(n_497),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_748),
.B(n_246),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_724),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_723),
.A2(n_359),
.B1(n_310),
.B2(n_311),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_827),
.A2(n_603),
.B(n_474),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_804),
.B(n_518),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_827),
.B(n_603),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_798),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_807),
.B(n_518),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_827),
.A2(n_476),
.B(n_503),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_846),
.A2(n_476),
.B(n_503),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_797),
.A2(n_519),
.B(n_503),
.C(n_497),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_699),
.B(n_352),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_846),
.A2(n_476),
.B(n_519),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_797),
.A2(n_356),
.B1(n_328),
.B2(n_343),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_798),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_849),
.Y(n_1010)
);

BUFx3_ASAP7_75t_L g1011 ( 
.A(n_720),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_814),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_695),
.Y(n_1013)
);

INVx4_ASAP7_75t_L g1014 ( 
.A(n_720),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_822),
.A2(n_519),
.B(n_360),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_846),
.A2(n_737),
.B(n_829),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_846),
.A2(n_476),
.B(n_512),
.Y(n_1017)
);

OR2x2_ASAP7_75t_L g1018 ( 
.A(n_780),
.B(n_350),
.Y(n_1018)
);

AOI21xp33_ASAP7_75t_L g1019 ( 
.A1(n_708),
.A2(n_825),
.B(n_830),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_818),
.A2(n_819),
.B(n_821),
.Y(n_1020)
);

INVxp67_ASAP7_75t_SL g1021 ( 
.A(n_849),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_834),
.A2(n_476),
.B(n_512),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_836),
.A2(n_476),
.B(n_518),
.Y(n_1023)
);

OAI21x1_ASAP7_75t_L g1024 ( 
.A1(n_763),
.A2(n_63),
.B(n_62),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_708),
.B(n_518),
.Y(n_1025)
);

CKINVDCx10_ASAP7_75t_R g1026 ( 
.A(n_698),
.Y(n_1026)
);

INVx3_ASAP7_75t_L g1027 ( 
.A(n_764),
.Y(n_1027)
);

INVxp67_ASAP7_75t_L g1028 ( 
.A(n_698),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_720),
.B(n_853),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_SL g1030 ( 
.A(n_765),
.B(n_269),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_808),
.Y(n_1031)
);

OA22x2_ASAP7_75t_L g1032 ( 
.A1(n_784),
.A2(n_691),
.B1(n_361),
.B2(n_351),
.Y(n_1032)
);

AND2x4_ASAP7_75t_L g1033 ( 
.A(n_852),
.B(n_123),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_843),
.B(n_246),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_839),
.A2(n_476),
.B(n_518),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_815),
.B(n_518),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_843),
.B(n_246),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_852),
.A2(n_269),
.B(n_246),
.C(n_15),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_839),
.A2(n_137),
.B(n_182),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_767),
.A2(n_119),
.B(n_163),
.Y(n_1040)
);

NOR2x1_ASAP7_75t_R g1041 ( 
.A(n_844),
.B(n_269),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_817),
.B(n_12),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_824),
.B(n_14),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_838),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_774),
.B(n_14),
.Y(n_1045)
);

NAND2xp33_ASAP7_75t_L g1046 ( 
.A(n_774),
.B(n_155),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_767),
.A2(n_153),
.B(n_151),
.Y(n_1047)
);

OAI21xp33_ASAP7_75t_L g1048 ( 
.A1(n_862),
.A2(n_952),
.B(n_977),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_931),
.B(n_774),
.Y(n_1049)
);

O2A1O1Ixp5_ASAP7_75t_L g1050 ( 
.A1(n_945),
.A2(n_775),
.B(n_782),
.C(n_837),
.Y(n_1050)
);

CKINVDCx20_ASAP7_75t_R g1051 ( 
.A(n_1001),
.Y(n_1051)
);

OAI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_863),
.A2(n_775),
.B(n_837),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_R g1053 ( 
.A(n_860),
.B(n_844),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_R g1054 ( 
.A(n_914),
.B(n_774),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_884),
.A2(n_823),
.B(n_786),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_1026),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_912),
.A2(n_774),
.B1(n_854),
.B2(n_786),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_867),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_987),
.B(n_823),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_960),
.A2(n_782),
.B(n_736),
.C(n_732),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_870),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_882),
.B(n_917),
.Y(n_1062)
);

NOR2xp33_ASAP7_75t_L g1063 ( 
.A(n_879),
.B(n_736),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_913),
.A2(n_732),
.B(n_728),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_L g1065 ( 
.A1(n_933),
.A2(n_881),
.B1(n_971),
.B2(n_994),
.Y(n_1065)
);

BUFx12f_ASAP7_75t_L g1066 ( 
.A(n_973),
.Y(n_1066)
);

OAI22xp5_ASAP7_75t_L g1067 ( 
.A1(n_960),
.A2(n_866),
.B1(n_873),
.B2(n_868),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_908),
.B(n_854),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_L g1069 ( 
.A1(n_980),
.A2(n_728),
.B(n_715),
.C(n_854),
.Y(n_1069)
);

AOI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_859),
.A2(n_864),
.B1(n_891),
.B2(n_996),
.Y(n_1070)
);

AND2x2_ASAP7_75t_L g1071 ( 
.A(n_963),
.B(n_854),
.Y(n_1071)
);

O2A1O1Ixp5_ASAP7_75t_SL g1072 ( 
.A1(n_1019),
.A2(n_715),
.B(n_16),
.C(n_21),
.Y(n_1072)
);

NOR2xp33_ASAP7_75t_L g1073 ( 
.A(n_905),
.B(n_15),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_877),
.Y(n_1074)
);

CKINVDCx16_ASAP7_75t_R g1075 ( 
.A(n_1011),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_892),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_SL g1077 ( 
.A(n_1014),
.B(n_148),
.Y(n_1077)
);

BUFx6f_ASAP7_75t_L g1078 ( 
.A(n_966),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_1009),
.B(n_146),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_16),
.B(n_22),
.C(n_23),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_948),
.B(n_22),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_922),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_SL g1083 ( 
.A(n_1014),
.B(n_139),
.Y(n_1083)
);

AOI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_1016),
.A2(n_103),
.B(n_99),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_956),
.B(n_24),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_921),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_966),
.Y(n_1087)
);

INVx3_ASAP7_75t_L g1088 ( 
.A(n_949),
.Y(n_1088)
);

OR2x6_ASAP7_75t_L g1089 ( 
.A(n_872),
.B(n_98),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_861),
.A2(n_97),
.B(n_92),
.Y(n_1090)
);

BUFx12f_ASAP7_75t_L g1091 ( 
.A(n_946),
.Y(n_1091)
);

O2A1O1Ixp33_ASAP7_75t_L g1092 ( 
.A1(n_890),
.A2(n_907),
.B(n_1008),
.C(n_997),
.Y(n_1092)
);

OAI21xp33_ASAP7_75t_L g1093 ( 
.A1(n_907),
.A2(n_27),
.B(n_30),
.Y(n_1093)
);

O2A1O1Ixp5_ASAP7_75t_L g1094 ( 
.A1(n_904),
.A2(n_89),
.B(n_88),
.C(n_78),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1012),
.B(n_27),
.Y(n_1095)
);

BUFx2_ASAP7_75t_SL g1096 ( 
.A(n_921),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_873),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_1097)
);

NOR2xp67_ASAP7_75t_L g1098 ( 
.A(n_1028),
.B(n_31),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_875),
.A2(n_60),
.B(n_37),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_878),
.A2(n_59),
.B(n_38),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_994),
.B(n_35),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1025),
.A2(n_40),
.B(n_45),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_900),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_876),
.A2(n_40),
.B1(n_48),
.B2(n_50),
.Y(n_1104)
);

INVxp67_ASAP7_75t_SL g1105 ( 
.A(n_966),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_997),
.A2(n_48),
.B(n_56),
.C(n_58),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_933),
.Y(n_1107)
);

O2A1O1Ixp5_ASAP7_75t_L g1108 ( 
.A1(n_886),
.A2(n_56),
.B(n_983),
.C(n_1015),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_901),
.Y(n_1109)
);

AO22x1_ASAP7_75t_L g1110 ( 
.A1(n_893),
.A2(n_995),
.B1(n_887),
.B2(n_1037),
.Y(n_1110)
);

AND3x1_ASAP7_75t_SL g1111 ( 
.A(n_1018),
.B(n_1041),
.C(n_1006),
.Y(n_1111)
);

O2A1O1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1008),
.A2(n_961),
.B(n_968),
.C(n_881),
.Y(n_1112)
);

OAI22x1_ASAP7_75t_L g1113 ( 
.A1(n_1034),
.A2(n_989),
.B1(n_872),
.B2(n_1033),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_869),
.B(n_984),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_986),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_874),
.A2(n_909),
.B(n_888),
.Y(n_1116)
);

A2O1A1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_874),
.A2(n_1015),
.B(n_975),
.C(n_876),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_976),
.B(n_982),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_869),
.A2(n_880),
.B1(n_926),
.B2(n_950),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_926),
.B(n_976),
.Y(n_1120)
);

OAI22xp5_ASAP7_75t_L g1121 ( 
.A1(n_925),
.A2(n_939),
.B1(n_928),
.B2(n_944),
.Y(n_1121)
);

HB1xp67_ASAP7_75t_L g1122 ( 
.A(n_921),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_949),
.B(n_1029),
.Y(n_1123)
);

O2A1O1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_961),
.A2(n_968),
.B(n_1030),
.C(n_1038),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1033),
.A2(n_865),
.B1(n_902),
.B2(n_896),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_982),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_R g1127 ( 
.A(n_955),
.B(n_1010),
.Y(n_1127)
);

O2A1O1Ixp5_ASAP7_75t_L g1128 ( 
.A1(n_1019),
.A2(n_958),
.B(n_938),
.C(n_932),
.Y(n_1128)
);

O2A1O1Ixp5_ASAP7_75t_L g1129 ( 
.A1(n_1020),
.A2(n_1000),
.B(n_941),
.C(n_981),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1042),
.A2(n_1043),
.B(n_974),
.C(n_1045),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_910),
.Y(n_1131)
);

A2O1A1Ixp33_ASAP7_75t_SL g1132 ( 
.A1(n_981),
.A2(n_871),
.B(n_955),
.C(n_1046),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_984),
.B(n_915),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_974),
.B(n_1010),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_L g1135 ( 
.A(n_986),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_986),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_954),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_979),
.B(n_1027),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_906),
.A2(n_1021),
.B1(n_871),
.B2(n_957),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_959),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_964),
.B(n_1027),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1031),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_898),
.B(n_957),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_894),
.A2(n_895),
.B(n_885),
.Y(n_1144)
);

O2A1O1Ixp33_ASAP7_75t_L g1145 ( 
.A1(n_929),
.A2(n_911),
.B(n_965),
.C(n_916),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_993),
.B(n_1013),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1044),
.Y(n_1147)
);

BUFx12f_ASAP7_75t_L g1148 ( 
.A(n_991),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_889),
.A2(n_972),
.B(n_998),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_1024),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_1036),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_991),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_951),
.A2(n_1032),
.B1(n_969),
.B2(n_899),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_918),
.B(n_947),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_972),
.A2(n_920),
.B(n_883),
.Y(n_1155)
);

BUFx12f_ASAP7_75t_L g1156 ( 
.A(n_991),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_L g1157 ( 
.A(n_923),
.B(n_930),
.Y(n_1157)
);

NOR2xp33_ASAP7_75t_L g1158 ( 
.A(n_937),
.B(n_985),
.Y(n_1158)
);

AO32x2_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_969),
.A3(n_897),
.B1(n_940),
.B2(n_970),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_919),
.A2(n_990),
.B(n_999),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_990),
.B(n_999),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1036),
.Y(n_1162)
);

A2O1A1Ixp33_ASAP7_75t_L g1163 ( 
.A1(n_934),
.A2(n_924),
.B(n_943),
.C(n_936),
.Y(n_1163)
);

BUFx2_ASAP7_75t_L g1164 ( 
.A(n_991),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1002),
.A2(n_992),
.B(n_953),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_991),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_903),
.Y(n_1167)
);

A2O1A1Ixp33_ASAP7_75t_SL g1168 ( 
.A1(n_927),
.A2(n_1005),
.B(n_942),
.C(n_1039),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_SL g1169 ( 
.A1(n_1040),
.A2(n_1047),
.B1(n_935),
.B2(n_962),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1003),
.A2(n_1007),
.B(n_1004),
.C(n_1035),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_967),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_978),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_988),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1022),
.A2(n_1023),
.B(n_1017),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1175)
);

AO32x2_ASAP7_75t_L g1176 ( 
.A1(n_881),
.A2(n_792),
.A3(n_989),
.B1(n_907),
.B2(n_890),
.Y(n_1176)
);

A2O1A1Ixp33_ASAP7_75t_SL g1177 ( 
.A1(n_862),
.A2(n_696),
.B(n_542),
.C(n_553),
.Y(n_1177)
);

NAND2x1p5_ASAP7_75t_L g1178 ( 
.A(n_1014),
.B(n_872),
.Y(n_1178)
);

BUFx12f_ASAP7_75t_L g1179 ( 
.A(n_914),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_862),
.B(n_711),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_SL g1181 ( 
.A(n_862),
.B(n_539),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_914),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_966),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_879),
.A2(n_699),
.B1(n_552),
.B2(n_637),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_862),
.B(n_542),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_862),
.B(n_711),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_865),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_SL g1189 ( 
.A(n_862),
.B(n_539),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_945),
.A2(n_711),
.B(n_862),
.C(n_696),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_917),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_862),
.B(n_539),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_867),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_966),
.Y(n_1195)
);

AOI22xp5_ASAP7_75t_L g1196 ( 
.A1(n_862),
.A2(n_700),
.B1(n_696),
.B2(n_987),
.Y(n_1196)
);

AOI21xp5_ASAP7_75t_L g1197 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_945),
.A2(n_711),
.B(n_696),
.C(n_862),
.Y(n_1198)
);

BUFx2_ASAP7_75t_L g1199 ( 
.A(n_870),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_966),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_862),
.B(n_539),
.Y(n_1203)
);

HB1xp67_ASAP7_75t_L g1204 ( 
.A(n_870),
.Y(n_1204)
);

OAI21xp33_ASAP7_75t_SL g1205 ( 
.A1(n_960),
.A2(n_700),
.B(n_862),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_884),
.A2(n_913),
.B(n_1016),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1192),
.Y(n_1207)
);

AO31x2_ASAP7_75t_L g1208 ( 
.A1(n_1191),
.A2(n_1067),
.A3(n_1139),
.B(n_1153),
.Y(n_1208)
);

OA21x2_ASAP7_75t_L g1209 ( 
.A1(n_1128),
.A2(n_1108),
.B(n_1129),
.Y(n_1209)
);

AO31x2_ASAP7_75t_L g1210 ( 
.A1(n_1067),
.A2(n_1139),
.A3(n_1153),
.B(n_1163),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1186),
.B(n_1181),
.Y(n_1211)
);

AO22x1_ASAP7_75t_L g1212 ( 
.A1(n_1118),
.A2(n_1126),
.B1(n_1063),
.B2(n_1120),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1051),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_SL g1215 ( 
.A1(n_1177),
.A2(n_1198),
.B(n_1187),
.C(n_1180),
.Y(n_1215)
);

AOI22xp5_ASAP7_75t_L g1216 ( 
.A1(n_1205),
.A2(n_1048),
.B1(n_1196),
.B2(n_1093),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1149),
.A2(n_1116),
.B(n_1144),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1189),
.B(n_1193),
.Y(n_1218)
);

AO31x2_ASAP7_75t_L g1219 ( 
.A1(n_1197),
.A2(n_1202),
.A3(n_1201),
.B(n_1206),
.Y(n_1219)
);

OAI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1117),
.A2(n_1092),
.B(n_1112),
.Y(n_1220)
);

AO22x2_ASAP7_75t_L g1221 ( 
.A1(n_1104),
.A2(n_1097),
.B1(n_1119),
.B2(n_1125),
.Y(n_1221)
);

AND2x2_ASAP7_75t_L g1222 ( 
.A(n_1203),
.B(n_1192),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1065),
.A2(n_1070),
.B1(n_1134),
.B2(n_1059),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1174),
.A2(n_1155),
.B(n_1165),
.Y(n_1224)
);

AOI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1101),
.A2(n_1110),
.B1(n_1082),
.B2(n_1095),
.Y(n_1225)
);

BUFx2_ASAP7_75t_L g1226 ( 
.A(n_1061),
.Y(n_1226)
);

BUFx2_ASAP7_75t_R g1227 ( 
.A(n_1056),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1204),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1124),
.A2(n_1130),
.B(n_1158),
.C(n_1069),
.Y(n_1229)
);

AOI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1091),
.A2(n_1125),
.B1(n_1113),
.B2(n_1083),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1199),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1133),
.B(n_1114),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1160),
.A2(n_1055),
.B(n_1064),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1170),
.A2(n_1145),
.B(n_1052),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1143),
.B(n_1107),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1052),
.A2(n_1050),
.B(n_1121),
.Y(n_1236)
);

AND2x4_ASAP7_75t_L g1237 ( 
.A(n_1167),
.B(n_1122),
.Y(n_1237)
);

OAI21x1_ASAP7_75t_L g1238 ( 
.A1(n_1121),
.A2(n_1084),
.B(n_1161),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_R g1239 ( 
.A(n_1179),
.B(n_1182),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1062),
.B(n_1185),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1146),
.B(n_1151),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1162),
.B(n_1142),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1086),
.B(n_1053),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1171),
.A2(n_1172),
.B(n_1090),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1140),
.B(n_1081),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1074),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1123),
.B(n_1088),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1085),
.B(n_1088),
.Y(n_1248)
);

BUFx2_ASAP7_75t_L g1249 ( 
.A(n_1075),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1073),
.B(n_1147),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1060),
.A2(n_1068),
.B(n_1100),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1132),
.A2(n_1169),
.B(n_1154),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1157),
.A2(n_1168),
.B(n_1049),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1138),
.A2(n_1173),
.B(n_1083),
.Y(n_1254)
);

INVx2_ASAP7_75t_L g1255 ( 
.A(n_1076),
.Y(n_1255)
);

NOR2x1_ASAP7_75t_R g1256 ( 
.A(n_1066),
.B(n_1096),
.Y(n_1256)
);

INVx2_ASAP7_75t_SL g1257 ( 
.A(n_1136),
.Y(n_1257)
);

AOI21xp33_ASAP7_75t_L g1258 ( 
.A1(n_1080),
.A2(n_1106),
.B(n_1097),
.Y(n_1258)
);

AND2x2_ASAP7_75t_L g1259 ( 
.A(n_1071),
.B(n_1188),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_1127),
.Y(n_1260)
);

OAI22x1_ASAP7_75t_L g1261 ( 
.A1(n_1103),
.A2(n_1194),
.B1(n_1109),
.B2(n_1123),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1078),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1166),
.Y(n_1263)
);

A2O1A1Ixp33_ASAP7_75t_L g1264 ( 
.A1(n_1099),
.A2(n_1057),
.B(n_1094),
.C(n_1077),
.Y(n_1264)
);

A2O1A1Ixp33_ASAP7_75t_L g1265 ( 
.A1(n_1077),
.A2(n_1131),
.B(n_1141),
.C(n_1152),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1164),
.A2(n_1150),
.B(n_1105),
.Y(n_1266)
);

OA21x2_ASAP7_75t_L g1267 ( 
.A1(n_1102),
.A2(n_1159),
.B(n_1104),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1072),
.A2(n_1178),
.B(n_1150),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1089),
.A2(n_1159),
.B(n_1098),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1078),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1178),
.B(n_1079),
.Y(n_1271)
);

BUFx2_ASAP7_75t_L g1272 ( 
.A(n_1087),
.Y(n_1272)
);

OAI21x1_ASAP7_75t_L g1273 ( 
.A1(n_1150),
.A2(n_1159),
.B(n_1176),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1166),
.A2(n_1089),
.B(n_1087),
.Y(n_1274)
);

A2O1A1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1176),
.A2(n_1166),
.B(n_1087),
.C(n_1195),
.Y(n_1275)
);

INVx4_ASAP7_75t_L g1276 ( 
.A(n_1115),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1089),
.A2(n_1200),
.B(n_1195),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1115),
.A2(n_1195),
.B(n_1135),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1115),
.Y(n_1279)
);

AOI21xp5_ASAP7_75t_L g1280 ( 
.A1(n_1135),
.A2(n_1184),
.B(n_1200),
.Y(n_1280)
);

OAI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1148),
.A2(n_1156),
.B1(n_1176),
.B2(n_1184),
.Y(n_1281)
);

AO21x1_ASAP7_75t_L g1282 ( 
.A1(n_1111),
.A2(n_1184),
.B(n_1200),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1054),
.A2(n_1183),
.B(n_1175),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1192),
.Y(n_1284)
);

OR2x2_ASAP7_75t_L g1285 ( 
.A(n_1192),
.B(n_539),
.Y(n_1285)
);

AO32x2_ASAP7_75t_L g1286 ( 
.A1(n_1067),
.A2(n_1139),
.A3(n_1104),
.B1(n_1097),
.B2(n_1153),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1191),
.A2(n_886),
.A3(n_1067),
.B(n_1139),
.Y(n_1287)
);

BUFx4f_ASAP7_75t_L g1288 ( 
.A(n_1179),
.Y(n_1288)
);

INVx3_ASAP7_75t_L g1289 ( 
.A(n_1166),
.Y(n_1289)
);

AO22x2_ASAP7_75t_L g1290 ( 
.A1(n_1104),
.A2(n_1097),
.B1(n_1067),
.B2(n_1119),
.Y(n_1290)
);

AOI21xp5_ASAP7_75t_L g1291 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1058),
.Y(n_1292)
);

AOI21xp5_ASAP7_75t_L g1293 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1058),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1186),
.A2(n_1205),
.B(n_1198),
.C(n_1048),
.Y(n_1297)
);

AOI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1166),
.Y(n_1299)
);

BUFx6f_ASAP7_75t_L g1300 ( 
.A(n_1086),
.Y(n_1300)
);

NOR2x1_ASAP7_75t_SL g1301 ( 
.A(n_1136),
.B(n_1125),
.Y(n_1301)
);

AO32x2_ASAP7_75t_L g1302 ( 
.A1(n_1067),
.A2(n_1139),
.A3(n_1104),
.B1(n_1097),
.B2(n_1153),
.Y(n_1302)
);

A2O1A1Ixp33_ASAP7_75t_L g1303 ( 
.A1(n_1186),
.A2(n_1205),
.B(n_1198),
.C(n_1048),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1304)
);

NOR4xp25_ASAP7_75t_L g1305 ( 
.A(n_1092),
.B(n_1198),
.C(n_1112),
.D(n_1205),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1186),
.B(n_539),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1307)
);

CKINVDCx12_ASAP7_75t_R g1308 ( 
.A(n_1062),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1309)
);

OAI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1186),
.A2(n_696),
.B(n_542),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1311)
);

BUFx4f_ASAP7_75t_L g1312 ( 
.A(n_1179),
.Y(n_1312)
);

AOI31xp67_ASAP7_75t_L g1313 ( 
.A1(n_1180),
.A2(n_1032),
.A3(n_1187),
.B(n_1196),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1161),
.A2(n_1025),
.B(n_1116),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1186),
.A2(n_1205),
.B(n_1198),
.C(n_1048),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1058),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1186),
.B(n_539),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1191),
.A2(n_886),
.A3(n_1067),
.B(n_1139),
.Y(n_1319)
);

OA21x2_ASAP7_75t_L g1320 ( 
.A1(n_1128),
.A2(n_1108),
.B(n_1129),
.Y(n_1320)
);

AOI221xp5_ASAP7_75t_L g1321 ( 
.A1(n_1186),
.A2(n_542),
.B1(n_696),
.B2(n_1118),
.C(n_1092),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1186),
.B(n_539),
.Y(n_1322)
);

O2A1O1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1048),
.C(n_945),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1149),
.A2(n_1116),
.B(n_1144),
.Y(n_1324)
);

OAI221xp5_ASAP7_75t_L g1325 ( 
.A1(n_1186),
.A2(n_1048),
.B1(n_542),
.B2(n_1177),
.C(n_862),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1186),
.A2(n_700),
.B1(n_1196),
.B2(n_711),
.Y(n_1326)
);

A2O1A1Ixp33_ASAP7_75t_L g1327 ( 
.A1(n_1186),
.A2(n_1205),
.B(n_1198),
.C(n_1048),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1167),
.B(n_1011),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1136),
.Y(n_1329)
);

OR2x6_ASAP7_75t_L g1330 ( 
.A(n_1096),
.B(n_720),
.Y(n_1330)
);

O2A1O1Ixp5_ASAP7_75t_SL g1331 ( 
.A1(n_1097),
.A2(n_1104),
.B(n_755),
.C(n_690),
.Y(n_1331)
);

OAI21x1_ASAP7_75t_L g1332 ( 
.A1(n_1149),
.A2(n_1116),
.B(n_1144),
.Y(n_1332)
);

OAI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1186),
.A2(n_1196),
.B1(n_806),
.B2(n_539),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1186),
.B(n_539),
.Y(n_1334)
);

O2A1O1Ixp33_ASAP7_75t_L g1335 ( 
.A1(n_1177),
.A2(n_1186),
.B(n_1048),
.C(n_945),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1336)
);

BUFx2_ASAP7_75t_L g1337 ( 
.A(n_1192),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1338)
);

AO31x2_ASAP7_75t_L g1339 ( 
.A1(n_1191),
.A2(n_886),
.A3(n_1067),
.B(n_1139),
.Y(n_1339)
);

O2A1O1Ixp5_ASAP7_75t_L g1340 ( 
.A1(n_1186),
.A2(n_1177),
.B(n_945),
.C(n_862),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1341)
);

INVx2_ASAP7_75t_L g1342 ( 
.A(n_1137),
.Y(n_1342)
);

BUFx6f_ASAP7_75t_L g1343 ( 
.A(n_1086),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1179),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1149),
.A2(n_1116),
.B(n_1144),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1058),
.Y(n_1347)
);

AOI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1348)
);

NAND2xp5_ASAP7_75t_L g1349 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1349)
);

NAND2xp5_ASAP7_75t_L g1350 ( 
.A(n_1186),
.B(n_1180),
.Y(n_1350)
);

INVx5_ASAP7_75t_L g1351 ( 
.A(n_1078),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1186),
.A2(n_1118),
.B1(n_1048),
.B2(n_700),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1186),
.B(n_1048),
.Y(n_1354)
);

AO32x2_ASAP7_75t_L g1355 ( 
.A1(n_1067),
.A2(n_1139),
.A3(n_1104),
.B1(n_1097),
.B2(n_1153),
.Y(n_1355)
);

OAI21xp5_ASAP7_75t_L g1356 ( 
.A1(n_1205),
.A2(n_1191),
.B(n_1198),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_SL g1358 ( 
.A1(n_1092),
.A2(n_1112),
.B(n_886),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1175),
.A2(n_1190),
.B(n_1183),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1186),
.A2(n_1118),
.B1(n_1048),
.B2(n_700),
.Y(n_1360)
);

CKINVDCx20_ASAP7_75t_R g1361 ( 
.A(n_1051),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1321),
.A2(n_1310),
.B1(n_1360),
.B2(n_1352),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1300),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1310),
.A2(n_1326),
.B1(n_1325),
.B2(n_1309),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_1361),
.Y(n_1365)
);

CKINVDCx6p67_ASAP7_75t_R g1366 ( 
.A(n_1344),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1326),
.A2(n_1341),
.B1(n_1349),
.B2(n_1354),
.Y(n_1367)
);

BUFx4_ASAP7_75t_R g1368 ( 
.A(n_1227),
.Y(n_1368)
);

BUFx3_ASAP7_75t_L g1369 ( 
.A(n_1207),
.Y(n_1369)
);

BUFx2_ASAP7_75t_SL g1370 ( 
.A(n_1300),
.Y(n_1370)
);

INVx1_ASAP7_75t_SL g1371 ( 
.A(n_1285),
.Y(n_1371)
);

OAI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1307),
.A2(n_1346),
.B1(n_1338),
.B2(n_1336),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_SL g1373 ( 
.A1(n_1290),
.A2(n_1356),
.B1(n_1211),
.B2(n_1221),
.Y(n_1373)
);

BUFx12f_ASAP7_75t_L g1374 ( 
.A(n_1213),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1333),
.A2(n_1220),
.B1(n_1290),
.B2(n_1216),
.Y(n_1375)
);

INVx11_ASAP7_75t_L g1376 ( 
.A(n_1308),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1343),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1249),
.Y(n_1378)
);

INVx11_ASAP7_75t_L g1379 ( 
.A(n_1256),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1284),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1356),
.A2(n_1221),
.B1(n_1220),
.B2(n_1350),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_L g1382 ( 
.A1(n_1216),
.A2(n_1258),
.B1(n_1223),
.B2(n_1358),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1223),
.A2(n_1225),
.B1(n_1318),
.B2(n_1322),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1258),
.A2(n_1334),
.B1(n_1218),
.B2(n_1240),
.Y(n_1384)
);

CKINVDCx6p67_ASAP7_75t_R g1385 ( 
.A(n_1343),
.Y(n_1385)
);

BUFx10_ASAP7_75t_L g1386 ( 
.A(n_1328),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1234),
.Y(n_1387)
);

AOI21xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1297),
.A2(n_1303),
.B(n_1316),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1225),
.A2(n_1250),
.B1(n_1222),
.B2(n_1230),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1342),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1269),
.A2(n_1245),
.B1(n_1337),
.B2(n_1259),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1246),
.Y(n_1392)
);

AOI22xp33_ASAP7_75t_L g1393 ( 
.A1(n_1230),
.A2(n_1269),
.B1(n_1235),
.B2(n_1241),
.Y(n_1393)
);

INVx1_ASAP7_75t_SL g1394 ( 
.A(n_1226),
.Y(n_1394)
);

BUFx8_ASAP7_75t_SL g1395 ( 
.A(n_1288),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1292),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1295),
.Y(n_1397)
);

BUFx8_ASAP7_75t_L g1398 ( 
.A(n_1272),
.Y(n_1398)
);

BUFx2_ASAP7_75t_R g1399 ( 
.A(n_1243),
.Y(n_1399)
);

INVx3_ASAP7_75t_SL g1400 ( 
.A(n_1260),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_1288),
.Y(n_1401)
);

INVx6_ASAP7_75t_L g1402 ( 
.A(n_1351),
.Y(n_1402)
);

BUFx8_ASAP7_75t_SL g1403 ( 
.A(n_1312),
.Y(n_1403)
);

INVx1_ASAP7_75t_SL g1404 ( 
.A(n_1231),
.Y(n_1404)
);

CKINVDCx11_ASAP7_75t_R g1405 ( 
.A(n_1260),
.Y(n_1405)
);

OAI22xp5_ASAP7_75t_SL g1406 ( 
.A1(n_1271),
.A2(n_1212),
.B1(n_1305),
.B2(n_1228),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1281),
.A2(n_1301),
.B1(n_1327),
.B2(n_1305),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1232),
.A2(n_1282),
.B1(n_1347),
.B2(n_1317),
.Y(n_1408)
);

BUFx2_ASAP7_75t_L g1409 ( 
.A(n_1262),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1242),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1261),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1270),
.Y(n_1412)
);

INVx8_ASAP7_75t_L g1413 ( 
.A(n_1351),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1281),
.A2(n_1320),
.B1(n_1209),
.B2(n_1302),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1237),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1247),
.Y(n_1416)
);

CKINVDCx11_ASAP7_75t_R g1417 ( 
.A(n_1330),
.Y(n_1417)
);

BUFx2_ASAP7_75t_L g1418 ( 
.A(n_1279),
.Y(n_1418)
);

CKINVDCx14_ASAP7_75t_R g1419 ( 
.A(n_1312),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1248),
.A2(n_1330),
.B1(n_1254),
.B2(n_1252),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1209),
.A2(n_1320),
.B1(n_1302),
.B2(n_1286),
.Y(n_1421)
);

BUFx10_ASAP7_75t_L g1422 ( 
.A(n_1257),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1215),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1229),
.A2(n_1264),
.B1(n_1265),
.B2(n_1323),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1267),
.A2(n_1247),
.B1(n_1251),
.B2(n_1253),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1274),
.A2(n_1267),
.B1(n_1277),
.B2(n_1286),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1286),
.A2(n_1302),
.B1(n_1355),
.B2(n_1273),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1251),
.A2(n_1340),
.B1(n_1236),
.B2(n_1355),
.Y(n_1428)
);

BUFx12f_ASAP7_75t_L g1429 ( 
.A(n_1329),
.Y(n_1429)
);

BUFx12f_ASAP7_75t_L g1430 ( 
.A(n_1329),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1335),
.B(n_1208),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1276),
.Y(n_1432)
);

BUFx10_ASAP7_75t_L g1433 ( 
.A(n_1256),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1355),
.A2(n_1238),
.B1(n_1331),
.B2(n_1283),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_L g1435 ( 
.A1(n_1263),
.A2(n_1299),
.B1(n_1289),
.B2(n_1244),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1275),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1263),
.A2(n_1299),
.B1(n_1289),
.B2(n_1208),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1266),
.A2(n_1276),
.B1(n_1278),
.B2(n_1280),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1208),
.A2(n_1298),
.B1(n_1214),
.B2(n_1357),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1291),
.A2(n_1304),
.B1(n_1353),
.B2(n_1348),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1239),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1313),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1293),
.A2(n_1296),
.B1(n_1315),
.B2(n_1311),
.Y(n_1443)
);

OAI22x1_ASAP7_75t_SL g1444 ( 
.A1(n_1239),
.A2(n_1339),
.B1(n_1319),
.B2(n_1287),
.Y(n_1444)
);

INVx3_ASAP7_75t_L g1445 ( 
.A(n_1268),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1287),
.Y(n_1446)
);

BUFx2_ASAP7_75t_L g1447 ( 
.A(n_1287),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1294),
.A2(n_1359),
.B1(n_1319),
.B2(n_1339),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1219),
.Y(n_1449)
);

BUFx2_ASAP7_75t_SL g1450 ( 
.A(n_1219),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1339),
.A2(n_1210),
.B1(n_1233),
.B2(n_1224),
.Y(n_1451)
);

BUFx6f_ASAP7_75t_L g1452 ( 
.A(n_1314),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1210),
.A2(n_1217),
.B1(n_1324),
.B2(n_1332),
.Y(n_1453)
);

BUFx4f_ASAP7_75t_SL g1454 ( 
.A(n_1219),
.Y(n_1454)
);

CKINVDCx11_ASAP7_75t_R g1455 ( 
.A(n_1345),
.Y(n_1455)
);

BUFx3_ASAP7_75t_L g1456 ( 
.A(n_1207),
.Y(n_1456)
);

BUFx12f_ASAP7_75t_L g1457 ( 
.A(n_1344),
.Y(n_1457)
);

INVx8_ASAP7_75t_L g1458 ( 
.A(n_1351),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1255),
.Y(n_1459)
);

CKINVDCx11_ASAP7_75t_R g1460 ( 
.A(n_1344),
.Y(n_1460)
);

NAND2xp33_ASAP7_75t_R g1461 ( 
.A(n_1213),
.B(n_756),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1255),
.Y(n_1462)
);

BUFx2_ASAP7_75t_SL g1463 ( 
.A(n_1361),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1321),
.A2(n_1186),
.B1(n_1310),
.B2(n_1352),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_SL g1465 ( 
.A(n_1300),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1255),
.Y(n_1466)
);

OAI22xp5_ASAP7_75t_L g1467 ( 
.A1(n_1352),
.A2(n_1186),
.B1(n_1360),
.B2(n_1196),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1255),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1344),
.Y(n_1469)
);

INVx6_ASAP7_75t_L g1470 ( 
.A(n_1300),
.Y(n_1470)
);

BUFx3_ASAP7_75t_L g1471 ( 
.A(n_1207),
.Y(n_1471)
);

CKINVDCx16_ASAP7_75t_R g1472 ( 
.A(n_1361),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1310),
.A2(n_1186),
.B1(n_1048),
.B2(n_879),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1350),
.B(n_1186),
.Y(n_1474)
);

BUFx3_ASAP7_75t_L g1475 ( 
.A(n_1207),
.Y(n_1475)
);

INVx6_ASAP7_75t_L g1476 ( 
.A(n_1300),
.Y(n_1476)
);

INVx6_ASAP7_75t_L g1477 ( 
.A(n_1300),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1344),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1321),
.A2(n_1186),
.B1(n_1310),
.B2(n_1352),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1321),
.A2(n_1186),
.B1(n_1310),
.B2(n_1352),
.Y(n_1480)
);

AOI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1310),
.A2(n_1186),
.B1(n_1048),
.B2(n_879),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1306),
.B(n_1318),
.Y(n_1482)
);

CKINVDCx11_ASAP7_75t_R g1483 ( 
.A(n_1344),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_SL g1484 ( 
.A1(n_1326),
.A2(n_1186),
.B1(n_700),
.B2(n_1205),
.Y(n_1484)
);

INVx3_ASAP7_75t_L g1485 ( 
.A(n_1300),
.Y(n_1485)
);

INVx4_ASAP7_75t_L g1486 ( 
.A(n_1300),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1255),
.Y(n_1487)
);

OR2x6_ASAP7_75t_L g1488 ( 
.A(n_1274),
.B(n_1110),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1352),
.A2(n_1186),
.B1(n_1360),
.B2(n_1196),
.Y(n_1489)
);

INVx8_ASAP7_75t_L g1490 ( 
.A(n_1413),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1453),
.A2(n_1439),
.B(n_1440),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1453),
.A2(n_1439),
.B(n_1440),
.Y(n_1493)
);

AO21x2_ASAP7_75t_L g1494 ( 
.A1(n_1426),
.A2(n_1420),
.B(n_1442),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1452),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1467),
.A2(n_1489),
.B1(n_1464),
.B2(n_1479),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1431),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1387),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1387),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1452),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1448),
.Y(n_1501)
);

OAI21x1_ASAP7_75t_L g1502 ( 
.A1(n_1443),
.A2(n_1445),
.B(n_1448),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1411),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1436),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1449),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1402),
.Y(n_1506)
);

INVx1_ASAP7_75t_L g1507 ( 
.A(n_1426),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1449),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1473),
.A2(n_1481),
.B(n_1479),
.Y(n_1509)
);

OAI21x1_ASAP7_75t_L g1510 ( 
.A1(n_1451),
.A2(n_1434),
.B(n_1435),
.Y(n_1510)
);

OA21x2_ASAP7_75t_L g1511 ( 
.A1(n_1434),
.A2(n_1428),
.B(n_1425),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1373),
.B(n_1484),
.Y(n_1512)
);

NAND2x1p5_ASAP7_75t_L g1513 ( 
.A(n_1423),
.B(n_1438),
.Y(n_1513)
);

INVx3_ASAP7_75t_L g1514 ( 
.A(n_1454),
.Y(n_1514)
);

INVx2_ASAP7_75t_SL g1515 ( 
.A(n_1402),
.Y(n_1515)
);

BUFx12f_ASAP7_75t_L g1516 ( 
.A(n_1460),
.Y(n_1516)
);

O2A1O1Ixp5_ASAP7_75t_L g1517 ( 
.A1(n_1424),
.A2(n_1420),
.B(n_1372),
.C(n_1383),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1428),
.A2(n_1425),
.B(n_1451),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1392),
.Y(n_1519)
);

INVx2_ASAP7_75t_SL g1520 ( 
.A(n_1402),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1396),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1444),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1427),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1421),
.Y(n_1524)
);

AOI21x1_ASAP7_75t_L g1525 ( 
.A1(n_1488),
.A2(n_1397),
.B(n_1412),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_L g1526 ( 
.A(n_1371),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1450),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1446),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1455),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1414),
.Y(n_1530)
);

OR2x2_ASAP7_75t_L g1531 ( 
.A(n_1375),
.B(n_1391),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1435),
.A2(n_1437),
.B(n_1388),
.Y(n_1532)
);

OAI21x1_ASAP7_75t_L g1533 ( 
.A1(n_1437),
.A2(n_1382),
.B(n_1364),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1459),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1381),
.Y(n_1535)
);

AO21x2_ASAP7_75t_L g1536 ( 
.A1(n_1372),
.A2(n_1468),
.B(n_1487),
.Y(n_1536)
);

INVx2_ASAP7_75t_SL g1537 ( 
.A(n_1413),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1482),
.B(n_1474),
.Y(n_1538)
);

OAI21x1_ASAP7_75t_L g1539 ( 
.A1(n_1382),
.A2(n_1364),
.B(n_1408),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1381),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1413),
.Y(n_1541)
);

INVx1_ASAP7_75t_SL g1542 ( 
.A(n_1400),
.Y(n_1542)
);

INVxp67_ASAP7_75t_L g1543 ( 
.A(n_1369),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1462),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1466),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1375),
.A2(n_1393),
.B(n_1408),
.Y(n_1546)
);

OAI21x1_ASAP7_75t_L g1547 ( 
.A1(n_1393),
.A2(n_1362),
.B(n_1367),
.Y(n_1547)
);

NOR2xp33_ASAP7_75t_L g1548 ( 
.A(n_1400),
.B(n_1472),
.Y(n_1548)
);

OR2x6_ASAP7_75t_L g1549 ( 
.A(n_1488),
.B(n_1406),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1373),
.B(n_1389),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_SL g1551 ( 
.A(n_1384),
.B(n_1367),
.Y(n_1551)
);

BUFx3_ASAP7_75t_L g1552 ( 
.A(n_1417),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1458),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1407),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1407),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1484),
.B(n_1384),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1389),
.B(n_1362),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1418),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1464),
.A2(n_1480),
.B(n_1390),
.Y(n_1559)
);

INVx2_ASAP7_75t_L g1560 ( 
.A(n_1410),
.Y(n_1560)
);

AND2x2_ASAP7_75t_L g1561 ( 
.A(n_1480),
.B(n_1416),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1415),
.B(n_1409),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1380),
.B(n_1475),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1404),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1394),
.B(n_1456),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1471),
.Y(n_1566)
);

OAI21x1_ASAP7_75t_L g1567 ( 
.A1(n_1485),
.A2(n_1465),
.B(n_1430),
.Y(n_1567)
);

OA21x2_ASAP7_75t_L g1568 ( 
.A1(n_1432),
.A2(n_1441),
.B(n_1401),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1485),
.A2(n_1465),
.B(n_1429),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1422),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1398),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1399),
.A2(n_1419),
.B1(n_1376),
.B2(n_1385),
.Y(n_1572)
);

OAI21x1_ASAP7_75t_L g1573 ( 
.A1(n_1422),
.A2(n_1370),
.B(n_1398),
.Y(n_1573)
);

AO21x1_ASAP7_75t_SL g1574 ( 
.A1(n_1379),
.A2(n_1433),
.B(n_1395),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1386),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1463),
.B(n_1363),
.Y(n_1576)
);

CKINVDCx8_ASAP7_75t_R g1577 ( 
.A(n_1368),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1503),
.Y(n_1578)
);

AND2x4_ASAP7_75t_SL g1579 ( 
.A(n_1558),
.B(n_1433),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1524),
.B(n_1378),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1503),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1526),
.B(n_1486),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1491),
.A2(n_1470),
.B(n_1476),
.Y(n_1583)
);

INVx5_ASAP7_75t_L g1584 ( 
.A(n_1549),
.Y(n_1584)
);

OR2x2_ASAP7_75t_L g1585 ( 
.A(n_1519),
.B(n_1366),
.Y(n_1585)
);

BUFx4f_ASAP7_75t_SL g1586 ( 
.A(n_1516),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1530),
.B(n_1377),
.Y(n_1587)
);

AOI211xp5_ASAP7_75t_L g1588 ( 
.A1(n_1509),
.A2(n_1461),
.B(n_1405),
.C(n_1403),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1538),
.B(n_1377),
.Y(n_1589)
);

AOI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1496),
.A2(n_1365),
.B1(n_1457),
.B2(n_1374),
.Y(n_1590)
);

OR2x2_ASAP7_75t_L g1591 ( 
.A(n_1519),
.B(n_1483),
.Y(n_1591)
);

A2O1A1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1517),
.A2(n_1470),
.B(n_1476),
.C(n_1477),
.Y(n_1592)
);

NAND4xp25_ASAP7_75t_L g1593 ( 
.A(n_1551),
.B(n_1478),
.C(n_1469),
.D(n_1470),
.Y(n_1593)
);

OAI21x1_ASAP7_75t_SL g1594 ( 
.A1(n_1529),
.A2(n_1525),
.B(n_1528),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1501),
.A2(n_1502),
.B(n_1493),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1516),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1523),
.B(n_1507),
.Y(n_1597)
);

AOI221xp5_ASAP7_75t_L g1598 ( 
.A1(n_1556),
.A2(n_1512),
.B1(n_1557),
.B2(n_1555),
.C(n_1554),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_L g1599 ( 
.A1(n_1557),
.A2(n_1550),
.B(n_1555),
.C(n_1554),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1507),
.B(n_1497),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1497),
.B(n_1519),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_L g1602 ( 
.A(n_1564),
.B(n_1560),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1556),
.B(n_1513),
.Y(n_1603)
);

NAND4xp25_ASAP7_75t_L g1604 ( 
.A(n_1535),
.B(n_1540),
.C(n_1522),
.D(n_1542),
.Y(n_1604)
);

BUFx2_ASAP7_75t_L g1605 ( 
.A(n_1566),
.Y(n_1605)
);

BUFx3_ASAP7_75t_L g1606 ( 
.A(n_1552),
.Y(n_1606)
);

O2A1O1Ixp33_ASAP7_75t_SL g1607 ( 
.A1(n_1550),
.A2(n_1529),
.B(n_1522),
.C(n_1531),
.Y(n_1607)
);

BUFx12f_ASAP7_75t_L g1608 ( 
.A(n_1516),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1563),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_L g1610 ( 
.A1(n_1513),
.A2(n_1510),
.B(n_1527),
.Y(n_1610)
);

OAI21xp5_ASAP7_75t_L g1611 ( 
.A1(n_1547),
.A2(n_1539),
.B(n_1559),
.Y(n_1611)
);

AOI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1549),
.A2(n_1529),
.B1(n_1546),
.B2(n_1547),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1549),
.A2(n_1546),
.B1(n_1528),
.B2(n_1512),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1492),
.Y(n_1614)
);

INVx2_ASAP7_75t_L g1615 ( 
.A(n_1521),
.Y(n_1615)
);

CKINVDCx5p33_ASAP7_75t_R g1616 ( 
.A(n_1577),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1540),
.B(n_1494),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1494),
.B(n_1528),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1534),
.B(n_1544),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1518),
.B(n_1534),
.Y(n_1620)
);

OR2x2_ASAP7_75t_L g1621 ( 
.A(n_1498),
.B(n_1499),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1534),
.Y(n_1622)
);

OA21x2_ASAP7_75t_L g1623 ( 
.A1(n_1532),
.A2(n_1533),
.B(n_1527),
.Y(n_1623)
);

NOR2xp67_ASAP7_75t_SL g1624 ( 
.A(n_1577),
.B(n_1552),
.Y(n_1624)
);

AOI221xp5_ASAP7_75t_L g1625 ( 
.A1(n_1561),
.A2(n_1531),
.B1(n_1504),
.B2(n_1562),
.C(n_1543),
.Y(n_1625)
);

BUFx3_ASAP7_75t_L g1626 ( 
.A(n_1552),
.Y(n_1626)
);

AOI211xp5_ASAP7_75t_L g1627 ( 
.A1(n_1572),
.A2(n_1548),
.B(n_1575),
.C(n_1576),
.Y(n_1627)
);

A2O1A1Ixp33_ASAP7_75t_L g1628 ( 
.A1(n_1532),
.A2(n_1546),
.B(n_1561),
.C(n_1514),
.Y(n_1628)
);

BUFx2_ASAP7_75t_L g1629 ( 
.A(n_1566),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1518),
.B(n_1545),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1518),
.B(n_1545),
.Y(n_1631)
);

AO21x2_ASAP7_75t_L g1632 ( 
.A1(n_1505),
.A2(n_1508),
.B(n_1499),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1622),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1620),
.B(n_1511),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1615),
.Y(n_1635)
);

BUFx3_ASAP7_75t_L g1636 ( 
.A(n_1594),
.Y(n_1636)
);

AND2x2_ASAP7_75t_L g1637 ( 
.A(n_1620),
.B(n_1511),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1630),
.B(n_1498),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_SL g1639 ( 
.A(n_1612),
.B(n_1513),
.Y(n_1639)
);

INVxp67_ASAP7_75t_SL g1640 ( 
.A(n_1614),
.Y(n_1640)
);

AND2x2_ASAP7_75t_L g1641 ( 
.A(n_1630),
.B(n_1511),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1536),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1631),
.Y(n_1643)
);

BUFx2_ASAP7_75t_L g1644 ( 
.A(n_1583),
.Y(n_1644)
);

NOR2xp33_ASAP7_75t_L g1645 ( 
.A(n_1604),
.B(n_1566),
.Y(n_1645)
);

INVx4_ASAP7_75t_L g1646 ( 
.A(n_1584),
.Y(n_1646)
);

HB1xp67_ASAP7_75t_L g1647 ( 
.A(n_1632),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1601),
.B(n_1536),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1623),
.B(n_1495),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1595),
.B(n_1495),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1632),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1623),
.B(n_1500),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1617),
.B(n_1500),
.Y(n_1653)
);

HB1xp67_ASAP7_75t_L g1654 ( 
.A(n_1621),
.Y(n_1654)
);

AOI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1598),
.A2(n_1549),
.B1(n_1562),
.B2(n_1504),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1583),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1618),
.B(n_1611),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1634),
.B(n_1618),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1635),
.Y(n_1659)
);

AOI22xp33_ASAP7_75t_L g1660 ( 
.A1(n_1655),
.A2(n_1593),
.B1(n_1613),
.B2(n_1625),
.Y(n_1660)
);

INVx2_ASAP7_75t_L g1661 ( 
.A(n_1649),
.Y(n_1661)
);

NAND4xp25_ASAP7_75t_L g1662 ( 
.A(n_1655),
.B(n_1599),
.C(n_1590),
.D(n_1588),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1634),
.B(n_1628),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1634),
.B(n_1628),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1647),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1648),
.B(n_1597),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1634),
.B(n_1610),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1637),
.B(n_1610),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1633),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1643),
.B(n_1605),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1637),
.B(n_1597),
.Y(n_1671)
);

BUFx2_ASAP7_75t_L g1672 ( 
.A(n_1650),
.Y(n_1672)
);

INVx3_ASAP7_75t_L g1673 ( 
.A(n_1650),
.Y(n_1673)
);

HB1xp67_ASAP7_75t_L g1674 ( 
.A(n_1647),
.Y(n_1674)
);

OAI21xp33_ASAP7_75t_L g1675 ( 
.A1(n_1655),
.A2(n_1603),
.B(n_1592),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1650),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVx4_ASAP7_75t_L g1678 ( 
.A(n_1646),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1648),
.B(n_1578),
.Y(n_1679)
);

O2A1O1Ixp33_ASAP7_75t_L g1680 ( 
.A1(n_1639),
.A2(n_1592),
.B(n_1607),
.C(n_1603),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1654),
.B(n_1581),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1638),
.B(n_1629),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1651),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1654),
.B(n_1602),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1642),
.B(n_1621),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1638),
.B(n_1619),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1652),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1665),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1663),
.B(n_1664),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1661),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1679),
.B(n_1657),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1662),
.A2(n_1639),
.B1(n_1584),
.B2(n_1580),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1663),
.B(n_1641),
.Y(n_1695)
);

INVxp67_ASAP7_75t_L g1696 ( 
.A(n_1681),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1664),
.B(n_1641),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1659),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1659),
.Y(n_1699)
);

INVx3_ASAP7_75t_L g1700 ( 
.A(n_1673),
.Y(n_1700)
);

AND2x2_ASAP7_75t_SL g1701 ( 
.A(n_1660),
.B(n_1646),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1664),
.B(n_1672),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_SL g1703 ( 
.A(n_1680),
.B(n_1636),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1672),
.B(n_1657),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1661),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1685),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1657),
.Y(n_1707)
);

AND2x4_ASAP7_75t_L g1708 ( 
.A(n_1678),
.B(n_1656),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1676),
.B(n_1656),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1681),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1686),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1656),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1662),
.A2(n_1584),
.B1(n_1580),
.B2(n_1608),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1666),
.B(n_1640),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1665),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1676),
.B(n_1644),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1644),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1685),
.B(n_1640),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1669),
.Y(n_1720)
);

INVx1_ASAP7_75t_SL g1721 ( 
.A(n_1670),
.Y(n_1721)
);

INVx3_ASAP7_75t_L g1722 ( 
.A(n_1673),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1687),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1669),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1689),
.B(n_1658),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1721),
.B(n_1670),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1699),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1699),
.Y(n_1728)
);

OAI211xp5_ASAP7_75t_L g1729 ( 
.A1(n_1703),
.A2(n_1675),
.B(n_1660),
.C(n_1680),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1699),
.Y(n_1730)
);

NOR2xp67_ASAP7_75t_SL g1731 ( 
.A(n_1703),
.B(n_1608),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1696),
.B(n_1645),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1689),
.B(n_1658),
.Y(n_1733)
);

INVx2_ASAP7_75t_SL g1734 ( 
.A(n_1708),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1696),
.B(n_1645),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1689),
.B(n_1658),
.Y(n_1736)
);

INVx2_ASAP7_75t_L g1737 ( 
.A(n_1709),
.Y(n_1737)
);

OR2x2_ASAP7_75t_L g1738 ( 
.A(n_1721),
.B(n_1670),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1698),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1698),
.Y(n_1740)
);

OR2x2_ASAP7_75t_L g1741 ( 
.A(n_1690),
.B(n_1686),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1690),
.B(n_1684),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1693),
.B(n_1684),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1708),
.Y(n_1744)
);

INVxp67_ASAP7_75t_SL g1745 ( 
.A(n_1716),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1693),
.B(n_1682),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1711),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1702),
.B(n_1671),
.Y(n_1748)
);

A2O1A1Ixp33_ASAP7_75t_L g1749 ( 
.A1(n_1701),
.A2(n_1675),
.B(n_1624),
.C(n_1627),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1711),
.Y(n_1750)
);

OR2x2_ASAP7_75t_L g1751 ( 
.A(n_1706),
.B(n_1682),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1713),
.B(n_1682),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1709),
.Y(n_1754)
);

OR2x2_ASAP7_75t_L g1755 ( 
.A(n_1706),
.B(n_1653),
.Y(n_1755)
);

AND2x4_ASAP7_75t_L g1756 ( 
.A(n_1702),
.B(n_1678),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1702),
.B(n_1671),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

OAI22xp5_ASAP7_75t_SL g1759 ( 
.A1(n_1714),
.A2(n_1586),
.B1(n_1596),
.B2(n_1616),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1720),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1691),
.B(n_1695),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1720),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1724),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1701),
.B(n_1607),
.C(n_1678),
.Y(n_1764)
);

INVx2_ASAP7_75t_L g1765 ( 
.A(n_1709),
.Y(n_1765)
);

NOR2x1_ASAP7_75t_L g1766 ( 
.A(n_1708),
.B(n_1606),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1715),
.B(n_1719),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1745),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1727),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1728),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1766),
.B(n_1708),
.Y(n_1772)
);

AOI211xp5_ASAP7_75t_L g1773 ( 
.A1(n_1729),
.A2(n_1701),
.B(n_1708),
.C(n_1688),
.Y(n_1773)
);

INVxp67_ASAP7_75t_SL g1774 ( 
.A(n_1731),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1732),
.B(n_1596),
.Y(n_1775)
);

AOI211x1_ASAP7_75t_L g1776 ( 
.A1(n_1764),
.A2(n_1707),
.B(n_1704),
.C(n_1719),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1725),
.B(n_1691),
.Y(n_1777)
);

AND4x1_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1714),
.C(n_1694),
.D(n_1701),
.Y(n_1778)
);

OR2x2_ASAP7_75t_L g1779 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1779)
);

AND2x2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.B(n_1736),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1761),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1761),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1749),
.A2(n_1759),
.B1(n_1694),
.B2(n_1735),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1730),
.Y(n_1784)
);

NAND2x1_ASAP7_75t_L g1785 ( 
.A(n_1756),
.B(n_1704),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1756),
.Y(n_1786)
);

OR2x2_ASAP7_75t_L g1787 ( 
.A(n_1726),
.B(n_1710),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1739),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1740),
.Y(n_1789)
);

AND2x4_ASAP7_75t_L g1790 ( 
.A(n_1756),
.B(n_1708),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1733),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1758),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1736),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1734),
.B(n_1606),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1747),
.B(n_1695),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1760),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1750),
.B(n_1695),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1752),
.B(n_1697),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1755),
.B(n_1697),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1748),
.Y(n_1800)
);

NAND4xp25_ASAP7_75t_L g1801 ( 
.A(n_1744),
.B(n_1591),
.C(n_1626),
.D(n_1589),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1751),
.B(n_1697),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1748),
.B(n_1704),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1774),
.B(n_1757),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1785),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1769),
.B(n_1757),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1792),
.Y(n_1808)
);

OAI32xp33_ASAP7_75t_L g1809 ( 
.A1(n_1782),
.A2(n_1765),
.A3(n_1737),
.B1(n_1754),
.B2(n_1726),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1775),
.B(n_1742),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1796),
.Y(n_1811)
);

AOI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1783),
.A2(n_1584),
.B1(n_1765),
.B2(n_1754),
.Y(n_1812)
);

NAND2xp5_ASAP7_75t_L g1813 ( 
.A(n_1776),
.B(n_1743),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1770),
.Y(n_1814)
);

AOI22xp33_ASAP7_75t_L g1815 ( 
.A1(n_1778),
.A2(n_1584),
.B1(n_1737),
.B2(n_1626),
.Y(n_1815)
);

AOI32xp33_ASAP7_75t_L g1816 ( 
.A1(n_1773),
.A2(n_1744),
.A3(n_1712),
.B1(n_1717),
.B2(n_1718),
.Y(n_1816)
);

AOI21xp33_ASAP7_75t_L g1817 ( 
.A1(n_1785),
.A2(n_1734),
.B(n_1738),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1771),
.Y(n_1818)
);

INVxp67_ASAP7_75t_L g1819 ( 
.A(n_1786),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1790),
.B(n_1707),
.Y(n_1820)
);

AOI22xp5_ASAP7_75t_L g1821 ( 
.A1(n_1801),
.A2(n_1678),
.B1(n_1707),
.B2(n_1636),
.Y(n_1821)
);

AOI31xp33_ASAP7_75t_L g1822 ( 
.A1(n_1786),
.A2(n_1616),
.A3(n_1738),
.B(n_1576),
.Y(n_1822)
);

AND2x2_ASAP7_75t_L g1823 ( 
.A(n_1790),
.B(n_1753),
.Y(n_1823)
);

INVx1_ASAP7_75t_SL g1824 ( 
.A(n_1790),
.Y(n_1824)
);

INVx1_ASAP7_75t_SL g1825 ( 
.A(n_1772),
.Y(n_1825)
);

O2A1O1Ixp33_ASAP7_75t_L g1826 ( 
.A1(n_1788),
.A2(n_1688),
.B(n_1716),
.C(n_1753),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1789),
.B(n_1715),
.Y(n_1827)
);

AOI32xp33_ASAP7_75t_L g1828 ( 
.A1(n_1772),
.A2(n_1717),
.A3(n_1712),
.B1(n_1718),
.B2(n_1668),
.Y(n_1828)
);

INVx2_ASAP7_75t_SL g1829 ( 
.A(n_1794),
.Y(n_1829)
);

OAI31xp33_ASAP7_75t_L g1830 ( 
.A1(n_1815),
.A2(n_1772),
.A3(n_1781),
.B(n_1800),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1807),
.B(n_1802),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1806),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1808),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1815),
.A2(n_1794),
.B(n_1787),
.Y(n_1834)
);

AOI22xp5_ASAP7_75t_L g1835 ( 
.A1(n_1804),
.A2(n_1781),
.B1(n_1800),
.B2(n_1793),
.Y(n_1835)
);

INVxp67_ASAP7_75t_L g1836 ( 
.A(n_1804),
.Y(n_1836)
);

AOI22xp5_ASAP7_75t_L g1837 ( 
.A1(n_1824),
.A2(n_1793),
.B1(n_1791),
.B2(n_1798),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1823),
.B(n_1780),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1825),
.B(n_1678),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1805),
.Y(n_1840)
);

NOR2x1_ASAP7_75t_SL g1841 ( 
.A(n_1805),
.B(n_1794),
.Y(n_1841)
);

AOI322xp5_ASAP7_75t_L g1842 ( 
.A1(n_1813),
.A2(n_1803),
.A3(n_1791),
.B1(n_1780),
.B2(n_1768),
.C1(n_1777),
.C2(n_1799),
.Y(n_1842)
);

AOI221xp5_ASAP7_75t_L g1843 ( 
.A1(n_1816),
.A2(n_1784),
.B1(n_1797),
.B2(n_1795),
.C(n_1779),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1823),
.B(n_1768),
.Y(n_1844)
);

O2A1O1Ixp33_ASAP7_75t_L g1845 ( 
.A1(n_1826),
.A2(n_1794),
.B(n_1779),
.C(n_1787),
.Y(n_1845)
);

INVx2_ASAP7_75t_SL g1846 ( 
.A(n_1820),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1809),
.A2(n_1803),
.B1(n_1763),
.B2(n_1762),
.C(n_1777),
.Y(n_1847)
);

AOI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1812),
.A2(n_1718),
.B1(n_1712),
.B2(n_1717),
.C(n_1683),
.Y(n_1848)
);

AOI21xp33_ASAP7_75t_SL g1849 ( 
.A1(n_1822),
.A2(n_1568),
.B(n_1573),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1811),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1836),
.Y(n_1851)
);

INVxp67_ASAP7_75t_L g1852 ( 
.A(n_1841),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1838),
.Y(n_1853)
);

OAI222xp33_ASAP7_75t_L g1854 ( 
.A1(n_1845),
.A2(n_1812),
.B1(n_1828),
.B2(n_1819),
.C1(n_1810),
.C2(n_1821),
.Y(n_1854)
);

CKINVDCx14_ASAP7_75t_R g1855 ( 
.A(n_1832),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1843),
.A2(n_1817),
.B1(n_1820),
.B2(n_1829),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1843),
.A2(n_1829),
.B1(n_1827),
.B2(n_1818),
.Y(n_1857)
);

AOI221xp5_ASAP7_75t_L g1858 ( 
.A1(n_1848),
.A2(n_1814),
.B1(n_1668),
.B2(n_1667),
.C(n_1683),
.Y(n_1858)
);

XNOR2xp5_ASAP7_75t_L g1859 ( 
.A(n_1837),
.B(n_1571),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1840),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1835),
.Y(n_1861)
);

INVxp67_ASAP7_75t_L g1862 ( 
.A(n_1839),
.Y(n_1862)
);

NOR2x1_ASAP7_75t_L g1863 ( 
.A(n_1833),
.B(n_1571),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1853),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1860),
.Y(n_1865)
);

OAI211xp5_ASAP7_75t_L g1866 ( 
.A1(n_1856),
.A2(n_1830),
.B(n_1848),
.C(n_1834),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1852),
.B(n_1846),
.Y(n_1867)
);

NAND2xp5_ASAP7_75t_L g1868 ( 
.A(n_1855),
.B(n_1831),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1861),
.B(n_1844),
.Y(n_1869)
);

NAND3xp33_ASAP7_75t_SL g1870 ( 
.A(n_1857),
.B(n_1858),
.C(n_1862),
.Y(n_1870)
);

AND4x1_ASAP7_75t_L g1871 ( 
.A(n_1851),
.B(n_1847),
.C(n_1850),
.D(n_1574),
.Y(n_1871)
);

NAND4xp75_ASAP7_75t_L g1872 ( 
.A(n_1863),
.B(n_1847),
.C(n_1568),
.D(n_1849),
.Y(n_1872)
);

OAI211xp5_ASAP7_75t_SL g1873 ( 
.A1(n_1866),
.A2(n_1842),
.B(n_1854),
.C(n_1859),
.Y(n_1873)
);

AOI221xp5_ASAP7_75t_L g1874 ( 
.A1(n_1870),
.A2(n_1854),
.B1(n_1570),
.B2(n_1565),
.C(n_1579),
.Y(n_1874)
);

O2A1O1Ixp5_ASAP7_75t_L g1875 ( 
.A1(n_1868),
.A2(n_1700),
.B(n_1722),
.C(n_1692),
.Y(n_1875)
);

OAI211xp5_ASAP7_75t_L g1876 ( 
.A1(n_1868),
.A2(n_1571),
.B(n_1568),
.C(n_1570),
.Y(n_1876)
);

AOI211xp5_ASAP7_75t_L g1877 ( 
.A1(n_1867),
.A2(n_1573),
.B(n_1567),
.C(n_1569),
.Y(n_1877)
);

OAI211xp5_ASAP7_75t_L g1878 ( 
.A1(n_1873),
.A2(n_1874),
.B(n_1864),
.C(n_1869),
.Y(n_1878)
);

O2A1O1Ixp33_ASAP7_75t_L g1879 ( 
.A1(n_1876),
.A2(n_1865),
.B(n_1871),
.C(n_1872),
.Y(n_1879)
);

OAI211xp5_ASAP7_75t_L g1880 ( 
.A1(n_1877),
.A2(n_1574),
.B(n_1569),
.C(n_1567),
.Y(n_1880)
);

AOI211xp5_ASAP7_75t_SL g1881 ( 
.A1(n_1875),
.A2(n_1575),
.B(n_1582),
.C(n_1700),
.Y(n_1881)
);

AOI222xp33_ASAP7_75t_L g1882 ( 
.A1(n_1873),
.A2(n_1579),
.B1(n_1636),
.B2(n_1674),
.C1(n_1609),
.C2(n_1667),
.Y(n_1882)
);

AOI22xp33_ASAP7_75t_L g1883 ( 
.A1(n_1873),
.A2(n_1636),
.B1(n_1646),
.B2(n_1587),
.Y(n_1883)
);

OR2x2_ASAP7_75t_L g1884 ( 
.A(n_1883),
.B(n_1741),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1881),
.Y(n_1885)
);

NOR2x1_ASAP7_75t_L g1886 ( 
.A(n_1878),
.B(n_1563),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1882),
.B(n_1879),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1880),
.B(n_1700),
.Y(n_1888)
);

XOR2xp5_ASAP7_75t_L g1889 ( 
.A(n_1886),
.B(n_1585),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_SL g1890 ( 
.A(n_1885),
.B(n_1741),
.Y(n_1890)
);

OAI22xp5_ASAP7_75t_SL g1891 ( 
.A1(n_1884),
.A2(n_1553),
.B1(n_1537),
.B2(n_1541),
.Y(n_1891)
);

AND2x4_ASAP7_75t_L g1892 ( 
.A(n_1890),
.B(n_1887),
.Y(n_1892)
);

OAI22x1_ASAP7_75t_L g1893 ( 
.A1(n_1892),
.A2(n_1889),
.B1(n_1888),
.B2(n_1891),
.Y(n_1893)
);

OA21x2_ASAP7_75t_L g1894 ( 
.A1(n_1893),
.A2(n_1705),
.B(n_1692),
.Y(n_1894)
);

CKINVDCx20_ASAP7_75t_R g1895 ( 
.A(n_1893),
.Y(n_1895)
);

NOR3xp33_ASAP7_75t_L g1896 ( 
.A(n_1895),
.B(n_1541),
.C(n_1537),
.Y(n_1896)
);

AOI22x1_ASAP7_75t_L g1897 ( 
.A1(n_1894),
.A2(n_1553),
.B1(n_1746),
.B2(n_1520),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1896),
.B(n_1897),
.Y(n_1898)
);

OAI22xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1896),
.A2(n_1553),
.B1(n_1520),
.B2(n_1506),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1898),
.B(n_1692),
.Y(n_1900)
);

OAI21xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1899),
.B(n_1705),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1901),
.Y(n_1902)
);

OAI221xp5_ASAP7_75t_R g1903 ( 
.A1(n_1902),
.A2(n_1490),
.B1(n_1700),
.B2(n_1722),
.C(n_1723),
.Y(n_1903)
);

AOI211xp5_ASAP7_75t_L g1904 ( 
.A1(n_1903),
.A2(n_1553),
.B(n_1515),
.C(n_1506),
.Y(n_1904)
);


endmodule