module fake_jpeg_29557_n_170 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_170);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_47),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_36),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_11),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_42),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_18),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g60 ( 
.A(n_38),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_14),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_9),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_13),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_16),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_11),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_17),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_32),
.B(n_40),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_SL g73 ( 
.A(n_69),
.Y(n_73)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

BUFx5_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_50),
.B(n_0),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_81),
.Y(n_83)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_79),
.Y(n_85)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_68),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_87),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_66),
.Y(n_87)
);

NOR2x1_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_68),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_83),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_81),
.B(n_60),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_90),
.B(n_94),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_60),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_62),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_71),
.B(n_65),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_86),
.A2(n_72),
.B1(n_57),
.B2(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_98),
.A2(n_100),
.B1(n_112),
.B2(n_114),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_83),
.A2(n_72),
.B1(n_64),
.B2(n_67),
.Y(n_100)
);

AND2x6_ASAP7_75t_L g101 ( 
.A(n_94),
.B(n_55),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_102),
.Y(n_120)
);

INVx13_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVxp33_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_95),
.B(n_54),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_107),
.Y(n_126)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_63),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_70),
.B(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_115),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_89),
.A2(n_61),
.B(n_59),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_109),
.B(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_1),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_111),
.B(n_113),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_64),
.B1(n_52),
.B2(n_49),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_93),
.B(n_48),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g114 ( 
.A1(n_90),
.A2(n_21),
.B1(n_45),
.B2(n_44),
.Y(n_114)
);

O2A1O1Ixp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_20),
.B(n_41),
.C(n_37),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_94),
.B(n_1),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_7),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_15),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_104),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_123),
.B(n_127),
.Y(n_148)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_129),
.B(n_132),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_115),
.B(n_5),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_5),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_133),
.B(n_134),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_114),
.B(n_6),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_136),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_101),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_7),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_137),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_130),
.A2(n_46),
.B(n_25),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_142),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_118),
.A2(n_8),
.B(n_9),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_145),
.B(n_147),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_29),
.C(n_34),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_128),
.B(n_23),
.C(n_33),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_130),
.A2(n_8),
.B1(n_10),
.B2(n_12),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_151),
.A2(n_127),
.B1(n_131),
.B2(n_10),
.Y(n_154)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_118),
.B(n_121),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_152),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_155),
.Y(n_160)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_149),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_120),
.B(n_126),
.Y(n_157)
);

NOR3xp33_ASAP7_75t_L g161 ( 
.A(n_157),
.B(n_138),
.C(n_139),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_141),
.A2(n_119),
.B1(n_22),
.B2(n_30),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_147),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g163 ( 
.A(n_162),
.B(n_145),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_163),
.A2(n_148),
.B(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_165),
.Y(n_166)
);

AOI322xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_156),
.A3(n_159),
.B1(n_164),
.B2(n_142),
.C1(n_160),
.C2(n_151),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_159),
.C(n_150),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_169),
.A2(n_143),
.B(n_144),
.Y(n_170)
);


endmodule