module fake_jpeg_31373_n_416 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_416);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_416;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_45),
.Y(n_99)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g47 ( 
.A(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_47),
.B(n_66),
.Y(n_97)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_18),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_51),
.Y(n_106)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVx6_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_57),
.Y(n_133)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_58),
.Y(n_127)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_60),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_62),
.Y(n_102)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_64),
.Y(n_140)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_44),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g67 ( 
.A(n_39),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_71),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_20),
.B(n_31),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_68),
.B(n_86),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_20),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_82),
.Y(n_90)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_73),
.Y(n_138)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_76),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_75),
.Y(n_137)
);

BUFx12_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_16),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_79),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_83),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_15),
.B(n_0),
.Y(n_82)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_85),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_38),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_19),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_19),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_87),
.B(n_23),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_88),
.B(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_73),
.A2(n_27),
.B1(n_36),
.B2(n_34),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_91),
.A2(n_114),
.B1(n_122),
.B2(n_42),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g101 ( 
.A1(n_69),
.A2(n_82),
.B(n_24),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_101),
.B(n_10),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_104),
.B(n_116),
.Y(n_168)
);

INVx2_ASAP7_75t_R g108 ( 
.A(n_76),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_108),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_50),
.A2(n_27),
.B1(n_43),
.B2(n_24),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_110),
.A2(n_111),
.B1(n_118),
.B2(n_128),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_58),
.A2(n_40),
.B1(n_43),
.B2(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_15),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_112),
.B(n_119),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_60),
.A2(n_30),
.B1(n_33),
.B2(n_32),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_74),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_75),
.A2(n_27),
.B1(n_17),
.B2(n_33),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_32),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_54),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_135),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_72),
.A2(n_62),
.B1(n_67),
.B2(n_66),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_47),
.A2(n_31),
.B1(n_30),
.B2(n_23),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_71),
.B(n_17),
.Y(n_135)
);

OAI21xp33_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_90),
.B(n_108),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_141),
.B(n_142),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_118),
.A2(n_42),
.B1(n_21),
.B2(n_10),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_90),
.B(n_89),
.Y(n_144)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_144),
.Y(n_208)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_145),
.Y(n_199)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_146),
.Y(n_198)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_103),
.Y(n_147)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_147),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_105),
.A2(n_56),
.B1(n_71),
.B2(n_21),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_148),
.A2(n_150),
.B1(n_172),
.B2(n_187),
.Y(n_213)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_138),
.Y(n_149)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_137),
.A2(n_56),
.B1(n_84),
.B2(n_85),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_41),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_163),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_153),
.A2(n_156),
.B1(n_170),
.B2(n_171),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_162),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_119),
.A2(n_42),
.B1(n_41),
.B2(n_25),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_158),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_98),
.B(n_42),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_160),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_161),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_109),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_41),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_164),
.B(n_169),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_93),
.A2(n_42),
.B1(n_14),
.B2(n_11),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_14),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_107),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_91),
.A2(n_41),
.B1(n_25),
.B2(n_10),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_122),
.A2(n_41),
.B1(n_25),
.B2(n_9),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_107),
.A2(n_25),
.B1(n_9),
.B2(n_2),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_25),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_173),
.B(n_183),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_93),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_174),
.Y(n_212)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_117),
.Y(n_176)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_177),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_1),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_182),
.Y(n_205)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_95),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_180),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_95),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_181),
.Y(n_223)
);

AO22x1_ASAP7_75t_SL g182 ( 
.A1(n_124),
.A2(n_8),
.B1(n_102),
.B2(n_127),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_100),
.B(n_8),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_93),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_184),
.B(n_185),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_115),
.Y(n_185)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_115),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_186),
.A2(n_120),
.B1(n_99),
.B2(n_92),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_96),
.A2(n_8),
.B1(n_139),
.B2(n_132),
.Y(n_187)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_124),
.Y(n_188)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_188),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_168),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_194),
.B(n_201),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_120),
.C(n_100),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_196),
.B(n_227),
.C(n_208),
.Y(n_264)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_200),
.B(n_179),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_168),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_149),
.Y(n_210)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_210),
.Y(n_234)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_211),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_163),
.A2(n_134),
.B1(n_131),
.B2(n_126),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_214),
.Y(n_251)
);

A2O1A1Ixp33_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_125),
.B(n_102),
.C(n_99),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_225),
.Y(n_235)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_161),
.Y(n_222)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_222),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

MAJx2_ASAP7_75t_L g227 ( 
.A(n_144),
.B(n_126),
.C(n_94),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_154),
.A2(n_127),
.B1(n_106),
.B2(n_139),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_228),
.A2(n_171),
.B1(n_213),
.B2(n_170),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_177),
.Y(n_229)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_229),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_159),
.B1(n_185),
.B2(n_155),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_230),
.A2(n_245),
.B1(n_265),
.B2(n_212),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_231),
.B(n_241),
.Y(n_279)
);

AOI32xp33_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_175),
.A3(n_162),
.B1(n_166),
.B2(n_178),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_233),
.B(n_250),
.Y(n_278)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_174),
.Y(n_236)
);

OR2x2_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_238),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_218),
.A2(n_152),
.B1(n_145),
.B2(n_131),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_237),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_204),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_192),
.B(n_169),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_264),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g242 ( 
.A(n_226),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_242),
.B(n_248),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_226),
.A2(n_153),
.B1(n_156),
.B2(n_155),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_244),
.A2(n_246),
.B1(n_231),
.B2(n_236),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_220),
.A2(n_142),
.B1(n_160),
.B2(n_165),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_172),
.B1(n_182),
.B2(n_143),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_203),
.Y(n_247)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_247),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_183),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_218),
.A2(n_126),
.B1(n_94),
.B2(n_188),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_249),
.A2(n_251),
.B1(n_229),
.B2(n_190),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_193),
.B(n_176),
.Y(n_250)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_203),
.Y(n_252)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_252),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_216),
.B(n_158),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_222),
.Y(n_254)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_254),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_255),
.A2(n_259),
.B(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_195),
.Y(n_256)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_256),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_224),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_197),
.A2(n_182),
.B1(n_167),
.B2(n_147),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_192),
.B(n_146),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_261),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_215),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_198),
.Y(n_262)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_205),
.B(n_182),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_263),
.B(n_196),
.Y(n_267)
);

OAI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_221),
.A2(n_212),
.B1(n_223),
.B2(n_205),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_267),
.B(n_270),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_211),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_234),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_271),
.B(n_287),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_227),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_272),
.B(n_256),
.C(n_243),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g315 ( 
.A1(n_273),
.A2(n_191),
.B(n_130),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_230),
.B(n_202),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_276),
.B(n_290),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_232),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_280),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_241),
.B1(n_236),
.B2(n_247),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_234),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g288 ( 
.A(n_239),
.B(n_202),
.C(n_210),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_283),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_251),
.B1(n_255),
.B2(n_213),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_235),
.B(n_238),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_246),
.B1(n_244),
.B2(n_259),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_258),
.B(n_189),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_293),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_240),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_233),
.B(n_189),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_294),
.B(n_296),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g295 ( 
.A(n_245),
.B(n_228),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_106),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_255),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g339 ( 
.A(n_297),
.B(n_314),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_266),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_298),
.B(n_280),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_300),
.A2(n_305),
.B1(n_310),
.B2(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_303),
.B(n_309),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_304),
.B(n_283),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_295),
.A2(n_254),
.B1(n_243),
.B2(n_252),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_306),
.B(n_319),
.C(n_288),
.Y(n_330)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_266),
.Y(n_307)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_307),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_286),
.A2(n_240),
.B1(n_261),
.B2(n_257),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_291),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_276),
.A2(n_206),
.B1(n_207),
.B2(n_209),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_285),
.A2(n_257),
.B1(n_199),
.B2(n_262),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_315),
.A2(n_321),
.B(n_289),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_268),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_316),
.Y(n_345)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_274),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_317),
.B(n_320),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_199),
.B(n_217),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_279),
.B1(n_293),
.B2(n_287),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_272),
.B(n_198),
.C(n_217),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_274),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_275),
.A2(n_130),
.B(n_190),
.Y(n_321)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_323),
.Y(n_337)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_324),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_325),
.B(n_306),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_322),
.A2(n_270),
.B(n_278),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_326),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_301),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_332),
.Y(n_355)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_329),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_330),
.B(n_300),
.C(n_312),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_331),
.A2(n_315),
.B1(n_323),
.B2(n_314),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_311),
.Y(n_332)
);

OAI32xp33_ASAP7_75t_L g335 ( 
.A1(n_312),
.A2(n_296),
.A3(n_267),
.B1(n_275),
.B2(n_279),
.Y(n_335)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_335),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_336),
.A2(n_271),
.B1(n_282),
.B2(n_269),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_302),
.B(n_281),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_338),
.B(n_316),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_273),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_343),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_299),
.B(n_277),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_302),
.B(n_284),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_344),
.A2(n_299),
.B1(n_308),
.B2(n_275),
.Y(n_346)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_346),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_347),
.B(n_350),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_341),
.B(n_319),
.Y(n_350)
);

NOR2x1_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_303),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_358),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_352),
.B(n_361),
.C(n_362),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_L g353 ( 
.A1(n_327),
.A2(n_297),
.B1(n_309),
.B2(n_285),
.Y(n_353)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_325),
.B(n_330),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_357),
.B(n_269),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_327),
.A2(n_279),
.B1(n_320),
.B2(n_317),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g372 ( 
.A(n_359),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_343),
.B(n_321),
.C(n_310),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_340),
.B(n_305),
.C(n_313),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_364),
.A2(n_334),
.B1(n_335),
.B2(n_282),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_348),
.A2(n_339),
.B(n_336),
.Y(n_366)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_366),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_370),
.B(n_356),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_352),
.B(n_340),
.C(n_339),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_371),
.B(n_374),
.C(n_375),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_354),
.B(n_339),
.C(n_333),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_347),
.B(n_324),
.C(n_337),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_348),
.A2(n_345),
.B(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_376),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_377),
.A2(n_378),
.B1(n_351),
.B2(n_363),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_360),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_379),
.B(n_359),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_388),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_381),
.B(n_390),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_350),
.C(n_356),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_384),
.B(n_386),
.C(n_373),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_385),
.Y(n_392)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_361),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_372),
.A2(n_355),
.B(n_362),
.Y(n_387)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_387),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_365),
.B(n_364),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_372),
.B(n_349),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_384),
.C(n_373),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_388),
.B(n_375),
.C(n_371),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_396),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_367),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_389),
.B(n_369),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_398),
.B(n_380),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_383),
.B(n_368),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_386),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_392),
.A2(n_382),
.B1(n_370),
.B2(n_377),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_400),
.B(n_403),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_402),
.B(n_391),
.C(n_395),
.Y(n_408)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_404),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g405 ( 
.A1(n_397),
.A2(n_393),
.B(n_394),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_405),
.A2(n_401),
.B(n_403),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_408),
.B(n_177),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_409),
.Y(n_411)
);

INVxp33_ASAP7_75t_L g412 ( 
.A(n_410),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_411),
.A2(n_407),
.B(n_406),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_413),
.B(n_130),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_414),
.B(n_412),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_415),
.B(n_132),
.Y(n_416)
);


endmodule