module fake_jpeg_3625_n_638 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_638);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_638;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_3),
.B(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_5),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g52 ( 
.A(n_16),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_7),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_7),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_0),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_62),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_63),
.Y(n_183)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_64),
.Y(n_196)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_65),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g142 ( 
.A(n_68),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_55),
.Y(n_69)
);

INVx6_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_71),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_72),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_10),
.B1(n_17),
.B2(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_73),
.A2(n_45),
.B1(n_43),
.B2(n_40),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_9),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_74),
.B(n_61),
.Y(n_165)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_75),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_76),
.Y(n_172)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_77),
.Y(n_176)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_78),
.Y(n_137)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_79),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_80),
.Y(n_212)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_34),
.Y(n_81)
);

INVx5_ASAP7_75t_L g207 ( 
.A(n_81),
.Y(n_207)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_82),
.Y(n_140)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_23),
.Y(n_83)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_83),
.Y(n_143)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_59),
.Y(n_87)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_87),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_32),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_88),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_89),
.Y(n_150)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_92),
.Y(n_156)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_93),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_94),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_58),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_96),
.B(n_99),
.Y(n_133)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_20),
.Y(n_98)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_58),
.B(n_8),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g100 ( 
.A(n_32),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_100),
.Y(n_171)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_101),
.Y(n_164)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_39),
.Y(n_102)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_26),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_38),
.A2(n_8),
.B(n_15),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_104),
.B(n_112),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_26),
.Y(n_105)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_105),
.Y(n_153)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_60),
.Y(n_106)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_106),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_107),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_44),
.B(n_14),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_108),
.B(n_33),
.Y(n_189)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_109),
.Y(n_180)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_32),
.Y(n_110)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_111),
.Y(n_192)
);

BUFx12f_ASAP7_75t_SL g112 ( 
.A(n_29),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_36),
.Y(n_114)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_114),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_60),
.Y(n_116)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_116),
.Y(n_151)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_50),
.Y(n_118)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_118),
.Y(n_178)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

BUFx24_ASAP7_75t_L g120 ( 
.A(n_29),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_121),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_30),
.B(n_18),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_122),
.Y(n_198)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_51),
.Y(n_123)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_123),
.Y(n_201)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_47),
.Y(n_124)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_124),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_51),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_53),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_127),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_51),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g128 ( 
.A(n_37),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_37),
.Y(n_162)
);

INVx11_ASAP7_75t_L g129 ( 
.A(n_39),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

OA22x2_ASAP7_75t_L g138 ( 
.A1(n_123),
.A2(n_57),
.B1(n_53),
.B2(n_49),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g257 ( 
.A1(n_138),
.A2(n_144),
.B1(n_204),
.B2(n_28),
.Y(n_257)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_74),
.A2(n_31),
.B(n_56),
.C(n_35),
.Y(n_139)
);

OAI21xp33_ASAP7_75t_L g271 ( 
.A1(n_139),
.A2(n_165),
.B(n_189),
.Y(n_271)
);

OA22x2_ASAP7_75t_L g144 ( 
.A1(n_128),
.A2(n_57),
.B1(n_53),
.B2(n_49),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_61),
.B(n_44),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_161),
.A2(n_4),
.B(n_130),
.Y(n_284)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_91),
.A2(n_57),
.B1(n_30),
.B2(n_27),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_163),
.A2(n_177),
.B1(n_182),
.B2(n_191),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_56),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_166),
.B(n_167),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_96),
.B(n_54),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_99),
.B(n_31),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_173),
.B(n_181),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_94),
.A2(n_22),
.B1(n_46),
.B2(n_27),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_95),
.A2(n_22),
.B1(n_46),
.B2(n_41),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_184),
.B1(n_64),
.B2(n_65),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_100),
.B(n_40),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_125),
.A2(n_41),
.B1(n_33),
.B2(n_43),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_88),
.B(n_45),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_186),
.B(n_199),
.Y(n_288)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_122),
.A2(n_35),
.B1(n_54),
.B2(n_21),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_105),
.B(n_12),
.Y(n_197)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_197),
.B(n_1),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_77),
.B(n_12),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_107),
.A2(n_39),
.B1(n_21),
.B2(n_25),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_200),
.A2(n_4),
.B1(n_159),
.B2(n_131),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_81),
.B(n_120),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_202),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g204 ( 
.A(n_80),
.B(n_28),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_62),
.B(n_11),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_210),
.Y(n_276)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_136),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_214),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_216),
.B(n_228),
.Y(n_312)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_212),
.Y(n_217)
);

INVx3_ASAP7_75t_SL g294 ( 
.A(n_217),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_204),
.A2(n_118),
.B1(n_115),
.B2(n_114),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g298 ( 
.A1(n_218),
.A2(n_246),
.B1(n_264),
.B2(n_149),
.Y(n_298)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_212),
.Y(n_219)
);

INVx3_ASAP7_75t_SL g296 ( 
.A(n_219),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_171),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_220),
.B(n_258),
.Y(n_301)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_146),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_221),
.B(n_224),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_183),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_222),
.Y(n_346)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_204),
.B(n_0),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_225),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_151),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_201),
.Y(n_227)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_227),
.Y(n_315)
);

NAND2xp33_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_0),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g229 ( 
.A1(n_141),
.A2(n_161),
.B(n_139),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_229),
.A2(n_285),
.B(n_250),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g230 ( 
.A1(n_163),
.A2(n_111),
.B1(n_89),
.B2(n_87),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_230),
.A2(n_260),
.B1(n_277),
.B2(n_244),
.Y(n_319)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_174),
.Y(n_232)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_232),
.Y(n_343)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_192),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g292 ( 
.A(n_233),
.Y(n_292)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

OAI22xp33_ASAP7_75t_L g235 ( 
.A1(n_200),
.A2(n_86),
.B1(n_76),
.B2(n_72),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_235),
.A2(n_248),
.B1(n_254),
.B2(n_267),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_236),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_144),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_237),
.B(n_240),
.Y(n_325)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_203),
.Y(n_238)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_238),
.Y(n_289)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_205),
.Y(n_239)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_239),
.Y(n_293)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_169),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_144),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_242),
.B(n_247),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_133),
.B(n_0),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_243),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_191),
.A2(n_71),
.B1(n_69),
.B2(n_66),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_244),
.A2(n_211),
.B1(n_170),
.B2(n_193),
.Y(n_333)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_245),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_177),
.A2(n_63),
.B1(n_21),
.B2(n_25),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_179),
.A2(n_28),
.B1(n_25),
.B2(n_11),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_180),
.Y(n_249)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_155),
.B(n_1),
.Y(n_250)
);

AND2x2_ASAP7_75t_SL g326 ( 
.A(n_250),
.B(n_282),
.Y(n_326)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_131),
.Y(n_251)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_251),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_170),
.Y(n_252)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_252),
.Y(n_332)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_140),
.Y(n_253)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_138),
.A2(n_28),
.B1(n_25),
.B2(n_11),
.Y(n_254)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_158),
.Y(n_256)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_256),
.Y(n_342)
);

NAND2xp33_ASAP7_75t_SL g345 ( 
.A(n_257),
.B(n_284),
.Y(n_345)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_194),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_176),
.Y(n_259)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_259),
.B(n_261),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_138),
.A2(n_28),
.B1(n_25),
.B2(n_13),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_143),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_266),
.Y(n_311)
);

OAI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_152),
.A2(n_18),
.B1(n_14),
.B2(n_13),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_L g299 ( 
.A1(n_263),
.A2(n_172),
.B1(n_154),
.B2(n_195),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_182),
.A2(n_13),
.B1(n_18),
.B2(n_3),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g267 ( 
.A1(n_198),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_150),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_268),
.B(n_273),
.Y(n_340)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_185),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_269),
.Y(n_317)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_176),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_270),
.B(n_272),
.Y(n_328)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_145),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_153),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_274),
.B(n_278),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_135),
.B(n_1),
.C(n_3),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_275),
.B(n_164),
.C(n_148),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g277 ( 
.A1(n_153),
.A2(n_5),
.B1(n_1),
.B2(n_4),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_207),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_279),
.Y(n_318)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_132),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_280),
.Y(n_322)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_207),
.Y(n_281)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_281),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_137),
.B(n_4),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_172),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_283),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_150),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g329 ( 
.A(n_286),
.B(n_195),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_287),
.A2(n_149),
.B1(n_157),
.B2(n_188),
.Y(n_306)
);

OA22x2_ASAP7_75t_L g295 ( 
.A1(n_223),
.A2(n_190),
.B1(n_159),
.B2(n_132),
.Y(n_295)
);

O2A1O1Ixp33_ASAP7_75t_SL g388 ( 
.A1(n_295),
.A2(n_335),
.B(n_289),
.C(n_293),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_298),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_299),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_255),
.A2(n_142),
.B1(n_190),
.B2(n_188),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g392 ( 
.A1(n_300),
.A2(n_313),
.B1(n_290),
.B2(n_324),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_160),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_303),
.B(n_327),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_304),
.B(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_271),
.B(n_156),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_305),
.B(n_329),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_306),
.A2(n_333),
.B1(n_235),
.B2(n_283),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_255),
.A2(n_287),
.B1(n_276),
.B2(n_225),
.Y(n_313)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_319),
.B(n_211),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_229),
.B(n_208),
.C(n_175),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_175),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_282),
.B(n_196),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_338),
.B(n_339),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_196),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_257),
.A2(n_208),
.B1(n_213),
.B2(n_158),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_341),
.A2(n_347),
.B1(n_219),
.B2(n_217),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_L g357 ( 
.A1(n_344),
.A2(n_275),
.B(n_269),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_223),
.A2(n_213),
.B1(n_134),
.B2(n_193),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_243),
.B(n_273),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_348),
.B(n_251),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_349),
.B(n_354),
.Y(n_396)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_302),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_352),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_312),
.A2(n_225),
.B1(n_288),
.B2(n_250),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_353),
.A2(n_358),
.B1(n_380),
.B2(n_382),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_325),
.A2(n_215),
.B1(n_243),
.B2(n_228),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_290),
.Y(n_355)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_355),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_SL g356 ( 
.A(n_305),
.B(n_265),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_356),
.B(n_370),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_357),
.Y(n_413)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g419 ( 
.A(n_359),
.Y(n_419)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_292),
.Y(n_360)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_360),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_267),
.B1(n_231),
.B2(n_274),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_361),
.A2(n_364),
.B1(n_376),
.B2(n_379),
.Y(n_428)
);

AO22x1_ASAP7_75t_SL g362 ( 
.A1(n_312),
.A2(n_261),
.B1(n_253),
.B2(n_272),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_389),
.Y(n_417)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_292),
.Y(n_363)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_347),
.A2(n_239),
.B1(n_238),
.B2(n_233),
.Y(n_364)
);

MAJx2_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_227),
.C(n_280),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g425 ( 
.A(n_365),
.B(n_366),
.C(n_330),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_325),
.A2(n_278),
.B1(n_270),
.B2(n_259),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_345),
.A2(n_334),
.B(n_327),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_367),
.A2(n_375),
.B(n_328),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g369 ( 
.A(n_342),
.Y(n_369)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_369),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g370 ( 
.A(n_340),
.B(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_314),
.Y(n_371)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_371),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_SL g372 ( 
.A(n_303),
.B(n_281),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_372),
.B(n_386),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_345),
.A2(n_234),
.B(n_232),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_334),
.A2(n_245),
.B1(n_241),
.B2(n_252),
.Y(n_376)
);

INVx4_ASAP7_75t_L g377 ( 
.A(n_302),
.Y(n_377)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_377),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_378),
.B(n_395),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_297),
.A2(n_222),
.B1(n_236),
.B2(n_134),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g382 ( 
.A1(n_297),
.A2(n_256),
.B1(n_209),
.B2(n_4),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_341),
.A2(n_209),
.B1(n_308),
.B2(n_306),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g430 ( 
.A1(n_384),
.A2(n_385),
.B1(n_387),
.B2(n_388),
.Y(n_430)
);

OAI22xp33_ASAP7_75t_L g385 ( 
.A1(n_295),
.A2(n_209),
.B1(n_318),
.B2(n_291),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_320),
.B(n_301),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_333),
.A2(n_323),
.B1(n_295),
.B2(n_337),
.Y(n_387)
);

AOI22xp33_ASAP7_75t_L g389 ( 
.A1(n_295),
.A2(n_318),
.B1(n_291),
.B2(n_342),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_320),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_390),
.B(n_315),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_337),
.A2(n_308),
.B1(n_339),
.B2(n_338),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_391),
.B(n_393),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_296),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_326),
.B(n_304),
.Y(n_393)
);

BUFx2_ASAP7_75t_L g394 ( 
.A(n_294),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_394),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_326),
.B(n_329),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_326),
.C(n_311),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_401),
.B(n_406),
.C(n_407),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_403),
.A2(n_409),
.B(n_418),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_404),
.A2(n_368),
.B1(n_374),
.B2(n_384),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_350),
.B(n_326),
.Y(n_406)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_393),
.B(n_309),
.C(n_322),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_367),
.A2(n_322),
.B(n_317),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_395),
.B(n_321),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_410),
.B(n_414),
.C(n_415),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_390),
.B(n_331),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g437 ( 
.A(n_412),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g414 ( 
.A(n_365),
.B(n_335),
.C(n_331),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g415 ( 
.A(n_357),
.B(n_328),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_375),
.A2(n_317),
.B(n_330),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_372),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_420),
.B(n_383),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_391),
.B(n_321),
.C(n_328),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_421),
.B(n_423),
.C(n_427),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_370),
.B(n_321),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_315),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_424),
.B(n_381),
.Y(n_454)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_425),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_353),
.B(n_330),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_368),
.A2(n_324),
.B(n_336),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_431),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_SL g432 ( 
.A(n_387),
.B(n_332),
.C(n_307),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_432),
.B(n_362),
.C(n_376),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_363),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_435),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_445),
.Y(n_472)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_416),
.Y(n_438)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_438),
.Y(n_496)
);

CKINVDCx14_ASAP7_75t_R g473 ( 
.A(n_439),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_373),
.Y(n_440)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_416),
.Y(n_441)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_441),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g479 ( 
.A1(n_442),
.A2(n_460),
.B(n_431),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_430),
.A2(n_351),
.B1(n_379),
.B2(n_380),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_443),
.A2(n_451),
.B1(n_458),
.B2(n_468),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_398),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_430),
.A2(n_351),
.B1(n_382),
.B2(n_380),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_446),
.A2(n_413),
.B1(n_417),
.B2(n_396),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_401),
.B(n_378),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_447),
.B(n_448),
.C(n_467),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g448 ( 
.A(n_406),
.B(n_354),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_429),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_449),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_409),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_450),
.B(n_470),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_422),
.A2(n_361),
.B1(n_349),
.B2(n_388),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_429),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_452),
.B(n_454),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_455),
.Y(n_490)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_426),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_457),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_422),
.A2(n_388),
.B1(n_366),
.B2(n_374),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_373),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_462),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_418),
.B(n_362),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_426),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_SL g463 ( 
.A(n_403),
.B(n_371),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_SL g499 ( 
.A(n_463),
.B(n_355),
.C(n_377),
.Y(n_499)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_464),
.B(n_359),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g500 ( 
.A(n_465),
.B(n_447),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_433),
.B(n_362),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_433),
.A2(n_364),
.B1(n_358),
.B2(n_369),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_399),
.B(n_289),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_417),
.A2(n_428),
.B1(n_396),
.B2(n_399),
.Y(n_471)
);

INVxp33_ASAP7_75t_SL g488 ( 
.A(n_471),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_407),
.C(n_415),
.Y(n_477)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_477),
.B(n_484),
.C(n_487),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_478),
.A2(n_486),
.B1(n_501),
.B2(n_468),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_479),
.A2(n_480),
.B(n_441),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_466),
.A2(n_413),
.B(n_396),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_451),
.A2(n_428),
.B1(n_414),
.B2(n_410),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_481),
.A2(n_482),
.B1(n_442),
.B2(n_438),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_458),
.A2(n_432),
.B1(n_427),
.B2(n_423),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g483 ( 
.A(n_448),
.B(n_402),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g531 ( 
.A(n_483),
.B(n_316),
.C(n_343),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_453),
.B(n_421),
.C(n_402),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_446),
.A2(n_425),
.B1(n_411),
.B2(n_408),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_425),
.C(n_411),
.Y(n_487)
);

FAx1_ASAP7_75t_L g489 ( 
.A(n_469),
.B(n_419),
.CI(n_397),
.CON(n_489),
.SN(n_489)
);

AOI211xp5_ASAP7_75t_SL g507 ( 
.A1(n_489),
.A2(n_469),
.B(n_460),
.C(n_465),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_405),
.C(n_400),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_493),
.C(n_495),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g493 ( 
.A(n_461),
.B(n_405),
.C(n_400),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_461),
.B(n_369),
.C(n_293),
.Y(n_495)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g526 ( 
.A(n_500),
.B(n_457),
.Y(n_526)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_440),
.A2(n_397),
.B1(n_352),
.B2(n_360),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_444),
.B(n_467),
.C(n_459),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_502),
.B(n_439),
.C(n_437),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_504),
.B(n_462),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_473),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_505),
.B(n_517),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_507),
.A2(n_394),
.B(n_310),
.Y(n_555)
);

OAI22xp5_ASAP7_75t_SL g508 ( 
.A1(n_474),
.A2(n_444),
.B1(n_466),
.B2(n_460),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g559 ( 
.A1(n_508),
.A2(n_519),
.B1(n_294),
.B2(n_346),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g509 ( 
.A(n_483),
.B(n_455),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_509),
.B(n_531),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_511),
.B(n_516),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_455),
.C(n_445),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_512),
.B(n_530),
.C(n_475),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g536 ( 
.A1(n_513),
.A2(n_494),
.B1(n_515),
.B2(n_528),
.Y(n_536)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_476),
.Y(n_514)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_514),
.Y(n_537)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_497),
.Y(n_515)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_515),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_443),
.Y(n_516)
);

CKINVDCx16_ASAP7_75t_R g517 ( 
.A(n_472),
.Y(n_517)
);

XOR2xp5_ASAP7_75t_L g538 ( 
.A(n_518),
.B(n_526),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_474),
.A2(n_488),
.B1(n_481),
.B2(n_482),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_SL g535 ( 
.A1(n_520),
.A2(n_480),
.B(n_489),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_493),
.B(n_436),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_521),
.B(n_523),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_522),
.B(n_528),
.Y(n_539)
);

CKINVDCx16_ASAP7_75t_R g523 ( 
.A(n_472),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g525 ( 
.A1(n_490),
.A2(n_452),
.B1(n_449),
.B2(n_464),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g556 ( 
.A1(n_525),
.A2(n_534),
.B1(n_394),
.B2(n_296),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_487),
.B(n_495),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_533),
.Y(n_544)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_503),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_529),
.B(n_532),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g530 ( 
.A(n_491),
.B(n_332),
.C(n_307),
.Y(n_530)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_485),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_500),
.B(n_310),
.Y(n_533)
);

CKINVDCx14_ASAP7_75t_R g534 ( 
.A(n_485),
.Y(n_534)
);

OAI21xp5_ASAP7_75t_L g565 ( 
.A1(n_535),
.A2(n_551),
.B(n_555),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_536),
.A2(n_508),
.B1(n_519),
.B2(n_522),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_541),
.B(n_530),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_510),
.B(n_475),
.C(n_502),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_546),
.B(n_549),
.Y(n_571)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_512),
.B(n_486),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g561 ( 
.A(n_548),
.B(n_526),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_510),
.B(n_489),
.C(n_478),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g550 ( 
.A(n_527),
.B(n_479),
.C(n_494),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_550),
.B(n_553),
.C(n_554),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_L g551 ( 
.A1(n_520),
.A2(n_492),
.B(n_501),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_506),
.B(n_498),
.C(n_504),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_506),
.B(n_503),
.C(n_496),
.Y(n_554)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_556),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_516),
.B(n_316),
.C(n_343),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_557),
.B(n_336),
.C(n_544),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g558 ( 
.A1(n_513),
.A2(n_346),
.B1(n_296),
.B2(n_294),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_L g564 ( 
.A1(n_558),
.A2(n_559),
.B1(n_514),
.B2(n_529),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_560),
.A2(n_569),
.B1(n_537),
.B2(n_535),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g584 ( 
.A(n_561),
.B(n_538),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g562 ( 
.A(n_538),
.B(n_533),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g581 ( 
.A(n_562),
.B(n_563),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_536),
.A2(n_507),
.B1(n_524),
.B2(n_509),
.Y(n_563)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_564),
.A2(n_550),
.B1(n_540),
.B2(n_546),
.Y(n_586)
);

AND2x2_ASAP7_75t_SL g566 ( 
.A(n_549),
.B(n_511),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_566),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_567),
.B(n_570),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g569 ( 
.A1(n_551),
.A2(n_531),
.B1(n_346),
.B2(n_336),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_545),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_573),
.B(n_574),
.Y(n_588)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_541),
.B(n_544),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_543),
.B(n_542),
.Y(n_575)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_575),
.Y(n_583)
);

OAI22xp5_ASAP7_75t_L g576 ( 
.A1(n_547),
.A2(n_559),
.B1(n_555),
.B2(n_545),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_576),
.B(n_577),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_554),
.B(n_552),
.C(n_548),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_552),
.B(n_557),
.C(n_553),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_578),
.B(n_574),
.Y(n_597)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_539),
.Y(n_579)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_579),
.Y(n_585)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_539),
.Y(n_580)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_580),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g601 ( 
.A1(n_582),
.A2(n_586),
.B1(n_565),
.B2(n_560),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_584),
.B(n_590),
.Y(n_598)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_567),
.B(n_540),
.C(n_578),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_587),
.B(n_595),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g590 ( 
.A(n_562),
.B(n_561),
.Y(n_590)
);

HB1xp67_ASAP7_75t_L g594 ( 
.A(n_575),
.Y(n_594)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_594),
.Y(n_610)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_569),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_577),
.B(n_568),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_596),
.B(n_597),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_596),
.B(n_568),
.C(n_571),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_599),
.B(n_603),
.Y(n_613)
);

INVx6_ASAP7_75t_L g600 ( 
.A(n_593),
.Y(n_600)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_600),
.Y(n_614)
);

INVxp67_ASAP7_75t_L g612 ( 
.A(n_601),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g603 ( 
.A(n_588),
.B(n_566),
.C(n_573),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_591),
.B(n_572),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_605),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g605 ( 
.A(n_588),
.B(n_566),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g606 ( 
.A(n_583),
.B(n_565),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_606),
.B(n_608),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_592),
.B(n_563),
.Y(n_607)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_607),
.Y(n_621)
);

AOI21xp5_ASAP7_75t_L g608 ( 
.A1(n_582),
.A2(n_585),
.B(n_589),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_SL g611 ( 
.A1(n_586),
.A2(n_581),
.B1(n_587),
.B2(n_584),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_611),
.B(n_581),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_616),
.B(n_617),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_599),
.B(n_590),
.C(n_609),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_603),
.C(n_602),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_618),
.Y(n_623)
);

NOR2x1_ASAP7_75t_L g619 ( 
.A(n_601),
.B(n_610),
.Y(n_619)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_619),
.Y(n_622)
);

INVxp67_ASAP7_75t_L g624 ( 
.A(n_613),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_624),
.B(n_627),
.Y(n_631)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_615),
.Y(n_625)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_625),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g627 ( 
.A(n_617),
.B(n_600),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_614),
.Y(n_628)
);

AOI21xp5_ASAP7_75t_L g629 ( 
.A1(n_628),
.A2(n_618),
.B(n_620),
.Y(n_629)
);

NAND3xp33_ASAP7_75t_SL g633 ( 
.A(n_629),
.B(n_632),
.C(n_626),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g632 ( 
.A1(n_622),
.A2(n_621),
.B(n_612),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_633),
.A2(n_634),
.B(n_630),
.Y(n_635)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_631),
.B(n_623),
.C(n_612),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g636 ( 
.A1(n_635),
.A2(n_619),
.B(n_608),
.Y(n_636)
);

OAI211xp5_ASAP7_75t_L g637 ( 
.A1(n_636),
.A2(n_598),
.B(n_611),
.C(n_635),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_637),
.Y(n_638)
);


endmodule