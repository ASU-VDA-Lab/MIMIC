module fake_netlist_1_3497_n_788 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_93, n_51, n_96, n_39, n_788);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_93;
input n_51;
input n_96;
input n_39;
output n_788;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_755;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_760;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_650;
wire n_625;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g98 ( .A(n_49), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_30), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_92), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_19), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_57), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_25), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_86), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_58), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_7), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_94), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_63), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_3), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_1), .Y(n_110) );
INVx2_ASAP7_75t_SL g111 ( .A(n_69), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_38), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_75), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_61), .Y(n_114) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_43), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_50), .Y(n_116) );
BUFx3_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_24), .Y(n_118) );
BUFx10_ASAP7_75t_L g119 ( .A(n_33), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_72), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_21), .Y(n_122) );
INVx1_ASAP7_75t_SL g123 ( .A(n_47), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_73), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_39), .Y(n_125) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_6), .B(n_1), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_16), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_83), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_22), .Y(n_129) );
BUFx2_ASAP7_75t_SL g130 ( .A(n_41), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_23), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_91), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_46), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_88), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_108), .B(n_0), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_129), .Y(n_136) );
XNOR2xp5_ASAP7_75t_L g137 ( .A(n_109), .B(n_0), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_99), .Y(n_138) );
NOR2x1_ASAP7_75t_L g139 ( .A(n_98), .B(n_2), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_100), .Y(n_140) );
INVx5_ASAP7_75t_L g141 ( .A(n_129), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_111), .B(n_2), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_119), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_129), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_111), .B(n_3), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_101), .Y(n_147) );
AOI22xp5_ASAP7_75t_SL g148 ( .A1(n_109), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_102), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_117), .Y(n_150) );
NOR2x1_ASAP7_75t_L g151 ( .A(n_103), .B(n_105), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_114), .B(n_4), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_106), .B(n_5), .Y(n_154) );
INVx2_ASAP7_75t_SL g155 ( .A(n_119), .Y(n_155) );
NOR2xp33_ASAP7_75t_SL g156 ( .A(n_104), .B(n_53), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_136), .Y(n_157) );
INVx2_ASAP7_75t_SL g158 ( .A(n_144), .Y(n_158) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_144), .B(n_119), .Y(n_159) );
INVx4_ASAP7_75t_L g160 ( .A(n_146), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_136), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_138), .Y(n_162) );
INVx3_ASAP7_75t_L g163 ( .A(n_146), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_136), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_144), .B(n_106), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_135), .B(n_104), .Y(n_167) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_136), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_145), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
OR2x2_ASAP7_75t_L g171 ( .A(n_135), .B(n_110), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_140), .B(n_131), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_145), .Y(n_175) );
INVx4_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
NAND3xp33_ASAP7_75t_L g177 ( .A(n_142), .B(n_127), .C(n_133), .Y(n_177) );
INVxp67_ASAP7_75t_SL g178 ( .A(n_154), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_138), .Y(n_179) );
INVx1_ASAP7_75t_L g180 ( .A(n_143), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_143), .Y(n_182) );
INVx8_ASAP7_75t_L g183 ( .A(n_141), .Y(n_183) );
CKINVDCx5p33_ASAP7_75t_R g184 ( .A(n_137), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_155), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_141), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_139), .B(n_117), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g188 ( .A(n_151), .B(n_134), .C(n_133), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_155), .B(n_124), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_140), .B(n_131), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_150), .Y(n_191) );
INVx1_ASAP7_75t_SL g192 ( .A(n_137), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_147), .B(n_134), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_147), .B(n_130), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_173), .Y(n_195) );
INVx3_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
INVxp67_ASAP7_75t_L g197 ( .A(n_167), .Y(n_197) );
AND2x6_ASAP7_75t_SL g198 ( .A(n_184), .B(n_152), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_178), .B(n_149), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_163), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_185), .B(n_149), .Y(n_201) );
NOR2xp33_ASAP7_75t_L g202 ( .A(n_166), .B(n_153), .Y(n_202) );
AOI22xp5_ASAP7_75t_L g203 ( .A1(n_173), .A2(n_115), .B1(n_116), .B2(n_153), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g204 ( .A1(n_163), .A2(n_151), .B(n_148), .C(n_139), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_162), .Y(n_205) );
A2O1A1Ixp33_ASAP7_75t_L g206 ( .A1(n_163), .A2(n_150), .B(n_126), .C(n_132), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_160), .B(n_156), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_158), .B(n_107), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_158), .B(n_112), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_194), .B(n_113), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_194), .B(n_118), .Y(n_211) );
NOR2xp33_ASAP7_75t_SL g212 ( .A(n_160), .B(n_115), .Y(n_212) );
AOI22xp5_ASAP7_75t_L g213 ( .A1(n_167), .A2(n_116), .B1(n_128), .B2(n_120), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_162), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_192), .Y(n_215) );
INVxp67_ASAP7_75t_L g216 ( .A(n_190), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_159), .B(n_123), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
NAND2x1p5_ASAP7_75t_L g219 ( .A(n_160), .B(n_129), .Y(n_219) );
NAND2xp33_ASAP7_75t_L g220 ( .A(n_163), .B(n_125), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_189), .B(n_176), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_171), .B(n_122), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_170), .A2(n_141), .B(n_54), .Y(n_223) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_176), .A2(n_141), .B1(n_8), .B2(n_9), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_176), .B(n_141), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_176), .B(n_141), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_179), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_170), .Y(n_228) );
NOR2xp67_ASAP7_75t_SL g229 ( .A(n_170), .B(n_52), .Y(n_229) );
NOR3xp33_ASAP7_75t_L g230 ( .A(n_188), .B(n_7), .C(n_8), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_193), .B(n_9), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_170), .B(n_56), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_171), .B(n_10), .Y(n_233) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_177), .B(n_59), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_180), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_191), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_180), .B(n_10), .Y(n_237) );
NAND2xp5_ASAP7_75t_SL g238 ( .A(n_191), .B(n_60), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_195), .A2(n_187), .B1(n_191), .B2(n_182), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_221), .A2(n_182), .B(n_183), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g241 ( .A1(n_200), .A2(n_183), .B(n_191), .Y(n_241) );
BUFx2_ASAP7_75t_L g242 ( .A(n_215), .Y(n_242) );
NOR2x1_ASAP7_75t_L g243 ( .A(n_233), .B(n_186), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_200), .A2(n_183), .B(n_186), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_228), .A2(n_183), .B(n_186), .Y(n_245) );
AOI21x1_ASAP7_75t_L g246 ( .A1(n_229), .A2(n_164), .B(n_157), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_196), .B(n_183), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_L g248 ( .A1(n_202), .A2(n_187), .B(n_181), .C(n_175), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_212), .B(n_165), .Y(n_249) );
OAI21xp5_ASAP7_75t_L g250 ( .A1(n_228), .A2(n_187), .B(n_164), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g251 ( .A1(n_225), .A2(n_169), .B(n_181), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_199), .B(n_187), .Y(n_252) );
OAI21xp5_ASAP7_75t_L g253 ( .A1(n_206), .A2(n_187), .B(n_181), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_222), .B(n_187), .Y(n_254) );
OAI21xp5_ASAP7_75t_L g255 ( .A1(n_206), .A2(n_187), .B(n_175), .Y(n_255) );
BUFx6f_ASAP7_75t_L g256 ( .A(n_219), .Y(n_256) );
INVx2_ASAP7_75t_SL g257 ( .A(n_231), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_201), .B(n_11), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_207), .A2(n_175), .B(n_174), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_226), .A2(n_174), .B(n_172), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_196), .Y(n_261) );
NAND2x1_ASAP7_75t_L g262 ( .A(n_196), .B(n_174), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_210), .B(n_11), .Y(n_263) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_205), .A2(n_172), .B(n_169), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_211), .B(n_12), .Y(n_265) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_219), .A2(n_172), .B(n_169), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_204), .B(n_161), .C(n_157), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g268 ( .A1(n_214), .A2(n_161), .B(n_157), .C(n_168), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_197), .B(n_12), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_207), .A2(n_161), .B(n_168), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_223), .A2(n_168), .B(n_165), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_213), .B(n_13), .Y(n_272) );
INVx6_ASAP7_75t_L g273 ( .A(n_237), .Y(n_273) );
AO31x2_ASAP7_75t_L g274 ( .A1(n_248), .A2(n_204), .A3(n_234), .B(n_235), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_272), .B(n_203), .Y(n_275) );
BUFx2_ASAP7_75t_L g276 ( .A(n_242), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_266), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_271), .A2(n_232), .B(n_238), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_269), .B(n_216), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_257), .B(n_227), .Y(n_280) );
OAI22xp33_ASAP7_75t_L g281 ( .A1(n_273), .A2(n_215), .B1(n_224), .B2(n_218), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_240), .A2(n_230), .B(n_236), .C(n_232), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_240), .A2(n_236), .B(n_220), .C(n_217), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_273), .B(n_220), .Y(n_284) );
OR2x2_ASAP7_75t_L g285 ( .A(n_258), .B(n_208), .Y(n_285) );
NOR4xp25_ASAP7_75t_L g286 ( .A(n_263), .B(n_238), .C(n_209), .D(n_15), .Y(n_286) );
AO32x2_ASAP7_75t_L g287 ( .A1(n_253), .A2(n_198), .A3(n_14), .B1(n_15), .B2(n_16), .Y(n_287) );
AO31x2_ASAP7_75t_L g288 ( .A1(n_268), .A2(n_13), .A3(n_14), .B(n_17), .Y(n_288) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_273), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_265), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_246), .A2(n_66), .B(n_18), .Y(n_291) );
AO21x2_ASAP7_75t_L g292 ( .A1(n_255), .A2(n_168), .B(n_165), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_254), .B(n_17), .Y(n_293) );
AO21x1_ASAP7_75t_L g294 ( .A1(n_249), .A2(n_20), .B(n_26), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_261), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_252), .B(n_27), .Y(n_296) );
AOI221x1_ASAP7_75t_L g297 ( .A1(n_259), .A2(n_168), .B1(n_165), .B2(n_31), .C(n_34), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_277), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_280), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_275), .B(n_239), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_277), .Y(n_301) );
AOI21x1_ASAP7_75t_L g302 ( .A1(n_297), .A2(n_270), .B(n_259), .Y(n_302) );
BUFx4f_ASAP7_75t_SL g303 ( .A(n_276), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_280), .B(n_256), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_288), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_286), .A2(n_250), .B(n_267), .Y(n_306) );
AOI21x1_ASAP7_75t_L g307 ( .A1(n_278), .A2(n_243), .B(n_260), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_278), .A2(n_264), .B(n_241), .Y(n_308) );
OA21x2_ASAP7_75t_L g309 ( .A1(n_291), .A2(n_241), .B(n_244), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_291), .A2(n_251), .B(n_244), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_290), .B(n_256), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_295), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_288), .Y(n_313) );
INVx1_ASAP7_75t_L g314 ( .A(n_288), .Y(n_314) );
INVx4_ASAP7_75t_L g315 ( .A(n_289), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_294), .A2(n_245), .B(n_262), .Y(n_316) );
AO21x2_ASAP7_75t_L g317 ( .A1(n_292), .A2(n_256), .B(n_168), .Y(n_317) );
OAI21x1_ASAP7_75t_L g318 ( .A1(n_294), .A2(n_247), .B(n_165), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_292), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_292), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_282), .A2(n_247), .B(n_165), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_274), .B(n_28), .Y(n_322) );
BUFx10_ASAP7_75t_L g323 ( .A(n_299), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_298), .Y(n_324) );
INVx6_ASAP7_75t_L g325 ( .A(n_315), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_305), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_305), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g328 ( .A(n_303), .B(n_281), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_304), .B(n_287), .Y(n_329) );
HB1xp67_ASAP7_75t_L g330 ( .A(n_303), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_298), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_304), .B(n_287), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
OR2x2_ASAP7_75t_L g334 ( .A(n_299), .B(n_274), .Y(n_334) );
OAI21x1_ASAP7_75t_L g335 ( .A1(n_321), .A2(n_302), .B(n_318), .Y(n_335) );
BUFx6f_ASAP7_75t_L g336 ( .A(n_298), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_305), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_313), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
OR2x2_ASAP7_75t_L g341 ( .A(n_304), .B(n_274), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_314), .Y(n_342) );
AND2x2_ASAP7_75t_L g343 ( .A(n_311), .B(n_287), .Y(n_343) );
INVx2_ASAP7_75t_SL g344 ( .A(n_311), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_312), .Y(n_345) );
INVx2_ASAP7_75t_R g346 ( .A(n_322), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_298), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_312), .Y(n_348) );
BUFx10_ASAP7_75t_L g349 ( .A(n_315), .Y(n_349) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_315), .B(n_285), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_321), .A2(n_296), .B(n_293), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_301), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_300), .A2(n_285), .B1(n_284), .B2(n_279), .Y(n_353) );
AND2x2_ASAP7_75t_L g354 ( .A(n_322), .B(n_287), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_315), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_322), .B(n_287), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_315), .B(n_283), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_301), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_301), .Y(n_359) );
BUFx3_ASAP7_75t_L g360 ( .A(n_301), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_306), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_319), .Y(n_362) );
INVx3_ASAP7_75t_L g363 ( .A(n_360), .Y(n_363) );
OAI221xp5_ASAP7_75t_L g364 ( .A1(n_353), .A2(n_300), .B1(n_282), .B2(n_283), .C(n_320), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_341), .B(n_319), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_324), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_328), .A2(n_306), .B1(n_320), .B2(n_319), .Y(n_367) );
BUFx3_ASAP7_75t_L g368 ( .A(n_349), .Y(n_368) );
AND2x4_ASAP7_75t_L g369 ( .A(n_338), .B(n_320), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_341), .B(n_319), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_329), .B(n_306), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_324), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_345), .B(n_274), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_349), .Y(n_374) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_350), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_338), .Y(n_376) );
AOI21xp5_ASAP7_75t_SL g377 ( .A1(n_350), .A2(n_309), .B(n_306), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_331), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_329), .B(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_332), .B(n_320), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_339), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_330), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g383 ( .A(n_345), .B(n_29), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_332), .B(n_320), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_348), .B(n_288), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_348), .B(n_317), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_355), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_362), .B(n_317), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_331), .Y(n_390) );
OR2x2_ASAP7_75t_L g391 ( .A(n_334), .B(n_317), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_343), .B(n_317), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_339), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_344), .B(n_317), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_343), .B(n_308), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_347), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_354), .B(n_308), .Y(n_397) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_346), .A2(n_309), .B1(n_308), .B2(n_316), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_347), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_349), .Y(n_400) );
OR2x2_ASAP7_75t_L g401 ( .A(n_334), .B(n_309), .Y(n_401) );
OR2x6_ASAP7_75t_L g402 ( .A(n_357), .B(n_318), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_340), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_344), .B(n_309), .Y(n_404) );
CKINVDCx8_ASAP7_75t_R g405 ( .A(n_336), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_354), .B(n_307), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_362), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_356), .B(n_307), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_340), .Y(n_409) );
BUFx6f_ASAP7_75t_L g410 ( .A(n_336), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_360), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_352), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
NAND2x1p5_ASAP7_75t_L g414 ( .A(n_333), .B(n_309), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_356), .B(n_307), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_333), .B(n_318), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_342), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_333), .A2(n_309), .B1(n_310), .B2(n_316), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_342), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_358), .Y(n_420) );
BUFx3_ASAP7_75t_L g421 ( .A(n_325), .Y(n_421) );
INVx3_ASAP7_75t_L g422 ( .A(n_336), .Y(n_422) );
INVxp67_ASAP7_75t_SL g423 ( .A(n_358), .Y(n_423) );
BUFx2_ASAP7_75t_L g424 ( .A(n_325), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_325), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_325), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_326), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_326), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_359), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_359), .Y(n_430) );
AND2x4_ASAP7_75t_SL g431 ( .A(n_375), .B(n_323), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_407), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_376), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_423), .B(n_327), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_371), .B(n_337), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_407), .Y(n_436) );
INVx2_ASAP7_75t_SL g437 ( .A(n_368), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_392), .B(n_327), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_368), .Y(n_439) );
HB1xp67_ASAP7_75t_L g440 ( .A(n_388), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_368), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_376), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_392), .B(n_337), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_381), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_381), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_365), .B(n_336), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_393), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_374), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_371), .B(n_361), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_382), .B(n_323), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_379), .B(n_323), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_391), .B(n_346), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_407), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_412), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_393), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_379), .B(n_323), .Y(n_456) );
BUFx2_ASAP7_75t_L g457 ( .A(n_374), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_380), .B(n_346), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_412), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_380), .B(n_384), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_384), .B(n_336), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_397), .B(n_357), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_391), .B(n_357), .Y(n_463) );
NAND2x1_ASAP7_75t_L g464 ( .A(n_400), .B(n_335), .Y(n_464) );
AND2x4_ASAP7_75t_L g465 ( .A(n_369), .B(n_335), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_427), .B(n_351), .Y(n_466) );
AND2x4_ASAP7_75t_L g467 ( .A(n_369), .B(n_351), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_403), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_403), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_397), .B(n_310), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_412), .Y(n_471) );
AND2x4_ASAP7_75t_L g472 ( .A(n_369), .B(n_310), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_395), .B(n_302), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_395), .B(n_302), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_406), .B(n_316), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_406), .B(n_35), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_408), .B(n_36), .Y(n_478) );
HB1xp67_ASAP7_75t_L g479 ( .A(n_374), .Y(n_479) );
INVx1_ASAP7_75t_SL g480 ( .A(n_400), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_405), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_427), .B(n_37), .Y(n_482) );
INVx2_ASAP7_75t_L g483 ( .A(n_413), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_387), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_409), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_408), .B(n_40), .Y(n_486) );
AND2x4_ASAP7_75t_L g487 ( .A(n_369), .B(n_42), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_417), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_417), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_413), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_419), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_419), .Y(n_492) );
INVx2_ASAP7_75t_L g493 ( .A(n_413), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_415), .B(n_44), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_420), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_415), .B(n_45), .Y(n_496) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_389), .B(n_48), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_428), .B(n_51), .Y(n_498) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_420), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_428), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_420), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_365), .B(n_370), .Y(n_502) );
BUFx2_ASAP7_75t_L g503 ( .A(n_424), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_429), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_429), .Y(n_505) );
INVx3_ASAP7_75t_L g506 ( .A(n_405), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_429), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_430), .Y(n_508) );
NOR2xp67_ASAP7_75t_L g509 ( .A(n_363), .B(n_55), .Y(n_509) );
OR2x2_ASAP7_75t_L g510 ( .A(n_370), .B(n_62), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_430), .B(n_64), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_430), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_401), .B(n_65), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_390), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_401), .B(n_67), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_416), .B(n_68), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_366), .B(n_70), .Y(n_517) );
INVx3_ASAP7_75t_L g518 ( .A(n_363), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_416), .B(n_71), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_373), .B(n_74), .Y(n_520) );
AND2x2_ASAP7_75t_SL g521 ( .A(n_424), .B(n_76), .Y(n_521) );
AND2x4_ASAP7_75t_SL g522 ( .A(n_426), .B(n_78), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_389), .B(n_79), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_386), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_414), .B(n_80), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g526 ( .A(n_480), .B(n_425), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_524), .B(n_385), .Y(n_527) );
HB1xp67_ASAP7_75t_L g528 ( .A(n_499), .Y(n_528) );
BUFx2_ASAP7_75t_L g529 ( .A(n_457), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_460), .B(n_411), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_440), .Y(n_531) );
AND2x4_ASAP7_75t_L g532 ( .A(n_437), .B(n_363), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_433), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_460), .B(n_411), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_502), .B(n_394), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_450), .B(n_425), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_442), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_438), .B(n_367), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_445), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_447), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_455), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_468), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_438), .B(n_390), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_469), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_443), .B(n_390), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_502), .B(n_363), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_473), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_435), .B(n_411), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_443), .B(n_411), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_504), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_488), .Y(n_553) );
AND2x2_ASAP7_75t_SL g554 ( .A(n_521), .B(n_383), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_489), .Y(n_555) );
OR2x2_ASAP7_75t_L g556 ( .A(n_449), .B(n_372), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_491), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_434), .B(n_372), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_484), .B(n_425), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_500), .B(n_366), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_492), .B(n_378), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_501), .B(n_378), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_437), .B(n_421), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_462), .B(n_421), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_432), .Y(n_565) );
INVxp33_ASAP7_75t_L g566 ( .A(n_448), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_396), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_451), .B(n_396), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_479), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_507), .B(n_508), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_462), .B(n_421), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_512), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_432), .Y(n_573) );
OR2x6_ASAP7_75t_L g574 ( .A(n_439), .B(n_377), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g575 ( .A(n_450), .B(n_364), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_436), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_470), .B(n_399), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_456), .B(n_399), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_503), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_461), .B(n_414), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_470), .B(n_418), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_461), .B(n_414), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_439), .B(n_402), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_441), .B(n_402), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_436), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_446), .B(n_404), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_453), .B(n_418), .Y(n_587) );
INVx2_ASAP7_75t_SL g588 ( .A(n_441), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_463), .B(n_454), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_458), .B(n_402), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_453), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_454), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_458), .B(n_402), .Y(n_593) );
OR2x2_ASAP7_75t_L g594 ( .A(n_463), .B(n_377), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_513), .B(n_402), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_459), .B(n_398), .Y(n_596) );
INVxp67_ASAP7_75t_SL g597 ( .A(n_464), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_513), .B(n_422), .Y(n_598) );
OR2x2_ASAP7_75t_L g599 ( .A(n_459), .B(n_422), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_471), .B(n_422), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_471), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_483), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_515), .B(n_422), .Y(n_603) );
AND2x2_ASAP7_75t_SL g604 ( .A(n_521), .B(n_410), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_515), .B(n_410), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_519), .B(n_410), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_519), .B(n_410), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_483), .B(n_410), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_490), .B(n_410), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_490), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_493), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_477), .B(n_81), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_493), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_495), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_495), .B(n_82), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_477), .B(n_84), .Y(n_616) );
NOR2x1p5_ASAP7_75t_L g617 ( .A(n_481), .B(n_85), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_514), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_478), .B(n_87), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_474), .B(n_89), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_474), .B(n_90), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_478), .B(n_93), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_530), .B(n_476), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_534), .B(n_476), .Y(n_624) );
NAND2x1p5_ASAP7_75t_L g625 ( .A(n_604), .B(n_487), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_531), .B(n_475), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g627 ( .A(n_566), .B(n_481), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_529), .B(n_481), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_528), .Y(n_629) );
AND2x4_ASAP7_75t_SL g630 ( .A(n_564), .B(n_506), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_581), .B(n_475), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g632 ( .A1(n_554), .A2(n_431), .B1(n_510), .B2(n_452), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_575), .B(n_506), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_533), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_539), .B(n_496), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_547), .B(n_518), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_528), .Y(n_637) );
OR2x2_ASAP7_75t_L g638 ( .A(n_535), .B(n_452), .Y(n_638) );
INVx1_ASAP7_75t_SL g639 ( .A(n_588), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_539), .B(n_486), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_579), .B(n_523), .C(n_497), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_581), .B(n_486), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_527), .B(n_496), .Y(n_643) );
O2A1O1Ixp33_ASAP7_75t_L g644 ( .A1(n_579), .A2(n_497), .B(n_523), .C(n_520), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_537), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_544), .B(n_514), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_538), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_527), .B(n_494), .Y(n_648) );
OR2x6_ASAP7_75t_L g649 ( .A(n_574), .B(n_487), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_540), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_551), .B(n_518), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_544), .B(n_466), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_546), .B(n_465), .Y(n_653) );
NAND2xp33_ASAP7_75t_L g654 ( .A(n_617), .B(n_525), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_541), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_552), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_542), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_543), .Y(n_658) );
NOR5xp2_ASAP7_75t_L g659 ( .A(n_597), .B(n_522), .C(n_509), .D(n_487), .E(n_516), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_546), .B(n_494), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_545), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_589), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_577), .B(n_472), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_548), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_532), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_577), .B(n_472), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_590), .B(n_518), .Y(n_667) );
AND2x2_ASAP7_75t_L g668 ( .A(n_593), .B(n_465), .Y(n_668) );
AND2x2_ASAP7_75t_L g669 ( .A(n_571), .B(n_465), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_550), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_553), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_555), .Y(n_672) );
INVx2_ASAP7_75t_SL g673 ( .A(n_563), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_557), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
NOR2xp67_ASAP7_75t_SL g676 ( .A(n_612), .B(n_616), .Y(n_676) );
NAND2x1_ASAP7_75t_SL g677 ( .A(n_532), .B(n_506), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_569), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_570), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_570), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_556), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_587), .B(n_472), .Y(n_682) );
AND2x2_ASAP7_75t_L g683 ( .A(n_580), .B(n_467), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_572), .Y(n_684) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_619), .B(n_525), .Y(n_685) );
INVx1_ASAP7_75t_SL g686 ( .A(n_563), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_587), .B(n_516), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_582), .B(n_467), .Y(n_688) );
AND2x2_ASAP7_75t_L g689 ( .A(n_559), .B(n_467), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_573), .B(n_516), .Y(n_690) );
CKINVDCx14_ASAP7_75t_R g691 ( .A(n_526), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_583), .B(n_431), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_560), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_679), .Y(n_694) );
NAND2x2_ASAP7_75t_L g695 ( .A(n_673), .B(n_594), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_685), .A2(n_574), .B1(n_549), .B2(n_536), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_680), .Y(n_697) );
O2A1O1Ixp5_ASAP7_75t_L g698 ( .A1(n_676), .A2(n_597), .B(n_596), .C(n_584), .Y(n_698) );
INVx2_ASAP7_75t_L g699 ( .A(n_629), .Y(n_699) );
O2A1O1Ixp33_ASAP7_75t_L g700 ( .A1(n_633), .A2(n_621), .B(n_620), .C(n_596), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_693), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_684), .Y(n_702) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_637), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_668), .B(n_574), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_631), .B(n_681), .Y(n_705) );
INVx1_ASAP7_75t_L g706 ( .A(n_634), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_645), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_647), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_632), .A2(n_595), .B1(n_603), .B2(n_598), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_631), .B(n_586), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g711 ( .A1(n_641), .A2(n_622), .B(n_621), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_654), .A2(n_567), .B(n_562), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_638), .B(n_568), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_691), .B(n_578), .Y(n_714) );
OR2x2_ASAP7_75t_L g715 ( .A(n_626), .B(n_592), .Y(n_715) );
INVx4_ASAP7_75t_L g716 ( .A(n_649), .Y(n_716) );
O2A1O1Ixp33_ASAP7_75t_SL g717 ( .A1(n_639), .A2(n_620), .B(n_561), .C(n_560), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_650), .Y(n_718) );
OAI211xp5_ASAP7_75t_L g719 ( .A1(n_677), .A2(n_600), .B(n_561), .C(n_606), .Y(n_719) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_656), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_632), .A2(n_607), .B1(n_605), .B2(n_613), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_655), .Y(n_722) );
INVxp67_ASAP7_75t_SL g723 ( .A(n_659), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_657), .Y(n_724) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_639), .B(n_600), .Y(n_725) );
A2O1A1Ixp33_ASAP7_75t_L g726 ( .A1(n_644), .A2(n_522), .B(n_511), .C(n_562), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_652), .B(n_602), .Y(n_727) );
O2A1O1Ixp33_ASAP7_75t_L g728 ( .A1(n_678), .A2(n_498), .B(n_482), .C(n_615), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_652), .B(n_585), .Y(n_729) );
NAND4xp25_ASAP7_75t_L g730 ( .A(n_641), .B(n_567), .C(n_599), .D(n_608), .Y(n_730) );
NAND2x1_ASAP7_75t_L g731 ( .A(n_649), .B(n_614), .Y(n_731) );
INVx1_ASAP7_75t_L g732 ( .A(n_658), .Y(n_732) );
HB1xp67_ASAP7_75t_L g733 ( .A(n_653), .Y(n_733) );
AND2x2_ASAP7_75t_L g734 ( .A(n_669), .B(n_611), .Y(n_734) );
AOI322xp5_ASAP7_75t_L g735 ( .A1(n_723), .A2(n_653), .A3(n_686), .B1(n_642), .B2(n_635), .C1(n_640), .C2(n_628), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g736 ( .A1(n_730), .A2(n_682), .B(n_663), .Y(n_736) );
OAI222xp33_ASAP7_75t_L g737 ( .A1(n_716), .A2(n_649), .B1(n_686), .B2(n_665), .C1(n_625), .C2(n_685), .Y(n_737) );
INVx1_ASAP7_75t_L g738 ( .A(n_701), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_727), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_696), .A2(n_627), .B1(n_665), .B2(n_666), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g741 ( .A1(n_696), .A2(n_695), .B1(n_716), .B2(n_721), .Y(n_741) );
AOI211xp5_ASAP7_75t_L g742 ( .A1(n_711), .A2(n_643), .B(n_648), .C(n_687), .Y(n_742) );
AOI322xp5_ASAP7_75t_L g743 ( .A1(n_714), .A2(n_624), .A3(n_623), .B1(n_660), .B2(n_662), .C1(n_675), .C2(n_636), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g744 ( .A1(n_698), .A2(n_625), .B(n_630), .Y(n_744) );
O2A1O1Ixp33_ASAP7_75t_L g745 ( .A1(n_711), .A2(n_674), .B(n_664), .C(n_661), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_729), .Y(n_746) );
NOR2xp67_ASAP7_75t_L g747 ( .A(n_719), .B(n_646), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_733), .B(n_670), .Y(n_748) );
AOI221x1_ASAP7_75t_SL g749 ( .A1(n_730), .A2(n_671), .B1(n_672), .B2(n_690), .C(n_576), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_705), .B(n_689), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_731), .A2(n_688), .B1(n_683), .B2(n_651), .Y(n_751) );
OA22x2_ASAP7_75t_L g752 ( .A1(n_709), .A2(n_692), .B1(n_667), .B2(n_690), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_725), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_712), .B(n_591), .Y(n_754) );
INVx1_ASAP7_75t_SL g755 ( .A(n_720), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_694), .B(n_601), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_749), .B(n_697), .Y(n_757) );
AOI31xp33_ASAP7_75t_L g758 ( .A1(n_744), .A2(n_726), .A3(n_717), .B(n_704), .Y(n_758) );
AOI21xp5_ASAP7_75t_SL g759 ( .A1(n_745), .A2(n_700), .B(n_728), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_755), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_752), .A2(n_702), .B1(n_732), .B2(n_724), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_748), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_741), .B(n_699), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_740), .A2(n_706), .B1(n_722), .B2(n_718), .C(n_707), .Y(n_764) );
NOR3xp33_ASAP7_75t_SL g765 ( .A(n_737), .B(n_708), .C(n_608), .Y(n_765) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_752), .A2(n_703), .B(n_715), .Y(n_766) );
OAI211xp5_ASAP7_75t_L g767 ( .A1(n_735), .A2(n_710), .B(n_713), .C(n_734), .Y(n_767) );
AOI221xp5_ASAP7_75t_L g768 ( .A1(n_759), .A2(n_753), .B1(n_736), .B2(n_739), .C(n_746), .Y(n_768) );
OAI21xp5_ASAP7_75t_L g769 ( .A1(n_766), .A2(n_747), .B(n_743), .Y(n_769) );
NOR2xp33_ASAP7_75t_SL g770 ( .A(n_760), .B(n_751), .Y(n_770) );
AND5x1_ASAP7_75t_L g771 ( .A(n_761), .B(n_742), .C(n_750), .D(n_754), .E(n_738), .Y(n_771) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_762), .B(n_756), .Y(n_772) );
XOR2x2_ASAP7_75t_L g773 ( .A(n_763), .B(n_517), .Y(n_773) );
NAND4xp25_ASAP7_75t_L g774 ( .A(n_768), .B(n_757), .C(n_767), .D(n_764), .Y(n_774) );
NOR2x1_ASAP7_75t_L g775 ( .A(n_769), .B(n_758), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_772), .Y(n_776) );
NAND2xp5_ASAP7_75t_SL g777 ( .A(n_775), .B(n_770), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_776), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_778), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_777), .B(n_774), .Y(n_780) );
OAI22x1_ASAP7_75t_L g781 ( .A1(n_780), .A2(n_771), .B1(n_765), .B2(n_773), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_779), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_782), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_783), .B(n_781), .Y(n_784) );
AOI21xp33_ASAP7_75t_SL g785 ( .A1(n_784), .A2(n_765), .B(n_96), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_785), .B(n_95), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g787 ( .A1(n_786), .A2(n_97), .B(n_565), .Y(n_787) );
AOI22xp33_ASAP7_75t_SL g788 ( .A1(n_787), .A2(n_610), .B1(n_618), .B2(n_609), .Y(n_788) );
endmodule