module real_jpeg_17072_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_0),
.B(n_70),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_0),
.B(n_127),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_0),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_0),
.B(n_279),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_0),
.B(n_385),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_0),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_0),
.B(n_406),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_1),
.B(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_1),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_1),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_2),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_2),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_2),
.B(n_350),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_2),
.B(n_374),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_2),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_2),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_2),
.B(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_3),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_3),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_4),
.Y(n_106)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_4),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_4),
.Y(n_236)
);

BUFx5_ASAP7_75t_L g377 ( 
.A(n_4),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_5),
.B(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_5),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_5),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_5),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_28),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_5),
.A2(n_12),
.B1(n_212),
.B2(n_215),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g315 ( 
.A(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_6),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_6),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_6),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_6),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_6),
.B(n_52),
.Y(n_183)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_7),
.Y(n_214)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_7),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g328 ( 
.A(n_7),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

NAND2x1_ASAP7_75t_L g91 ( 
.A(n_8),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_8),
.B(n_176),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g190 ( 
.A(n_8),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g225 ( 
.A(n_8),
.B(n_226),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_8),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_8),
.B(n_323),
.Y(n_322)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_8),
.B(n_52),
.Y(n_392)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_9),
.Y(n_76)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_9),
.Y(n_125)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_9),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_9),
.Y(n_228)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_9),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_10),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_10),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_10),
.B(n_221),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_10),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_10),
.B(n_52),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_11),
.B(n_78),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_11),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_11),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_11),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_11),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_232),
.Y(n_231)
);

INVxp33_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_11),
.B(n_326),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_12),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_12),
.B(n_166),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_12),
.B(n_275),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_12),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_12),
.B(n_353),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_12),
.B(n_377),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_12),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_12),
.B(n_413),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_13),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_13),
.Y(n_111)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_13),
.Y(n_334)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_14),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_14),
.Y(n_118)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g187 ( 
.A(n_15),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_15),
.Y(n_391)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_16),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_198),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_196),
.Y(n_18)
);

INVxp67_ASAP7_75t_SL g19 ( 
.A(n_20),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_154),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_22),
.B(n_154),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_97),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_67),
.C(n_89),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g155 ( 
.A(n_25),
.B(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_43),
.C(n_53),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_26),
.B(n_43),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_31),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_27),
.B(n_32),
.C(n_39),
.Y(n_149)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_30),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_39),
.Y(n_31)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_51),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_44),
.B(n_162),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_47),
.A2(n_51),
.B1(n_65),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_47),
.Y(n_163)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_49),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_50),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_51),
.A2(n_61),
.B1(n_65),
.B2(n_66),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_51),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_55),
.C(n_61),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_53),
.B(n_251),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_54),
.B(n_219),
.C(n_220),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_54),
.A2(n_55),
.B1(n_220),
.B2(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_57),
.Y(n_55)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_57),
.Y(n_121)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_61),
.A2(n_66),
.B1(n_103),
.B2(n_104),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_62),
.B(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_64),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_64),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_66),
.B(n_104),
.C(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_67),
.B(n_89),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.C(n_84),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_68),
.B(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_73),
.C(n_77),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_69),
.B(n_77),
.Y(n_180)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_73),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_79),
.Y(n_144)
);

BUFx5_ASAP7_75t_L g275 ( 
.A(n_79),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_80),
.Y(n_195)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_82),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_83),
.Y(n_93)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_SL g90 ( 
.A(n_85),
.B(n_91),
.Y(n_90)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_85),
.B(n_91),
.C(n_96),
.Y(n_131)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_88),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_89)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_91),
.B(n_183),
.C(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx5_ASAP7_75t_L g136 ( 
.A(n_93),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_94),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_129),
.B1(n_152),
.B2(n_153),
.Y(n_97)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_98),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_112),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_100),
.B(n_108),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_104),
.B2(n_107),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_101),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g103 ( 
.A(n_104),
.Y(n_103)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_106),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_119),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_118),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_118),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.C(n_126),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_120),
.B(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_126),
.Y(n_148)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_129),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_146),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_132),
.Y(n_130)
);

XNOR2x1_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_141),
.B1(n_142),
.B2(n_145),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_138),
.Y(n_145)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx5_ASAP7_75t_L g375 ( 
.A(n_144),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_149),
.C(n_150),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_149),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_158),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.C(n_159),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_155),
.B(n_157),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_159),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_181),
.C(n_193),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_160),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_164),
.C(n_179),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_161),
.B(n_164),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_174),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_165),
.A2(n_174),
.B1(n_175),
.B2(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_169),
.B(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_173),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_174),
.B(n_349),
.C(n_352),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_174),
.A2(n_175),
.B1(n_349),
.B2(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2x2_ASAP7_75t_SL g260 ( 
.A(n_179),
.B(n_261),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_181),
.B(n_193),
.Y(n_249)
);

MAJx2_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.C(n_189),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_182),
.B(n_245),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_183),
.B(n_184),
.Y(n_209)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_188),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_189),
.A2(n_190),
.B1(n_330),
.B2(n_331),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_190),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_192),
.Y(n_313)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

AO21x2_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_293),
.B(n_468),
.Y(n_199)
);

NOR2xp67_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_287),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_254),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g469 ( 
.A(n_202),
.B(n_254),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_247),
.Y(n_202)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_203),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_223),
.C(n_242),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_205),
.B(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_210),
.C(n_218),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_206),
.B(n_336),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_210),
.A2(n_211),
.B1(n_218),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_211),
.A2(n_309),
.B(n_314),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_213),
.Y(n_386)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

BUFx3_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_218),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_219),
.B(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_222),
.B(n_271),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_223),
.A2(n_243),
.B1(n_244),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_223),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_234),
.C(n_237),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_224),
.B(n_282),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.C(n_231),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_225),
.A2(n_231),
.B1(n_306),
.B2(n_307),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_225),
.B(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_229),
.B(n_305),
.Y(n_304)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_231),
.Y(n_307)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_234),
.A2(n_235),
.B1(n_237),
.B2(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_237),
.Y(n_283)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_247)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_248),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_250),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_252),
.B(n_291),
.C(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_260),
.C(n_262),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_256),
.A2(n_257),
.B1(n_260),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g262 ( 
.A(n_263),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_263),
.B(n_297),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_281),
.C(n_284),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_264),
.B(n_302),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.C(n_273),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_266),
.B(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_269),
.B(n_273),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_270),
.B(n_272),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_276),
.C(n_278),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_274),
.A2(n_276),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_274),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_276),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_276),
.A2(n_346),
.B1(n_422),
.B2(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_276),
.B(n_418),
.C(n_422),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_278),
.B(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_284),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_287),
.A2(n_469),
.B(n_470),
.Y(n_468)
);

AND2x2_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_290),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g470 ( 
.A(n_288),
.B(n_290),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_364),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_299),
.C(n_338),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_296),
.B(n_300),
.Y(n_467)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_303),
.C(n_335),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_301),
.B(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g363 ( 
.A(n_303),
.B(n_335),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_308),
.C(n_320),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_308),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_306),
.B(n_373),
.C(n_376),
.Y(n_397)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_316),
.Y(n_314)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx4_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g340 ( 
.A(n_320),
.B(n_341),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_329),
.C(n_330),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_321),
.B(n_454),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_325),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_322),
.B(n_325),
.Y(n_404)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_322),
.A2(n_411),
.B1(n_412),
.B2(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2x1_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_362),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_362),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.C(n_359),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_340),
.B(n_465),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_342),
.B(n_360),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_347),
.C(n_357),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_343),
.B(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_348),
.B(n_358),
.Y(n_459)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

XOR2x2_ASAP7_75t_L g398 ( 
.A(n_352),
.B(n_399),
.Y(n_398)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

NAND3xp33_ASAP7_75t_SL g364 ( 
.A(n_365),
.B(n_366),
.C(n_467),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_462),
.B(n_466),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_368),
.A2(n_448),
.B(n_461),
.Y(n_367)
);

OAI21x1_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_407),
.B(n_447),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_395),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g447 ( 
.A(n_370),
.B(n_395),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_378),
.C(n_387),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_371),
.B(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_377),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_378),
.A2(n_379),
.B1(n_387),
.B2(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_384),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_SL g419 ( 
.A(n_380),
.B(n_384),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx4_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx6_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

AO22x1_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_392),
.B1(n_393),
.B2(n_394),
.Y(n_387)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_388),
.Y(n_393)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_392),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_393),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_394),
.B(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_397),
.B(n_398),
.C(n_401),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_403),
.Y(n_401)
);

MAJx2_ASAP7_75t_L g456 ( 
.A(n_402),
.B(n_404),
.C(n_405),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_405),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_408),
.A2(n_441),
.B(n_446),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_409),
.A2(n_425),
.B(n_440),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_417),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_410),
.B(n_417),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_412),
.Y(n_433)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_SL g414 ( 
.A(n_415),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_420),
.B2(n_421),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_426),
.A2(n_434),
.B(n_439),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_432),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_427),
.B(n_432),
.Y(n_439)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_442),
.B(n_445),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_449),
.B(n_460),
.Y(n_448)
);

NOR2xp67_ASAP7_75t_SL g461 ( 
.A(n_449),
.B(n_460),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_450),
.A2(n_451),
.B1(n_457),
.B2(n_458),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_455),
.B2(n_456),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_452),
.B(n_456),
.C(n_457),
.Y(n_463)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

NOR2x1_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_464),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_463),
.B(n_464),
.Y(n_466)
);


endmodule