module fake_netlist_1_2878_n_1384 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_336, n_348, n_252, n_152, n_113, n_353, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_334, n_275, n_0, n_131, n_112, n_205, n_330, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_351, n_83, n_28, n_48, n_100, n_305, n_228, n_345, n_236, n_340, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_333, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_354, n_32, n_235, n_243, n_331, n_352, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_338, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_342, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_344, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_349, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_339, n_240, n_346, n_103, n_180, n_104, n_74, n_335, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_343, n_127, n_291, n_170, n_281, n_341, n_58, n_122, n_187, n_138, n_323, n_347, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_355, n_226, n_159, n_337, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_332, n_350, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1384);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_336;
input n_348;
input n_252;
input n_152;
input n_113;
input n_353;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_334;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_330;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_351;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_345;
input n_236;
input n_340;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_333;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_354;
input n_32;
input n_235;
input n_243;
input n_331;
input n_352;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_338;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_342;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_344;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_349;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_339;
input n_240;
input n_346;
input n_103;
input n_180;
input n_104;
input n_74;
input n_335;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_343;
input n_127;
input n_291;
input n_170;
input n_281;
input n_341;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_347;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_355;
input n_226;
input n_159;
input n_337;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_332;
input n_350;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1384;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_545;
wire n_896;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1209;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1240;
wire n_1139;
wire n_577;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1102;
wire n_723;
wire n_972;
wire n_997;
wire n_1244;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_359;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_930;
wire n_994;
wire n_410;
wire n_774;
wire n_1207;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_382;
wire n_658;
wire n_691;
wire n_444;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_1306;
wire n_958;
wire n_468;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_796;
wire n_1216;
wire n_927;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_799;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_1157;
wire n_806;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1117;
wire n_1007;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_834;
wire n_901;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_1292;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_1087;
wire n_662;
wire n_1372;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_882;
wire n_871;
wire n_803;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1058;
wire n_388;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_615;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_397;
wire n_1109;
wire n_1008;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_458;
wire n_1084;
wire n_618;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_538;
wire n_492;
wire n_1150;
wire n_1327;
wire n_368;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_1022;
wire n_802;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_401;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_955;
wire n_1275;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_455;
wire n_529;
wire n_1025;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1160;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_374;
wire n_718;
wire n_1238;
wire n_1114;
wire n_1304;
wire n_948;
wire n_1286;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1021;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_700;
wire n_534;
wire n_1296;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_967;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_695;
wire n_1104;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g356 ( .A(n_244), .Y(n_356) );
CKINVDCx5p33_ASAP7_75t_R g357 ( .A(n_234), .Y(n_357) );
INVx1_ASAP7_75t_SL g358 ( .A(n_31), .Y(n_358) );
CKINVDCx5p33_ASAP7_75t_R g359 ( .A(n_343), .Y(n_359) );
CKINVDCx16_ASAP7_75t_R g360 ( .A(n_183), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_107), .Y(n_361) );
INVx4_ASAP7_75t_R g362 ( .A(n_200), .Y(n_362) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_235), .B(n_82), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_325), .Y(n_364) );
NOR2xp67_ASAP7_75t_L g365 ( .A(n_48), .B(n_148), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_96), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_310), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_100), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_216), .Y(n_369) );
CKINVDCx5p33_ASAP7_75t_R g370 ( .A(n_91), .Y(n_370) );
INVx1_ASAP7_75t_SL g371 ( .A(n_340), .Y(n_371) );
CKINVDCx20_ASAP7_75t_R g372 ( .A(n_2), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_38), .Y(n_373) );
BUFx3_ASAP7_75t_L g374 ( .A(n_85), .Y(n_374) );
INVx1_ASAP7_75t_SL g375 ( .A(n_88), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_35), .Y(n_376) );
INVx1_ASAP7_75t_SL g377 ( .A(n_156), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_184), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_321), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_220), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_113), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_140), .Y(n_382) );
CKINVDCx5p33_ASAP7_75t_R g383 ( .A(n_329), .Y(n_383) );
CKINVDCx5p33_ASAP7_75t_R g384 ( .A(n_162), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_192), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_294), .Y(n_386) );
BUFx6f_ASAP7_75t_L g387 ( .A(n_127), .Y(n_387) );
INVxp67_ASAP7_75t_SL g388 ( .A(n_304), .Y(n_388) );
CKINVDCx5p33_ASAP7_75t_R g389 ( .A(n_178), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_324), .Y(n_390) );
CKINVDCx5p33_ASAP7_75t_R g391 ( .A(n_223), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_204), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_328), .Y(n_393) );
CKINVDCx20_ASAP7_75t_R g394 ( .A(n_277), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g395 ( .A(n_99), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g396 ( .A(n_303), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_188), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_335), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_14), .Y(n_399) );
INVxp67_ASAP7_75t_L g400 ( .A(n_5), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_39), .Y(n_401) );
CKINVDCx5p33_ASAP7_75t_R g402 ( .A(n_172), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_222), .Y(n_403) );
INVxp67_ASAP7_75t_L g404 ( .A(n_142), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_215), .Y(n_405) );
CKINVDCx16_ASAP7_75t_R g406 ( .A(n_225), .Y(n_406) );
CKINVDCx20_ASAP7_75t_R g407 ( .A(n_259), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_334), .Y(n_408) );
INVx1_ASAP7_75t_SL g409 ( .A(n_344), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g410 ( .A(n_289), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_147), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g412 ( .A(n_70), .Y(n_412) );
CKINVDCx20_ASAP7_75t_R g413 ( .A(n_106), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_152), .Y(n_414) );
CKINVDCx5p33_ASAP7_75t_R g415 ( .A(n_133), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_240), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_137), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_266), .Y(n_418) );
BUFx5_ASAP7_75t_L g419 ( .A(n_231), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_213), .Y(n_420) );
CKINVDCx16_ASAP7_75t_R g421 ( .A(n_168), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_296), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_59), .Y(n_423) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_70), .B(n_115), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_330), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_336), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_252), .Y(n_427) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_275), .Y(n_428) );
CKINVDCx5p33_ASAP7_75t_R g429 ( .A(n_260), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_278), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_43), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_122), .Y(n_432) );
INVx2_ASAP7_75t_SL g433 ( .A(n_108), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_238), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_268), .B(n_158), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_273), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_239), .B(n_152), .Y(n_437) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_115), .Y(n_438) );
CKINVDCx5p33_ASAP7_75t_R g439 ( .A(n_122), .Y(n_439) );
INVxp67_ASAP7_75t_L g440 ( .A(n_311), .Y(n_440) );
BUFx6f_ASAP7_75t_L g441 ( .A(n_263), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_124), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_104), .Y(n_443) );
CKINVDCx5p33_ASAP7_75t_R g444 ( .A(n_14), .Y(n_444) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_298), .Y(n_445) );
CKINVDCx16_ASAP7_75t_R g446 ( .A(n_265), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_341), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_144), .Y(n_448) );
INVx2_ASAP7_75t_SL g449 ( .A(n_209), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_136), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_3), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_320), .B(n_288), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_46), .Y(n_453) );
CKINVDCx5p33_ASAP7_75t_R g454 ( .A(n_241), .Y(n_454) );
CKINVDCx5p33_ASAP7_75t_R g455 ( .A(n_194), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_138), .Y(n_456) );
BUFx6f_ASAP7_75t_L g457 ( .A(n_164), .Y(n_457) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_269), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_51), .Y(n_459) );
BUFx6f_ASAP7_75t_L g460 ( .A(n_312), .Y(n_460) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_196), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_295), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_89), .Y(n_463) );
NOR2xp67_ASAP7_75t_L g464 ( .A(n_339), .B(n_224), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_270), .Y(n_465) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_208), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_337), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_332), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_313), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_267), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_202), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_86), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_205), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_354), .Y(n_474) );
BUFx3_ASAP7_75t_L g475 ( .A(n_319), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_258), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_195), .Y(n_477) );
CKINVDCx5p33_ASAP7_75t_R g478 ( .A(n_22), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_127), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_148), .Y(n_480) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_93), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_217), .Y(n_482) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_232), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_9), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_249), .Y(n_485) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_153), .Y(n_486) );
CKINVDCx5p33_ASAP7_75t_R g487 ( .A(n_80), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_101), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_170), .Y(n_489) );
INVxp67_ASAP7_75t_SL g490 ( .A(n_307), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_250), .Y(n_491) );
CKINVDCx5p33_ASAP7_75t_R g492 ( .A(n_24), .Y(n_492) );
CKINVDCx5p33_ASAP7_75t_R g493 ( .A(n_233), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_246), .Y(n_494) );
CKINVDCx5p33_ASAP7_75t_R g495 ( .A(n_163), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g496 ( .A(n_128), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_54), .Y(n_497) );
CKINVDCx5p33_ASAP7_75t_R g498 ( .A(n_64), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_17), .Y(n_499) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_345), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_26), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_284), .Y(n_502) );
BUFx5_ASAP7_75t_L g503 ( .A(n_112), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_186), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_82), .Y(n_505) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_218), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_228), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_134), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_212), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_306), .Y(n_510) );
CKINVDCx5p33_ASAP7_75t_R g511 ( .A(n_141), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_103), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_65), .Y(n_513) );
INVxp33_ASAP7_75t_L g514 ( .A(n_77), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_80), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_56), .Y(n_516) );
CKINVDCx5p33_ASAP7_75t_R g517 ( .A(n_333), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g518 ( .A(n_37), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_226), .Y(n_519) );
CKINVDCx5p33_ASAP7_75t_R g520 ( .A(n_261), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_120), .Y(n_521) );
BUFx2_ASAP7_75t_SL g522 ( .A(n_146), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_198), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_179), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_352), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_176), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_227), .Y(n_527) );
INVx2_ASAP7_75t_L g528 ( .A(n_274), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_264), .Y(n_529) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_33), .Y(n_530) );
CKINVDCx5p33_ASAP7_75t_R g531 ( .A(n_297), .Y(n_531) );
INVxp33_ASAP7_75t_SL g532 ( .A(n_104), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_36), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_120), .Y(n_534) );
CKINVDCx5p33_ASAP7_75t_R g535 ( .A(n_64), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_24), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_124), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_193), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_281), .Y(n_539) );
CKINVDCx5p33_ASAP7_75t_R g540 ( .A(n_43), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_342), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g542 ( .A(n_129), .Y(n_542) );
CKINVDCx5p33_ASAP7_75t_R g543 ( .A(n_22), .Y(n_543) );
INVx1_ASAP7_75t_L g544 ( .A(n_79), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g545 ( .A(n_256), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_315), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_242), .Y(n_547) );
BUFx2_ASAP7_75t_L g548 ( .A(n_138), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_126), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g550 ( .A(n_280), .Y(n_550) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_309), .Y(n_551) );
NOR2xp67_ASAP7_75t_L g552 ( .A(n_121), .B(n_301), .Y(n_552) );
INVxp67_ASAP7_75t_L g553 ( .A(n_54), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_203), .Y(n_554) );
CKINVDCx5p33_ASAP7_75t_R g555 ( .A(n_350), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_420), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_503), .Y(n_557) );
NOR2x1_ASAP7_75t_L g558 ( .A(n_374), .B(n_0), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_503), .Y(n_559) );
NOR2xp33_ASAP7_75t_SL g560 ( .A(n_360), .B(n_355), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_419), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_394), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_503), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_433), .B(n_0), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_481), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_548), .B(n_534), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_419), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_514), .B(n_1), .Y(n_568) );
OA21x2_ASAP7_75t_L g569 ( .A1(n_364), .A2(n_159), .B(n_157), .Y(n_569) );
OAI22xp5_ASAP7_75t_SL g570 ( .A1(n_372), .A2(n_6), .B1(n_4), .B2(n_5), .Y(n_570) );
BUFx6f_ASAP7_75t_L g571 ( .A(n_420), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_374), .B(n_4), .Y(n_572) );
INVx6_ASAP7_75t_L g573 ( .A(n_419), .Y(n_573) );
CKINVDCx11_ASAP7_75t_R g574 ( .A(n_372), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_514), .B(n_6), .Y(n_575) );
OA21x2_ASAP7_75t_L g576 ( .A1(n_364), .A2(n_161), .B(n_160), .Y(n_576) );
INVx2_ASAP7_75t_L g577 ( .A(n_419), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_419), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_419), .Y(n_579) );
OAI22xp5_ASAP7_75t_L g580 ( .A1(n_407), .A2(n_9), .B1(n_7), .B2(n_8), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_503), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_420), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_406), .B(n_10), .Y(n_583) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_420), .Y(n_584) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_426), .B(n_10), .Y(n_585) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_552), .B(n_11), .Y(n_586) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_428), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_449), .B(n_11), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_428), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_503), .Y(n_590) );
INVx3_ASAP7_75t_L g591 ( .A(n_503), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_399), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_399), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_428), .Y(n_594) );
OAI22xp5_ASAP7_75t_SL g595 ( .A1(n_413), .A2(n_15), .B1(n_12), .B2(n_13), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_524), .B(n_12), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_591), .B(n_425), .Y(n_597) );
BUFx3_ASAP7_75t_L g598 ( .A(n_591), .Y(n_598) );
BUFx10_ASAP7_75t_L g599 ( .A(n_573), .Y(n_599) );
INVx3_ASAP7_75t_L g600 ( .A(n_591), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_560), .B(n_421), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_591), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_561), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_556), .Y(n_604) );
BUFx3_ASAP7_75t_L g605 ( .A(n_573), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_566), .B(n_368), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_556), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_575), .B(n_446), .Y(n_608) );
OR2x6_ASAP7_75t_L g609 ( .A(n_570), .B(n_522), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_575), .B(n_482), .Y(n_610) );
BUFx10_ASAP7_75t_L g611 ( .A(n_573), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_583), .B(n_500), .Y(n_612) );
INVx2_ASAP7_75t_SL g613 ( .A(n_573), .Y(n_613) );
INVxp67_ASAP7_75t_SL g614 ( .A(n_568), .Y(n_614) );
AND2x6_ASAP7_75t_L g615 ( .A(n_572), .B(n_475), .Y(n_615) );
INVx2_ASAP7_75t_L g616 ( .A(n_556), .Y(n_616) );
NAND2xp5_ASAP7_75t_SL g617 ( .A(n_560), .B(n_523), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_557), .B(n_369), .Y(n_618) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_557), .B(n_378), .C(n_356), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_561), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_561), .Y(n_621) );
BUFx10_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
INVx4_ASAP7_75t_L g623 ( .A(n_572), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_559), .B(n_369), .Y(n_624) );
INVx5_ASAP7_75t_L g625 ( .A(n_556), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_567), .Y(n_626) );
NAND2xp33_ASAP7_75t_L g627 ( .A(n_588), .B(n_357), .Y(n_627) );
HB1xp67_ASAP7_75t_L g628 ( .A(n_583), .Y(n_628) );
INVxp67_ASAP7_75t_L g629 ( .A(n_562), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_592), .B(n_593), .Y(n_630) );
INVx5_ASAP7_75t_L g631 ( .A(n_556), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_559), .B(n_385), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_556), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_572), .A2(n_361), .B1(n_373), .B2(n_366), .Y(n_634) );
CKINVDCx5p33_ASAP7_75t_R g635 ( .A(n_574), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_571), .Y(n_636) );
INVx2_ASAP7_75t_SL g637 ( .A(n_623), .Y(n_637) );
OAI221xp5_ASAP7_75t_L g638 ( .A1(n_634), .A2(n_564), .B1(n_588), .B2(n_596), .C(n_565), .Y(n_638) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_614), .A2(n_580), .B1(n_585), .B2(n_410), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_606), .B(n_546), .Y(n_640) );
NAND2xp5_ASAP7_75t_SL g641 ( .A(n_623), .B(n_567), .Y(n_641) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_623), .B(n_567), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_597), .B(n_596), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_630), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_608), .B(n_558), .Y(n_645) );
BUFx6f_ASAP7_75t_L g646 ( .A(n_599), .Y(n_646) );
BUFx2_ASAP7_75t_L g647 ( .A(n_628), .Y(n_647) );
BUFx4f_ASAP7_75t_L g648 ( .A(n_615), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_610), .B(n_563), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_618), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_623), .B(n_563), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_618), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_615), .Y(n_653) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_615), .A2(n_581), .B1(n_590), .B2(n_532), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_606), .B(n_581), .Y(n_655) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_612), .A2(n_565), .B1(n_580), .B2(n_595), .C(n_570), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_615), .A2(n_590), .B1(n_578), .B2(n_579), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_603), .Y(n_658) );
NAND2xp33_ASAP7_75t_L g659 ( .A(n_615), .B(n_577), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_615), .B(n_592), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_615), .A2(n_578), .B1(n_579), .B2(n_577), .Y(n_661) );
INVx2_ASAP7_75t_SL g662 ( .A(n_615), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_603), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_627), .B(n_593), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_600), .B(n_359), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g666 ( .A1(n_624), .A2(n_578), .B(n_579), .C(n_577), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_600), .B(n_367), .Y(n_667) );
NAND2x1_ASAP7_75t_L g668 ( .A(n_600), .B(n_362), .Y(n_668) );
NAND2xp33_ASAP7_75t_L g669 ( .A(n_602), .B(n_428), .Y(n_669) );
INVx2_ASAP7_75t_SL g670 ( .A(n_599), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_629), .B(n_370), .Y(n_671) );
INVx2_ASAP7_75t_SL g672 ( .A(n_601), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_620), .B(n_379), .Y(n_673) );
NAND2xp5_ASAP7_75t_SL g674 ( .A(n_620), .B(n_390), .Y(n_674) );
NOR3xp33_ASAP7_75t_L g675 ( .A(n_617), .B(n_595), .C(n_404), .Y(n_675) );
BUFx3_ASAP7_75t_L g676 ( .A(n_599), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g677 ( .A1(n_619), .A2(n_410), .B1(n_447), .B2(n_407), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_600), .B(n_380), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_598), .B(n_383), .Y(n_679) );
AOI22xp5_ASAP7_75t_L g680 ( .A1(n_619), .A2(n_461), .B1(n_467), .B2(n_447), .Y(n_680) );
AOI22xp5_ASAP7_75t_SL g681 ( .A1(n_635), .A2(n_438), .B1(n_496), .B2(n_413), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_621), .A2(n_381), .B1(n_382), .B2(n_376), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_626), .B(n_392), .Y(n_683) );
OR2x2_ASAP7_75t_L g684 ( .A(n_609), .B(n_358), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_624), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_626), .B(n_393), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_598), .B(n_384), .Y(n_687) );
OAI22xp33_ASAP7_75t_L g688 ( .A1(n_609), .A2(n_496), .B1(n_501), .B2(n_438), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_598), .B(n_386), .Y(n_689) );
AOI22xp33_ASAP7_75t_SL g690 ( .A1(n_609), .A2(n_530), .B1(n_501), .B2(n_512), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_602), .B(n_389), .Y(n_691) );
INVx3_ASAP7_75t_L g692 ( .A(n_599), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_632), .B(n_391), .Y(n_693) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_609), .A2(n_530), .B1(n_467), .B2(n_483), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_632), .B(n_375), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_605), .B(n_396), .Y(n_696) );
BUFx2_ASAP7_75t_L g697 ( .A(n_605), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_604), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_611), .B(n_402), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g700 ( .A(n_611), .B(n_416), .Y(n_700) );
BUFx3_ASAP7_75t_L g701 ( .A(n_611), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_604), .Y(n_702) );
NAND2xp5_ASAP7_75t_SL g703 ( .A(n_611), .B(n_397), .Y(n_703) );
AND2x6_ASAP7_75t_SL g704 ( .A(n_625), .B(n_401), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_622), .B(n_429), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_622), .B(n_395), .Y(n_706) );
NAND2xp5_ASAP7_75t_SL g707 ( .A(n_613), .B(n_398), .Y(n_707) );
BUFx6f_ASAP7_75t_SL g708 ( .A(n_625), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_625), .B(n_440), .Y(n_709) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_625), .A2(n_417), .B1(n_423), .B2(n_411), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g711 ( .A1(n_604), .A2(n_576), .B(n_569), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_625), .B(n_436), .Y(n_712) );
NAND2xp5_ASAP7_75t_SL g713 ( .A(n_625), .B(n_403), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_631), .B(n_445), .Y(n_714) );
OR2x6_ASAP7_75t_L g715 ( .A(n_647), .B(n_365), .Y(n_715) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_640), .B(n_461), .Y(n_716) );
BUFx8_ASAP7_75t_L g717 ( .A(n_708), .Y(n_717) );
A2O1A1Ixp33_ASAP7_75t_L g718 ( .A1(n_650), .A2(n_431), .B(n_442), .C(n_432), .Y(n_718) );
NAND2xp5_ASAP7_75t_SL g719 ( .A(n_646), .B(n_483), .Y(n_719) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_641), .A2(n_576), .B(n_569), .Y(n_720) );
INVx4_ASAP7_75t_L g721 ( .A(n_708), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_643), .B(n_400), .Y(n_722) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_646), .B(n_539), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_658), .Y(n_724) );
AOI21xp5_ASAP7_75t_L g725 ( .A1(n_641), .A2(n_576), .B(n_569), .Y(n_725) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_638), .B(n_539), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_652), .A2(n_550), .B1(n_509), .B2(n_424), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g728 ( .A(n_646), .B(n_550), .Y(n_728) );
BUFx6f_ASAP7_75t_L g729 ( .A(n_646), .Y(n_729) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_642), .A2(n_490), .B(n_388), .Y(n_730) );
BUFx3_ASAP7_75t_L g731 ( .A(n_658), .Y(n_731) );
NAND2xp5_ASAP7_75t_SL g732 ( .A(n_676), .B(n_454), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_685), .A2(n_448), .B1(n_451), .B2(n_443), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_663), .Y(n_734) );
AND2x2_ASAP7_75t_L g735 ( .A(n_695), .B(n_412), .Y(n_735) );
O2A1O1Ixp33_ASAP7_75t_L g736 ( .A1(n_655), .A2(n_553), .B(n_459), .C(n_463), .Y(n_736) );
NOR2xp33_ASAP7_75t_SL g737 ( .A(n_648), .B(n_455), .Y(n_737) );
NOR2xp33_ASAP7_75t_L g738 ( .A(n_671), .B(n_415), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_644), .B(n_439), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_645), .B(n_444), .Y(n_740) );
A2O1A1Ixp33_ASAP7_75t_L g741 ( .A1(n_649), .A2(n_472), .B(n_479), .C(n_456), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_672), .B(n_450), .Y(n_742) );
O2A1O1Ixp5_ASAP7_75t_L g743 ( .A1(n_703), .A2(n_437), .B(n_363), .C(n_435), .Y(n_743) );
NAND2xp5_ASAP7_75t_SL g744 ( .A(n_676), .B(n_458), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g745 ( .A(n_648), .B(n_414), .Y(n_745) );
A2O1A1Ixp33_ASAP7_75t_L g746 ( .A1(n_666), .A2(n_488), .B(n_497), .C(n_480), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g747 ( .A(n_666), .B(n_586), .C(n_387), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_681), .Y(n_748) );
O2A1O1Ixp33_ASAP7_75t_L g749 ( .A1(n_675), .A2(n_505), .B(n_513), .C(n_499), .Y(n_749) );
AOI21xp5_ASAP7_75t_L g750 ( .A1(n_651), .A2(n_408), .B(n_405), .Y(n_750) );
O2A1O1Ixp33_ASAP7_75t_SL g751 ( .A1(n_668), .A2(n_430), .B(n_434), .C(n_427), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g752 ( .A1(n_663), .A2(n_521), .B(n_533), .C(n_516), .Y(n_752) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_684), .B(n_478), .Y(n_753) );
O2A1O1Ixp33_ASAP7_75t_L g754 ( .A1(n_660), .A2(n_544), .B(n_549), .C(n_537), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_706), .B(n_484), .Y(n_755) );
OAI21x1_ASAP7_75t_L g756 ( .A1(n_711), .A2(n_616), .B(n_607), .Y(n_756) );
INVx1_ASAP7_75t_L g757 ( .A(n_664), .Y(n_757) );
BUFx3_ASAP7_75t_L g758 ( .A(n_677), .Y(n_758) );
NAND2xp5_ASAP7_75t_SL g759 ( .A(n_701), .B(n_466), .Y(n_759) );
NAND2xp5_ASAP7_75t_SL g760 ( .A(n_701), .B(n_493), .Y(n_760) );
NAND2xp5_ASAP7_75t_SL g761 ( .A(n_670), .B(n_495), .Y(n_761) );
BUFx6f_ASAP7_75t_L g762 ( .A(n_662), .Y(n_762) );
NAND2x1p5_ASAP7_75t_L g763 ( .A(n_653), .B(n_453), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_639), .A2(n_508), .B1(n_536), .B2(n_453), .Y(n_764) );
INVxp67_ASAP7_75t_L g765 ( .A(n_680), .Y(n_765) );
NOR2x1_ASAP7_75t_L g766 ( .A(n_707), .B(n_586), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_690), .B(n_486), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_659), .A2(n_465), .B(n_462), .Y(n_768) );
AND2x2_ASAP7_75t_L g769 ( .A(n_682), .B(n_487), .Y(n_769) );
AOI21xp5_ASAP7_75t_L g770 ( .A1(n_659), .A2(n_469), .B(n_468), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g771 ( .A(n_670), .B(n_504), .Y(n_771) );
AOI21xp5_ASAP7_75t_L g772 ( .A1(n_637), .A2(n_473), .B(n_470), .Y(n_772) );
NOR3xp33_ASAP7_75t_L g773 ( .A(n_694), .B(n_498), .C(n_492), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_654), .A2(n_511), .B1(n_518), .B2(n_515), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_657), .A2(n_535), .B1(n_542), .B2(n_540), .Y(n_775) );
NAND2xp5_ASAP7_75t_SL g776 ( .A(n_637), .B(n_506), .Y(n_776) );
BUFx2_ASAP7_75t_L g777 ( .A(n_704), .Y(n_777) );
OAI22xp5_ASAP7_75t_L g778 ( .A1(n_693), .A2(n_543), .B1(n_536), .B2(n_387), .Y(n_778) );
NOR2xp33_ASAP7_75t_L g779 ( .A(n_653), .B(n_371), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_689), .B(n_363), .Y(n_780) );
BUFx2_ASAP7_75t_L g781 ( .A(n_688), .Y(n_781) );
O2A1O1Ixp33_ASAP7_75t_L g782 ( .A1(n_673), .A2(n_474), .B(n_477), .C(n_476), .Y(n_782) );
NAND2xp5_ASAP7_75t_SL g783 ( .A(n_692), .B(n_517), .Y(n_783) );
INVx2_ASAP7_75t_L g784 ( .A(n_708), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_697), .Y(n_785) );
AND2x2_ASAP7_75t_L g786 ( .A(n_710), .B(n_387), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g787 ( .A(n_661), .B(n_437), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_692), .B(n_520), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_673), .Y(n_789) );
BUFx4f_ASAP7_75t_L g790 ( .A(n_692), .Y(n_790) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_674), .B(n_529), .Y(n_791) );
NOR2xp33_ASAP7_75t_L g792 ( .A(n_691), .B(n_377), .Y(n_792) );
AOI221xp5_ASAP7_75t_L g793 ( .A1(n_674), .A2(n_387), .B1(n_489), .B2(n_494), .C(n_485), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g794 ( .A(n_699), .B(n_531), .Y(n_794) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_665), .B(n_409), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_683), .B(n_545), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_686), .B(n_551), .Y(n_797) );
AOI21x1_ASAP7_75t_L g798 ( .A1(n_713), .A2(n_616), .B(n_607), .Y(n_798) );
AOI21xp33_ASAP7_75t_L g799 ( .A1(n_700), .A2(n_502), .B(n_471), .Y(n_799) );
OAI21xp33_ASAP7_75t_L g800 ( .A1(n_679), .A2(n_687), .B(n_678), .Y(n_800) );
OAI22xp5_ASAP7_75t_L g801 ( .A1(n_705), .A2(n_510), .B1(n_519), .B2(n_507), .Y(n_801) );
NOR2xp67_ASAP7_75t_SL g802 ( .A(n_703), .B(n_555), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_686), .B(n_525), .Y(n_803) );
OAI21xp33_ASAP7_75t_L g804 ( .A1(n_667), .A2(n_527), .B(n_526), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_709), .Y(n_805) );
NAND2xp5_ASAP7_75t_SL g806 ( .A(n_696), .B(n_541), .Y(n_806) );
AOI21xp5_ASAP7_75t_L g807 ( .A1(n_713), .A2(n_554), .B(n_547), .Y(n_807) );
OAI22xp5_ASAP7_75t_L g808 ( .A1(n_712), .A2(n_418), .B1(n_422), .B2(n_385), .Y(n_808) );
AOI21xp5_ASAP7_75t_L g809 ( .A1(n_698), .A2(n_422), .B(n_418), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_714), .B(n_475), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_698), .A2(n_528), .B1(n_538), .B2(n_491), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_702), .B(n_15), .Y(n_812) );
NOR2xp33_ASAP7_75t_L g813 ( .A(n_702), .B(n_16), .Y(n_813) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_669), .A2(n_528), .B1(n_538), .B2(n_491), .Y(n_814) );
BUFx6f_ASAP7_75t_L g815 ( .A(n_646), .Y(n_815) );
CKINVDCx10_ASAP7_75t_R g816 ( .A(n_681), .Y(n_816) );
INVx1_ASAP7_75t_L g817 ( .A(n_644), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_644), .Y(n_818) );
CKINVDCx10_ASAP7_75t_R g819 ( .A(n_681), .Y(n_819) );
BUFx6f_ASAP7_75t_L g820 ( .A(n_646), .Y(n_820) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_640), .A2(n_452), .B1(n_435), .B2(n_464), .Y(n_821) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_640), .A2(n_452), .B1(n_457), .B2(n_441), .Y(n_822) );
AOI21xp5_ASAP7_75t_L g823 ( .A1(n_641), .A2(n_636), .B(n_633), .Y(n_823) );
NOR3xp33_ASAP7_75t_L g824 ( .A(n_656), .B(n_589), .C(n_582), .Y(n_824) );
NAND2xp33_ASAP7_75t_L g825 ( .A(n_646), .B(n_441), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g826 ( .A1(n_641), .A2(n_636), .B(n_633), .Y(n_826) );
AOI21x1_ASAP7_75t_L g827 ( .A1(n_711), .A2(n_594), .B(n_582), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_658), .Y(n_828) );
OAI22xp5_ASAP7_75t_L g829 ( .A1(n_650), .A2(n_457), .B1(n_460), .B2(n_441), .Y(n_829) );
OR2x6_ASAP7_75t_L g830 ( .A(n_647), .B(n_441), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_650), .A2(n_460), .B1(n_457), .B2(n_571), .Y(n_831) );
OR2x6_ASAP7_75t_L g832 ( .A(n_647), .B(n_457), .Y(n_832) );
AOI22xp5_ASAP7_75t_L g833 ( .A1(n_640), .A2(n_460), .B1(n_584), .B2(n_571), .Y(n_833) );
AOI21xp5_ASAP7_75t_L g834 ( .A1(n_641), .A2(n_631), .B(n_460), .Y(n_834) );
AOI21xp5_ASAP7_75t_L g835 ( .A1(n_720), .A2(n_587), .B(n_584), .Y(n_835) );
OAI22xp33_ASAP7_75t_L g836 ( .A1(n_781), .A2(n_20), .B1(n_18), .B2(n_19), .Y(n_836) );
O2A1O1Ixp33_ASAP7_75t_L g837 ( .A1(n_764), .A2(n_20), .B(n_18), .C(n_19), .Y(n_837) );
OAI21x1_ASAP7_75t_L g838 ( .A1(n_756), .A2(n_584), .B(n_571), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_817), .B(n_21), .Y(n_839) );
OAI21x1_ASAP7_75t_L g840 ( .A1(n_827), .A2(n_584), .B(n_571), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_818), .Y(n_841) );
OA21x2_ASAP7_75t_L g842 ( .A1(n_725), .A2(n_587), .B(n_165), .Y(n_842) );
O2A1O1Ixp33_ASAP7_75t_L g843 ( .A1(n_764), .A2(n_25), .B(n_21), .C(n_23), .Y(n_843) );
BUFx6f_ASAP7_75t_L g844 ( .A(n_729), .Y(n_844) );
O2A1O1Ixp5_ASAP7_75t_SL g845 ( .A1(n_811), .A2(n_587), .B(n_166), .C(n_167), .Y(n_845) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_735), .B(n_23), .Y(n_846) );
AO32x2_ASAP7_75t_L g847 ( .A1(n_811), .A2(n_587), .A3(n_27), .B1(n_25), .B2(n_26), .Y(n_847) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_800), .A2(n_30), .B(n_28), .C(n_29), .Y(n_848) );
AOI221xp5_ASAP7_75t_SL g849 ( .A1(n_736), .A2(n_28), .B1(n_29), .B2(n_30), .C(n_32), .Y(n_849) );
INVx2_ASAP7_75t_L g850 ( .A(n_731), .Y(n_850) );
OAI21xp33_ASAP7_75t_L g851 ( .A1(n_753), .A2(n_32), .B(n_33), .Y(n_851) );
O2A1O1Ixp33_ASAP7_75t_L g852 ( .A1(n_718), .A2(n_36), .B(n_34), .C(n_35), .Y(n_852) );
AO32x2_ASAP7_75t_L g853 ( .A1(n_808), .A2(n_34), .A3(n_37), .B1(n_38), .B2(n_39), .Y(n_853) );
OAI21x1_ASAP7_75t_L g854 ( .A1(n_798), .A2(n_171), .B(n_169), .Y(n_854) );
AND2x4_ASAP7_75t_L g855 ( .A(n_721), .B(n_40), .Y(n_855) );
INVx5_ASAP7_75t_L g856 ( .A(n_830), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_716), .B(n_40), .Y(n_857) );
INVx2_ASAP7_75t_L g858 ( .A(n_724), .Y(n_858) );
A2O1A1Ixp33_ASAP7_75t_L g859 ( .A1(n_754), .A2(n_44), .B(n_41), .C(n_42), .Y(n_859) );
AO31x2_ASAP7_75t_L g860 ( .A1(n_746), .A2(n_47), .A3(n_45), .B(n_46), .Y(n_860) );
AOI221xp5_ASAP7_75t_SL g861 ( .A1(n_749), .A2(n_45), .B1(n_47), .B2(n_48), .C(n_49), .Y(n_861) );
NAND3x1_ASAP7_75t_L g862 ( .A(n_816), .B(n_49), .C(n_50), .Y(n_862) );
O2A1O1Ixp33_ASAP7_75t_L g863 ( .A1(n_741), .A2(n_52), .B(n_50), .C(n_51), .Y(n_863) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_830), .A2(n_55), .B1(n_52), .B2(n_53), .Y(n_864) );
AOI21xp5_ASAP7_75t_L g865 ( .A1(n_810), .A2(n_174), .B(n_173), .Y(n_865) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_757), .A2(n_177), .B(n_175), .Y(n_866) );
OR2x2_ASAP7_75t_L g867 ( .A(n_727), .B(n_53), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_765), .B(n_55), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_772), .A2(n_181), .B(n_180), .Y(n_869) );
CKINVDCx6p67_ASAP7_75t_R g870 ( .A(n_819), .Y(n_870) );
INVx2_ASAP7_75t_L g871 ( .A(n_734), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_717), .Y(n_872) );
CKINVDCx20_ASAP7_75t_R g873 ( .A(n_717), .Y(n_873) );
AOI21xp5_ASAP7_75t_L g874 ( .A1(n_823), .A2(n_185), .B(n_182), .Y(n_874) );
OAI21xp5_ASAP7_75t_L g875 ( .A1(n_747), .A2(n_189), .B(n_187), .Y(n_875) );
BUFx10_ASAP7_75t_L g876 ( .A(n_830), .Y(n_876) );
OAI21x1_ASAP7_75t_L g877 ( .A1(n_826), .A2(n_191), .B(n_190), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_828), .Y(n_878) );
OAI21x1_ASAP7_75t_L g879 ( .A1(n_834), .A2(n_199), .B(n_197), .Y(n_879) );
AOI31xp67_ASAP7_75t_L g880 ( .A1(n_821), .A2(n_206), .A3(n_207), .B(n_201), .Y(n_880) );
NOR2x1_ASAP7_75t_SL g881 ( .A(n_832), .B(n_56), .Y(n_881) );
AO31x2_ASAP7_75t_L g882 ( .A1(n_813), .A2(n_59), .A3(n_57), .B(n_58), .Y(n_882) );
O2A1O1Ixp33_ASAP7_75t_SL g883 ( .A1(n_805), .A2(n_211), .B(n_214), .C(n_210), .Y(n_883) );
AO31x2_ASAP7_75t_L g884 ( .A1(n_831), .A2(n_60), .A3(n_57), .B(n_58), .Y(n_884) );
AND2x2_ASAP7_75t_L g885 ( .A(n_726), .B(n_61), .Y(n_885) );
A2O1A1Ixp33_ASAP7_75t_L g886 ( .A1(n_782), .A2(n_63), .B(n_61), .C(n_62), .Y(n_886) );
O2A1O1Ixp33_ASAP7_75t_L g887 ( .A1(n_752), .A2(n_65), .B(n_62), .C(n_63), .Y(n_887) );
BUFx8_ASAP7_75t_L g888 ( .A(n_777), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_739), .Y(n_889) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_832), .Y(n_890) );
INVx3_ASAP7_75t_L g891 ( .A(n_721), .Y(n_891) );
AOI221xp5_ASAP7_75t_L g892 ( .A1(n_733), .A2(n_66), .B1(n_67), .B2(n_68), .C(n_69), .Y(n_892) );
NAND3x1_ASAP7_75t_L g893 ( .A(n_773), .B(n_66), .C(n_67), .Y(n_893) );
OAI22xp5_ASAP7_75t_L g894 ( .A1(n_832), .A2(n_69), .B1(n_71), .B2(n_72), .Y(n_894) );
INVx5_ASAP7_75t_L g895 ( .A(n_729), .Y(n_895) );
AOI21xp5_ASAP7_75t_L g896 ( .A1(n_806), .A2(n_221), .B(n_219), .Y(n_896) );
A2O1A1Ixp33_ASAP7_75t_L g897 ( .A1(n_747), .A2(n_71), .B(n_72), .C(n_73), .Y(n_897) );
OAI21xp33_ASAP7_75t_L g898 ( .A1(n_738), .A2(n_73), .B(n_74), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_824), .Y(n_899) );
A2O1A1Ixp33_ASAP7_75t_L g900 ( .A1(n_750), .A2(n_74), .B(n_75), .C(n_76), .Y(n_900) );
CKINVDCx5p33_ASAP7_75t_R g901 ( .A(n_748), .Y(n_901) );
A2O1A1Ixp33_ASAP7_75t_L g902 ( .A1(n_804), .A2(n_768), .B(n_770), .C(n_743), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_829), .A2(n_75), .A3(n_76), .B(n_77), .Y(n_903) );
INVx2_ASAP7_75t_SL g904 ( .A(n_719), .Y(n_904) );
BUFx6f_ASAP7_75t_L g905 ( .A(n_815), .Y(n_905) );
INVxp67_ASAP7_75t_SL g906 ( .A(n_815), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_722), .B(n_78), .Y(n_907) );
AND2x6_ASAP7_75t_L g908 ( .A(n_784), .B(n_78), .Y(n_908) );
O2A1O1Ixp33_ASAP7_75t_L g909 ( .A1(n_780), .A2(n_79), .B(n_81), .C(n_83), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g910 ( .A(n_758), .B(n_81), .Y(n_910) );
NAND2x1p5_ASAP7_75t_L g911 ( .A(n_815), .B(n_83), .Y(n_911) );
AO31x2_ASAP7_75t_L g912 ( .A1(n_787), .A2(n_84), .A3(n_85), .B(n_86), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_769), .B(n_84), .Y(n_913) );
OAI21xp5_ASAP7_75t_L g914 ( .A1(n_789), .A2(n_230), .B(n_229), .Y(n_914) );
AOI21xp5_ASAP7_75t_SL g915 ( .A1(n_820), .A2(n_237), .B(n_236), .Y(n_915) );
INVxp67_ASAP7_75t_SL g916 ( .A(n_820), .Y(n_916) );
AO31x2_ASAP7_75t_L g917 ( .A1(n_809), .A2(n_87), .A3(n_88), .B(n_89), .Y(n_917) );
O2A1O1Ixp33_ASAP7_75t_L g918 ( .A1(n_778), .A2(n_87), .B(n_90), .C(n_91), .Y(n_918) );
AND2x2_ASAP7_75t_L g919 ( .A(n_767), .B(n_90), .Y(n_919) );
AND2x4_ASAP7_75t_L g920 ( .A(n_785), .B(n_92), .Y(n_920) );
BUFx3_ASAP7_75t_L g921 ( .A(n_820), .Y(n_921) );
AO32x2_ASAP7_75t_L g922 ( .A1(n_801), .A2(n_814), .A3(n_775), .B1(n_774), .B2(n_751), .Y(n_922) );
BUFx3_ASAP7_75t_L g923 ( .A(n_715), .Y(n_923) );
OAI21x1_ASAP7_75t_L g924 ( .A1(n_763), .A2(n_245), .B(n_243), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_740), .B(n_92), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g926 ( .A1(n_788), .A2(n_248), .B(n_247), .Y(n_926) );
OAI21xp5_ASAP7_75t_L g927 ( .A1(n_730), .A2(n_253), .B(n_251), .Y(n_927) );
OAI21xp5_ASAP7_75t_L g928 ( .A1(n_807), .A2(n_255), .B(n_254), .Y(n_928) );
OAI21x1_ASAP7_75t_L g929 ( .A1(n_745), .A2(n_262), .B(n_257), .Y(n_929) );
A2O1A1Ixp33_ASAP7_75t_L g930 ( .A1(n_795), .A2(n_93), .B(n_94), .C(n_95), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_755), .B(n_94), .Y(n_931) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_822), .B(n_95), .C(n_96), .Y(n_932) );
AO21x2_ASAP7_75t_L g933 ( .A1(n_799), .A2(n_285), .B(n_351), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_792), .B(n_97), .Y(n_934) );
AOI22xp5_ASAP7_75t_L g935 ( .A1(n_723), .A2(n_97), .B1(n_98), .B2(n_99), .Y(n_935) );
BUFx3_ASAP7_75t_L g936 ( .A(n_715), .Y(n_936) );
AO31x2_ASAP7_75t_L g937 ( .A1(n_803), .A2(n_98), .A3(n_100), .B(n_101), .Y(n_937) );
OAI21xp5_ASAP7_75t_L g938 ( .A1(n_833), .A2(n_287), .B(n_349), .Y(n_938) );
INVx2_ASAP7_75t_L g939 ( .A(n_812), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g940 ( .A(n_790), .B(n_102), .Y(n_940) );
INVx1_ASAP7_75t_L g941 ( .A(n_786), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g942 ( .A1(n_790), .A2(n_105), .B1(n_106), .B2(n_107), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_728), .B(n_108), .Y(n_943) );
NOR2xp67_ASAP7_75t_L g944 ( .A(n_742), .B(n_109), .Y(n_944) );
AND2x2_ASAP7_75t_L g945 ( .A(n_715), .B(n_109), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_766), .B(n_110), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g947 ( .A1(n_793), .A2(n_110), .B1(n_111), .B2(n_112), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_791), .Y(n_948) );
OAI22x1_ASAP7_75t_L g949 ( .A1(n_761), .A2(n_111), .B1(n_113), .B2(n_114), .Y(n_949) );
BUFx3_ASAP7_75t_L g950 ( .A(n_762), .Y(n_950) );
AO31x2_ASAP7_75t_L g951 ( .A1(n_779), .A2(n_114), .A3(n_116), .B(n_117), .Y(n_951) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_794), .Y(n_952) );
BUFx10_ASAP7_75t_L g953 ( .A(n_762), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_796), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_797), .Y(n_955) );
AOI21xp5_ASAP7_75t_L g956 ( .A1(n_783), .A2(n_293), .B(n_348), .Y(n_956) );
A2O1A1Ixp33_ASAP7_75t_L g957 ( .A1(n_802), .A2(n_116), .B(n_117), .C(n_118), .Y(n_957) );
A2O1A1Ixp33_ASAP7_75t_L g958 ( .A1(n_771), .A2(n_119), .B(n_121), .C(n_123), .Y(n_958) );
NAND2xp5_ASAP7_75t_SL g959 ( .A(n_737), .B(n_119), .Y(n_959) );
AO31x2_ASAP7_75t_L g960 ( .A1(n_825), .A2(n_123), .A3(n_125), .B(n_126), .Y(n_960) );
AND2x4_ASAP7_75t_L g961 ( .A(n_732), .B(n_125), .Y(n_961) );
INVx2_ASAP7_75t_SL g962 ( .A(n_744), .Y(n_962) );
INVx1_ASAP7_75t_L g963 ( .A(n_776), .Y(n_963) );
OAI21xp5_ASAP7_75t_L g964 ( .A1(n_759), .A2(n_299), .B(n_347), .Y(n_964) );
AO31x2_ASAP7_75t_L g965 ( .A1(n_737), .A2(n_128), .A3(n_129), .B(n_130), .Y(n_965) );
HB1xp67_ASAP7_75t_L g966 ( .A(n_760), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_762), .Y(n_967) );
AO21x2_ASAP7_75t_L g968 ( .A1(n_827), .A2(n_300), .B(n_346), .Y(n_968) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_716), .B(n_130), .Y(n_969) );
INVx2_ASAP7_75t_L g970 ( .A(n_817), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_817), .B(n_131), .Y(n_971) );
BUFx2_ASAP7_75t_L g972 ( .A(n_717), .Y(n_972) );
OR2x6_ASAP7_75t_L g973 ( .A(n_830), .B(n_131), .Y(n_973) );
HB1xp67_ASAP7_75t_L g974 ( .A(n_830), .Y(n_974) );
AND2x2_ASAP7_75t_L g975 ( .A(n_735), .B(n_132), .Y(n_975) );
BUFx6f_ASAP7_75t_L g976 ( .A(n_729), .Y(n_976) );
OR2x2_ASAP7_75t_L g977 ( .A(n_727), .B(n_132), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g978 ( .A(n_817), .B(n_133), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_817), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_L g980 ( .A1(n_800), .A2(n_135), .B(n_136), .C(n_137), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g981 ( .A1(n_817), .A2(n_135), .B1(n_139), .B2(n_140), .Y(n_981) );
OAI21x1_ASAP7_75t_L g982 ( .A1(n_756), .A2(n_302), .B(n_338), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g983 ( .A1(n_727), .A2(n_139), .B1(n_141), .B2(n_142), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_817), .B(n_143), .Y(n_984) );
OAI22xp5_ASAP7_75t_L g985 ( .A1(n_973), .A2(n_143), .B1(n_144), .B2(n_145), .Y(n_985) );
INVx1_ASAP7_75t_L g986 ( .A(n_970), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_841), .Y(n_987) );
INVxp67_ASAP7_75t_SL g988 ( .A(n_920), .Y(n_988) );
NAND2xp5_ASAP7_75t_L g989 ( .A(n_889), .B(n_145), .Y(n_989) );
OAI21xp5_ASAP7_75t_L g990 ( .A1(n_899), .A2(n_146), .B(n_147), .Y(n_990) );
OAI21xp5_ASAP7_75t_L g991 ( .A1(n_902), .A2(n_149), .B(n_150), .Y(n_991) );
AOI21xp5_ASAP7_75t_L g992 ( .A1(n_835), .A2(n_308), .B(n_331), .Y(n_992) );
NAND2x1_ASAP7_75t_L g993 ( .A(n_973), .B(n_305), .Y(n_993) );
AND2x4_ASAP7_75t_L g994 ( .A(n_979), .B(n_150), .Y(n_994) );
OR2x2_ASAP7_75t_L g995 ( .A(n_867), .B(n_151), .Y(n_995) );
AO31x2_ASAP7_75t_L g996 ( .A1(n_848), .A2(n_151), .A3(n_153), .B(n_154), .Y(n_996) );
INVx2_ASAP7_75t_L g997 ( .A(n_858), .Y(n_997) );
INVx2_ASAP7_75t_L g998 ( .A(n_871), .Y(n_998) );
INVx2_ASAP7_75t_SL g999 ( .A(n_873), .Y(n_999) );
AND2x4_ASAP7_75t_L g1000 ( .A(n_856), .B(n_155), .Y(n_1000) );
OR2x2_ASAP7_75t_L g1001 ( .A(n_977), .B(n_271), .Y(n_1001) );
INVx1_ASAP7_75t_L g1002 ( .A(n_839), .Y(n_1002) );
NAND3xp33_ASAP7_75t_L g1003 ( .A(n_849), .B(n_272), .C(n_276), .Y(n_1003) );
BUFx12f_ASAP7_75t_L g1004 ( .A(n_888), .Y(n_1004) );
INVx2_ASAP7_75t_L g1005 ( .A(n_878), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_856), .B(n_279), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_971), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1008 ( .A1(n_885), .A2(n_282), .B1(n_283), .B2(n_286), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_948), .B(n_290), .Y(n_1009) );
INVx1_ASAP7_75t_L g1010 ( .A(n_978), .Y(n_1010) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_975), .B(n_291), .Y(n_1011) );
NAND2x1p5_ASAP7_75t_L g1012 ( .A(n_856), .B(n_292), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_984), .Y(n_1013) );
INVxp33_ASAP7_75t_L g1014 ( .A(n_919), .Y(n_1014) );
OA21x2_ASAP7_75t_L g1015 ( .A1(n_982), .A2(n_314), .B(n_316), .Y(n_1015) );
OAI21xp5_ASAP7_75t_L g1016 ( .A1(n_941), .A2(n_317), .B(n_318), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_954), .B(n_322), .Y(n_1017) );
INVx1_ASAP7_75t_L g1018 ( .A(n_908), .Y(n_1018) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_955), .B(n_323), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_939), .B(n_326), .Y(n_1020) );
INVx8_ASAP7_75t_L g1021 ( .A(n_895), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_925), .A2(n_327), .B(n_353), .Y(n_1022) );
OAI21xp5_ASAP7_75t_L g1023 ( .A1(n_845), .A2(n_932), .B(n_875), .Y(n_1023) );
AOI21xp5_ASAP7_75t_L g1024 ( .A1(n_842), .A2(n_883), .B(n_934), .Y(n_1024) );
OAI21x1_ASAP7_75t_L g1025 ( .A1(n_854), .A2(n_842), .B(n_877), .Y(n_1025) );
NAND2xp5_ASAP7_75t_L g1026 ( .A(n_913), .B(n_907), .Y(n_1026) );
AO31x2_ASAP7_75t_L g1027 ( .A1(n_980), .A2(n_897), .A3(n_859), .B(n_886), .Y(n_1027) );
CKINVDCx5p33_ASAP7_75t_R g1028 ( .A(n_888), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_908), .Y(n_1029) );
AO31x2_ASAP7_75t_L g1030 ( .A1(n_874), .A2(n_949), .A3(n_900), .B(n_881), .Y(n_1030) );
AO21x2_ASAP7_75t_L g1031 ( .A1(n_914), .A2(n_938), .B(n_968), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1032 ( .A(n_901), .B(n_846), .Y(n_1032) );
NAND2xp5_ASAP7_75t_L g1033 ( .A(n_931), .B(n_868), .Y(n_1033) );
AND2x2_ASAP7_75t_L g1034 ( .A(n_945), .B(n_904), .Y(n_1034) );
NAND2xp5_ASAP7_75t_L g1035 ( .A(n_850), .B(n_963), .Y(n_1035) );
OA21x2_ASAP7_75t_L g1036 ( .A1(n_879), .A2(n_927), .B(n_861), .Y(n_1036) );
AO31x2_ASAP7_75t_L g1037 ( .A1(n_930), .A2(n_926), .A3(n_865), .B(n_866), .Y(n_1037) );
AOI21xp33_ASAP7_75t_SL g1038 ( .A1(n_836), .A2(n_855), .B(n_969), .Y(n_1038) );
OA21x2_ASAP7_75t_L g1039 ( .A1(n_928), .A2(n_929), .B(n_924), .Y(n_1039) );
BUFx2_ASAP7_75t_L g1040 ( .A(n_872), .Y(n_1040) );
NOR2x1_ASAP7_75t_SL g1041 ( .A(n_895), .B(n_844), .Y(n_1041) );
AO21x2_ASAP7_75t_L g1042 ( .A1(n_933), .A2(n_964), .B(n_946), .Y(n_1042) );
INVx1_ASAP7_75t_L g1043 ( .A(n_908), .Y(n_1043) );
AND2x4_ASAP7_75t_L g1044 ( .A(n_891), .B(n_962), .Y(n_1044) );
CKINVDCx20_ASAP7_75t_R g1045 ( .A(n_870), .Y(n_1045) );
NAND2x1p5_ASAP7_75t_L g1046 ( .A(n_855), .B(n_921), .Y(n_1046) );
INVx3_ASAP7_75t_L g1047 ( .A(n_953), .Y(n_1047) );
AOI211xp5_ASAP7_75t_L g1048 ( .A1(n_942), .A2(n_857), .B(n_864), .C(n_894), .Y(n_1048) );
INVx2_ASAP7_75t_SL g1049 ( .A(n_876), .Y(n_1049) );
INVx2_ASAP7_75t_L g1050 ( .A(n_911), .Y(n_1050) );
OR2x2_ASAP7_75t_L g1051 ( .A(n_910), .B(n_923), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_981), .Y(n_1052) );
A2O1A1Ixp33_ASAP7_75t_L g1053 ( .A1(n_851), .A2(n_918), .B(n_898), .C(n_863), .Y(n_1053) );
CKINVDCx5p33_ASAP7_75t_R g1054 ( .A(n_936), .Y(n_1054) );
NOR2xp33_ASAP7_75t_L g1055 ( .A(n_952), .B(n_966), .Y(n_1055) );
NAND2xp5_ASAP7_75t_L g1056 ( .A(n_961), .B(n_943), .Y(n_1056) );
AOI22xp5_ASAP7_75t_L g1057 ( .A1(n_983), .A2(n_892), .B1(n_961), .B2(n_935), .Y(n_1057) );
AO21x2_ASAP7_75t_L g1058 ( .A1(n_944), .A2(n_869), .B(n_957), .Y(n_1058) );
OR2x2_ASAP7_75t_L g1059 ( .A(n_890), .B(n_974), .Y(n_1059) );
OA21x2_ASAP7_75t_L g1060 ( .A1(n_956), .A2(n_958), .B(n_896), .Y(n_1060) );
OAI21x1_ASAP7_75t_L g1061 ( .A1(n_906), .A2(n_916), .B(n_915), .Y(n_1061) );
AND2x2_ASAP7_75t_L g1062 ( .A(n_847), .B(n_853), .Y(n_1062) );
AOI222xp33_ASAP7_75t_L g1063 ( .A1(n_940), .A2(n_947), .B1(n_862), .B2(n_959), .C1(n_893), .C2(n_967), .Y(n_1063) );
A2O1A1Ixp33_ASAP7_75t_L g1064 ( .A1(n_852), .A2(n_837), .B(n_843), .C(n_887), .Y(n_1064) );
NOR2x1_ASAP7_75t_L g1065 ( .A(n_909), .B(n_950), .Y(n_1065) );
A2O1A1Ixp33_ASAP7_75t_L g1066 ( .A1(n_922), .A2(n_976), .B(n_905), .C(n_860), .Y(n_1066) );
OAI22xp5_ASAP7_75t_L g1067 ( .A1(n_905), .A2(n_976), .B1(n_922), .B2(n_847), .Y(n_1067) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_860), .B(n_905), .Y(n_1068) );
OAI21x1_ASAP7_75t_L g1069 ( .A1(n_880), .A2(n_922), .B(n_917), .Y(n_1069) );
OAI21x1_ASAP7_75t_L g1070 ( .A1(n_917), .A2(n_912), .B(n_882), .Y(n_1070) );
AND2x2_ASAP7_75t_L g1071 ( .A(n_853), .B(n_937), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1072 ( .A(n_882), .B(n_951), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_882), .A2(n_951), .B(n_917), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_937), .Y(n_1074) );
NAND2x1p5_ASAP7_75t_L g1075 ( .A(n_965), .B(n_960), .Y(n_1075) );
HB1xp67_ASAP7_75t_L g1076 ( .A(n_960), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_951), .B(n_912), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g1078 ( .A(n_912), .B(n_937), .Y(n_1078) );
NAND2xp5_ASAP7_75t_L g1079 ( .A(n_903), .B(n_884), .Y(n_1079) );
OAI21x1_ASAP7_75t_L g1080 ( .A1(n_965), .A2(n_884), .B(n_903), .Y(n_1080) );
INVx2_ASAP7_75t_L g1081 ( .A(n_884), .Y(n_1081) );
OR2x2_ASAP7_75t_L g1082 ( .A(n_903), .B(n_727), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_889), .B(n_817), .Y(n_1083) );
AND2x2_ASAP7_75t_L g1084 ( .A(n_889), .B(n_735), .Y(n_1084) );
INVx3_ASAP7_75t_L g1085 ( .A(n_953), .Y(n_1085) );
AOI21xp5_ASAP7_75t_L g1086 ( .A1(n_835), .A2(n_725), .B(n_720), .Y(n_1086) );
AOI21xp5_ASAP7_75t_L g1087 ( .A1(n_835), .A2(n_725), .B(n_720), .Y(n_1087) );
NAND2xp5_ASAP7_75t_L g1088 ( .A(n_889), .B(n_817), .Y(n_1088) );
INVx1_ASAP7_75t_L g1089 ( .A(n_970), .Y(n_1089) );
AND2x2_ASAP7_75t_L g1090 ( .A(n_889), .B(n_735), .Y(n_1090) );
INVx2_ASAP7_75t_SL g1091 ( .A(n_972), .Y(n_1091) );
AOI21xp5_ASAP7_75t_L g1092 ( .A1(n_835), .A2(n_725), .B(n_720), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1093 ( .A1(n_889), .A2(n_781), .B1(n_716), .B2(n_758), .Y(n_1093) );
NAND2xp5_ASAP7_75t_L g1094 ( .A(n_899), .B(n_817), .Y(n_1094) );
AOI22xp33_ASAP7_75t_SL g1095 ( .A1(n_881), .A2(n_681), .B1(n_781), .B2(n_748), .Y(n_1095) );
AND2x4_ASAP7_75t_L g1096 ( .A(n_889), .B(n_817), .Y(n_1096) );
NOR2xp33_ASAP7_75t_L g1097 ( .A(n_889), .B(n_716), .Y(n_1097) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_889), .A2(n_656), .B1(n_690), .B2(n_716), .C(n_639), .Y(n_1098) );
NAND2xp5_ASAP7_75t_L g1099 ( .A(n_889), .B(n_817), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1100 ( .A1(n_973), .A2(n_920), .B1(n_856), .B2(n_830), .Y(n_1100) );
OAI21xp5_ASAP7_75t_L g1101 ( .A1(n_899), .A2(n_747), .B(n_902), .Y(n_1101) );
INVx2_ASAP7_75t_L g1102 ( .A(n_970), .Y(n_1102) );
BUFx3_ASAP7_75t_L g1103 ( .A(n_873), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_899), .B(n_817), .Y(n_1104) );
INVx2_ASAP7_75t_L g1105 ( .A(n_970), .Y(n_1105) );
OA21x2_ASAP7_75t_L g1106 ( .A1(n_838), .A2(n_835), .B(n_840), .Y(n_1106) );
INVx3_ASAP7_75t_L g1107 ( .A(n_953), .Y(n_1107) );
AND2x4_ASAP7_75t_L g1108 ( .A(n_889), .B(n_817), .Y(n_1108) );
INVx1_ASAP7_75t_L g1109 ( .A(n_970), .Y(n_1109) );
AND2x4_ASAP7_75t_L g1110 ( .A(n_889), .B(n_817), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_970), .Y(n_1111) );
INVx2_ASAP7_75t_L g1112 ( .A(n_970), .Y(n_1112) );
INVx1_ASAP7_75t_L g1113 ( .A(n_970), .Y(n_1113) );
NAND2xp5_ASAP7_75t_L g1114 ( .A(n_899), .B(n_817), .Y(n_1114) );
AND2x4_ASAP7_75t_L g1115 ( .A(n_889), .B(n_817), .Y(n_1115) );
AND2x6_ASAP7_75t_L g1116 ( .A(n_855), .B(n_920), .Y(n_1116) );
INVx2_ASAP7_75t_L g1117 ( .A(n_970), .Y(n_1117) );
AND2x4_ASAP7_75t_L g1118 ( .A(n_1116), .B(n_1018), .Y(n_1118) );
BUFx12f_ASAP7_75t_L g1119 ( .A(n_1004), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1120 ( .A(n_1084), .B(n_1090), .Y(n_1120) );
OR2x2_ASAP7_75t_L g1121 ( .A(n_1082), .B(n_988), .Y(n_1121) );
AND2x2_ASAP7_75t_L g1122 ( .A(n_1102), .B(n_1105), .Y(n_1122) );
OR2x6_ASAP7_75t_L g1123 ( .A(n_1100), .B(n_1046), .Y(n_1123) );
AND2x2_ASAP7_75t_L g1124 ( .A(n_1112), .B(n_1117), .Y(n_1124) );
NOR2x1_ASAP7_75t_R g1125 ( .A(n_1028), .B(n_1103), .Y(n_1125) );
INVx1_ASAP7_75t_L g1126 ( .A(n_987), .Y(n_1126) );
BUFx6f_ASAP7_75t_L g1127 ( .A(n_1061), .Y(n_1127) );
BUFx3_ASAP7_75t_L g1128 ( .A(n_1021), .Y(n_1128) );
BUFx2_ASAP7_75t_L g1129 ( .A(n_1116), .Y(n_1129) );
INVx2_ASAP7_75t_SL g1130 ( .A(n_1021), .Y(n_1130) );
INVx1_ASAP7_75t_L g1131 ( .A(n_986), .Y(n_1131) );
BUFx2_ASAP7_75t_L g1132 ( .A(n_1116), .Y(n_1132) );
INVx4_ASAP7_75t_L g1133 ( .A(n_1021), .Y(n_1133) );
AO21x2_ASAP7_75t_L g1134 ( .A1(n_1073), .A2(n_1078), .B(n_1077), .Y(n_1134) );
AND2x2_ASAP7_75t_L g1135 ( .A(n_997), .B(n_998), .Y(n_1135) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1089), .Y(n_1136) );
NAND2xp5_ASAP7_75t_L g1137 ( .A(n_1097), .B(n_1093), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1005), .B(n_1109), .Y(n_1138) );
AO21x2_ASAP7_75t_L g1139 ( .A1(n_1078), .A2(n_1077), .B(n_1066), .Y(n_1139) );
OR2x2_ASAP7_75t_L g1140 ( .A(n_1056), .B(n_1072), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1111), .B(n_1113), .Y(n_1141) );
OAI21x1_ASAP7_75t_L g1142 ( .A1(n_1025), .A2(n_1087), .B(n_1086), .Y(n_1142) );
NAND2xp5_ASAP7_75t_L g1143 ( .A(n_1096), .B(n_1108), .Y(n_1143) );
INVx4_ASAP7_75t_L g1144 ( .A(n_1116), .Y(n_1144) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1096), .B(n_1108), .Y(n_1145) );
AO21x2_ASAP7_75t_L g1146 ( .A1(n_1079), .A2(n_1072), .B(n_1024), .Y(n_1146) );
INVx1_ASAP7_75t_L g1147 ( .A(n_1110), .Y(n_1147) );
AND2x4_ASAP7_75t_L g1148 ( .A(n_1029), .B(n_1043), .Y(n_1148) );
INVx1_ASAP7_75t_L g1149 ( .A(n_1110), .Y(n_1149) );
AO21x2_ASAP7_75t_L g1150 ( .A1(n_1079), .A2(n_1101), .B(n_1092), .Y(n_1150) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1115), .B(n_1002), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_1064), .A2(n_1053), .B(n_1057), .Y(n_1152) );
AO21x2_ASAP7_75t_L g1153 ( .A1(n_1101), .A2(n_991), .B(n_1069), .Y(n_1153) );
INVx1_ASAP7_75t_L g1154 ( .A(n_1115), .Y(n_1154) );
AND2x4_ASAP7_75t_L g1155 ( .A(n_1041), .B(n_1006), .Y(n_1155) );
OA21x2_ASAP7_75t_L g1156 ( .A1(n_1070), .A2(n_1080), .B(n_1068), .Y(n_1156) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_1095), .A2(n_1098), .B1(n_1063), .B2(n_1052), .Y(n_1157) );
NAND2xp5_ASAP7_75t_L g1158 ( .A(n_1083), .B(n_1088), .Y(n_1158) );
AND2x2_ASAP7_75t_L g1159 ( .A(n_1007), .B(n_1010), .Y(n_1159) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1013), .B(n_1094), .Y(n_1160) );
HB1xp67_ASAP7_75t_L g1161 ( .A(n_1040), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1099), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1035), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_1035), .Y(n_1164) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1106), .Y(n_1165) );
AND2x2_ASAP7_75t_L g1166 ( .A(n_1094), .B(n_1104), .Y(n_1166) );
AND2x2_ASAP7_75t_L g1167 ( .A(n_1104), .B(n_1114), .Y(n_1167) );
AOI21x1_ASAP7_75t_L g1168 ( .A1(n_1067), .A2(n_1074), .B(n_1076), .Y(n_1168) );
OAI21xp5_ASAP7_75t_L g1169 ( .A1(n_1057), .A2(n_1003), .B(n_1033), .Y(n_1169) );
AO21x2_ASAP7_75t_L g1170 ( .A1(n_1081), .A2(n_1023), .B(n_1071), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1114), .B(n_990), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1172 ( .A(n_990), .B(n_1062), .Y(n_1172) );
INVx3_ASAP7_75t_L g1173 ( .A(n_1012), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_994), .Y(n_1174) );
AO21x2_ASAP7_75t_L g1175 ( .A1(n_1031), .A2(n_1042), .B(n_1016), .Y(n_1175) );
OAI211xp5_ASAP7_75t_SL g1176 ( .A1(n_1032), .A2(n_1063), .B(n_1051), .C(n_995), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1026), .B(n_1033), .Y(n_1177) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_1100), .Y(n_1178) );
INVx2_ASAP7_75t_SL g1179 ( .A(n_1047), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_989), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1034), .B(n_1014), .Y(n_1181) );
AO21x2_ASAP7_75t_L g1182 ( .A1(n_1031), .A2(n_1042), .B(n_1058), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1000), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1026), .B(n_1011), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_985), .B(n_1001), .Y(n_1185) );
OR2x6_ASAP7_75t_L g1186 ( .A(n_993), .B(n_1012), .Y(n_1186) );
AND2x2_ASAP7_75t_L g1187 ( .A(n_985), .B(n_996), .Y(n_1187) );
INVx2_ASAP7_75t_SL g1188 ( .A(n_1085), .Y(n_1188) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_1075), .Y(n_1189) );
INVx1_ASAP7_75t_L g1190 ( .A(n_1059), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1191 ( .A(n_996), .B(n_1017), .Y(n_1191) );
HB1xp67_ASAP7_75t_L g1192 ( .A(n_1107), .Y(n_1192) );
INVxp67_ASAP7_75t_L g1193 ( .A(n_1055), .Y(n_1193) );
AND2x2_ASAP7_75t_L g1194 ( .A(n_996), .B(n_1019), .Y(n_1194) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_1048), .A2(n_1038), .B1(n_1019), .B2(n_1009), .Y(n_1195) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1009), .B(n_1017), .Y(n_1196) );
INVx1_ASAP7_75t_L g1197 ( .A(n_1044), .Y(n_1197) );
BUFx2_ASAP7_75t_L g1198 ( .A(n_1075), .Y(n_1198) );
INVx4_ASAP7_75t_L g1199 ( .A(n_1049), .Y(n_1199) );
OR2x6_ASAP7_75t_L g1200 ( .A(n_1050), .B(n_1065), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1201 ( .A(n_1048), .B(n_1030), .Y(n_1201) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_1008), .A2(n_1020), .B1(n_1091), .B2(n_1054), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_999), .A2(n_1020), .B1(n_1036), .B2(n_1060), .Y(n_1203) );
INVx1_ASAP7_75t_SL g1204 ( .A(n_1045), .Y(n_1204) );
HB1xp67_ASAP7_75t_L g1205 ( .A(n_1030), .Y(n_1205) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1027), .Y(n_1206) );
INVx1_ASAP7_75t_L g1207 ( .A(n_1027), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1037), .B(n_1015), .Y(n_1208) );
AND2x4_ASAP7_75t_L g1209 ( .A(n_1022), .B(n_992), .Y(n_1209) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1039), .Y(n_1210) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_1116), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1212 ( .A(n_1102), .B(n_1105), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1201), .B(n_1172), .Y(n_1213) );
BUFx3_ASAP7_75t_L g1214 ( .A(n_1155), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1201), .B(n_1172), .Y(n_1215) );
OR2x2_ASAP7_75t_L g1216 ( .A(n_1140), .B(n_1121), .Y(n_1216) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1140), .B(n_1121), .Y(n_1217) );
HB1xp67_ASAP7_75t_L g1218 ( .A(n_1161), .Y(n_1218) );
AND2x4_ASAP7_75t_SL g1219 ( .A(n_1144), .B(n_1155), .Y(n_1219) );
AND2x2_ASAP7_75t_L g1220 ( .A(n_1187), .B(n_1166), .Y(n_1220) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1206), .Y(n_1221) );
BUFx6f_ASAP7_75t_L g1222 ( .A(n_1127), .Y(n_1222) );
INVx2_ASAP7_75t_L g1223 ( .A(n_1165), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1207), .Y(n_1224) );
NAND2x1p5_ASAP7_75t_L g1225 ( .A(n_1144), .B(n_1173), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1167), .B(n_1177), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1167), .B(n_1177), .Y(n_1227) );
AND2x4_ASAP7_75t_SL g1228 ( .A(n_1144), .B(n_1123), .Y(n_1228) );
OR2x2_ASAP7_75t_L g1229 ( .A(n_1178), .B(n_1152), .Y(n_1229) );
INVxp67_ASAP7_75t_SL g1230 ( .A(n_1174), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1141), .B(n_1160), .Y(n_1231) );
AND2x2_ASAP7_75t_L g1232 ( .A(n_1122), .B(n_1124), .Y(n_1232) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1122), .B(n_1124), .Y(n_1233) );
OAI22xp5_ASAP7_75t_L g1234 ( .A1(n_1157), .A2(n_1185), .B1(n_1123), .B2(n_1178), .Y(n_1234) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1134), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1212), .B(n_1138), .Y(n_1236) );
HB1xp67_ASAP7_75t_L g1237 ( .A(n_1151), .Y(n_1237) );
AND2x4_ASAP7_75t_L g1238 ( .A(n_1189), .B(n_1198), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1212), .B(n_1138), .Y(n_1239) );
NAND2xp5_ASAP7_75t_L g1240 ( .A(n_1162), .B(n_1159), .Y(n_1240) );
INVx1_ASAP7_75t_L g1241 ( .A(n_1134), .Y(n_1241) );
NAND2xp5_ASAP7_75t_L g1242 ( .A(n_1159), .B(n_1163), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1135), .B(n_1184), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1190), .B(n_1120), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1135), .B(n_1184), .Y(n_1245) );
AND2x2_ASAP7_75t_L g1246 ( .A(n_1171), .B(n_1191), .Y(n_1246) );
NAND2xp5_ASAP7_75t_L g1247 ( .A(n_1164), .B(n_1137), .Y(n_1247) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_1185), .A2(n_1123), .B1(n_1132), .B2(n_1129), .Y(n_1248) );
AND2x2_ASAP7_75t_L g1249 ( .A(n_1171), .B(n_1191), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1194), .B(n_1170), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1194), .B(n_1170), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1145), .B(n_1126), .Y(n_1252) );
HB1xp67_ASAP7_75t_L g1253 ( .A(n_1192), .Y(n_1253) );
NAND2x1p5_ASAP7_75t_SL g1254 ( .A(n_1196), .B(n_1130), .Y(n_1254) );
OR2x2_ASAP7_75t_L g1255 ( .A(n_1143), .B(n_1158), .Y(n_1255) );
INVx2_ASAP7_75t_SL g1256 ( .A(n_1128), .Y(n_1256) );
AND2x4_ASAP7_75t_L g1257 ( .A(n_1123), .B(n_1118), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1150), .B(n_1131), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1150), .B(n_1136), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1260 ( .A(n_1139), .B(n_1169), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1139), .B(n_1205), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1153), .B(n_1148), .Y(n_1262) );
AND2x2_ASAP7_75t_L g1263 ( .A(n_1153), .B(n_1148), .Y(n_1263) );
NAND2xp5_ASAP7_75t_L g1264 ( .A(n_1147), .B(n_1149), .Y(n_1264) );
OR2x2_ASAP7_75t_L g1265 ( .A(n_1181), .B(n_1132), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1266 ( .A(n_1154), .B(n_1180), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1221), .Y(n_1267) );
AND2x2_ASAP7_75t_L g1268 ( .A(n_1246), .B(n_1156), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1269 ( .A(n_1249), .B(n_1208), .Y(n_1269) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1221), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1224), .Y(n_1271) );
AND2x4_ASAP7_75t_L g1272 ( .A(n_1262), .B(n_1127), .Y(n_1272) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1249), .B(n_1146), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1231), .B(n_1197), .Y(n_1274) );
BUFx2_ASAP7_75t_L g1275 ( .A(n_1254), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1220), .B(n_1153), .Y(n_1276) );
INVx2_ASAP7_75t_L g1277 ( .A(n_1223), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1258), .Y(n_1278) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1258), .Y(n_1279) );
INVx3_ASAP7_75t_L g1280 ( .A(n_1222), .Y(n_1280) );
AND2x2_ASAP7_75t_L g1281 ( .A(n_1220), .B(n_1210), .Y(n_1281) );
NAND2x1p5_ASAP7_75t_L g1282 ( .A(n_1214), .B(n_1211), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1259), .Y(n_1283) );
AND2x4_ASAP7_75t_L g1284 ( .A(n_1262), .B(n_1127), .Y(n_1284) );
HB1xp67_ASAP7_75t_L g1285 ( .A(n_1253), .Y(n_1285) );
INVxp67_ASAP7_75t_L g1286 ( .A(n_1218), .Y(n_1286) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1263), .B(n_1127), .Y(n_1287) );
OR2x2_ASAP7_75t_L g1288 ( .A(n_1216), .B(n_1203), .Y(n_1288) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1213), .B(n_1168), .Y(n_1289) );
INVx2_ASAP7_75t_SL g1290 ( .A(n_1228), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1215), .B(n_1182), .Y(n_1291) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1236), .B(n_1148), .Y(n_1292) );
NAND2xp5_ASAP7_75t_SL g1293 ( .A(n_1256), .B(n_1199), .Y(n_1293) );
NAND2x1p5_ASAP7_75t_L g1294 ( .A(n_1214), .B(n_1133), .Y(n_1294) );
NAND2xp5_ASAP7_75t_L g1295 ( .A(n_1239), .B(n_1195), .Y(n_1295) );
BUFx2_ASAP7_75t_L g1296 ( .A(n_1254), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1297 ( .A(n_1232), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1298 ( .A(n_1226), .B(n_1183), .Y(n_1298) );
INVx2_ASAP7_75t_SL g1299 ( .A(n_1228), .Y(n_1299) );
HB1xp67_ASAP7_75t_L g1300 ( .A(n_1232), .Y(n_1300) );
HB1xp67_ASAP7_75t_L g1301 ( .A(n_1233), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1250), .B(n_1175), .Y(n_1302) );
HB1xp67_ASAP7_75t_L g1303 ( .A(n_1233), .Y(n_1303) );
OR2x2_ASAP7_75t_L g1304 ( .A(n_1217), .B(n_1193), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1251), .B(n_1142), .Y(n_1305) );
NOR2x1_ASAP7_75t_L g1306 ( .A(n_1238), .B(n_1186), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1267), .Y(n_1307) );
INVx2_ASAP7_75t_L g1308 ( .A(n_1277), .Y(n_1308) );
OR2x2_ASAP7_75t_L g1309 ( .A(n_1297), .B(n_1217), .Y(n_1309) );
NAND2xp5_ASAP7_75t_L g1310 ( .A(n_1300), .B(n_1227), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1311 ( .A(n_1268), .B(n_1261), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1273), .B(n_1261), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1301), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1273), .B(n_1260), .Y(n_1314) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1303), .Y(n_1315) );
INVx2_ASAP7_75t_L g1316 ( .A(n_1277), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1270), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_1281), .B(n_1243), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1281), .B(n_1243), .Y(n_1319) );
NAND2xp5_ASAP7_75t_L g1320 ( .A(n_1295), .B(n_1245), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1285), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1291), .B(n_1235), .Y(n_1322) );
INVx1_ASAP7_75t_SL g1323 ( .A(n_1304), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g1324 ( .A(n_1286), .B(n_1237), .Y(n_1324) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1304), .B(n_1204), .Y(n_1325) );
AND2x2_ASAP7_75t_SL g1326 ( .A(n_1275), .B(n_1228), .Y(n_1326) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1278), .B(n_1229), .Y(n_1327) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1271), .Y(n_1328) );
OR2x2_ASAP7_75t_L g1329 ( .A(n_1279), .B(n_1229), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1276), .B(n_1241), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1276), .B(n_1241), .Y(n_1331) );
NAND2x1_ASAP7_75t_SL g1332 ( .A(n_1306), .B(n_1257), .Y(n_1332) );
NAND2x1p5_ASAP7_75t_L g1333 ( .A(n_1306), .B(n_1133), .Y(n_1333) );
OAI31xp33_ASAP7_75t_L g1334 ( .A1(n_1296), .A2(n_1176), .A3(n_1234), .B(n_1248), .Y(n_1334) );
NAND2xp5_ASAP7_75t_L g1335 ( .A(n_1298), .B(n_1240), .Y(n_1335) );
NAND3xp33_ASAP7_75t_L g1336 ( .A(n_1334), .B(n_1288), .C(n_1296), .Y(n_1336) );
INVx1_ASAP7_75t_L g1337 ( .A(n_1309), .Y(n_1337) );
OR2x2_ASAP7_75t_L g1338 ( .A(n_1318), .B(n_1283), .Y(n_1338) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1309), .Y(n_1339) );
INVx2_ASAP7_75t_L g1340 ( .A(n_1308), .Y(n_1340) );
AND2x2_ASAP7_75t_L g1341 ( .A(n_1311), .B(n_1289), .Y(n_1341) );
INVx1_ASAP7_75t_L g1342 ( .A(n_1307), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1343 ( .A(n_1311), .B(n_1289), .Y(n_1343) );
NAND2xp5_ASAP7_75t_L g1344 ( .A(n_1314), .B(n_1283), .Y(n_1344) );
OAI21xp5_ASAP7_75t_L g1345 ( .A1(n_1333), .A2(n_1293), .B(n_1294), .Y(n_1345) );
INVx2_ASAP7_75t_L g1346 ( .A(n_1308), .Y(n_1346) );
OAI22xp5_ASAP7_75t_L g1347 ( .A1(n_1326), .A2(n_1294), .B1(n_1290), .B2(n_1299), .Y(n_1347) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1317), .Y(n_1348) );
INVx1_ASAP7_75t_L g1349 ( .A(n_1328), .Y(n_1349) );
INVx2_ASAP7_75t_L g1350 ( .A(n_1316), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1351 ( .A1(n_1333), .A2(n_1294), .B1(n_1299), .B2(n_1282), .Y(n_1351) );
NOR4xp25_ASAP7_75t_L g1352 ( .A(n_1321), .B(n_1244), .C(n_1247), .D(n_1266), .Y(n_1352) );
OR2x2_ASAP7_75t_L g1353 ( .A(n_1319), .B(n_1288), .Y(n_1353) );
OR2x2_ASAP7_75t_L g1354 ( .A(n_1310), .B(n_1269), .Y(n_1354) );
NAND4xp25_ASAP7_75t_L g1355 ( .A(n_1325), .B(n_1265), .C(n_1255), .D(n_1242), .Y(n_1355) );
INVx1_ASAP7_75t_L g1356 ( .A(n_1342), .Y(n_1356) );
AOI222xp33_ASAP7_75t_L g1357 ( .A1(n_1336), .A2(n_1323), .B1(n_1324), .B2(n_1320), .C1(n_1315), .C2(n_1313), .Y(n_1357) );
NAND2xp5_ASAP7_75t_L g1358 ( .A(n_1352), .B(n_1312), .Y(n_1358) );
AOI22xp5_ASAP7_75t_L g1359 ( .A1(n_1355), .A2(n_1330), .B1(n_1331), .B2(n_1322), .Y(n_1359) );
CKINVDCx16_ASAP7_75t_R g1360 ( .A(n_1347), .Y(n_1360) );
OAI21xp5_ASAP7_75t_SL g1361 ( .A1(n_1345), .A2(n_1219), .B(n_1225), .Y(n_1361) );
OAI221xp5_ASAP7_75t_L g1362 ( .A1(n_1351), .A2(n_1332), .B1(n_1329), .B2(n_1327), .C(n_1335), .Y(n_1362) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_1340), .Y(n_1363) );
OAI31xp33_ASAP7_75t_L g1364 ( .A1(n_1337), .A2(n_1219), .A3(n_1202), .B(n_1327), .Y(n_1364) );
OAI221xp5_ASAP7_75t_L g1365 ( .A1(n_1339), .A2(n_1329), .B1(n_1292), .B2(n_1230), .C(n_1274), .Y(n_1365) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_1360), .A2(n_1362), .B1(n_1359), .B2(n_1361), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1367 ( .A1(n_1358), .A2(n_1341), .B1(n_1343), .B2(n_1344), .C(n_1353), .Y(n_1367) );
OAI221xp5_ASAP7_75t_L g1368 ( .A1(n_1364), .A2(n_1338), .B1(n_1354), .B2(n_1349), .C(n_1348), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1369 ( .A1(n_1357), .A2(n_1252), .B1(n_1265), .B2(n_1305), .Y(n_1369) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1356), .Y(n_1370) );
NOR3xp33_ASAP7_75t_L g1371 ( .A(n_1365), .B(n_1125), .C(n_1199), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1372 ( .A(n_1363), .B(n_1302), .Y(n_1372) );
A2O1A1Ixp33_ASAP7_75t_SL g1373 ( .A1(n_1364), .A2(n_1350), .B(n_1346), .C(n_1280), .Y(n_1373) );
NAND3xp33_ASAP7_75t_L g1374 ( .A(n_1366), .B(n_1369), .C(n_1367), .Y(n_1374) );
NOR3xp33_ASAP7_75t_L g1375 ( .A(n_1373), .B(n_1371), .C(n_1368), .Y(n_1375) );
AOI221x1_ASAP7_75t_L g1376 ( .A1(n_1375), .A2(n_1199), .B1(n_1370), .B2(n_1119), .C(n_1372), .Y(n_1376) );
AND2x4_ASAP7_75t_L g1377 ( .A(n_1376), .B(n_1374), .Y(n_1377) );
NAND2x1_ASAP7_75t_L g1378 ( .A(n_1377), .B(n_1376), .Y(n_1378) );
OAI21xp5_ASAP7_75t_L g1379 ( .A1(n_1378), .A2(n_1179), .B(n_1188), .Y(n_1379) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1379), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1380), .Y(n_1381) );
OAI21xp5_ASAP7_75t_L g1382 ( .A1(n_1381), .A2(n_1200), .B(n_1264), .Y(n_1382) );
AOI21xp5_ASAP7_75t_L g1383 ( .A1(n_1382), .A2(n_1200), .B(n_1209), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1384 ( .A1(n_1383), .A2(n_1272), .B1(n_1284), .B2(n_1287), .Y(n_1384) );
endmodule