module fake_jpeg_2098_n_163 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_163);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_163;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_1),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_56),
.Y(n_65)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

AO22x1_ASAP7_75t_L g66 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_44),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g60 ( 
.A(n_47),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

BUFx4f_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_59),
.A2(n_38),
.B1(n_49),
.B2(n_51),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_64),
.B1(n_52),
.B2(n_56),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_61),
.A2(n_49),
.B1(n_44),
.B2(n_51),
.Y(n_64)
);

INVxp67_ASAP7_75t_SL g87 ( 
.A(n_66),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_67),
.B(n_69),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_37),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_60),
.A2(n_51),
.B1(n_44),
.B2(n_53),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_72),
.A2(n_57),
.B1(n_58),
.B2(n_47),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_81),
.B1(n_86),
.B2(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_74),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_76),
.B(n_79),
.Y(n_96)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_58),
.B(n_57),
.C(n_54),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_1),
.B(n_2),
.Y(n_93)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_41),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_61),
.B1(n_56),
.B2(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_45),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_85),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_83),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_62),
.B(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_64),
.A2(n_53),
.B1(n_48),
.B2(n_58),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_83),
.B(n_53),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_91),
.C(n_23),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_65),
.C(n_70),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_70),
.B1(n_65),
.B2(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_92),
.A2(n_99),
.B1(n_5),
.B2(n_6),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_7),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_75),
.B(n_4),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_104),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_77),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_78),
.Y(n_103)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_103),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_4),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_102),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_105),
.A2(n_111),
.B1(n_13),
.B2(n_14),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_114),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_110),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_112),
.B(n_113),
.Y(n_128)
);

NAND3xp33_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_8),
.C(n_9),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_25),
.B1(n_30),
.B2(n_29),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_95),
.B1(n_88),
.B2(n_90),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_116),
.A2(n_120),
.B(n_18),
.Y(n_132)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_117),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_97),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_118),
.B(n_119),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_11),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_91),
.A2(n_24),
.B1(n_28),
.B2(n_27),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_13),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_96),
.B(n_12),
.Y(n_122)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_122),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_97),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_123),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_125),
.B(n_126),
.Y(n_143)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_109),
.Y(n_130)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_132),
.B(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_106),
.Y(n_133)
);

INVx13_ASAP7_75t_L g134 ( 
.A(n_123),
.Y(n_134)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_107),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_137),
.B(n_138),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_110),
.A2(n_14),
.B(n_32),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_127),
.A2(n_108),
.B1(n_121),
.B2(n_119),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_140),
.A2(n_144),
.B1(n_131),
.B2(n_126),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_129),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_130),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_127),
.A2(n_108),
.B1(n_120),
.B2(n_115),
.Y(n_144)
);

XNOR2x1_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_152),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_142),
.A2(n_132),
.B(n_124),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_150),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_143),
.B(n_135),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_144),
.B(n_137),
.CI(n_128),
.CON(n_152),
.SN(n_152)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_156),
.B(n_154),
.Y(n_157)
);

FAx1_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_155),
.CI(n_152),
.CON(n_158),
.SN(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_147),
.B(n_141),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_159),
.A2(n_140),
.B(n_146),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_160),
.A2(n_145),
.B(n_124),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_161),
.B(n_134),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_162),
.B(n_125),
.Y(n_163)
);


endmodule