module fake_jpeg_31332_n_184 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_184);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_184;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_2),
.B(n_5),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx6_ASAP7_75t_SL g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_8),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_28),
.Y(n_41)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_8),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

BUFx8_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_44),
.A2(n_32),
.B1(n_15),
.B2(n_24),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_51),
.A2(n_46),
.B1(n_34),
.B2(n_33),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_29),
.B1(n_18),
.B2(n_15),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_52),
.A2(n_30),
.B1(n_17),
.B2(n_3),
.Y(n_92)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_37),
.B(n_22),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_59),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_25),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_60),
.B(n_61),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_25),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_71),
.Y(n_93)
);

OA22x2_ASAP7_75t_L g66 ( 
.A1(n_36),
.A2(n_30),
.B1(n_20),
.B2(n_24),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_24),
.B1(n_15),
.B2(n_23),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_22),
.Y(n_68)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_10),
.C(n_14),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_35),
.B(n_16),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_73),
.A2(n_76),
.B1(n_67),
.B2(n_56),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g75 ( 
.A(n_65),
.B(n_30),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g98 ( 
.A1(n_75),
.A2(n_63),
.B(n_48),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_79),
.Y(n_100)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_66),
.B(n_21),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_80),
.B(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_81),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_52),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_95),
.Y(n_101)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_89),
.Y(n_104)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_69),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_88),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_16),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_53),
.B(n_30),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_94),
.Y(n_112)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_63),
.Y(n_91)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_92),
.A2(n_67),
.B1(n_50),
.B2(n_64),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_30),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_72),
.B(n_17),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_102),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_74),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_109),
.B(n_110),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_93),
.B(n_70),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_64),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_87),
.C(n_76),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g127 ( 
.A(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_86),
.B(n_11),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_89),
.B(n_11),
.Y(n_117)
);

NOR2x1_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_80),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_118),
.B(n_124),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_120),
.B(n_128),
.Y(n_137)
);

XOR2x2_ASAP7_75t_SL g121 ( 
.A(n_112),
.B(n_75),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_114),
.C(n_78),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_123),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_101),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_125),
.B(n_129),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_90),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_108),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_104),
.B(n_94),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_133),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_104),
.A2(n_48),
.B(n_74),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_132),
.A2(n_109),
.B(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_88),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_105),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_138),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_126),
.A2(n_111),
.B(n_114),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_121),
.A2(n_118),
.A3(n_126),
.B1(n_131),
.B2(n_130),
.C1(n_120),
.C2(n_128),
.Y(n_139)
);

OA21x2_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_141),
.B(n_127),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_122),
.B(n_100),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g153 ( 
.A1(n_140),
.A2(n_134),
.B(n_129),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_100),
.C(n_103),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_144),
.B(n_145),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_111),
.B(n_107),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_148),
.A2(n_132),
.B1(n_127),
.B2(n_133),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_145),
.B(n_138),
.Y(n_164)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_142),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_151),
.B(n_152),
.Y(n_160)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_143),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_153),
.A2(n_155),
.B1(n_157),
.B2(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AOI322xp5_ASAP7_75t_L g165 ( 
.A1(n_158),
.A2(n_91),
.A3(n_50),
.B1(n_106),
.B2(n_85),
.C1(n_54),
.C2(n_9),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_150),
.A2(n_148),
.B1(n_147),
.B2(n_136),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_161),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_150),
.A2(n_157),
.B1(n_137),
.B2(n_156),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_151),
.A2(n_137),
.B1(n_144),
.B2(n_146),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_163),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_164),
.A2(n_54),
.B(n_17),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_165),
.B(n_166),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_152),
.B2(n_73),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_164),
.A2(n_154),
.B1(n_77),
.B2(n_83),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_168),
.A2(n_170),
.B(n_172),
.Y(n_174)
);

AOI31xp67_ASAP7_75t_L g169 ( 
.A1(n_161),
.A2(n_12),
.A3(n_17),
.B(n_3),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_169),
.B(n_160),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_173),
.B(n_176),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_174),
.A2(n_175),
.B(n_168),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_167),
.A2(n_162),
.B(n_159),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_171),
.B(n_166),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_0),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_179),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_1),
.C(n_3),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_1),
.C(n_4),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_182),
.A2(n_181),
.B1(n_5),
.B2(n_48),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_183),
.Y(n_184)
);


endmodule