module fake_jpeg_28988_n_112 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_112);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_112;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_5),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_29),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_17),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_41),
.Y(n_57)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_51),
.B(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_39),
.B(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_53),
.Y(n_59)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_0),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_42),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_63),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_43),
.B1(n_41),
.B2(n_40),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_2),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_49),
.B(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_66),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_54),
.B(n_44),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_68),
.B(n_20),
.Y(n_79)
);

INVxp33_ASAP7_75t_L g69 ( 
.A(n_67),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_71),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_65),
.A2(n_48),
.B1(n_1),
.B2(n_2),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_70),
.A2(n_78),
.B(n_12),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_58),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_57),
.A2(n_35),
.B1(n_15),
.B2(n_18),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_63),
.B(n_0),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_74),
.B(n_75),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_1),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_76),
.B(n_79),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_59),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_80),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_64),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_9),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_83),
.B(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_77),
.B(n_25),
.C(n_32),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_72),
.A2(n_7),
.B(n_8),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_87),
.A2(n_92),
.B(n_93),
.Y(n_101)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_9),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_91),
.B(n_31),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_70),
.B(n_10),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_14),
.C(n_19),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_94),
.B(n_23),
.C(n_28),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_77),
.B(n_34),
.C(n_26),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_95),
.B(n_92),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_97),
.B(n_100),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_99),
.A2(n_95),
.B(n_85),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_104),
.B(n_105),
.Y(n_107)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_103),
.A2(n_82),
.B(n_98),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_101),
.Y(n_108)
);

NOR3xp33_ASAP7_75t_SL g109 ( 
.A(n_108),
.B(n_107),
.C(n_102),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_109),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_97),
.C(n_89),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_111),
.B(n_86),
.Y(n_112)
);


endmodule