module real_jpeg_16015_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_166;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_148;
wire n_373;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_0),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_1),
.A2(n_15),
.B(n_378),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_1),
.B(n_379),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g23 ( 
.A1(n_2),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_2),
.A2(n_24),
.B1(n_115),
.B2(n_118),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_2),
.A2(n_24),
.B1(n_123),
.B2(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_2),
.A2(n_24),
.B1(n_59),
.B2(n_250),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g290 ( 
.A(n_3),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_3),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_4),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_5),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_58)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_5),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_6),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_6),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_6),
.A2(n_76),
.B1(n_201),
.B2(n_204),
.Y(n_200)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_7),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_7),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_7),
.Y(n_175)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_8),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_8),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_8),
.Y(n_268)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_9),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_9),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_9),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_9),
.Y(n_235)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_10),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_10),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_10),
.A2(n_145),
.B1(n_147),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_10),
.A2(n_49),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

OAI32xp33_ASAP7_75t_L g263 ( 
.A1(n_10),
.A2(n_88),
.A3(n_264),
.B1(n_266),
.B2(n_269),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_10),
.B(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_10),
.B(n_308),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_10),
.B(n_335),
.Y(n_334)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_11),
.Y(n_379)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_13),
.Y(n_127)
);

BUFx8_ASAP7_75t_L g150 ( 
.A(n_13),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_216),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_215),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_194),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_19),
.B(n_194),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_152),
.C(n_177),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_20),
.B(n_152),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_83),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_21),
.B(n_85),
.C(n_121),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_57),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_22),
.A2(n_57),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_22),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_22),
.B(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_22),
.A2(n_229),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

AO22x1_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_42),
.B2(n_48),
.Y(n_22)
);

AO22x2_ASAP7_75t_L g188 ( 
.A1(n_23),
.A2(n_32),
.B1(n_42),
.B2(n_48),
.Y(n_188)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_31),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_32),
.Y(n_347)
);

NOR2x1p5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_42),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_36),
.Y(n_164)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_36),
.Y(n_283)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AO22x2_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_43),
.B1(n_45),
.B2(n_46),
.Y(n_42)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_42),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_42),
.A2(n_167),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_42),
.B(n_315),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_45),
.Y(n_185)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_45),
.Y(n_251)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_48),
.B(n_167),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_48),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_50),
.B(n_53),
.Y(n_48)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI32xp33_ASAP7_75t_L g279 ( 
.A1(n_53),
.A2(n_280),
.A3(n_284),
.B1(n_286),
.B2(n_291),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_54),
.B(n_159),
.Y(n_269)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_57),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_65),
.B1(n_73),
.B2(n_80),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_58),
.A2(n_180),
.B(n_183),
.Y(n_179)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_63),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_64),
.A2(n_157),
.B1(n_159),
.B2(n_162),
.Y(n_156)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_64),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_65),
.A2(n_249),
.B1(n_252),
.B2(n_254),
.Y(n_248)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_66),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_66),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_70),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_68),
.Y(n_253)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_69),
.Y(n_311)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_70),
.Y(n_285)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_72),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g296 ( 
.A(n_72),
.Y(n_296)
);

NOR2x1_ASAP7_75t_L g169 ( 
.A(n_73),
.B(n_170),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_84),
.A2(n_85),
.B1(n_121),
.B2(n_151),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_84),
.A2(n_85),
.B1(n_188),
.B2(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_84),
.B(n_188),
.C(n_262),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_84),
.A2(n_85),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_84),
.B(n_346),
.C(n_367),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_85),
.Y(n_84)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_102),
.B1(n_107),
.B2(n_114),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_86),
.A2(n_102),
.B(n_107),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_86),
.A2(n_102),
.B1(n_107),
.B2(n_114),
.Y(n_206)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_102),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_95),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_89),
.A2(n_103),
.B1(n_104),
.B2(n_105),
.Y(n_102)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_94),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_98),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_100),
.Y(n_141)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_101),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_101),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_101),
.Y(n_241)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_102),
.Y(n_275)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx2_ASAP7_75t_SL g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_120),
.Y(n_246)
);

INVx2_ASAP7_75t_SL g151 ( 
.A(n_121),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_121),
.B(n_206),
.C(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_121),
.A2(n_151),
.B1(n_206),
.B2(n_336),
.Y(n_360)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B1(n_137),
.B2(n_144),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g191 ( 
.A1(n_122),
.A2(n_128),
.B1(n_137),
.B2(n_144),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_126),
.B(n_130),
.Y(n_129)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_127),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_127),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_128),
.B(n_137),
.Y(n_213)
);

OAI21x1_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_133),
.B(n_137),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_129),
.Y(n_245)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_132),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_137),
.Y(n_335)
);

OA22x2_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_141),
.B2(n_142),
.Y(n_137)
);

INVx6_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_147),
.B(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_147),
.Y(n_315)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_168),
.B2(n_176),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_155),
.B(n_176),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_165),
.B(n_166),
.Y(n_155)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_165),
.A2(n_347),
.B(n_348),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g176 ( 
.A(n_168),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_169),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_170),
.B(n_254),
.Y(n_270)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OA21x2_ASAP7_75t_L g312 ( 
.A1(n_172),
.A2(n_183),
.B(n_249),
.Y(n_312)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_175),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_177),
.B(n_221),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.C(n_192),
.Y(n_177)
);

XNOR2x1_ASAP7_75t_L g223 ( 
.A(n_178),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_188),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_179),
.A2(n_188),
.B1(n_272),
.B2(n_364),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_179),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_184),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g272 ( 
.A(n_188),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_188),
.B(n_279),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_188),
.A2(n_272),
.B1(n_279),
.B2(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_191),
.A2(n_192),
.B1(n_193),
.B2(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_191),
.Y(n_225)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_191),
.Y(n_367)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_208),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_206),
.B(n_207),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_198),
.B(n_206),
.Y(n_207)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_206),
.A2(n_331),
.B1(n_332),
.B2(n_336),
.Y(n_330)
);

INVx1_ASAP7_75t_SL g336 ( 
.A(n_206),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_206),
.B(n_312),
.C(n_334),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_255),
.B(n_377),
.Y(n_216)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_222),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_220),
.B(n_222),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_226),
.C(n_230),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_223),
.B(n_227),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_SL g343 ( 
.A(n_225),
.B(n_344),
.Y(n_343)
);

HB1xp67_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_229),
.B(n_248),
.C(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_229),
.B(n_327),
.C(n_329),
.Y(n_341)
);

XNOR2x1_ASAP7_75t_L g369 ( 
.A(n_230),
.B(n_370),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_231),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_247),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_232),
.A2(n_247),
.B1(n_248),
.B2(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_232),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_242),
.B1(n_245),
.B2(n_246),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_247),
.A2(n_248),
.B1(n_298),
.B2(n_299),
.Y(n_297)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_248),
.B(n_314),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_248),
.B(n_314),
.Y(n_316)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_354),
.B(n_372),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_340),
.B(n_353),
.Y(n_257)
);

AOI21x1_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_324),
.B(n_339),
.Y(n_258)
);

OAI21x1_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_276),
.B(n_323),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_273),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_261),
.B(n_273),
.Y(n_323)
);

XOR2x2_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_271),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_270),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_263),
.B(n_270),
.Y(n_327)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

AOI21x1_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_300),
.B(n_322),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_297),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_SL g322 ( 
.A(n_278),
.B(n_297),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx4_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx5_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

INVx6_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_317),
.B(n_321),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_313),
.B(n_316),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_312),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_307),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_312),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_318),
.B1(n_333),
.B2(n_334),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_318),
.B(n_319),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_338),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_338),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_329),
.B1(n_330),
.B2(n_337),
.Y(n_325)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_327),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_341),
.B(n_342),
.Y(n_353)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_349),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_350),
.C(n_351),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_SL g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_368),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_357),
.B(n_358),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_359),
.B(n_363),
.C(n_365),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_365),
.B2(n_366),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

INVx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_368),
.B(n_375),
.Y(n_374)
);

NAND2x1_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g376 ( 
.A(n_369),
.B(n_371),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);


endmodule