module real_jpeg_5755_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_0),
.A2(n_68),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_0),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_0),
.A2(n_71),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_0),
.A2(n_71),
.B1(n_305),
.B2(n_306),
.Y(n_304)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_1),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_101),
.B1(n_110),
.B2(n_112),
.Y(n_109)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_2),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_2),
.A2(n_112),
.B1(n_147),
.B2(n_149),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_2),
.A2(n_112),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_2),
.A2(n_112),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_3),
.A2(n_29),
.B1(n_139),
.B2(n_140),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_3),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_3),
.A2(n_139),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_3),
.A2(n_139),
.B1(n_351),
.B2(n_352),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_L g368 ( 
.A1(n_3),
.A2(n_139),
.B1(n_363),
.B2(n_369),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_4),
.B(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_4),
.A2(n_40),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_4),
.B(n_142),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_4),
.B(n_329),
.C(n_331),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_L g333 ( 
.A1(n_4),
.A2(n_334),
.B1(n_335),
.B2(n_337),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_4),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_4),
.B(n_235),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_4),
.A2(n_44),
.B1(n_189),
.B2(n_380),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_5),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_5),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_5),
.A2(n_99),
.B1(n_118),
.B2(n_181),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g340 ( 
.A1(n_5),
.A2(n_118),
.B1(n_337),
.B2(n_341),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_5),
.A2(n_118),
.B1(n_369),
.B2(n_381),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_7),
.A2(n_54),
.B1(n_59),
.B2(n_60),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_7),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_7),
.A2(n_59),
.B1(n_153),
.B2(n_200),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_7),
.A2(n_59),
.B1(n_280),
.B2(n_282),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_SL g465 ( 
.A1(n_7),
.A2(n_59),
.B1(n_466),
.B2(n_467),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_8),
.A2(n_99),
.B1(n_103),
.B2(n_104),
.Y(n_98)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_8),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_8),
.A2(n_103),
.B1(n_121),
.B2(n_244),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_8),
.A2(n_103),
.B1(n_357),
.B2(n_360),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_8),
.A2(n_103),
.B1(n_337),
.B2(n_420),
.Y(n_419)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_9),
.Y(n_83)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_10),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_10),
.Y(n_190)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_10),
.Y(n_229)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_10),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_10),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_11),
.Y(n_131)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_11),
.Y(n_135)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_13),
.Y(n_117)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_13),
.Y(n_121)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_13),
.Y(n_125)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_13),
.Y(n_128)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_13),
.Y(n_469)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_14),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_169)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_14),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_L g192 ( 
.A1(n_14),
.A2(n_172),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_14),
.A2(n_172),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_14),
.A2(n_121),
.B1(n_172),
.B2(n_318),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g156 ( 
.A(n_15),
.Y(n_156)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_15),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_451),
.Y(n_16)
);

OA21x2_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_320),
.B(n_445),
.Y(n_17)
);

NAND3xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_262),
.C(n_297),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_247),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_20),
.A2(n_447),
.B(n_448),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_203),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_21),
.B(n_203),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_144),
.C(n_185),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_22),
.B(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_75),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_23),
.B(n_76),
.C(n_113),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_43),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_24),
.B(n_43),
.Y(n_250)
);

OAI32xp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_29),
.A3(n_31),
.B1(n_34),
.B2(n_39),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_27),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g281 ( 
.A(n_27),
.Y(n_281)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_28),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_28),
.Y(n_134)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_33),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_36),
.Y(n_89)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_36),
.Y(n_111)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_36),
.Y(n_182)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_36),
.Y(n_307)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_52),
.B1(n_63),
.B2(n_67),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_44),
.A2(n_67),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_44),
.B(n_192),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_44),
.A2(n_221),
.B(n_270),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_44),
.A2(n_219),
.B(n_356),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_44),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_44),
.A2(n_189),
.B1(n_368),
.B2(n_380),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_44),
.A2(n_187),
.B(n_221),
.Y(n_414)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_48),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_47),
.Y(n_363)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_47),
.Y(n_369)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_51),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_51),
.Y(n_389)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_53),
.A2(n_218),
.B(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_57),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_58),
.Y(n_227)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g331 ( 
.A(n_68),
.Y(n_331)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_69),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_70),
.Y(n_196)
);

INVx6_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_73),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_113),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_98),
.B(n_108),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g183 ( 
.A(n_77),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_77),
.B(n_236),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_77),
.A2(n_235),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_77),
.A2(n_235),
.B1(n_259),
.B2(n_417),
.Y(n_416)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_77),
.A2(n_304),
.B(n_461),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_78),
.B(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_78),
.A2(n_180),
.B1(n_183),
.B2(n_184),
.Y(n_179)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_78),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_78),
.A2(n_180),
.B1(n_183),
.B2(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_78),
.A2(n_279),
.B(n_285),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B1(n_84),
.B2(n_86),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_79),
.Y(n_201)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_80),
.Y(n_336)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g411 ( 
.A(n_82),
.Y(n_411)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_83),
.Y(n_92)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_84),
.Y(n_211)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_85),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_85),
.Y(n_339)
);

INVx6_ASAP7_75t_L g344 ( 
.A(n_85),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_85),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_90),
.B1(n_93),
.B2(n_96),
.Y(n_87)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_88),
.Y(n_237)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_91),
.Y(n_407)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_94),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_132)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_98),
.Y(n_184)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_102),
.Y(n_284)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_109),
.A2(n_183),
.B(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_122),
.B1(n_137),
.B2(n_142),
.Y(n_113)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_115),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_117),
.Y(n_292)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_121),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_122),
.A2(n_289),
.B(n_316),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_122),
.B(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_143),
.B1(n_176),
.B2(n_178),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_123),
.A2(n_138),
.B1(n_143),
.B2(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_123),
.A2(n_243),
.B(n_288),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_132),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_133),
.Y(n_181)
);

INVx6_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_142),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_143),
.B(n_317),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_143),
.A2(n_465),
.B(n_470),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_144),
.B(n_185),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_175),
.C(n_179),
.Y(n_144)
);

FAx1_ASAP7_75t_SL g249 ( 
.A(n_145),
.B(n_175),
.CI(n_179),
.CON(n_249),
.SN(n_249)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_150),
.B(n_167),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_146),
.B(n_202),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_146),
.A2(n_150),
.B(n_202),
.Y(n_459)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_148),
.Y(n_413)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_149),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_150),
.A2(n_198),
.B1(n_199),
.B2(n_202),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_150),
.A2(n_167),
.B(n_273),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g310 ( 
.A(n_150),
.B(n_198),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_150),
.A2(n_435),
.B(n_436),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_151),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_151),
.A2(n_168),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_151),
.A2(n_168),
.B1(n_333),
.B2(n_340),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_151),
.A2(n_168),
.B1(n_340),
.B2(n_350),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_151),
.A2(n_168),
.B1(n_350),
.B2(n_419),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_162),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_154),
.B1(n_157),
.B2(n_161),
.Y(n_152)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_153),
.Y(n_327)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_156),
.Y(n_163)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_160),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_161),
.Y(n_351)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_162),
.Y(n_168)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_168),
.Y(n_202)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_169),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_197),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_186),
.B(n_197),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

INVx3_ASAP7_75t_SL g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_202),
.B(n_334),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_204),
.B(n_206),
.C(n_230),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_230),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_215),
.B2(n_216),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_207),
.B(n_216),
.Y(n_276)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_219),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_220),
.B(n_228),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_226),
.Y(n_382)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_227),
.Y(n_359)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_227),
.Y(n_393)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_246),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_242),
.B2(n_245),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_232),
.B(n_245),
.C(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_234),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_239),
.B(n_334),
.Y(n_408)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx5_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_241),
.Y(n_305)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_260),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_248),
.B(n_260),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_249),
.B(n_443),
.Y(n_442)
);

BUFx24_ASAP7_75t_SL g476 ( 
.A(n_249),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_250),
.B(n_251),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_255),
.C(n_257),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_252),
.A2(n_253),
.B1(n_255),
.B2(n_256),
.Y(n_430)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g429 ( 
.A(n_257),
.B(n_430),
.Y(n_429)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

A2O1A1O1Ixp25_ASAP7_75t_L g445 ( 
.A1(n_262),
.A2(n_297),
.B(n_446),
.C(n_449),
.D(n_450),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_296),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_263),
.B(n_296),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_266),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_267),
.C(n_295),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_275),
.B1(n_294),
.B2(n_295),
.Y(n_266)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_269),
.B1(n_272),
.B2(n_274),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_269),
.B1(n_315),
.B2(n_319),
.Y(n_314)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_272),
.Y(n_313)
);

AOI21xp33_ASAP7_75t_L g473 ( 
.A1(n_269),
.A2(n_313),
.B(n_315),
.Y(n_473)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_275),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_277),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_286),
.C(n_293),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_286),
.B1(n_287),
.B2(n_293),
.Y(n_277)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_278),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

OAI32xp33_ASAP7_75t_L g401 ( 
.A1(n_280),
.A2(n_402),
.A3(n_405),
.B1(n_408),
.B2(n_409),
.Y(n_401)
);

INVx3_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

OAI21xp33_ASAP7_75t_SL g417 ( 
.A1(n_281),
.A2(n_334),
.B(n_408),
.Y(n_417)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_298),
.B(n_299),
.Y(n_450)
);

BUFx24_ASAP7_75t_SL g479 ( 
.A(n_299),
.Y(n_479)
);

FAx1_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.CI(n_312),
.CON(n_299),
.SN(n_299)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_300),
.B(n_301),
.C(n_312),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_308),
.B(n_311),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_302),
.B(n_308),
.Y(n_311)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_309),
.Y(n_436)
);

FAx1_ASAP7_75t_SL g455 ( 
.A(n_311),
.B(n_456),
.CI(n_473),
.CON(n_455),
.SN(n_455)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_315),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_317),
.Y(n_471)
);

INVx8_ASAP7_75t_L g466 ( 
.A(n_318),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_440),
.B(n_444),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_425),
.B(n_439),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_323),
.A2(n_397),
.B(n_424),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_324),
.A2(n_364),
.B(n_396),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_345),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_325),
.B(n_345),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_332),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_332),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_334),
.B(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx4_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_344),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_355),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_349),
.B2(n_354),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_347),
.B(n_354),
.C(n_355),
.Y(n_398)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_SL g354 ( 
.A(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_356),
.Y(n_371)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx6_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_376),
.B(n_395),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_375),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_366),
.B(n_375),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_367),
.A2(n_370),
.B1(n_371),
.B2(n_372),
.Y(n_366)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_383),
.B(n_394),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_378),
.B(n_379),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g394 ( 
.A(n_378),
.B(n_379),
.Y(n_394)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_390),
.Y(n_385)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx8_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx4_ASAP7_75t_SL g391 ( 
.A(n_392),
.Y(n_391)
);

INVx4_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_399),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_399),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_415),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_400),
.B(n_416),
.C(n_418),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g400 ( 
.A(n_401),
.B(n_414),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_401),
.B(n_414),
.Y(n_433)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx11_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g435 ( 
.A(n_419),
.Y(n_435)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_427),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_426),
.B(n_427),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g427 ( 
.A1(n_428),
.A2(n_429),
.B1(n_431),
.B2(n_432),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_428),
.B(n_434),
.C(n_437),
.Y(n_441)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_437),
.B2(n_438),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_433),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_434),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_441),
.B(n_442),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_474),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_454),
.B(n_455),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_455),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g477 ( 
.A(n_455),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_457),
.A2(n_458),
.B1(n_464),
.B2(n_472),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_459),
.A2(n_460),
.B1(n_462),
.B2(n_463),
.Y(n_458)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_459),
.Y(n_463)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_460),
.Y(n_462)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_464),
.Y(n_472)
);

INVx8_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx8_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);


endmodule