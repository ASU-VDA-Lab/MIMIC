module fake_jpeg_12184_n_79 (n_13, n_21, n_1, n_10, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_79);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_79;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_36)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_28),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_38),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_35),
.A2(n_24),
.B1(n_34),
.B2(n_26),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_35),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_39),
.B(n_41),
.Y(n_44)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_11),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_34),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_42),
.B(n_3),
.Y(n_51)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_45),
.B(n_51),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_32),
.B(n_43),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_56),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_39),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_58),
.C(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_33),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_49),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_25),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_48),
.B(n_31),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_6),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_61),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_55),
.B(n_54),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_65),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_54),
.A2(n_24),
.B1(n_23),
.B2(n_4),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_64),
.A2(n_7),
.B1(n_13),
.B2(n_17),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_52),
.C(n_8),
.Y(n_67)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_67),
.B(n_62),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_19),
.B1(n_21),
.B2(n_22),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_71),
.Y(n_73)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_70),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_66),
.C(n_69),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_73),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_77),
.B(n_78),
.Y(n_79)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);


endmodule