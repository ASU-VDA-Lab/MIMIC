module fake_jpeg_7425_n_90 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_90);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_90;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_24;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_22),
.B(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_4),
.B(n_9),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_16),
.B(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_3),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_27),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_48),
.B(n_50),
.Y(n_71)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_55),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_2),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_5),
.Y(n_51)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_14),
.B1(n_17),
.B2(n_7),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g53 ( 
.A1(n_43),
.A2(n_26),
.B(n_36),
.C(n_45),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_45),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_37),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

OA22x2_ASAP7_75t_L g57 ( 
.A1(n_24),
.A2(n_46),
.B1(n_35),
.B2(n_41),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_46),
.Y(n_58)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_59),
.C(n_62),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_34),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_28),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_25),
.B(n_31),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_69),
.A2(n_38),
.B1(n_57),
.B2(n_58),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_74),
.A2(n_69),
.B1(n_48),
.B2(n_72),
.Y(n_81)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_75),
.Y(n_79)
);

FAx1_ASAP7_75t_SL g76 ( 
.A(n_68),
.B(n_55),
.CI(n_59),
.CON(n_76),
.SN(n_76)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_76),
.A2(n_77),
.B1(n_78),
.B2(n_73),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_67),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_77),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_81),
.B(n_74),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_76),
.C(n_79),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_83),
.B(n_81),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_84),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_85),
.B(n_76),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_87),
.A2(n_54),
.B(n_65),
.Y(n_88)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_89),
.A3(n_29),
.B1(n_39),
.B2(n_61),
.C1(n_70),
.C2(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);


endmodule