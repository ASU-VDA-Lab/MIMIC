module real_jpeg_24278_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx3_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_1),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_1),
.B(n_106),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_1),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_85),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_1),
.B(n_60),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_1),
.B(n_48),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_1),
.B(n_36),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_1),
.B(n_51),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_2),
.B(n_48),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_85),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_2),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_2),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_36),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_51),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_2),
.B(n_24),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_3),
.B(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_3),
.B(n_98),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_3),
.B(n_85),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_3),
.B(n_36),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_3),
.B(n_51),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_3),
.B(n_24),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_4),
.B(n_17),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_4),
.B(n_98),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_4),
.B(n_85),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_4),
.B(n_60),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_48),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_4),
.B(n_36),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_4),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_4),
.B(n_333),
.Y(n_332)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_6),
.Y(n_99)
);

INVx8_ASAP7_75t_SL g30 ( 
.A(n_7),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_8),
.B(n_24),
.Y(n_23)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_8),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_8),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_8),
.B(n_85),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g238 ( 
.A(n_9),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_9),
.B(n_98),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_9),
.B(n_85),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_9),
.B(n_60),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_9),
.B(n_48),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_9),
.B(n_36),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_10),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_10),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_10),
.B(n_98),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_10),
.B(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_10),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_10),
.B(n_36),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_10),
.B(n_51),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_10),
.B(n_57),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_13),
.B(n_85),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_13),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_13),
.B(n_60),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_13),
.B(n_48),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_13),
.B(n_36),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_13),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_13),
.B(n_57),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_14),
.B(n_106),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_98),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_14),
.B(n_85),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_14),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_14),
.B(n_48),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_14),
.B(n_36),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_16),
.B(n_48),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_16),
.B(n_36),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_16),
.B(n_60),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_16),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_16),
.B(n_98),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_51),
.Y(n_169)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_17),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_21),
.B1(n_40),
.B2(n_41),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_34),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_25),
.B(n_140),
.Y(n_200)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_27),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_28),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g34 ( 
.A(n_28),
.B(n_35),
.C(n_39),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_28),
.A2(n_33),
.B1(n_35),
.B2(n_49),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_29),
.B(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_29),
.B(n_287),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_29),
.B(n_251),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_31),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_31),
.B(n_120),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_31),
.B(n_236),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_35),
.A2(n_46),
.B1(n_47),
.B2(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_62),
.C(n_63),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_42),
.B(n_391),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_53),
.C(n_54),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_43),
.B(n_389),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_45),
.B1(n_50),
.B2(n_52),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_46),
.A2(n_47),
.B1(n_58),
.B2(n_347),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_55),
.C(n_58),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_47),
.B(n_49),
.C(n_52),
.Y(n_62)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_48),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_50),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_53),
.B(n_54),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_55),
.A2(n_56),
.B1(n_379),
.B2(n_380),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_58),
.A2(n_318),
.B1(n_319),
.B2(n_347),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_58),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_SL g377 ( 
.A(n_58),
.B(n_319),
.C(n_345),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_59),
.B(n_214),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_59),
.B(n_251),
.Y(n_250)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_62),
.B(n_63),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_390),
.C(n_392),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_384),
.C(n_385),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_366),
.C(n_367),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_337),
.C(n_338),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_311),
.C(n_312),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_279),
.C(n_280),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_244),
.C(n_245),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_206),
.C(n_207),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_176),
.C(n_177),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_151),
.C(n_152),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_109),
.C(n_122),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_92),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_87),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_78),
.B(n_87),
.C(n_92),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_81),
.C(n_83),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_80),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_84),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_85),
.Y(n_141)
);

BUFx24_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_88),
.B(n_90),
.C(n_91),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_100),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_93),
.B(n_101),
.C(n_102),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_102),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_104),
.B1(n_105),
.B2(n_108),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_103),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_104),
.B(n_108),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_121),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_110),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_113),
.A2(n_114),
.B1(n_121),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_121),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_147),
.C(n_148),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_131),
.C(n_137),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_129),
.C(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_132),
.B(n_135),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_132),
.A2(n_133),
.B1(n_135),
.B2(n_136),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.C(n_142),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_165),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_166),
.C(n_175),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_161),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_160),
.C(n_161),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_159),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx24_ASAP7_75t_SL g394 ( 
.A(n_161),
.Y(n_394)
);

FAx1_ASAP7_75t_SL g161 ( 
.A(n_162),
.B(n_163),
.CI(n_164),
.CON(n_161),
.SN(n_161)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.C(n_164),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_175),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_173),
.B2(n_174),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_171),
.B2(n_172),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_169),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_173),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_180),
.B1(n_181),
.B2(n_182),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_180),
.B(n_181),
.C(n_192),
.Y(n_206)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_187),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_183),
.B(n_188),
.C(n_191),
.Y(n_210)
);

BUFx24_ASAP7_75t_SL g397 ( 
.A(n_183),
.Y(n_397)
);

FAx1_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.CI(n_186),
.CON(n_183),
.SN(n_183)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_184),
.B(n_185),
.C(n_186),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_199),
.C(n_204),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_199),
.B1(n_204),
.B2(n_205),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B(n_198),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_197),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_198),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_198),
.B(n_231),
.C(n_232),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_199),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_202),
.C(n_203),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_227),
.B2(n_243),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_208),
.B(n_228),
.C(n_229),
.Y(n_244)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_210),
.B(n_212),
.C(n_220),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_220),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_213),
.B(n_216),
.C(n_219),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_254),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_218),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_226),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_225),
.C(n_226),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_224),
.Y(n_225)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g232 ( 
.A(n_233),
.B(n_242),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_234),
.B(n_237),
.C(n_242),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_277),
.B2(n_278),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_247),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_248),
.B(n_268),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_268),
.C(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_257),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_249),
.B(n_258),
.C(n_259),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_250),
.B(n_253),
.C(n_255),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_255),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_260),
.A2(n_261),
.B1(n_262),
.B2(n_267),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_260),
.Y(n_267)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_265),
.B2(n_266),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_263),
.A2(n_264),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_266),
.C(n_267),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_263),
.B(n_286),
.C(n_289),
.Y(n_335)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_271),
.C(n_272),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_276),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_274),
.B(n_275),
.C(n_276),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_281),
.B(n_283),
.C(n_310),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_297),
.B2(n_310),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_291),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_285),
.B(n_292),
.C(n_293),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g290 ( 
.A(n_289),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g317 ( 
.A1(n_289),
.A2(n_290),
.B1(n_318),
.B2(n_319),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_SL g351 ( 
.A(n_289),
.B(n_316),
.C(n_319),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

BUFx24_ASAP7_75t_SL g395 ( 
.A(n_293),
.Y(n_395)
);

FAx1_ASAP7_75t_SL g293 ( 
.A(n_294),
.B(n_295),
.CI(n_296),
.CON(n_293),
.SN(n_293)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_294),
.B(n_295),
.C(n_296),
.Y(n_321)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_297),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_299),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_298),
.B(n_300),
.C(n_301),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_302),
.A2(n_303),
.B1(n_304),
.B2(n_309),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_302),
.B(n_305),
.C(n_307),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_307),
.B2(n_308),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_305),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g331 ( 
.A1(n_306),
.A2(n_307),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_334),
.C(n_335),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_336),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_326),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_326),
.C(n_336),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_320),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_321),
.C(n_322),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g393 ( 
.A(n_322),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g322 ( 
.A(n_323),
.B(n_324),
.CI(n_325),
.CON(n_322),
.SN(n_322)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_323),
.B(n_324),
.C(n_325),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_328),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_327),
.B(n_329),
.C(n_330),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_332),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_339),
.B(n_341),
.C(n_353),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_352),
.B2(n_353),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_343),
.A2(n_344),
.B1(n_348),
.B2(n_349),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_343),
.B(n_350),
.C(n_351),
.Y(n_369)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_346),
.Y(n_344)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_354),
.B(n_355),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_354),
.B(n_356),
.C(n_359),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_359),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_359),
.Y(n_358)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_360),
.B(n_362),
.C(n_365),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_363),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_364),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_381),
.B1(n_382),
.B2(n_383),
.Y(n_367)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_368),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_369),
.B(n_370),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_369),
.B(n_370),
.C(n_383),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_371),
.B(n_377),
.C(n_378),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_372),
.B(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_386),
.C(n_388),
.Y(n_392)
);

FAx1_ASAP7_75t_SL g372 ( 
.A(n_373),
.B(n_374),
.CI(n_375),
.CON(n_372),
.SN(n_372)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_378),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_379),
.Y(n_380)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_381),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);


endmodule