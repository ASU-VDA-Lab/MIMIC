module real_jpeg_17800_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_148;
wire n_373;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_358;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

BUFx3_ASAP7_75t_L g92 ( 
.A(n_0),
.Y(n_92)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_0),
.Y(n_101)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_1),
.A2(n_120),
.B1(n_123),
.B2(n_127),
.Y(n_119)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_1),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_1),
.A2(n_58),
.B1(n_127),
.B2(n_178),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_1),
.A2(n_127),
.B1(n_242),
.B2(n_306),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_1),
.A2(n_44),
.B1(n_127),
.B2(n_358),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_2),
.Y(n_205)
);

BUFx5_ASAP7_75t_L g211 ( 
.A(n_2),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_2),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_2),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_3),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_3),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_3),
.A2(n_143),
.B1(n_223),
.B2(n_227),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_4),
.A2(n_190),
.B1(n_191),
.B2(n_198),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_4),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_4),
.A2(n_144),
.B1(n_190),
.B2(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_5),
.Y(n_152)
);

BUFx5_ASAP7_75t_L g366 ( 
.A(n_5),
.Y(n_366)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_6),
.Y(n_108)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_6),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_6),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_6),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_6),
.Y(n_226)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_6),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_6),
.Y(n_331)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_7),
.A2(n_34),
.B1(n_38),
.B2(n_39),
.Y(n_33)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_8),
.A2(n_130),
.B1(n_133),
.B2(n_134),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_8),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_8),
.A2(n_133),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g337 ( 
.A1(n_8),
.A2(n_133),
.B1(n_316),
.B2(n_338),
.Y(n_337)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_9),
.B(n_154),
.Y(n_153)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_9),
.A2(n_97),
.A3(n_247),
.B1(n_251),
.B2(n_256),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_9),
.B(n_128),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_9),
.A2(n_23),
.B1(n_268),
.B2(n_357),
.Y(n_356)
);

AOI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_9),
.A2(n_57),
.B1(n_378),
.B2(n_381),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_10),
.A2(n_44),
.B1(n_51),
.B2(n_54),
.Y(n_43)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_11),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_11),
.Y(n_158)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_11),
.Y(n_175)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_12),
.A2(n_184),
.B1(n_185),
.B2(n_186),
.Y(n_183)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_12),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_12),
.A2(n_185),
.B1(n_240),
.B2(n_241),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_12),
.A2(n_185),
.B1(n_312),
.B2(n_315),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_13),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx4f_ASAP7_75t_L g146 ( 
.A(n_14),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_15),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g180 ( 
.A(n_15),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_272),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_270),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_232),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_19),
.B(n_232),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_164),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.Y(n_20)
);

XOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_55),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_32),
.B1(n_41),
.B2(n_43),
.Y(n_22)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_23),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_23),
.A2(n_311),
.B1(n_318),
.B2(n_319),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_23),
.A2(n_337),
.B1(n_357),
.B2(n_364),
.Y(n_363)
);

OR2x2_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_24),
.Y(n_318)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g355 ( 
.A(n_26),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_30),
.Y(n_266)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_31),
.Y(n_283)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_33),
.A2(n_138),
.B1(n_147),
.B2(n_148),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_37),
.Y(n_208)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx6_ASAP7_75t_L g341 ( 
.A(n_41),
.Y(n_341)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_49),
.Y(n_142)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_50),
.Y(n_209)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_50),
.Y(n_314)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_50),
.Y(n_340)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_61),
.B1(n_72),
.B2(n_78),
.Y(n_55)
);

OAI21xp33_ASAP7_75t_SL g166 ( 
.A1(n_56),
.A2(n_57),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_57),
.B(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_57),
.B(n_290),
.Y(n_289)
);

OAI21xp33_ASAP7_75t_SL g301 ( 
.A1(n_57),
.A2(n_289),
.B(n_302),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_57),
.B(n_354),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_57),
.B(n_231),
.Y(n_367)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_67),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_66),
.Y(n_163)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_71),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_71),
.Y(n_96)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_76),
.Y(n_122)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_76),
.Y(n_132)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_77),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OA21x2_ASAP7_75t_L g171 ( 
.A1(n_79),
.A2(n_155),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_83),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_81),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_82),
.Y(n_170)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_137),
.C(n_153),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_86),
.B(n_235),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_118),
.B1(n_128),
.B2(n_129),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_87),
.A2(n_128),
.B1(n_129),
.B2(n_183),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_88),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_88),
.A2(n_119),
.B1(n_377),
.B2(n_383),
.Y(n_376)
);

AO21x2_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_97),
.B(n_106),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_104),
.Y(n_255)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_104),
.Y(n_380)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_105),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_106)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_108),
.Y(n_281)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_112),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_113),
.Y(n_291)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_115),
.Y(n_220)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_115),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_123),
.Y(n_382)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_128),
.Y(n_383)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

BUFx2_ASAP7_75t_SL g134 ( 
.A(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_137),
.B(n_153),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_138),
.A2(n_147),
.B1(n_263),
.B2(n_267),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_145),
.Y(n_317)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_146),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_147),
.A2(n_336),
.B1(n_341),
.B2(n_342),
.Y(n_335)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_151),
.Y(n_269)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_154),
.A2(n_166),
.B1(n_171),
.B2(n_177),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22x1_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_159),
.B1(n_160),
.B2(n_162),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_181),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx12f_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_188),
.Y(n_181)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_201),
.B1(n_221),
.B2(n_230),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_189),
.Y(n_243)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_197),
.Y(n_229)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_200),
.Y(n_213)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_200),
.Y(n_308)
);

BUFx12f_ASAP7_75t_L g327 ( 
.A(n_200),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_201),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_201),
.A2(n_230),
.B1(n_301),
.B2(n_305),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_201),
.A2(n_230),
.B1(n_305),
.B2(n_324),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_201),
.A2(n_230),
.B1(n_239),
.B2(n_324),
.Y(n_385)
);

AND2x2_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_212),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_206),
.B1(n_209),
.B2(n_210),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_205),
.Y(n_218)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_208),
.Y(n_352)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

OAI22xp33_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_214),
.B1(n_216),
.B2(n_219),
.Y(n_212)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_213),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_218),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_231),
.A2(n_237),
.B1(n_238),
.B2(n_243),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_244),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_233),
.A2(n_234),
.B1(n_391),
.B2(n_392),
.Y(n_390)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_236),
.A2(n_244),
.B1(n_245),
.B2(n_393),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_236),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_261),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_246),
.A2(n_261),
.B1(n_262),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_246),
.Y(n_387)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_263),
.Y(n_319)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_389),
.B(n_395),
.Y(n_272)
);

AOI21x1_ASAP7_75t_SL g273 ( 
.A1(n_274),
.A2(n_371),
.B(n_388),
.Y(n_273)
);

OAI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_333),
.B(n_370),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_276),
.B(n_309),
.Y(n_275)
);

OR2x2_ASAP7_75t_L g370 ( 
.A(n_276),
.B(n_309),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_299),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_277),
.A2(n_299),
.B1(n_300),
.B2(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_277),
.Y(n_344)
);

OAI32xp33_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_282),
.A3(n_284),
.B1(n_289),
.B2(n_292),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_310),
.B(n_320),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_310),
.B(n_322),
.C(n_332),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_311),
.Y(n_342)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_321),
.A2(n_322),
.B1(n_323),
.B2(n_332),
.Y(n_320)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx3_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_334),
.A2(n_345),
.B(n_369),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_343),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_335),
.B(n_343),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_346),
.A2(n_362),
.B(n_368),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_356),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_353),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_367),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_363),
.B(n_367),
.Y(n_368)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_372),
.B(n_373),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_386),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_375),
.A2(n_376),
.B1(n_384),
.B2(n_385),
.Y(n_374)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_375),
.B(n_385),
.C(n_386),
.Y(n_394)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_394),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_390),
.B(n_394),
.Y(n_395)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);


endmodule