module real_aes_520_n_77 (n_17, n_28, n_76, n_56, n_34, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_43, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_44, n_7, n_4, n_6, n_12, n_68, n_69, n_46, n_59, n_25, n_73, n_48, n_37, n_70, n_50, n_26, n_13, n_24, n_2, n_55, n_62, n_67, n_33, n_14, n_11, n_16, n_39, n_5, n_45, n_60, n_38, n_0, n_63, n_1, n_53, n_36, n_77);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_43;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_44;
input n_7;
input n_4;
input n_6;
input n_12;
input n_68;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_48;
input n_37;
input n_70;
input n_50;
input n_26;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_67;
input n_33;
input n_14;
input n_11;
input n_16;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_0;
input n_63;
input n_1;
input n_53;
input n_36;
output n_77;
wire n_480;
wire n_113;
wire n_476;
wire n_187;
wire n_436;
wire n_90;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_522;
wire n_485;
wire n_222;
wire n_287;
wire n_357;
wire n_503;
wire n_386;
wire n_518;
wire n_254;
wire n_207;
wire n_469;
wire n_83;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_540;
wire n_299;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_341;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_260;
wire n_97;
wire n_186;
wire n_138;
wire n_379;
wire n_374;
wire n_453;
wire n_235;
wire n_399;
wire n_378;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_145;
wire n_415;
wire n_227;
wire n_92;
wire n_519;
wire n_510;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_94;
wire n_289;
wire n_462;
wire n_280;
wire n_333;
wire n_213;
wire n_356;
wire n_478;
wire n_408;
wire n_184;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_98;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_82;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_174;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_506;
wire n_513;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_119;
wire n_455;
wire n_504;
wire n_164;
wire n_231;
wire n_102;
wire n_454;
wire n_122;
wire n_443;
wire n_534;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_80;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_367;
wire n_267;
wire n_218;
wire n_204;
wire n_339;
wire n_398;
wire n_89;
wire n_277;
wire n_425;
wire n_331;
wire n_93;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_323;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_368;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_250;
wire n_85;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_402;
wire n_171;
wire n_87;
wire n_78;
wire n_531;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_391;
wire n_360;
wire n_165;
wire n_361;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_501;
wire n_488;
wire n_251;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_115;
wire n_96;
wire n_110;
wire n_392;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_95;
wire n_188;
wire n_269;
wire n_430;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_158;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_109;
wire n_536;
wire n_203;
wire n_470;
wire n_81;
wire n_133;
wire n_494;
wire n_377;
wire n_273;
wire n_114;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_486;
wire n_411;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_88;
wire n_159;
wire n_108;
wire n_373;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_526;
wire n_155;
wire n_243;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_446;
wire n_221;
wire n_156;
wire n_359;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_180;
wire n_212;
wire n_210;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_371;
wire n_103;
wire n_166;
wire n_224;
wire n_151;
wire n_130;
wire n_253;
wire n_459;
wire n_99;
wire n_440;
wire n_525;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_79;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_305;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_473;
wire n_465;
wire n_474;
wire n_170;
wire n_86;
wire n_375;
wire n_340;
wire n_483;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_105;
wire n_84;
wire n_294;
wire n_393;
wire n_258;
wire n_206;
wire n_307;
wire n_500;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_403;
wire n_194;
wire n_137;
wire n_424;
wire n_225;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_264;
wire n_237;
wire n_91;
AO22x2_ASAP7_75t_L g91 ( .A1(n_0), .A2(n_55), .B1(n_92), .B2(n_93), .Y(n_91) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_1), .B(n_197), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_2), .B(n_212), .Y(n_230) );
INVx1_ASAP7_75t_L g184 ( .A(n_3), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g169 ( .A1(n_4), .A2(n_49), .B1(n_170), .B2(n_171), .Y(n_169) );
INVx1_ASAP7_75t_L g171 ( .A(n_4), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g150 ( .A1(n_5), .A2(n_21), .B1(n_151), .B2(n_154), .Y(n_150) );
AO22x2_ASAP7_75t_L g95 ( .A1(n_6), .A2(n_16), .B1(n_92), .B2(n_96), .Y(n_95) );
AND2x2_ASAP7_75t_L g232 ( .A(n_7), .B(n_221), .Y(n_232) );
AND2x2_ASAP7_75t_L g241 ( .A(n_8), .B(n_242), .Y(n_241) );
INVx2_ASAP7_75t_L g218 ( .A(n_9), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g143 ( .A1(n_10), .A2(n_15), .B1(n_144), .B2(n_147), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_11), .B(n_212), .Y(n_251) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_12), .B(n_197), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_13), .A2(n_70), .B1(n_197), .B2(n_305), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g110 ( .A1(n_14), .A2(n_31), .B1(n_111), .B2(n_117), .Y(n_110) );
OAI221xp5_ASAP7_75t_L g176 ( .A1(n_16), .A2(n_55), .B1(n_59), .B2(n_177), .C(n_179), .Y(n_176) );
OR2x2_ASAP7_75t_L g219 ( .A(n_17), .B(n_69), .Y(n_219) );
OA21x2_ASAP7_75t_L g222 ( .A1(n_17), .A2(n_69), .B(n_218), .Y(n_222) );
INVx3_ASAP7_75t_L g92 ( .A(n_18), .Y(n_92) );
AOI22xp33_ASAP7_75t_L g135 ( .A1(n_19), .A2(n_27), .B1(n_136), .B2(n_140), .Y(n_135) );
AO21x2_ASAP7_75t_L g246 ( .A1(n_20), .A2(n_242), .B(n_247), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_22), .A2(n_205), .B(n_228), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_23), .B(n_212), .Y(n_261) );
OAI22xp5_ASAP7_75t_SL g166 ( .A1(n_24), .A2(n_64), .B1(n_167), .B2(n_168), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_24), .Y(n_167) );
INVx1_ASAP7_75t_SL g100 ( .A(n_25), .Y(n_100) );
INVx1_ASAP7_75t_L g186 ( .A(n_26), .Y(n_186) );
AND2x2_ASAP7_75t_L g203 ( .A(n_26), .B(n_184), .Y(n_203) );
AND2x2_ASAP7_75t_L g206 ( .A(n_26), .B(n_207), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_28), .B(n_197), .Y(n_231) );
AOI22xp33_ASAP7_75t_L g87 ( .A1(n_29), .A2(n_37), .B1(n_88), .B2(n_105), .Y(n_87) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_30), .B(n_212), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_32), .B(n_197), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_33), .A2(n_205), .B(n_237), .Y(n_236) );
AOI22xp5_ASAP7_75t_L g532 ( .A1(n_34), .A2(n_82), .B1(n_83), .B2(n_533), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_34), .Y(n_533) );
AO22x2_ASAP7_75t_L g103 ( .A1(n_35), .A2(n_59), .B1(n_92), .B2(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_36), .B(n_214), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_38), .B(n_197), .Y(n_248) );
AOI22xp33_ASAP7_75t_L g121 ( .A1(n_39), .A2(n_52), .B1(n_122), .B2(n_124), .Y(n_121) );
INVx1_ASAP7_75t_L g200 ( .A(n_40), .Y(n_200) );
INVx1_ASAP7_75t_L g209 ( .A(n_40), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_41), .B(n_212), .Y(n_239) );
AOI22xp5_ASAP7_75t_L g524 ( .A1(n_41), .A2(n_82), .B1(n_83), .B2(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_41), .Y(n_525) );
AND2x2_ASAP7_75t_L g277 ( .A(n_42), .B(n_216), .Y(n_277) );
INVx1_ASAP7_75t_L g101 ( .A(n_43), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_44), .B(n_214), .Y(n_238) );
INVx1_ASAP7_75t_L g540 ( .A(n_44), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_45), .B(n_214), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_46), .B(n_197), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g279 ( .A(n_47), .B(n_197), .Y(n_279) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_48), .A2(n_205), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g170 ( .A(n_49), .Y(n_170) );
AND2x2_ASAP7_75t_L g272 ( .A(n_50), .B(n_217), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_51), .B(n_214), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_53), .B(n_214), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g309 ( .A1(n_54), .A2(n_72), .B1(n_205), .B2(n_310), .Y(n_309) );
INVxp33_ASAP7_75t_L g181 ( .A(n_55), .Y(n_181) );
INVx1_ASAP7_75t_L g81 ( .A(n_56), .Y(n_81) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_56), .B(n_212), .Y(n_269) );
INVx1_ASAP7_75t_L g202 ( .A(n_57), .Y(n_202) );
INVx1_ASAP7_75t_L g207 ( .A(n_57), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_58), .B(n_214), .Y(n_229) );
INVxp67_ASAP7_75t_L g180 ( .A(n_59), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_60), .A2(n_76), .B1(n_158), .B2(n_162), .Y(n_157) );
AOI21xp5_ASAP7_75t_L g280 ( .A1(n_61), .A2(n_205), .B(n_281), .Y(n_280) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_62), .A2(n_205), .B(n_210), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_63), .A2(n_205), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g168 ( .A(n_64), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_65), .B(n_129), .Y(n_128) );
AND2x2_ASAP7_75t_L g263 ( .A(n_66), .B(n_217), .Y(n_263) );
NAND2xp5_ASAP7_75t_SL g302 ( .A(n_67), .B(n_216), .Y(n_302) );
AND2x2_ASAP7_75t_L g220 ( .A(n_68), .B(n_221), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_71), .A2(n_205), .B(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_73), .B(n_212), .Y(n_211) );
BUFx2_ASAP7_75t_L g271 ( .A(n_74), .Y(n_271) );
BUFx2_ASAP7_75t_SL g178 ( .A(n_75), .Y(n_178) );
AOI221xp5_ASAP7_75t_L g77 ( .A1(n_78), .A2(n_173), .B1(n_187), .B2(n_520), .C(n_523), .Y(n_77) );
XOR2xp5_ASAP7_75t_L g78 ( .A(n_79), .B(n_164), .Y(n_78) );
AOI22xp5_ASAP7_75t_L g79 ( .A1(n_80), .A2(n_81), .B1(n_82), .B2(n_83), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_81), .Y(n_80) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_83), .Y(n_82) );
HB1xp67_ASAP7_75t_L g83 ( .A(n_84), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_85), .Y(n_84) );
NOR2xp67_ASAP7_75t_L g85 ( .A(n_86), .B(n_134), .Y(n_85) );
NAND4xp25_ASAP7_75t_L g86 ( .A(n_87), .B(n_110), .C(n_121), .D(n_128), .Y(n_86) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_89), .Y(n_88) );
AND2x2_ASAP7_75t_L g89 ( .A(n_90), .B(n_97), .Y(n_89) );
AND2x2_ASAP7_75t_L g139 ( .A(n_90), .B(n_115), .Y(n_139) );
AND2x4_ASAP7_75t_L g156 ( .A(n_90), .B(n_149), .Y(n_156) );
AND2x2_ASAP7_75t_L g90 ( .A(n_91), .B(n_94), .Y(n_90) );
INVx2_ASAP7_75t_L g114 ( .A(n_91), .Y(n_114) );
AND2x2_ASAP7_75t_L g126 ( .A(n_91), .B(n_95), .Y(n_126) );
INVx1_ASAP7_75t_L g93 ( .A(n_92), .Y(n_93) );
INVx2_ASAP7_75t_L g96 ( .A(n_92), .Y(n_96) );
OAI22x1_ASAP7_75t_L g98 ( .A1(n_92), .A2(n_99), .B1(n_100), .B2(n_101), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_92), .Y(n_99) );
INVx1_ASAP7_75t_L g104 ( .A(n_92), .Y(n_104) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_94), .Y(n_109) );
INVx1_ASAP7_75t_L g94 ( .A(n_95), .Y(n_94) );
AND2x4_ASAP7_75t_L g113 ( .A(n_95), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g133 ( .A(n_95), .Y(n_133) );
AND2x2_ASAP7_75t_L g123 ( .A(n_97), .B(n_113), .Y(n_123) );
AND2x4_ASAP7_75t_L g146 ( .A(n_97), .B(n_132), .Y(n_146) );
AND2x2_ASAP7_75t_L g97 ( .A(n_98), .B(n_102), .Y(n_97) );
AND2x2_ASAP7_75t_L g107 ( .A(n_98), .B(n_103), .Y(n_107) );
INVx2_ASAP7_75t_L g116 ( .A(n_98), .Y(n_116) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
AND2x4_ASAP7_75t_L g149 ( .A(n_102), .B(n_116), .Y(n_149) );
INVx2_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
AND2x2_ASAP7_75t_L g115 ( .A(n_103), .B(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g142 ( .A(n_103), .Y(n_142) );
BUFx4f_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x4_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x4_ASAP7_75t_L g119 ( .A(n_107), .B(n_120), .Y(n_119) );
AND2x2_ASAP7_75t_L g131 ( .A(n_107), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_115), .Y(n_112) );
AND2x4_ASAP7_75t_L g148 ( .A(n_113), .B(n_149), .Y(n_148) );
INVxp67_ASAP7_75t_L g120 ( .A(n_114), .Y(n_120) );
AND2x4_ASAP7_75t_L g132 ( .A(n_114), .B(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g153 ( .A(n_115), .B(n_132), .Y(n_153) );
INVx2_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
INVx6_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
BUFx5_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
BUFx12f_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x4_ASAP7_75t_L g141 ( .A(n_126), .B(n_142), .Y(n_141) );
AND2x4_ASAP7_75t_L g163 ( .A(n_126), .B(n_149), .Y(n_163) );
INVx4_ASAP7_75t_SL g129 ( .A(n_130), .Y(n_129) );
INVx6_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AND2x4_ASAP7_75t_L g161 ( .A(n_132), .B(n_149), .Y(n_161) );
NAND4xp25_ASAP7_75t_L g134 ( .A(n_135), .B(n_143), .C(n_150), .D(n_157), .Y(n_134) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
BUFx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx6_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
BUFx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_SL g151 ( .A(n_152), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_153), .Y(n_152) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx8_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx4_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx8_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
BUFx2_ASAP7_75t_SL g162 ( .A(n_163), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_166), .B1(n_169), .B2(n_172), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g165 ( .A(n_166), .Y(n_165) );
CKINVDCx20_ASAP7_75t_R g172 ( .A(n_169), .Y(n_172) );
INVx1_ASAP7_75t_SL g173 ( .A(n_174), .Y(n_173) );
CKINVDCx20_ASAP7_75t_R g174 ( .A(n_175), .Y(n_174) );
AND3x1_ASAP7_75t_SL g175 ( .A(n_176), .B(n_182), .C(n_185), .Y(n_175) );
INVxp67_ASAP7_75t_L g531 ( .A(n_176), .Y(n_531) );
CKINVDCx8_ASAP7_75t_R g177 ( .A(n_178), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_180), .B(n_181), .Y(n_179) );
CKINVDCx16_ASAP7_75t_R g529 ( .A(n_182), .Y(n_529) );
AOI21xp33_ASAP7_75t_L g536 ( .A1(n_182), .A2(n_537), .B(n_538), .Y(n_536) );
INVx1_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AND2x2_ASAP7_75t_L g306 ( .A(n_183), .B(n_307), .Y(n_306) );
OR2x2_ASAP7_75t_SL g534 ( .A(n_183), .B(n_185), .Y(n_534) );
HB1xp67_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g208 ( .A(n_184), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_185), .B(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
NOR2x1p5_ASAP7_75t_L g311 ( .A(n_186), .B(n_312), .Y(n_311) );
INVx5_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
AND2x4_ASAP7_75t_L g188 ( .A(n_189), .B(n_424), .Y(n_188) );
NOR3xp33_ASAP7_75t_L g189 ( .A(n_190), .B(n_349), .C(n_385), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_191), .B(n_323), .Y(n_190) );
AOI211xp5_ASAP7_75t_L g191 ( .A1(n_192), .A2(n_243), .B(n_273), .C(n_298), .Y(n_191) );
AND2x2_ASAP7_75t_L g414 ( .A(n_192), .B(n_275), .Y(n_414) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_223), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_193), .B(n_396), .Y(n_395) );
AND2x2_ASAP7_75t_L g447 ( .A(n_193), .B(n_329), .Y(n_447) );
AND2x2_ASAP7_75t_L g463 ( .A(n_193), .B(n_290), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_193), .B(n_473), .Y(n_472) );
NAND2x1p5_ASAP7_75t_L g496 ( .A(n_193), .B(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AND2x4_ASAP7_75t_SL g285 ( .A(n_194), .B(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g318 ( .A(n_194), .Y(n_318) );
AND2x2_ASAP7_75t_L g365 ( .A(n_194), .B(n_300), .Y(n_365) );
AND2x2_ASAP7_75t_L g384 ( .A(n_194), .B(n_223), .Y(n_384) );
BUFx2_ASAP7_75t_L g389 ( .A(n_194), .Y(n_389) );
AND2x2_ASAP7_75t_L g433 ( .A(n_194), .B(n_233), .Y(n_433) );
AND2x4_ASAP7_75t_L g505 ( .A(n_194), .B(n_506), .Y(n_505) );
NOR2x1_ASAP7_75t_L g517 ( .A(n_194), .B(n_289), .Y(n_517) );
OR2x6_ASAP7_75t_L g194 ( .A(n_195), .B(n_220), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_204), .B(n_216), .Y(n_195) );
AND2x4_ASAP7_75t_L g197 ( .A(n_198), .B(n_203), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_199), .B(n_201), .Y(n_198) );
AND2x6_ASAP7_75t_L g214 ( .A(n_199), .B(n_207), .Y(n_214) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
AND2x4_ASAP7_75t_L g212 ( .A(n_201), .B(n_209), .Y(n_212) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx5_ASAP7_75t_L g215 ( .A(n_203), .Y(n_215) );
AND2x6_ASAP7_75t_L g205 ( .A(n_206), .B(n_208), .Y(n_205) );
BUFx3_ASAP7_75t_L g308 ( .A(n_206), .Y(n_308) );
INVx2_ASAP7_75t_L g313 ( .A(n_207), .Y(n_313) );
AND2x4_ASAP7_75t_L g310 ( .A(n_208), .B(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g307 ( .A(n_209), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_215), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_214), .B(n_271), .Y(n_270) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_215), .A2(n_229), .B(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_215), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_215), .A2(n_251), .B(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_215), .A2(n_260), .B(n_261), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_215), .A2(n_269), .B(n_270), .Y(n_268) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_215), .A2(n_282), .B(n_283), .Y(n_281) );
CKINVDCx5p33_ASAP7_75t_R g225 ( .A(n_216), .Y(n_225) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_216), .A2(n_304), .B(n_309), .Y(n_303) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_SL g217 ( .A(n_218), .B(n_219), .Y(n_217) );
AND2x4_ASAP7_75t_L g253 ( .A(n_218), .B(n_219), .Y(n_253) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_221), .A2(n_266), .B(n_267), .Y(n_265) );
BUFx4f_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx3_ASAP7_75t_L g234 ( .A(n_222), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_223), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g436 ( .A(n_223), .Y(n_436) );
BUFx2_ASAP7_75t_L g485 ( .A(n_223), .Y(n_485) );
INVx1_ASAP7_75t_L g507 ( .A(n_223), .Y(n_507) );
AND2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_233), .Y(n_223) );
INVx3_ASAP7_75t_L g286 ( .A(n_224), .Y(n_286) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_224), .Y(n_473) );
AOI21x1_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_232), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_231), .Y(n_226) );
INVx2_ASAP7_75t_L g289 ( .A(n_233), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_233), .B(n_286), .Y(n_290) );
INVx2_ASAP7_75t_L g373 ( .A(n_233), .Y(n_373) );
OR2x2_ASAP7_75t_L g380 ( .A(n_233), .B(n_329), .Y(n_380) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B(n_241), .Y(n_233) );
INVx4_ASAP7_75t_L g242 ( .A(n_234), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_240), .Y(n_235) );
INVx3_ASAP7_75t_L g256 ( .A(n_242), .Y(n_256) );
AND2x2_ASAP7_75t_L g335 ( .A(n_243), .B(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g369 ( .A(n_243), .B(n_332), .Y(n_369) );
AND2x2_ASAP7_75t_L g243 ( .A(n_244), .B(n_254), .Y(n_243) );
AND2x2_ASAP7_75t_L g405 ( .A(n_244), .B(n_296), .Y(n_405) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g362 ( .A(n_245), .B(n_255), .Y(n_362) );
AND2x2_ASAP7_75t_L g481 ( .A(n_245), .B(n_264), .Y(n_481) );
INVx2_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
INVx1_ASAP7_75t_L g295 ( .A(n_246), .Y(n_295) );
INVx1_ASAP7_75t_L g321 ( .A(n_246), .Y(n_321) );
AND2x2_ASAP7_75t_L g377 ( .A(n_246), .B(n_255), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_246), .B(n_276), .Y(n_382) );
OR2x2_ASAP7_75t_L g445 ( .A(n_246), .B(n_264), .Y(n_445) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_246), .Y(n_454) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_249), .B(n_253), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_253), .A2(n_279), .B(n_280), .Y(n_278) );
AND2x2_ASAP7_75t_L g275 ( .A(n_254), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
NOR2x1_ASAP7_75t_SL g254 ( .A(n_255), .B(n_264), .Y(n_254) );
AO21x1_ASAP7_75t_SL g255 ( .A1(n_256), .A2(n_257), .B(n_263), .Y(n_255) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_256), .A2(n_257), .B(n_263), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_262), .Y(n_257) );
AND2x2_ASAP7_75t_L g292 ( .A(n_264), .B(n_293), .Y(n_292) );
INVx2_ASAP7_75t_SL g348 ( .A(n_264), .Y(n_348) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_264), .B(n_276), .Y(n_358) );
OR2x2_ASAP7_75t_L g363 ( .A(n_264), .B(n_293), .Y(n_363) );
BUFx2_ASAP7_75t_L g419 ( .A(n_264), .Y(n_419) );
AND2x2_ASAP7_75t_L g455 ( .A(n_264), .B(n_334), .Y(n_455) );
AND2x2_ASAP7_75t_L g466 ( .A(n_264), .B(n_296), .Y(n_466) );
OR2x6_ASAP7_75t_L g264 ( .A(n_265), .B(n_272), .Y(n_264) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
AOI22xp5_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_284), .B1(n_290), .B2(n_291), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_275), .A2(n_463), .B1(n_513), .B2(n_518), .Y(n_512) );
INVx4_ASAP7_75t_L g293 ( .A(n_276), .Y(n_293) );
INVx2_ASAP7_75t_L g332 ( .A(n_276), .Y(n_332) );
HB1xp67_ASAP7_75t_L g403 ( .A(n_276), .Y(n_403) );
OR2x2_ASAP7_75t_L g418 ( .A(n_276), .B(n_296), .Y(n_418) );
OR2x2_ASAP7_75t_SL g444 ( .A(n_276), .B(n_445), .Y(n_444) );
OR2x6_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
AND2x2_ASAP7_75t_SL g284 ( .A(n_285), .B(n_287), .Y(n_284) );
INVx2_ASAP7_75t_SL g325 ( .A(n_285), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_285), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g393 ( .A(n_285), .B(n_341), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_285), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g315 ( .A(n_286), .Y(n_315) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_286), .Y(n_340) );
AND2x2_ASAP7_75t_L g396 ( .A(n_286), .B(n_373), .Y(n_396) );
INVx1_ASAP7_75t_L g506 ( .A(n_286), .Y(n_506) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g317 ( .A(n_288), .B(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_288), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g314 ( .A(n_289), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_290), .B(n_447), .Y(n_446) );
AOI321xp33_ASAP7_75t_L g468 ( .A1(n_291), .A2(n_370), .A3(n_438), .B1(n_469), .B2(n_470), .C(n_474), .Y(n_468) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVxp67_ASAP7_75t_SL g367 ( .A(n_292), .Y(n_367) );
AND2x2_ASAP7_75t_L g392 ( .A(n_292), .B(n_321), .Y(n_392) );
AND2x2_ASAP7_75t_L g467 ( .A(n_292), .B(n_377), .Y(n_467) );
INVx1_ASAP7_75t_L g336 ( .A(n_293), .Y(n_336) );
BUFx2_ASAP7_75t_L g346 ( .A(n_293), .Y(n_346) );
NOR2xp67_ASAP7_75t_L g453 ( .A(n_293), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_SL g391 ( .A(n_294), .Y(n_391) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
BUFx2_ASAP7_75t_L g398 ( .A(n_295), .Y(n_398) );
INVx2_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_296), .Y(n_357) );
INVx3_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AOI21xp33_ASAP7_75t_SL g298 ( .A1(n_299), .A2(n_316), .B(n_319), .Y(n_298) );
NOR2xp67_ASAP7_75t_L g450 ( .A(n_299), .B(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_314), .Y(n_300) );
INVx3_ASAP7_75t_L g341 ( .A(n_301), .Y(n_341) );
AND2x2_ASAP7_75t_L g372 ( .A(n_301), .B(n_373), .Y(n_372) );
AND2x4_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x4_ASAP7_75t_L g329 ( .A(n_302), .B(n_303), .Y(n_329) );
INVx1_ASAP7_75t_L g522 ( .A(n_305), .Y(n_522) );
AND2x4_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
HB1xp67_ASAP7_75t_L g537 ( .A(n_307), .Y(n_537) );
INVx1_ASAP7_75t_L g539 ( .A(n_308), .Y(n_539) );
INVx3_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g412 ( .A(n_314), .Y(n_412) );
INVx1_ASAP7_75t_SL g497 ( .A(n_315), .Y(n_497) );
INVxp33_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g371 ( .A(n_318), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g423 ( .A(n_318), .B(n_380), .Y(n_423) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_L g427 ( .A(n_320), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_320), .B(n_442), .Y(n_441) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_321), .B(n_358), .Y(n_413) );
NOR4xp25_ASAP7_75t_L g508 ( .A(n_321), .B(n_352), .C(n_509), .D(n_510), .Y(n_508) );
OR2x2_ASAP7_75t_L g476 ( .A(n_322), .B(n_477), .Y(n_476) );
AOI221xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_330), .B1(n_335), .B2(n_337), .C(n_342), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g351 ( .A(n_326), .B(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OR2x2_ASAP7_75t_L g388 ( .A(n_327), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g408 ( .A(n_328), .Y(n_408) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
BUFx3_ASAP7_75t_L g431 ( .A(n_329), .Y(n_431) );
AND2x2_ASAP7_75t_L g438 ( .A(n_329), .B(n_439), .Y(n_438) );
INVxp67_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
OR2x2_ASAP7_75t_L g375 ( .A(n_332), .B(n_376), .Y(n_375) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_334), .B(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx2_ASAP7_75t_L g352 ( .A(n_339), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_339), .B(n_422), .Y(n_421) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
INVx2_ASAP7_75t_L g344 ( .A(n_341), .Y(n_344) );
OAI321xp33_ASAP7_75t_L g456 ( .A1(n_341), .A2(n_449), .A3(n_457), .B1(n_462), .B2(n_464), .C(n_468), .Y(n_456) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
OR2x2_ASAP7_75t_L g411 ( .A(n_344), .B(n_412), .Y(n_411) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g511 ( .A(n_347), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_348), .B(n_391), .Y(n_390) );
NAND2xp33_ASAP7_75t_SL g491 ( .A(n_348), .B(n_362), .Y(n_491) );
OAI211xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B(n_364), .C(n_368), .Y(n_349) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_354), .B(n_359), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g355 ( .A(n_356), .B(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g460 ( .A(n_357), .Y(n_460) );
INVx3_ASAP7_75t_L g399 ( .A(n_358), .Y(n_399) );
OR2x2_ASAP7_75t_L g502 ( .A(n_358), .B(n_376), .Y(n_502) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_360), .A2(n_444), .B1(n_446), .B2(n_448), .Y(n_443) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_SL g442 ( .A(n_363), .Y(n_442) );
OR2x2_ASAP7_75t_L g519 ( .A(n_363), .B(n_376), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
AOI21xp5_ASAP7_75t_SL g368 ( .A1(n_369), .A2(n_370), .B(n_374), .Y(n_368) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_372), .B(n_389), .Y(n_488) );
AND2x2_ASAP7_75t_L g494 ( .A(n_372), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g439 ( .A(n_373), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g374 ( .A1(n_375), .A2(n_378), .B1(n_381), .B2(n_383), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g420 ( .A1(n_376), .A2(n_419), .B(n_421), .C(n_423), .Y(n_420) );
INVx2_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_379), .B(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_379), .B(n_471), .Y(n_493) );
INVx2_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g465 ( .A(n_382), .B(n_466), .Y(n_465) );
INVx2_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
A2O1A1Ixp33_ASAP7_75t_L g415 ( .A1(n_384), .A2(n_416), .B(n_419), .C(n_420), .Y(n_415) );
NAND3xp33_ASAP7_75t_SL g385 ( .A(n_386), .B(n_400), .C(n_415), .Y(n_385) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_390), .B1(n_392), .B2(n_393), .C1(n_394), .C2(n_397), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g449 ( .A(n_389), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_389), .B(n_422), .Y(n_475) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_SL g409 ( .A(n_396), .Y(n_409) );
AND2x2_ASAP7_75t_L g397 ( .A(n_398), .B(n_399), .Y(n_397) );
OR2x2_ASAP7_75t_L g514 ( .A(n_398), .B(n_431), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_399), .A2(n_490), .B1(n_492), .B2(n_494), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_406), .B1(n_410), .B2(n_413), .C(n_414), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI21xp5_ASAP7_75t_SL g474 ( .A1(n_407), .A2(n_475), .B(n_476), .Y(n_474) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx2_ASAP7_75t_L g422 ( .A(n_408), .Y(n_422) );
AND2x2_ASAP7_75t_L g516 ( .A(n_408), .B(n_517), .Y(n_516) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g500 ( .A(n_412), .Y(n_500) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OR2x2_ASAP7_75t_L g429 ( .A(n_418), .B(n_419), .Y(n_429) );
INVx1_ASAP7_75t_L g482 ( .A(n_418), .Y(n_482) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_456), .C(n_478), .Y(n_424) );
OAI211xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_430), .B(n_432), .C(n_437), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g432 ( .A1(n_427), .A2(n_433), .B(n_434), .Y(n_432) );
INVx1_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI211xp5_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_440), .B(n_443), .C(n_450), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g461 ( .A(n_444), .Y(n_461) );
INVxp67_ASAP7_75t_SL g486 ( .A(n_445), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_447), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g509 ( .A(n_447), .Y(n_509) );
AND2x2_ASAP7_75t_L g499 ( .A(n_449), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g469 ( .A(n_451), .Y(n_469) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_455), .Y(n_452) );
INVx1_ASAP7_75t_L g477 ( .A(n_453), .Y(n_477) );
INVx2_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_461), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g462 ( .A(n_463), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g498 ( .A1(n_465), .A2(n_499), .B1(n_501), .B2(n_503), .C(n_508), .Y(n_498) );
OAI21xp33_ASAP7_75t_SL g513 ( .A1(n_470), .A2(n_514), .B(n_515), .Y(n_513) );
INVx2_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND4xp25_ASAP7_75t_L g478 ( .A(n_479), .B(n_489), .C(n_498), .D(n_512), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B1(n_486), .B2(n_487), .Y(n_479) );
AND2x4_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
INVx1_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_SL g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_507), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_521), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
OAI222xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_526), .B1(n_532), .B2(n_534), .C1(n_535), .C2(n_540), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g526 ( .A(n_527), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_528), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_536), .Y(n_535) );
INVxp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
endmodule