module fake_jpeg_2113_n_647 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_647);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_647;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVxp33_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_9),
.B(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx4f_ASAP7_75t_SL g44 ( 
.A(n_4),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_14),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_7),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_59),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_61),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_36),
.A2(n_0),
.B1(n_2),
.B2(n_4),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_62),
.A2(n_30),
.B1(n_19),
.B2(n_26),
.Y(n_188)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_32),
.Y(n_63)
);

INVx3_ASAP7_75t_L g199 ( 
.A(n_63),
.Y(n_199)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_52),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_64),
.Y(n_177)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_65),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_18),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_66),
.B(n_79),
.Y(n_141)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_68),
.Y(n_175)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_69),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_70),
.Y(n_134)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_71),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_38),
.B(n_15),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_72),
.B(n_83),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_56),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_73),
.Y(n_202)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_74),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_76),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_77),
.Y(n_189)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_27),
.B(n_12),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_80),
.Y(n_213)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g147 ( 
.A(n_82),
.Y(n_147)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_42),
.B(n_15),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_24),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_84),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_24),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_85),
.Y(n_183)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_34),
.Y(n_86)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_49),
.Y(n_87)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_87),
.Y(n_208)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_88),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_33),
.B(n_43),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_89),
.B(n_128),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_90),
.Y(n_190)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_91),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_45),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_127),
.Y(n_148)
);

BUFx12_ASAP7_75t_L g93 ( 
.A(n_44),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_93),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_54),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_94),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_95),
.B(n_99),
.Y(n_150)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_51),
.Y(n_96)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_96),
.Y(n_184)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_97),
.Y(n_220)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_98),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_56),
.Y(n_99)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_100),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_55),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_101),
.Y(n_214)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_102),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_55),
.Y(n_103)
);

INVx6_ASAP7_75t_L g156 ( 
.A(n_103),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx6_ASAP7_75t_L g176 ( 
.A(n_104),
.Y(n_176)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_44),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g223 ( 
.A(n_105),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_106),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_20),
.Y(n_107)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_21),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_108),
.Y(n_154)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_58),
.Y(n_109)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_20),
.Y(n_110)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_20),
.Y(n_111)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_29),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_114),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_29),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_29),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_115),
.B(n_123),
.Y(n_160)
);

BUFx24_ASAP7_75t_L g116 ( 
.A(n_36),
.Y(n_116)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_116),
.Y(n_204)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_52),
.Y(n_118)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_118),
.Y(n_155)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_119),
.Y(n_157)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx8_ASAP7_75t_L g195 ( 
.A(n_120),
.Y(n_195)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_25),
.Y(n_121)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_121),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_31),
.Y(n_122)
);

INVx8_ASAP7_75t_L g200 ( 
.A(n_122),
.Y(n_200)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_31),
.Y(n_124)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_124),
.Y(n_162)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_23),
.Y(n_125)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_125),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_126),
.Y(n_163)
);

INVx2_ASAP7_75t_SL g127 ( 
.A(n_46),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_27),
.B(n_12),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_46),
.Y(n_129)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_129),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_83),
.B(n_53),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_149),
.B(n_153),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_105),
.Y(n_151)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_151),
.B(n_116),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_106),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_80),
.B(n_43),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_158),
.B(n_161),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_108),
.B(n_37),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_129),
.B(n_53),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_166),
.B(n_170),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_120),
.A2(n_124),
.B1(n_126),
.B2(n_122),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_167),
.A2(n_104),
.B1(n_103),
.B2(n_101),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g168 ( 
.A1(n_88),
.A2(n_19),
.B1(n_57),
.B2(n_26),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_168),
.A2(n_188),
.B1(n_205),
.B2(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_75),
.B(n_37),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_75),
.B(n_77),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_171),
.B(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_67),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_173),
.B(n_174),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_74),
.Y(n_174)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_100),
.Y(n_178)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_178),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_107),
.B(n_47),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_77),
.B(n_30),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_182),
.B(n_187),
.Y(n_251)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_185),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_111),
.B(n_47),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_70),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_192),
.B(n_197),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_76),
.B(n_41),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_194),
.B(n_198),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_84),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_98),
.B(n_41),
.Y(n_198)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_85),
.Y(n_201)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_201),
.Y(n_248)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_90),
.Y(n_203)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_203),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_112),
.A2(n_19),
.B1(n_57),
.B2(n_50),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_SL g207 ( 
.A(n_116),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_207),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_93),
.B(n_39),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_209),
.B(n_210),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_82),
.B(n_39),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_28),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_212),
.B(n_218),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_94),
.B(n_28),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_65),
.A2(n_50),
.B1(n_46),
.B2(n_48),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_226),
.A2(n_273),
.B1(n_285),
.B2(n_292),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_165),
.A2(n_50),
.B1(n_35),
.B2(n_48),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_227),
.A2(n_246),
.B1(n_274),
.B2(n_281),
.Y(n_363)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_217),
.Y(n_228)
);

INVx4_ASAP7_75t_L g339 ( 
.A(n_228),
.Y(n_339)
);

INVx4_ASAP7_75t_L g230 ( 
.A(n_155),
.Y(n_230)
);

INVx4_ASAP7_75t_L g343 ( 
.A(n_230),
.Y(n_343)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_181),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_231),
.Y(n_362)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_217),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g357 ( 
.A(n_233),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_134),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_234),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g346 ( 
.A(n_236),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx11_ASAP7_75t_L g304 ( 
.A(n_237),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_146),
.B(n_86),
.Y(n_238)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_238),
.Y(n_305)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_239),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_71),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_240),
.B(n_256),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_202),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_241),
.B(n_255),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_243),
.Y(n_319)
);

INVx5_ASAP7_75t_L g244 ( 
.A(n_217),
.Y(n_244)
);

INVx3_ASAP7_75t_L g322 ( 
.A(n_244),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_L g246 ( 
.A1(n_139),
.A2(n_48),
.B1(n_35),
.B2(n_62),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_184),
.Y(n_249)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_162),
.Y(n_250)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_250),
.Y(n_321)
);

A2O1A1O1Ixp25_ASAP7_75t_L g252 ( 
.A1(n_135),
.A2(n_102),
.B(n_21),
.C(n_15),
.D(n_12),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_252),
.B(n_291),
.Y(n_360)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_196),
.Y(n_253)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_253),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_148),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_220),
.B(n_2),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_148),
.B(n_4),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_257),
.Y(n_332)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_219),
.Y(n_259)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g262 ( 
.A(n_151),
.B(n_5),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g336 ( 
.A(n_262),
.Y(n_336)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_160),
.Y(n_263)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_263),
.Y(n_318)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_131),
.Y(n_264)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_264),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_204),
.B(n_5),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_150),
.B(n_5),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_266),
.B(n_267),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_159),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_175),
.B(n_147),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_268),
.B(n_272),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_205),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_269),
.A2(n_164),
.B1(n_140),
.B2(n_193),
.Y(n_353)
);

INVx3_ASAP7_75t_L g270 ( 
.A(n_204),
.Y(n_270)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_270),
.Y(n_342)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_172),
.Y(n_271)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_271),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_147),
.B(n_6),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_221),
.A2(n_143),
.B1(n_138),
.B2(n_211),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_156),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_136),
.Y(n_275)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_275),
.Y(n_344)
);

INVx4_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_276),
.Y(n_361)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_130),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_277),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_172),
.Y(n_278)
);

BUFx2_ASAP7_75t_SL g312 ( 
.A(n_278),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_142),
.Y(n_279)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_279),
.Y(n_334)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_213),
.Y(n_280)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_280),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_156),
.A2(n_6),
.B1(n_10),
.B2(n_176),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_130),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_283),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_133),
.Y(n_283)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_180),
.Y(n_284)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_176),
.A2(n_10),
.B1(n_191),
.B2(n_214),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_152),
.B(n_10),
.Y(n_286)
);

NOR2x1_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_288),
.Y(n_306)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_157),
.Y(n_287)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_287),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_186),
.B(n_199),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_154),
.B(n_10),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_290),
.B(n_293),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_208),
.B(n_169),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g292 ( 
.A1(n_168),
.A2(n_191),
.B1(n_163),
.B2(n_206),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_163),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_177),
.B(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_294),
.B(n_295),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_189),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_195),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_296),
.B(n_298),
.Y(n_354)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_180),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_297),
.Y(n_307)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_133),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_223),
.B(n_190),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_300),
.B(n_211),
.Y(n_314)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_131),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_301),
.Y(n_310)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_137),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_302),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_247),
.B(n_213),
.C(n_177),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_309),
.B(n_330),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_232),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_313),
.B(n_314),
.Y(n_364)
);

OA22x2_ASAP7_75t_L g315 ( 
.A1(n_229),
.A2(n_145),
.B1(n_222),
.B2(n_137),
.Y(n_315)
);

INVx3_ASAP7_75t_L g393 ( 
.A(n_315),
.Y(n_393)
);

OAI22xp33_ASAP7_75t_SL g316 ( 
.A1(n_246),
.A2(n_229),
.B1(n_227),
.B2(n_261),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_316),
.A2(n_305),
.B1(n_319),
.B2(n_363),
.Y(n_379)
);

OA22x2_ASAP7_75t_L g326 ( 
.A1(n_269),
.A2(n_145),
.B1(n_222),
.B2(n_164),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_253),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_235),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_329),
.B(n_338),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_238),
.B(n_132),
.C(n_214),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_273),
.A2(n_195),
.B1(n_206),
.B2(n_183),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_333),
.A2(n_341),
.B1(n_225),
.B2(n_271),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_291),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_243),
.A2(n_216),
.B(n_144),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g389 ( 
.A1(n_340),
.A2(n_233),
.B(n_239),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_292),
.A2(n_190),
.B1(n_183),
.B2(n_140),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_228),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_244),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_314),
.B(n_251),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_365),
.B(n_370),
.Y(n_419)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_337),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g438 ( 
.A(n_367),
.Y(n_438)
);

INVx13_ASAP7_75t_L g368 ( 
.A(n_304),
.Y(n_368)
);

BUFx8_ASAP7_75t_L g426 ( 
.A(n_368),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g369 ( 
.A(n_328),
.B(n_299),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g422 ( 
.A(n_369),
.B(n_381),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_306),
.B(n_258),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_371),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_354),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_377),
.Y(n_415)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_321),
.Y(n_374)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_374),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_306),
.B(n_260),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_376),
.Y(n_437)
);

A2O1A1Ixp33_ASAP7_75t_L g376 ( 
.A1(n_360),
.A2(n_257),
.B(n_252),
.C(n_262),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_323),
.Y(n_377)
);

INVx1_ASAP7_75t_SL g378 ( 
.A(n_340),
.Y(n_378)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_378),
.Y(n_429)
);

OAI22xp33_ASAP7_75t_SL g423 ( 
.A1(n_379),
.A2(n_382),
.B1(n_399),
.B2(n_403),
.Y(n_423)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_321),
.Y(n_380)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_380),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_351),
.B(n_303),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_356),
.Y(n_383)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_383),
.Y(n_441)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_298),
.B1(n_276),
.B2(n_277),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g439 ( 
.A(n_384),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_385),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_320),
.A2(n_264),
.B1(n_250),
.B2(n_224),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_386),
.A2(n_404),
.B1(n_359),
.B2(n_317),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_348),
.A2(n_265),
.B(n_270),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_326),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_349),
.B(n_348),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_388),
.B(n_396),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g449 ( 
.A(n_389),
.B(n_408),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_335),
.B(n_245),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_390),
.B(n_398),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_SL g391 ( 
.A1(n_307),
.A2(n_230),
.B1(n_280),
.B2(n_295),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_391),
.Y(n_424)
);

OR2x2_ASAP7_75t_L g392 ( 
.A(n_360),
.B(n_225),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_392),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g394 ( 
.A(n_344),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g420 ( 
.A(n_394),
.B(n_352),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_309),
.B(n_242),
.Y(n_396)
);

INVx6_ASAP7_75t_SL g397 ( 
.A(n_357),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_397),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_362),
.B(n_248),
.Y(n_398)
);

AOI22xp33_ASAP7_75t_SL g399 ( 
.A1(n_315),
.A2(n_279),
.B1(n_132),
.B2(n_223),
.Y(n_399)
);

INVx8_ASAP7_75t_L g400 ( 
.A(n_312),
.Y(n_400)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_400),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_401),
.A2(n_407),
.B1(n_342),
.B2(n_317),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_360),
.B(n_324),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_402),
.Y(n_421)
);

AOI22xp33_ASAP7_75t_L g403 ( 
.A1(n_320),
.A2(n_254),
.B1(n_278),
.B2(n_234),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_333),
.A2(n_193),
.B1(n_200),
.B2(n_236),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_297),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_405),
.B(n_406),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_284),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_341),
.A2(n_200),
.B1(n_132),
.B2(n_237),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_336),
.A2(n_237),
.B(n_332),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_358),
.B(n_308),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_409),
.B(n_342),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_339),
.Y(n_410)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_410),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_395),
.B(n_396),
.C(n_364),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_412),
.B(n_432),
.Y(n_467)
);

OAI32xp33_ASAP7_75t_L g413 ( 
.A1(n_375),
.A2(n_330),
.A3(n_355),
.B1(n_358),
.B2(n_344),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_413),
.B(n_392),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_414),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_395),
.B(n_345),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_SL g472 ( 
.A(n_416),
.B(n_433),
.Y(n_472)
);

AOI32xp33_ASAP7_75t_L g418 ( 
.A1(n_366),
.A2(n_310),
.A3(n_311),
.B1(n_343),
.B2(n_315),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_418),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_420),
.Y(n_485)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_427),
.A2(n_401),
.B1(n_444),
.B2(n_407),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_379),
.A2(n_393),
.B1(n_382),
.B2(n_386),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g456 ( 
.A1(n_428),
.A2(n_393),
.B1(n_382),
.B2(n_403),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_334),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_430),
.B(n_442),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_409),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_431),
.B(n_373),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_364),
.B(n_325),
.C(n_361),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_325),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_381),
.B(n_357),
.Y(n_442)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_444),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g453 ( 
.A(n_448),
.B(n_366),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g507 ( 
.A(n_453),
.B(n_455),
.Y(n_507)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_449),
.A2(n_414),
.B(n_429),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_454),
.A2(n_459),
.B(n_463),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_456),
.A2(n_468),
.B1(n_408),
.B2(n_434),
.Y(n_509)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_441),
.Y(n_457)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_438),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_458),
.B(n_460),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g459 ( 
.A1(n_449),
.A2(n_393),
.B(n_378),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_438),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_441),
.Y(n_461)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_461),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_429),
.A2(n_378),
.B(n_389),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g501 ( 
.A(n_462),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_421),
.A2(n_387),
.B(n_392),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_464),
.A2(n_476),
.B1(n_432),
.B2(n_411),
.Y(n_500)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_417),
.Y(n_465)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_465),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_L g466 ( 
.A1(n_436),
.A2(n_372),
.B(n_402),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_466),
.B(n_411),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_428),
.A2(n_402),
.B1(n_370),
.B2(n_404),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g470 ( 
.A(n_415),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_470),
.B(n_471),
.Y(n_490)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_439),
.A2(n_385),
.B(n_397),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_446),
.B(n_406),
.Y(n_473)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_473),
.Y(n_505)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_417),
.Y(n_474)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_474),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_445),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_478),
.Y(n_494)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_425),
.Y(n_477)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_477),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_446),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_433),
.B(n_405),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_479),
.B(n_480),
.Y(n_497)
);

NOR2x1_ASAP7_75t_L g480 ( 
.A(n_437),
.B(n_421),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_425),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_481),
.B(n_483),
.Y(n_502)
);

INVx13_ASAP7_75t_L g482 ( 
.A(n_426),
.Y(n_482)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_482),
.Y(n_506)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_435),
.Y(n_483)
);

INVx13_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_484),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_487),
.B(n_480),
.Y(n_529)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_467),
.B(n_412),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_491),
.B(n_514),
.C(n_519),
.Y(n_521)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_467),
.B(n_416),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_492),
.B(n_508),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_469),
.A2(n_437),
.B1(n_440),
.B2(n_427),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_493),
.A2(n_503),
.B1(n_509),
.B2(n_511),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g495 ( 
.A(n_455),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_495),
.B(n_498),
.Y(n_536)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_451),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_470),
.B(n_369),
.Y(n_499)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_499),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_500),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_464),
.A2(n_419),
.B1(n_423),
.B2(n_424),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_453),
.B(n_390),
.Y(n_504)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_504),
.Y(n_538)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_419),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_451),
.B(n_485),
.Y(n_510)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_510),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_450),
.A2(n_424),
.B1(n_439),
.B2(n_413),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_468),
.A2(n_435),
.B1(n_422),
.B2(n_443),
.Y(n_512)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_472),
.B(n_388),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_SL g515 ( 
.A1(n_450),
.A2(n_443),
.B1(n_315),
.B2(n_447),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_515),
.B(n_456),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_479),
.B(n_376),
.Y(n_519)
);

AOI22xp5_ASAP7_75t_SL g556 ( 
.A1(n_520),
.A2(n_511),
.B1(n_501),
.B2(n_515),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_494),
.B(n_460),
.Y(n_523)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_523),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_501),
.A2(n_459),
.B(n_454),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g570 ( 
.A(n_525),
.B(n_529),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_494),
.B(n_458),
.Y(n_526)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_526),
.Y(n_563)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_502),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_527),
.B(n_530),
.Y(n_555)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_502),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_507),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_532),
.B(n_533),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_507),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_488),
.Y(n_534)
);

AOI22xp33_ASAP7_75t_SL g562 ( 
.A1(n_534),
.A2(n_541),
.B1(n_545),
.B2(n_546),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_491),
.B(n_452),
.C(n_466),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_537),
.C(n_540),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_492),
.B(n_452),
.C(n_478),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_SL g540 ( 
.A(n_490),
.B(n_503),
.C(n_493),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_488),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_514),
.B(n_463),
.C(n_475),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_542),
.B(n_547),
.C(n_521),
.Y(n_553)
);

HB1xp67_ASAP7_75t_L g543 ( 
.A(n_506),
.Y(n_543)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_543),
.Y(n_564)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_505),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_505),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_473),
.C(n_462),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_480),
.Y(n_548)
);

CKINVDCx14_ASAP7_75t_R g569 ( 
.A(n_548),
.Y(n_569)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_486),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_549),
.A2(n_457),
.B1(n_461),
.B2(n_481),
.Y(n_566)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_544),
.A2(n_509),
.B1(n_512),
.B2(n_497),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g587 ( 
.A1(n_550),
.A2(n_552),
.B1(n_558),
.B2(n_561),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_524),
.A2(n_490),
.B1(n_476),
.B2(n_471),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g591 ( 
.A(n_553),
.B(n_559),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_SL g554 ( 
.A(n_542),
.B(n_519),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g575 ( 
.A(n_554),
.B(n_565),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_556),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g558 ( 
.A1(n_528),
.A2(n_517),
.B1(n_518),
.B2(n_489),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_531),
.B(n_517),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_R g560 ( 
.A(n_548),
.B(n_516),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_571),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_522),
.A2(n_513),
.B1(n_496),
.B2(n_474),
.Y(n_561)
);

XNOR2xp5_ASAP7_75t_SL g565 ( 
.A(n_535),
.B(n_376),
.Y(n_565)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_566),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g567 ( 
.A1(n_544),
.A2(n_522),
.B1(n_520),
.B2(n_534),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_567),
.A2(n_526),
.B1(n_549),
.B2(n_477),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_531),
.B(n_465),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_568),
.B(n_530),
.C(n_527),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_521),
.B(n_537),
.C(n_547),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_573),
.B(n_554),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g576 ( 
.A(n_551),
.B(n_540),
.C(n_525),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_576),
.B(n_579),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_564),
.B(n_539),
.Y(n_579)
);

BUFx12_ASAP7_75t_L g580 ( 
.A(n_568),
.Y(n_580)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_580),
.Y(n_593)
);

AOI21xp5_ASAP7_75t_SL g581 ( 
.A1(n_563),
.A2(n_572),
.B(n_523),
.Y(n_581)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_581),
.Y(n_601)
);

INVxp67_ASAP7_75t_L g582 ( 
.A(n_562),
.Y(n_582)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_582),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_560),
.B(n_536),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_583),
.B(n_585),
.Y(n_603)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_567),
.A2(n_550),
.B(n_555),
.Y(n_584)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_584),
.B(n_588),
.Y(n_599)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_557),
.Y(n_585)
);

CKINVDCx20_ASAP7_75t_R g586 ( 
.A(n_569),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_586),
.B(n_589),
.Y(n_606)
);

CKINVDCx16_ASAP7_75t_R g589 ( 
.A(n_570),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_551),
.B(n_483),
.C(n_447),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_590),
.B(n_559),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_538),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_592),
.B(n_594),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_591),
.B(n_571),
.C(n_553),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_584),
.A2(n_570),
.B1(n_558),
.B2(n_561),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_595),
.B(n_598),
.Y(n_610)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_597),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_SL g598 ( 
.A(n_574),
.B(n_383),
.Y(n_598)
);

BUFx24_ASAP7_75t_SL g600 ( 
.A(n_591),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_600),
.B(n_602),
.Y(n_608)
);

BUFx24_ASAP7_75t_SL g602 ( 
.A(n_581),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_604),
.B(n_605),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_576),
.B(n_556),
.C(n_565),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_594),
.B(n_584),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g624 ( 
.A(n_609),
.B(n_612),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g612 ( 
.A(n_596),
.B(n_606),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_603),
.B(n_607),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_613),
.B(n_614),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_593),
.B(n_573),
.C(n_587),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_599),
.B(n_605),
.C(n_582),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_615),
.B(n_410),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_L g616 ( 
.A(n_599),
.B(n_577),
.Y(n_616)
);

INVxp67_ASAP7_75t_L g629 ( 
.A(n_616),
.Y(n_629)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_601),
.A2(n_578),
.B1(n_575),
.B2(n_580),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g626 ( 
.A1(n_617),
.A2(n_380),
.B1(n_374),
.B2(n_484),
.Y(n_626)
);

OAI21xp5_ASAP7_75t_SL g619 ( 
.A1(n_596),
.A2(n_578),
.B(n_580),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g623 ( 
.A1(n_619),
.A2(n_426),
.B(n_484),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_618),
.B(n_506),
.C(n_359),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_622),
.B(n_623),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_398),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_625),
.B(n_624),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_626),
.B(n_627),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_620),
.A2(n_371),
.B(n_410),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_628),
.B(n_630),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_610),
.A2(n_482),
.B1(n_346),
.B2(n_367),
.Y(n_630)
);

AOI322xp5_ASAP7_75t_L g631 ( 
.A1(n_621),
.A2(n_611),
.A3(n_614),
.B1(n_615),
.B2(n_617),
.C1(n_616),
.C2(n_482),
.Y(n_631)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_631),
.A2(n_632),
.B(n_400),
.Y(n_640)
);

AOI322xp5_ASAP7_75t_L g632 ( 
.A1(n_629),
.A2(n_368),
.A3(n_400),
.B1(n_346),
.B2(n_326),
.C1(n_361),
.C2(n_327),
.Y(n_632)
);

NOR2x1_ASAP7_75t_L g638 ( 
.A(n_635),
.B(n_327),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g637 ( 
.A(n_633),
.B(n_629),
.C(n_622),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_637),
.B(n_638),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_636),
.B(n_634),
.Y(n_639)
);

AOI322xp5_ASAP7_75t_L g641 ( 
.A1(n_639),
.A2(n_640),
.A3(n_368),
.B1(n_326),
.B2(n_304),
.C1(n_322),
.C2(n_339),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g643 ( 
.A1(n_641),
.A2(n_642),
.B(n_322),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_643),
.B(n_331),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_644),
.B(n_331),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g646 ( 
.A(n_645),
.B(n_352),
.Y(n_646)
);

BUFx24_ASAP7_75t_SL g647 ( 
.A(n_646),
.Y(n_647)
);


endmodule