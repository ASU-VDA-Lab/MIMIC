module fake_netlist_6_2296_n_1845 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1845);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1845;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_1058;
wire n_854;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_L g170 ( 
.A(n_28),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_87),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g172 ( 
.A(n_117),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_84),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_141),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_79),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_152),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_149),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_30),
.Y(n_178)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_119),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_68),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_43),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_48),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_59),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_145),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_99),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_19),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_9),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_73),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_93),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_18),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_112),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_22),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_75),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_103),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_70),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_148),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_136),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_156),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_139),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_32),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_6),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_14),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_2),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_33),
.Y(n_209)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_137),
.Y(n_211)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_96),
.Y(n_213)
);

BUFx10_ASAP7_75t_L g214 ( 
.A(n_44),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g215 ( 
.A(n_22),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_77),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_54),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_165),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_33),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_46),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_60),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_31),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_52),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_126),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_124),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_95),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_157),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_45),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_160),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_19),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_82),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_18),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_39),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_83),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_36),
.Y(n_238)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_107),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_74),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_106),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_4),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_21),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_72),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_16),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_2),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_40),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_132),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_24),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_7),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_151),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_94),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_131),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_40),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_111),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g257 ( 
.A(n_110),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_109),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_11),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_143),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_146),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_127),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_80),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_42),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_64),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_32),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_58),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_108),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_92),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_125),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_28),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_101),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_9),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_150),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_105),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_42),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_70),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_8),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_159),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_166),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_61),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_27),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_102),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_43),
.Y(n_286)
);

BUFx3_ASAP7_75t_L g287 ( 
.A(n_133),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_67),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_29),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_34),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_121),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_56),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_5),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_16),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_27),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_46),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_114),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_29),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_15),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_6),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_69),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_63),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_7),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_65),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_71),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_24),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_57),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_155),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_104),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_13),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_45),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_154),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_60),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_26),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_21),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_8),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_13),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_163),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_169),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_12),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_135),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_89),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_20),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_0),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_116),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g328 ( 
.A(n_10),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_130),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_65),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_25),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_26),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_76),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_47),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_30),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_17),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_37),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_67),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_39),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_53),
.Y(n_340)
);

BUFx10_ASAP7_75t_L g341 ( 
.A(n_100),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_49),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_225),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_239),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_225),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_225),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_225),
.Y(n_347)
);

INVxp33_ASAP7_75t_L g348 ( 
.A(n_239),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_225),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_266),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_173),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_266),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_328),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_266),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_179),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_266),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_186),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_272),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_272),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_328),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g362 ( 
.A(n_192),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_272),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_272),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_272),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_171),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_178),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_267),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_267),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_314),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_267),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_170),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_175),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_177),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_170),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_180),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_180),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_191),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_194),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_197),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_314),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_172),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_172),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_209),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_253),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_174),
.B(n_0),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_182),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_209),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_310),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_184),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_183),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_310),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_196),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_210),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_184),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_337),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_205),
.Y(n_398)
);

INVxp33_ASAP7_75t_L g399 ( 
.A(n_205),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_255),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_208),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_282),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_208),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_221),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_187),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_174),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_285),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_210),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_224),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_261),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_224),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_212),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_198),
.Y(n_414)
);

CKINVDCx16_ASAP7_75t_R g415 ( 
.A(n_261),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_226),
.Y(n_416)
);

INVxp33_ASAP7_75t_L g417 ( 
.A(n_226),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_236),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_236),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_238),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_238),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_313),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_243),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_243),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_201),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_248),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_248),
.Y(n_427)
);

CKINVDCx16_ASAP7_75t_R g428 ( 
.A(n_199),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_202),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_203),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g431 ( 
.A(n_251),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_212),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_343),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_343),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_383),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_368),
.B(n_181),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_366),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_345),
.Y(n_438)
);

CKINVDCx9p33_ASAP7_75t_R g439 ( 
.A(n_354),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_373),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_354),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_391),
.A2(n_284),
.B1(n_259),
.B2(n_299),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_369),
.B(n_234),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_400),
.A2(n_330),
.B1(n_283),
.B2(n_339),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_374),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_346),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_346),
.Y(n_448)
);

INVxp33_ASAP7_75t_L g449 ( 
.A(n_405),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_347),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_347),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_349),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_367),
.B(n_211),
.Y(n_453)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_395),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_349),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_L g456 ( 
.A(n_378),
.B(n_379),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_350),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_350),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_344),
.A2(n_215),
.B1(n_293),
.B2(n_326),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_352),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_394),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_352),
.Y(n_462)
);

AND2x6_ASAP7_75t_L g463 ( 
.A(n_369),
.B(n_181),
.Y(n_463)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_408),
.B(n_234),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_353),
.Y(n_465)
);

INVx3_ASAP7_75t_L g466 ( 
.A(n_353),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_414),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_361),
.A2(n_342),
.B1(n_340),
.B2(n_336),
.Y(n_468)
);

AND2x4_ASAP7_75t_L g469 ( 
.A(n_371),
.B(n_287),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_355),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_355),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_425),
.Y(n_472)
);

BUFx3_ASAP7_75t_L g473 ( 
.A(n_357),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_387),
.B(n_245),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_351),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_357),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_413),
.B(n_213),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_359),
.Y(n_478)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_370),
.B(n_287),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_358),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_359),
.B(n_220),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_381),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g483 ( 
.A1(n_380),
.A2(n_342),
.B1(n_340),
.B2(n_336),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_360),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_348),
.A2(n_286),
.B1(n_188),
.B2(n_277),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_429),
.Y(n_486)
);

CKINVDCx20_ASAP7_75t_R g487 ( 
.A(n_402),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_360),
.Y(n_488)
);

OAI21x1_ASAP7_75t_L g489 ( 
.A1(n_406),
.A2(n_371),
.B(n_258),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_363),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_363),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_399),
.B(n_251),
.Y(n_492)
);

OAI21x1_ASAP7_75t_L g493 ( 
.A1(n_406),
.A2(n_258),
.B(n_219),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_407),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_422),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g496 ( 
.A(n_364),
.B(n_219),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_364),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_356),
.B(n_257),
.Y(n_498)
);

OA22x2_ASAP7_75t_SL g499 ( 
.A1(n_398),
.A2(n_264),
.B1(n_265),
.B2(n_332),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_430),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_365),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_365),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_372),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_362),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_398),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_401),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_386),
.B(n_227),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_401),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_385),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_229),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_442),
.Y(n_511)
);

NAND2xp33_ASAP7_75t_R g512 ( 
.A(n_504),
.B(n_189),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_435),
.B(n_232),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_435),
.B(n_372),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_464),
.B(n_375),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_483),
.A2(n_193),
.B1(n_250),
.B2(n_247),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_442),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_237),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_489),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_448),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_489),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_448),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_489),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_454),
.B(n_411),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_473),
.Y(n_525)
);

NAND3xp33_ASAP7_75t_L g526 ( 
.A(n_498),
.B(n_396),
.C(n_390),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_454),
.B(n_415),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_473),
.Y(n_528)
);

INVx1_ASAP7_75t_SL g529 ( 
.A(n_480),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_477),
.B(n_507),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_473),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_501),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_501),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_448),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_470),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_450),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_443),
.A2(n_428),
.B1(n_265),
.B2(n_264),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_450),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_450),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_501),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_433),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_507),
.B(n_240),
.Y(n_542)
);

BUFx6f_ASAP7_75t_L g543 ( 
.A(n_493),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_451),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_451),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_481),
.Y(n_546)
);

INVx4_ASAP7_75t_L g547 ( 
.A(n_470),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

INVx2_ASAP7_75t_SL g549 ( 
.A(n_479),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_432),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_451),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_452),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_452),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_453),
.B(n_417),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_438),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_437),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_479),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_432),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_470),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_482),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_452),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_447),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_460),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_481),
.B(n_241),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_474),
.B(n_419),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_460),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_470),
.Y(n_569)
);

INVx8_ASAP7_75t_L g570 ( 
.A(n_436),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_460),
.Y(n_571)
);

BUFx16f_ASAP7_75t_R g572 ( 
.A(n_439),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_449),
.B(n_431),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_464),
.B(n_242),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_434),
.Y(n_575)
);

INVx3_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_493),
.Y(n_577)
);

OAI22xp33_ASAP7_75t_SL g578 ( 
.A1(n_485),
.A2(n_269),
.B1(n_273),
.B2(n_319),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_440),
.B(n_249),
.Y(n_579)
);

OR2x2_ASAP7_75t_L g580 ( 
.A(n_482),
.B(n_416),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_464),
.B(n_252),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_446),
.Y(n_583)
);

BUFx6f_ASAP7_75t_SL g584 ( 
.A(n_432),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_461),
.B(n_249),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_455),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_434),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_455),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_457),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_457),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_434),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_432),
.B(n_254),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_493),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_467),
.B(n_249),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_503),
.Y(n_595)
);

INVx8_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

INVxp33_ASAP7_75t_L g597 ( 
.A(n_443),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_492),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_458),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_458),
.Y(n_600)
);

INVx3_ASAP7_75t_L g601 ( 
.A(n_488),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_465),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_465),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_444),
.B(n_176),
.Y(n_604)
);

OAI22xp33_ASAP7_75t_L g605 ( 
.A1(n_485),
.A2(n_246),
.B1(n_235),
.B2(n_338),
.Y(n_605)
);

INVx2_ASAP7_75t_SL g606 ( 
.A(n_492),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_503),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_471),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_503),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_488),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_503),
.Y(n_611)
);

NOR2x1p5_ASAP7_75t_L g612 ( 
.A(n_509),
.B(n_274),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_471),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_472),
.B(n_249),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_486),
.B(n_341),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_476),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_503),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_503),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_476),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_478),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_488),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_478),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_444),
.B(n_341),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_488),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_459),
.B(n_421),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_444),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_434),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_441),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_484),
.Y(n_629)
);

INVxp67_ASAP7_75t_SL g630 ( 
.A(n_488),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_441),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_484),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_441),
.Y(n_633)
);

BUFx6f_ASAP7_75t_L g634 ( 
.A(n_488),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_483),
.A2(n_292),
.B1(n_290),
.B2(n_335),
.Y(n_635)
);

AND2x2_ASAP7_75t_L g636 ( 
.A(n_469),
.B(n_375),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_490),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_469),
.B(n_341),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_441),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_469),
.B(n_490),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_496),
.B(n_176),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_L g642 ( 
.A(n_456),
.B(n_195),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_497),
.Y(n_643)
);

INVx3_ASAP7_75t_L g644 ( 
.A(n_462),
.Y(n_644)
);

INVx4_ASAP7_75t_L g645 ( 
.A(n_436),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_497),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_502),
.Y(n_648)
);

AOI22xp33_ASAP7_75t_L g649 ( 
.A1(n_468),
.A2(n_279),
.B1(n_288),
.B2(n_294),
.Y(n_649)
);

HB1xp67_ASAP7_75t_L g650 ( 
.A(n_480),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_475),
.Y(n_652)
);

OAI22xp33_ASAP7_75t_L g653 ( 
.A1(n_459),
.A2(n_298),
.B1(n_206),
.B2(n_207),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_462),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_462),
.Y(n_655)
);

OAI21xp33_ASAP7_75t_SL g656 ( 
.A1(n_505),
.A2(n_279),
.B(n_274),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_506),
.Y(n_657)
);

INVx2_ASAP7_75t_SL g658 ( 
.A(n_496),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_462),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_466),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_530),
.B(n_466),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_636),
.Y(n_662)
);

INVxp67_ASAP7_75t_L g663 ( 
.A(n_573),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_546),
.B(n_466),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_549),
.B(n_559),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_636),
.Y(n_666)
);

INVx2_ASAP7_75t_SL g667 ( 
.A(n_511),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_555),
.B(n_468),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_549),
.B(n_466),
.Y(n_669)
);

NAND2x1p5_ASAP7_75t_L g670 ( 
.A(n_550),
.B(n_185),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_559),
.B(n_491),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_567),
.B(n_491),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_550),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_550),
.Y(n_674)
);

OAI22xp5_ASAP7_75t_L g675 ( 
.A1(n_598),
.A2(n_275),
.B1(n_185),
.B2(n_204),
.Y(n_675)
);

BUFx8_ASAP7_75t_L g676 ( 
.A(n_511),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_606),
.B(n_658),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_606),
.A2(n_319),
.B1(n_276),
.B2(n_273),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_562),
.B(n_500),
.Y(n_679)
);

NOR3xp33_ASAP7_75t_L g680 ( 
.A(n_537),
.B(n_445),
.C(n_500),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_560),
.Y(n_681)
);

INVxp67_ASAP7_75t_L g682 ( 
.A(n_524),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_560),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_658),
.B(n_181),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_560),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_527),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_619),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_626),
.B(n_181),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_510),
.B(n_445),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g690 ( 
.A(n_558),
.B(n_487),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_542),
.B(n_491),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_513),
.B(n_218),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_626),
.B(n_181),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_518),
.B(n_491),
.Y(n_694)
);

AOI22xp33_ASAP7_75t_L g695 ( 
.A1(n_604),
.A2(n_217),
.B1(n_308),
.B2(n_305),
.Y(n_695)
);

AOI22xp33_ASAP7_75t_L g696 ( 
.A1(n_604),
.A2(n_217),
.B1(n_308),
.B2(n_305),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_566),
.B(n_190),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_525),
.B(n_190),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_651),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_525),
.B(n_200),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_528),
.B(n_200),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_657),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_528),
.B(n_204),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_519),
.B(n_256),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_619),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_531),
.B(n_216),
.Y(n_706)
);

NAND3x1_ASAP7_75t_L g707 ( 
.A(n_516),
.B(n_294),
.C(n_288),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_531),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_L g709 ( 
.A(n_574),
.B(n_223),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_620),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_532),
.B(n_216),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_532),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_519),
.B(n_260),
.Y(n_713)
);

INVx8_ASAP7_75t_L g714 ( 
.A(n_584),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_604),
.A2(n_309),
.B1(n_228),
.B2(n_269),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_533),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_620),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_581),
.B(n_231),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_642),
.B(n_580),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_580),
.B(n_233),
.Y(n_720)
);

AOI22xp33_ASAP7_75t_L g721 ( 
.A1(n_604),
.A2(n_323),
.B1(n_309),
.B2(n_320),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_533),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_519),
.B(n_262),
.Y(n_723)
);

INVx5_ASAP7_75t_L g724 ( 
.A(n_519),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_648),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_648),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_514),
.B(n_268),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_540),
.B(n_222),
.Y(n_728)
);

A2O1A1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_640),
.A2(n_222),
.B(n_228),
.C(n_230),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_517),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_541),
.Y(n_731)
);

OR2x6_ASAP7_75t_L g732 ( 
.A(n_650),
.B(n_439),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_514),
.B(n_278),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_541),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_540),
.Y(n_735)
);

NOR2xp67_ASAP7_75t_SL g736 ( 
.A(n_645),
.B(n_230),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_517),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_644),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_526),
.B(n_289),
.C(n_280),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_515),
.B(n_295),
.Y(n_740)
);

NOR3xp33_ASAP7_75t_L g741 ( 
.A(n_537),
.B(n_302),
.C(n_301),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_519),
.B(n_263),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_515),
.B(n_304),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_583),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_641),
.A2(n_322),
.B1(n_276),
.B2(n_320),
.Y(n_745)
);

BUFx6f_ASAP7_75t_SL g746 ( 
.A(n_583),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_529),
.B(n_508),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_553),
.B(n_275),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_SL g749 ( 
.A(n_583),
.B(n_494),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_516),
.B(n_635),
.C(n_649),
.Y(n_750)
);

O2A1O1Ixp33_ASAP7_75t_L g751 ( 
.A1(n_578),
.A2(n_508),
.B(n_331),
.C(n_303),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_553),
.B(n_322),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_583),
.B(n_199),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_543),
.B(n_270),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_543),
.B(n_271),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_556),
.B(n_323),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_556),
.B(n_333),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_557),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_557),
.B(n_333),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_612),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_564),
.B(n_436),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_564),
.Y(n_762)
);

NOR2xp67_ASAP7_75t_L g763 ( 
.A(n_579),
.B(n_281),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_582),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_625),
.B(n_403),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_543),
.B(n_291),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_586),
.B(n_436),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_543),
.B(n_297),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_543),
.B(n_324),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_577),
.B(n_327),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_586),
.Y(n_771)
);

AND2x2_ASAP7_75t_L g772 ( 
.A(n_625),
.B(n_199),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_588),
.B(n_436),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_577),
.B(n_329),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_588),
.B(n_436),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_641),
.B(n_403),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_577),
.B(n_341),
.Y(n_777)
);

INVxp33_ASAP7_75t_L g778 ( 
.A(n_635),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_589),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_589),
.B(n_436),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_612),
.B(n_199),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_641),
.A2(n_463),
.B1(n_316),
.B2(n_300),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_590),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_590),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_584),
.A2(n_592),
.B1(n_623),
.B2(n_638),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_599),
.Y(n_786)
);

BUFx6f_ASAP7_75t_L g787 ( 
.A(n_577),
.Y(n_787)
);

NOR3xp33_ASAP7_75t_L g788 ( 
.A(n_578),
.B(n_307),
.C(n_321),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_584),
.A2(n_334),
.B1(n_306),
.B2(n_325),
.Y(n_789)
);

NAND2xp33_ASAP7_75t_L g790 ( 
.A(n_577),
.B(n_593),
.Y(n_790)
);

OR2x2_ASAP7_75t_L g791 ( 
.A(n_652),
.B(n_404),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_512),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_593),
.B(n_311),
.Y(n_793)
);

INVx8_ASAP7_75t_L g794 ( 
.A(n_584),
.Y(n_794)
);

BUFx6f_ASAP7_75t_L g795 ( 
.A(n_593),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_600),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_602),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_603),
.B(n_463),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_603),
.B(n_463),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_585),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_608),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_644),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_608),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_594),
.B(n_312),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_613),
.Y(n_805)
);

INVx4_ASAP7_75t_L g806 ( 
.A(n_610),
.Y(n_806)
);

AO221x1_ASAP7_75t_L g807 ( 
.A1(n_605),
.A2(n_332),
.B1(n_331),
.B2(n_317),
.C(n_316),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_616),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_616),
.B(n_463),
.Y(n_809)
);

NOR3xp33_ASAP7_75t_L g810 ( 
.A(n_614),
.B(n_318),
.C(n_315),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_597),
.B(n_214),
.Y(n_811)
);

NOR2x1_ASAP7_75t_L g812 ( 
.A(n_615),
.B(n_495),
.Y(n_812)
);

INVxp67_ASAP7_75t_SL g813 ( 
.A(n_659),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_641),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_622),
.B(n_463),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_622),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_629),
.B(n_463),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_593),
.B(n_214),
.Y(n_818)
);

NOR3xp33_ASAP7_75t_L g819 ( 
.A(n_653),
.B(n_300),
.C(n_296),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_593),
.B(n_214),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_521),
.A2(n_303),
.B(n_317),
.C(n_296),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_724),
.B(n_645),
.Y(n_822)
);

AOI22xp5_ASAP7_75t_L g823 ( 
.A1(n_814),
.A2(n_632),
.B1(n_629),
.B2(n_637),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_772),
.B(n_632),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_672),
.B(n_637),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_731),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_668),
.A2(n_656),
.B(n_523),
.C(n_521),
.Y(n_827)
);

AOI22xp33_ASAP7_75t_L g828 ( 
.A1(n_750),
.A2(n_523),
.B1(n_656),
.B2(n_643),
.Y(n_828)
);

INVx5_ASAP7_75t_L g829 ( 
.A(n_787),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_689),
.A2(n_646),
.B1(n_643),
.B2(n_647),
.Y(n_830)
);

AND2x6_ASAP7_75t_SL g831 ( 
.A(n_668),
.B(n_572),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_731),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_734),
.Y(n_833)
);

BUFx2_ASAP7_75t_L g834 ( 
.A(n_679),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_787),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_734),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_692),
.B(n_646),
.Y(n_837)
);

NOR2xp33_ASAP7_75t_L g838 ( 
.A(n_663),
.B(n_647),
.Y(n_838)
);

AND2x6_ASAP7_75t_L g839 ( 
.A(n_787),
.B(n_644),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_692),
.B(n_644),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_724),
.B(n_645),
.Y(n_841)
);

BUFx12f_ASAP7_75t_L g842 ( 
.A(n_676),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_776),
.B(n_630),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_776),
.B(n_661),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_744),
.Y(n_845)
);

NAND3xp33_ASAP7_75t_SL g846 ( 
.A(n_778),
.B(n_409),
.C(n_404),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_682),
.B(n_686),
.Y(n_847)
);

NAND3xp33_ASAP7_75t_SL g848 ( 
.A(n_800),
.B(n_410),
.C(n_427),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_720),
.B(n_214),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_689),
.A2(n_595),
.B1(n_607),
.B2(n_609),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_764),
.Y(n_851)
);

BUFx3_ASAP7_75t_L g852 ( 
.A(n_714),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_776),
.B(n_709),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_SL g854 ( 
.A1(n_749),
.A2(n_244),
.B1(n_596),
.B2(n_570),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_662),
.B(n_595),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_719),
.B(n_654),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_819),
.A2(n_244),
.B1(n_575),
.B2(n_655),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_718),
.B(n_575),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_764),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_724),
.B(n_645),
.Y(n_860)
);

BUFx3_ASAP7_75t_L g861 ( 
.A(n_714),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_792),
.B(n_575),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_783),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_718),
.A2(n_617),
.B1(n_607),
.B2(n_609),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_783),
.Y(n_865)
);

AOI22xp33_ASAP7_75t_L g866 ( 
.A1(n_807),
.A2(n_244),
.B1(n_655),
.B2(n_639),
.Y(n_866)
);

BUFx2_ASAP7_75t_L g867 ( 
.A(n_667),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_784),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_720),
.B(n_244),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_730),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_784),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_699),
.B(n_587),
.Y(n_872)
);

OR2x2_ASAP7_75t_L g873 ( 
.A(n_791),
.B(n_409),
.Y(n_873)
);

OAI22xp33_ASAP7_75t_L g874 ( 
.A1(n_665),
.A2(n_631),
.B1(n_627),
.B2(n_655),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_724),
.B(n_659),
.Y(n_875)
);

BUFx3_ASAP7_75t_L g876 ( 
.A(n_714),
.Y(n_876)
);

INVx2_ASAP7_75t_SL g877 ( 
.A(n_747),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_803),
.Y(n_878)
);

INVx2_ASAP7_75t_SL g879 ( 
.A(n_765),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_803),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_683),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_805),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_787),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_805),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_SL g885 ( 
.A(n_680),
.B(n_426),
.C(n_424),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_SL g886 ( 
.A(n_795),
.B(n_659),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_790),
.A2(n_596),
.B(n_570),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_788),
.A2(n_627),
.B1(n_591),
.B2(n_639),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_795),
.B(n_659),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_781),
.Y(n_890)
);

INVx4_ASAP7_75t_L g891 ( 
.A(n_795),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_816),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_666),
.B(n_611),
.Y(n_893)
);

AND2x4_ASAP7_75t_SL g894 ( 
.A(n_732),
.B(n_683),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_795),
.B(n_683),
.Y(n_895)
);

INVx1_ASAP7_75t_SL g896 ( 
.A(n_753),
.Y(n_896)
);

NOR3xp33_ASAP7_75t_SL g897 ( 
.A(n_811),
.B(n_499),
.C(n_410),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_702),
.B(n_591),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_683),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_816),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_794),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_687),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_673),
.B(n_618),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_681),
.B(n_659),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_758),
.B(n_591),
.Y(n_905)
);

INVx2_ASAP7_75t_SL g906 ( 
.A(n_760),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_794),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_687),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_SL g909 ( 
.A1(n_811),
.A2(n_412),
.B1(n_427),
.B2(n_426),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_705),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_762),
.B(n_627),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_677),
.B(n_628),
.Y(n_912)
);

AOI22xp5_ASAP7_75t_L g913 ( 
.A1(n_793),
.A2(n_624),
.B1(n_576),
.B2(n_561),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_705),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_677),
.B(n_737),
.Y(n_915)
);

OR2x2_ASAP7_75t_L g916 ( 
.A(n_740),
.B(n_412),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_681),
.B(n_659),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_771),
.B(n_628),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_779),
.B(n_631),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_785),
.A2(n_639),
.B1(n_631),
.B2(n_633),
.Y(n_920)
);

OAI21xp5_ASAP7_75t_L g921 ( 
.A1(n_704),
.A2(n_633),
.B(n_551),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_786),
.B(n_633),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_727),
.B(n_733),
.Y(n_923)
);

AOI22xp33_ASAP7_75t_L g924 ( 
.A1(n_745),
.A2(n_544),
.B1(n_545),
.B2(n_539),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_710),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_676),
.Y(n_926)
);

OR2x6_ASAP7_75t_L g927 ( 
.A(n_794),
.B(n_570),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_738),
.Y(n_928)
);

NOR3xp33_ASAP7_75t_SL g929 ( 
.A(n_739),
.B(n_499),
.C(n_424),
.Y(n_929)
);

AND2x4_ASAP7_75t_SL g930 ( 
.A(n_732),
.B(n_660),
.Y(n_930)
);

AOI21xp33_ASAP7_75t_L g931 ( 
.A1(n_727),
.A2(n_570),
.B(n_596),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_710),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_717),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_796),
.B(n_660),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_797),
.B(n_660),
.Y(n_935)
);

NOR2x2_ASAP7_75t_L g936 ( 
.A(n_732),
.B(n_1),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_738),
.B(n_660),
.Y(n_937)
);

NOR3xp33_ASAP7_75t_SL g938 ( 
.A(n_789),
.B(n_423),
.C(n_420),
.Y(n_938)
);

AND2x2_ASAP7_75t_SL g939 ( 
.A(n_810),
.B(n_547),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_802),
.B(n_660),
.Y(n_940)
);

AOI22xp33_ASAP7_75t_L g941 ( 
.A1(n_777),
.A2(n_545),
.B1(n_544),
.B2(n_539),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_801),
.B(n_660),
.Y(n_942)
);

BUFx4f_ASAP7_75t_L g943 ( 
.A(n_670),
.Y(n_943)
);

INVx2_ASAP7_75t_L g944 ( 
.A(n_717),
.Y(n_944)
);

INVx3_ASAP7_75t_L g945 ( 
.A(n_802),
.Y(n_945)
);

NAND3xp33_ASAP7_75t_SL g946 ( 
.A(n_741),
.B(n_423),
.C(n_420),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_725),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_733),
.B(n_418),
.Y(n_948)
);

AND2x2_ASAP7_75t_SL g949 ( 
.A(n_697),
.B(n_547),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_676),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_808),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_725),
.Y(n_952)
);

BUFx3_ASAP7_75t_L g953 ( 
.A(n_708),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_674),
.B(n_535),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_806),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_685),
.B(n_535),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_726),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_746),
.Y(n_958)
);

A2O1A1Ixp33_ASAP7_75t_L g959 ( 
.A1(n_751),
.A2(n_376),
.B(n_377),
.C(n_384),
.Y(n_959)
);

AOI22xp5_ASAP7_75t_L g960 ( 
.A1(n_818),
.A2(n_569),
.B1(n_624),
.B2(n_621),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_726),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_743),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_712),
.B(n_548),
.Y(n_963)
);

INVx3_ASAP7_75t_L g964 ( 
.A(n_716),
.Y(n_964)
);

CKINVDCx5p33_ASAP7_75t_R g965 ( 
.A(n_746),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_722),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_690),
.B(n_376),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_735),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_L g969 ( 
.A(n_664),
.B(n_548),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_L g970 ( 
.A(n_669),
.B(n_671),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_698),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_806),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_818),
.B(n_548),
.Y(n_973)
);

AOI22xp5_ASAP7_75t_L g974 ( 
.A1(n_820),
.A2(n_601),
.B1(n_624),
.B2(n_621),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_700),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_701),
.Y(n_976)
);

INVxp33_ASAP7_75t_L g977 ( 
.A(n_812),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_703),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_706),
.Y(n_979)
);

NOR2xp33_ASAP7_75t_L g980 ( 
.A(n_820),
.B(n_561),
.Y(n_980)
);

INVx2_ASAP7_75t_SL g981 ( 
.A(n_748),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_691),
.B(n_561),
.Y(n_982)
);

BUFx12f_ASAP7_75t_L g983 ( 
.A(n_670),
.Y(n_983)
);

OR2x2_ASAP7_75t_L g984 ( 
.A(n_804),
.B(n_377),
.Y(n_984)
);

HB1xp67_ASAP7_75t_L g985 ( 
.A(n_707),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_694),
.B(n_561),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_711),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_813),
.B(n_569),
.Y(n_988)
);

AO22x1_ASAP7_75t_L g989 ( 
.A1(n_675),
.A2(n_384),
.B1(n_388),
.B2(n_389),
.Y(n_989)
);

AND2x2_ASAP7_75t_SL g990 ( 
.A(n_678),
.B(n_547),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_728),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_752),
.Y(n_992)
);

NAND2xp33_ASAP7_75t_L g993 ( 
.A(n_761),
.B(n_596),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_763),
.B(n_388),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_695),
.B(n_569),
.Y(n_995)
);

AOI22xp33_ASAP7_75t_L g996 ( 
.A1(n_777),
.A2(n_538),
.B1(n_520),
.B2(n_522),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_756),
.Y(n_997)
);

AND2x4_ASAP7_75t_L g998 ( 
.A(n_821),
.B(n_576),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_696),
.B(n_576),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_715),
.B(n_576),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_867),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_887),
.A2(n_742),
.B(n_723),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_845),
.Y(n_1003)
);

INVx5_ASAP7_75t_L g1004 ( 
.A(n_839),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_836),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_835),
.Y(n_1006)
);

INVxp67_ASAP7_75t_L g1007 ( 
.A(n_877),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_829),
.A2(n_742),
.B(n_723),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_962),
.B(n_713),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_853),
.A2(n_754),
.B1(n_755),
.B2(n_774),
.Y(n_1010)
);

AO21x1_ASAP7_75t_L g1011 ( 
.A1(n_980),
.A2(n_754),
.B(n_769),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_948),
.B(n_757),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_824),
.B(n_759),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_836),
.Y(n_1014)
);

AOI222xp33_ASAP7_75t_L g1015 ( 
.A1(n_849),
.A2(n_869),
.B1(n_885),
.B2(n_848),
.C1(n_846),
.C2(n_834),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_851),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_851),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_838),
.B(n_721),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_890),
.B(n_684),
.Y(n_1019)
);

AND2x2_ASAP7_75t_L g1020 ( 
.A(n_879),
.B(n_684),
.Y(n_1020)
);

BUFx2_ASAP7_75t_L g1021 ( 
.A(n_870),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_951),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_835),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_829),
.A2(n_768),
.B(n_770),
.Y(n_1024)
);

AO32x1_ASAP7_75t_L g1025 ( 
.A1(n_920),
.A2(n_389),
.A3(n_392),
.B1(n_393),
.B2(n_397),
.Y(n_1025)
);

A2O1A1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_837),
.A2(n_766),
.B(n_769),
.C(n_774),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_829),
.A2(n_755),
.B(n_766),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_835),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_847),
.A2(n_729),
.B(n_688),
.C(n_693),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_822),
.A2(n_688),
.B(n_693),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_896),
.B(n_767),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_915),
.A2(n_817),
.B1(n_815),
.B2(n_809),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_847),
.B(n_773),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_977),
.A2(n_985),
.B1(n_906),
.B2(n_842),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_822),
.A2(n_799),
.B(n_798),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_901),
.B(n_736),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_838),
.B(n_775),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_L g1038 ( 
.A(n_916),
.B(n_780),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_981),
.B(n_782),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_SL g1040 ( 
.A(n_943),
.B(n_610),
.Y(n_1040)
);

AOI22xp5_ASAP7_75t_L g1041 ( 
.A1(n_915),
.A2(n_624),
.B1(n_621),
.B2(n_601),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_997),
.B(n_534),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_841),
.A2(n_634),
.B(n_610),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_943),
.B(n_610),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_860),
.A2(n_634),
.B(n_621),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_971),
.B(n_534),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_977),
.B(n_601),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_823),
.B(n_953),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_SL g1049 ( 
.A(n_953),
.B(n_634),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_978),
.B(n_536),
.Y(n_1050)
);

HB1xp67_ASAP7_75t_L g1051 ( 
.A(n_899),
.Y(n_1051)
);

A2O1A1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_979),
.A2(n_601),
.B(n_536),
.C(n_568),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_SL g1053 ( 
.A(n_983),
.B(n_551),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_967),
.B(n_392),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_972),
.A2(n_571),
.B(n_568),
.Y(n_1055)
);

BUFx3_ASAP7_75t_L g1056 ( 
.A(n_842),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_868),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_987),
.B(n_970),
.Y(n_1058)
);

AND2x2_ASAP7_75t_L g1059 ( 
.A(n_873),
.B(n_393),
.Y(n_1059)
);

A2O1A1Ixp33_ASAP7_75t_L g1060 ( 
.A1(n_970),
.A2(n_571),
.B(n_568),
.C(n_565),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_856),
.A2(n_844),
.B(n_912),
.C(n_840),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_868),
.Y(n_1062)
);

INVx2_ASAP7_75t_L g1063 ( 
.A(n_871),
.Y(n_1063)
);

A2O1A1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_856),
.A2(n_565),
.B(n_563),
.C(n_554),
.Y(n_1064)
);

AO21x1_ASAP7_75t_L g1065 ( 
.A1(n_980),
.A2(n_571),
.B(n_565),
.Y(n_1065)
);

HB1xp67_ASAP7_75t_L g1066 ( 
.A(n_899),
.Y(n_1066)
);

AOI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_858),
.A2(n_563),
.B(n_554),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_871),
.Y(n_1068)
);

INVx1_ASAP7_75t_SL g1069 ( 
.A(n_936),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_830),
.B(n_1),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_966),
.B(n_3),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_946),
.B(n_397),
.C(n_554),
.Y(n_1072)
);

NAND2x1p5_ASAP7_75t_L g1073 ( 
.A(n_901),
.B(n_899),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_825),
.B(n_862),
.Y(n_1074)
);

INVxp67_ASAP7_75t_SL g1075 ( 
.A(n_835),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_862),
.B(n_563),
.Y(n_1076)
);

INVx4_ASAP7_75t_L g1077 ( 
.A(n_901),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_R g1078 ( 
.A(n_958),
.B(n_965),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_899),
.Y(n_1079)
);

INVx8_ASAP7_75t_L g1080 ( 
.A(n_839),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_880),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_827),
.A2(n_552),
.B(n_551),
.C(n_10),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_880),
.Y(n_1083)
);

A2O1A1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_912),
.A2(n_3),
.B(n_4),
.C(n_14),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_843),
.A2(n_162),
.B(n_161),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_955),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_900),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_900),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_826),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_910),
.Y(n_1090)
);

AND2x2_ASAP7_75t_L g1091 ( 
.A(n_909),
.B(n_17),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_SL g1092 ( 
.A(n_983),
.B(n_147),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_992),
.B(n_144),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_910),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_975),
.B(n_976),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_897),
.A2(n_23),
.B(n_25),
.C(n_31),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_990),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_1097)
);

AND2x2_ASAP7_75t_L g1098 ( 
.A(n_894),
.B(n_35),
.Y(n_1098)
);

OR2x2_ASAP7_75t_L g1099 ( 
.A(n_984),
.B(n_968),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_975),
.B(n_36),
.Y(n_1100)
);

INVx2_ASAP7_75t_SL g1101 ( 
.A(n_894),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_950),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_SL g1103 ( 
.A(n_968),
.B(n_142),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_990),
.A2(n_37),
.B1(n_38),
.B2(n_41),
.Y(n_1104)
);

NAND3xp33_ASAP7_75t_L g1105 ( 
.A(n_938),
.B(n_38),
.C(n_41),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_901),
.Y(n_1106)
);

NOR2xp33_ASAP7_75t_R g1107 ( 
.A(n_852),
.B(n_140),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_852),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_832),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_964),
.B(n_44),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_976),
.B(n_47),
.Y(n_1111)
);

AOI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_994),
.A2(n_138),
.B1(n_123),
.B2(n_122),
.Y(n_1112)
);

O2A1O1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_827),
.A2(n_959),
.B(n_991),
.C(n_929),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_964),
.B(n_118),
.Y(n_1114)
);

OAI21xp33_ASAP7_75t_SL g1115 ( 
.A1(n_828),
.A2(n_48),
.B(n_50),
.Y(n_1115)
);

INVx2_ASAP7_75t_L g1116 ( 
.A(n_914),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_991),
.B(n_115),
.Y(n_1117)
);

AOI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_828),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_L g1119 ( 
.A1(n_959),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_1119)
);

CKINVDCx20_ASAP7_75t_R g1120 ( 
.A(n_861),
.Y(n_1120)
);

AO21x1_ASAP7_75t_L g1121 ( 
.A1(n_973),
.A2(n_55),
.B(n_56),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_949),
.A2(n_883),
.B1(n_928),
.B2(n_945),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_883),
.Y(n_1123)
);

NOR2xp33_ASAP7_75t_L g1124 ( 
.A(n_831),
.B(n_855),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_833),
.A2(n_55),
.B(n_58),
.C(n_59),
.Y(n_1125)
);

A2O1A1Ixp33_ASAP7_75t_L g1126 ( 
.A1(n_859),
.A2(n_61),
.B(n_62),
.C(n_64),
.Y(n_1126)
);

BUFx2_ASAP7_75t_SL g1127 ( 
.A(n_861),
.Y(n_1127)
);

NOR2xp33_ASAP7_75t_L g1128 ( 
.A(n_855),
.B(n_62),
.Y(n_1128)
);

A2O1A1Ixp33_ASAP7_75t_L g1129 ( 
.A1(n_863),
.A2(n_66),
.B(n_68),
.C(n_69),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_865),
.Y(n_1130)
);

INVxp67_ASAP7_75t_L g1131 ( 
.A(n_855),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_926),
.Y(n_1132)
);

OAI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_949),
.A2(n_88),
.B1(n_78),
.B2(n_81),
.Y(n_1133)
);

OR2x6_ASAP7_75t_L g1134 ( 
.A(n_927),
.B(n_85),
.Y(n_1134)
);

AND2x2_ASAP7_75t_L g1135 ( 
.A(n_930),
.B(n_893),
.Y(n_1135)
);

INVx6_ASAP7_75t_L g1136 ( 
.A(n_876),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_931),
.A2(n_86),
.B(n_90),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_982),
.A2(n_986),
.B(n_969),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_883),
.B(n_91),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_L g1140 ( 
.A(n_893),
.B(n_66),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_955),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_914),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_SL g1143 ( 
.A1(n_930),
.A2(n_97),
.B1(n_98),
.B2(n_876),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_883),
.B(n_893),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_886),
.A2(n_889),
.B(n_904),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_850),
.A2(n_888),
.B(n_921),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_928),
.A2(n_945),
.B1(n_884),
.B2(n_882),
.Y(n_1147)
);

OR2x2_ASAP7_75t_L g1148 ( 
.A(n_878),
.B(n_892),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_904),
.A2(n_917),
.B(n_895),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_891),
.A2(n_1000),
.B1(n_995),
.B2(n_999),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_866),
.A2(n_993),
.B(n_881),
.C(n_888),
.Y(n_1151)
);

BUFx3_ASAP7_75t_L g1152 ( 
.A(n_907),
.Y(n_1152)
);

AO31x2_ASAP7_75t_L g1153 ( 
.A1(n_1065),
.A2(n_1011),
.A3(n_1026),
.B(n_1002),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1058),
.B(n_952),
.Y(n_1154)
);

OAI21xp33_ASAP7_75t_SL g1155 ( 
.A1(n_1097),
.A2(n_1104),
.B(n_1118),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1138),
.A2(n_891),
.B(n_895),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_SL g1157 ( 
.A1(n_1151),
.A2(n_875),
.B(n_917),
.C(n_937),
.Y(n_1157)
);

AO31x2_ASAP7_75t_L g1158 ( 
.A1(n_1061),
.A2(n_934),
.A3(n_942),
.B(n_935),
.Y(n_1158)
);

AOI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1012),
.A2(n_875),
.B(n_988),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1074),
.B(n_944),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_SL g1161 ( 
.A(n_1015),
.B(n_907),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1067),
.A2(n_941),
.B(n_996),
.Y(n_1162)
);

NOR2xp33_ASAP7_75t_L g1163 ( 
.A(n_1009),
.B(n_963),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1014),
.Y(n_1164)
);

AO21x1_ASAP7_75t_L g1165 ( 
.A1(n_1082),
.A2(n_973),
.B(n_998),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1095),
.B(n_944),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1148),
.Y(n_1167)
);

NAND2xp33_ASAP7_75t_L g1168 ( 
.A(n_1018),
.B(n_839),
.Y(n_1168)
);

AOI21x1_ASAP7_75t_SL g1169 ( 
.A1(n_1100),
.A2(n_998),
.B(n_973),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1146),
.A2(n_988),
.B(n_940),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_SL g1171 ( 
.A1(n_1113),
.A2(n_866),
.B(n_922),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_L g1172 ( 
.A(n_1004),
.B(n_839),
.Y(n_1172)
);

OAI21xp5_ASAP7_75t_SL g1173 ( 
.A1(n_1097),
.A2(n_854),
.B(n_857),
.Y(n_1173)
);

BUFx8_ASAP7_75t_L g1174 ( 
.A(n_1021),
.Y(n_1174)
);

OAI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1149),
.A2(n_996),
.B(n_941),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_L g1176 ( 
.A1(n_1145),
.A2(n_919),
.B(n_905),
.Y(n_1176)
);

AND2x4_ASAP7_75t_L g1177 ( 
.A(n_1101),
.B(n_881),
.Y(n_1177)
);

OR2x6_ASAP7_75t_L g1178 ( 
.A(n_1080),
.B(n_927),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1033),
.B(n_932),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1033),
.B(n_932),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1037),
.B(n_1038),
.Y(n_1181)
);

HB1xp67_ASAP7_75t_L g1182 ( 
.A(n_1022),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1008),
.A2(n_988),
.B(n_940),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1059),
.B(n_963),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1010),
.A2(n_864),
.B(n_874),
.Y(n_1185)
);

BUFx8_ASAP7_75t_SL g1186 ( 
.A(n_1003),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_SL g1187 ( 
.A(n_1070),
.B(n_911),
.C(n_872),
.Y(n_1187)
);

INVx2_ASAP7_75t_SL g1188 ( 
.A(n_1001),
.Y(n_1188)
);

NAND2xp33_ASAP7_75t_R g1189 ( 
.A(n_1078),
.B(n_956),
.Y(n_1189)
);

AOI221xp5_ASAP7_75t_L g1190 ( 
.A1(n_1070),
.A2(n_989),
.B1(n_957),
.B2(n_902),
.C(n_961),
.Y(n_1190)
);

AO31x2_ASAP7_75t_L g1191 ( 
.A1(n_1052),
.A2(n_1150),
.A3(n_1024),
.B(n_1027),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1030),
.A2(n_918),
.B(n_898),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1037),
.B(n_952),
.Y(n_1193)
);

HB1xp67_ASAP7_75t_L g1194 ( 
.A(n_1022),
.Y(n_1194)
);

OAI21x1_ASAP7_75t_L g1195 ( 
.A1(n_1043),
.A2(n_913),
.B(n_933),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1007),
.Y(n_1196)
);

NOR2xp67_ASAP7_75t_L g1197 ( 
.A(n_1007),
.B(n_908),
.Y(n_1197)
);

OR2x6_ASAP7_75t_L g1198 ( 
.A(n_1080),
.B(n_927),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_1135),
.B(n_963),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1009),
.A2(n_939),
.B(n_998),
.C(n_960),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1089),
.Y(n_1201)
);

INVx2_ASAP7_75t_L g1202 ( 
.A(n_1057),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1038),
.B(n_933),
.Y(n_1203)
);

BUFx2_ASAP7_75t_L g1204 ( 
.A(n_1120),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_1098),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1013),
.B(n_925),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1076),
.B(n_947),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1104),
.A2(n_924),
.B1(n_974),
.B2(n_939),
.Y(n_1208)
);

AND2x2_ASAP7_75t_L g1209 ( 
.A(n_1124),
.B(n_1099),
.Y(n_1209)
);

AO21x2_ASAP7_75t_L g1210 ( 
.A1(n_1060),
.A2(n_903),
.B(n_954),
.Y(n_1210)
);

O2A1O1Ixp5_ASAP7_75t_L g1211 ( 
.A1(n_1137),
.A2(n_1048),
.B(n_1040),
.C(n_1044),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1118),
.A2(n_924),
.B1(n_903),
.B2(n_956),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1080),
.Y(n_1213)
);

NOR2xp67_ASAP7_75t_L g1214 ( 
.A(n_1077),
.B(n_954),
.Y(n_1214)
);

OAI21x1_ASAP7_75t_L g1215 ( 
.A1(n_1045),
.A2(n_956),
.B(n_1035),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_L g1216 ( 
.A(n_1124),
.B(n_1069),
.Y(n_1216)
);

AOI22xp5_ASAP7_75t_L g1217 ( 
.A1(n_1034),
.A2(n_1092),
.B1(n_1140),
.B2(n_1128),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1062),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1042),
.B(n_1046),
.Y(n_1219)
);

AO31x2_ASAP7_75t_L g1220 ( 
.A1(n_1121),
.A2(n_1064),
.A3(n_1147),
.B(n_1122),
.Y(n_1220)
);

OAI21xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1091),
.A2(n_1143),
.B(n_1112),
.Y(n_1221)
);

AOI221xp5_ASAP7_75t_SL g1222 ( 
.A1(n_1096),
.A2(n_1084),
.B1(n_1115),
.B2(n_1071),
.C(n_1119),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1050),
.B(n_1131),
.Y(n_1223)
);

AOI21xp33_ASAP7_75t_L g1224 ( 
.A1(n_1029),
.A2(n_1111),
.B(n_1110),
.Y(n_1224)
);

OAI22xp5_ASAP7_75t_L g1225 ( 
.A1(n_1004),
.A2(n_1143),
.B1(n_1039),
.B2(n_1131),
.Y(n_1225)
);

AND2x4_ASAP7_75t_L g1226 ( 
.A(n_1108),
.B(n_1152),
.Y(n_1226)
);

O2A1O1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1125),
.A2(n_1129),
.B(n_1126),
.C(n_1031),
.Y(n_1227)
);

NAND3x1_ASAP7_75t_L g1228 ( 
.A(n_1020),
.B(n_1128),
.C(n_1140),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1019),
.A2(n_1085),
.B(n_1047),
.C(n_1105),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_L g1230 ( 
.A1(n_1004),
.A2(n_1109),
.B1(n_1130),
.B2(n_1134),
.Y(n_1230)
);

AO21x1_ASAP7_75t_L g1231 ( 
.A1(n_1093),
.A2(n_1117),
.B(n_1114),
.Y(n_1231)
);

AO31x2_ASAP7_75t_L g1232 ( 
.A1(n_1133),
.A2(n_1025),
.A3(n_1055),
.B(n_1016),
.Y(n_1232)
);

INVx2_ASAP7_75t_SL g1233 ( 
.A(n_1136),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1075),
.A2(n_1144),
.B(n_1049),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1005),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1017),
.B(n_1087),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1063),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1075),
.A2(n_1103),
.B(n_1025),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1068),
.Y(n_1239)
);

AOI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1081),
.A2(n_1088),
.B(n_1083),
.Y(n_1240)
);

INVx4_ASAP7_75t_L g1241 ( 
.A(n_1136),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1025),
.A2(n_1086),
.B(n_1141),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1090),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1094),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1116),
.B(n_1142),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1032),
.A2(n_1139),
.B(n_1053),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1051),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1086),
.A2(n_1141),
.B(n_1041),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_SL g1249 ( 
.A1(n_1132),
.A2(n_1127),
.B1(n_1023),
.B2(n_1028),
.C(n_1006),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1051),
.B(n_1079),
.Y(n_1250)
);

OAI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1072),
.A2(n_1036),
.B(n_1079),
.Y(n_1251)
);

INVxp67_ASAP7_75t_L g1252 ( 
.A(n_1102),
.Y(n_1252)
);

OAI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1072),
.A2(n_1036),
.B(n_1066),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1066),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1006),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1006),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1107),
.B(n_1077),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1073),
.A2(n_1134),
.B(n_1023),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1106),
.B(n_1028),
.Y(n_1259)
);

INVx4_ASAP7_75t_L g1260 ( 
.A(n_1136),
.Y(n_1260)
);

INVx2_ASAP7_75t_SL g1261 ( 
.A(n_1056),
.Y(n_1261)
);

OAI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1123),
.A2(n_1026),
.B(n_1061),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_1123),
.B(n_1058),
.Y(n_1263)
);

O2A1O1Ixp5_ASAP7_75t_L g1264 ( 
.A1(n_1123),
.A2(n_923),
.B(n_1011),
.C(n_1026),
.Y(n_1264)
);

AO31x2_ASAP7_75t_L g1265 ( 
.A1(n_1065),
.A2(n_1011),
.A3(n_1026),
.B(n_1002),
.Y(n_1265)
);

AOI21xp5_ASAP7_75t_L g1266 ( 
.A1(n_1002),
.A2(n_790),
.B(n_724),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1021),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1148),
.Y(n_1268)
);

NAND3xp33_ASAP7_75t_L g1269 ( 
.A(n_1015),
.B(n_567),
.C(n_555),
.Y(n_1269)
);

BUFx3_ASAP7_75t_L g1270 ( 
.A(n_1120),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1054),
.B(n_663),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1014),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1275)
);

O2A1O1Ixp5_ASAP7_75t_L g1276 ( 
.A1(n_1011),
.A2(n_923),
.B(n_1026),
.C(n_1002),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1026),
.A2(n_1061),
.B(n_1010),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1278)
);

INVx5_ASAP7_75t_L g1279 ( 
.A(n_1080),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1065),
.A2(n_1011),
.A3(n_1026),
.B(n_1002),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1004),
.B(n_829),
.Y(n_1281)
);

BUFx3_ASAP7_75t_L g1282 ( 
.A(n_1120),
.Y(n_1282)
);

AOI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1002),
.A2(n_790),
.B(n_724),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1002),
.A2(n_724),
.B(n_790),
.Y(n_1284)
);

AOI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1070),
.A2(n_668),
.B1(n_689),
.B2(n_597),
.C(n_778),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1287)
);

AND2x4_ASAP7_75t_L g1288 ( 
.A(n_1101),
.B(n_852),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1070),
.A2(n_668),
.B1(n_567),
.B2(n_555),
.Y(n_1289)
);

OAI22x1_ASAP7_75t_L g1290 ( 
.A1(n_1070),
.A2(n_668),
.B1(n_750),
.B2(n_516),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1014),
.Y(n_1291)
);

NAND3xp33_ASAP7_75t_L g1292 ( 
.A(n_1015),
.B(n_567),
.C(n_555),
.Y(n_1292)
);

NOR2xp33_ASAP7_75t_L g1293 ( 
.A(n_1058),
.B(n_663),
.Y(n_1293)
);

OR2x2_ASAP7_75t_L g1294 ( 
.A(n_1099),
.B(n_652),
.Y(n_1294)
);

AO21x2_ASAP7_75t_L g1295 ( 
.A1(n_1002),
.A2(n_1011),
.B(n_1146),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1148),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1054),
.B(n_663),
.Y(n_1297)
);

CKINVDCx8_ASAP7_75t_R g1298 ( 
.A(n_1127),
.Y(n_1298)
);

OA21x2_ASAP7_75t_L g1299 ( 
.A1(n_1146),
.A2(n_1065),
.B(n_1026),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_1003),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1058),
.B(n_1074),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1148),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1058),
.B(n_663),
.Y(n_1303)
);

INVx2_ASAP7_75t_SL g1304 ( 
.A(n_1241),
.Y(n_1304)
);

NOR2x1_ASAP7_75t_L g1305 ( 
.A(n_1241),
.B(n_1260),
.Y(n_1305)
);

BUFx2_ASAP7_75t_L g1306 ( 
.A(n_1182),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1196),
.Y(n_1307)
);

HB1xp67_ASAP7_75t_L g1308 ( 
.A(n_1194),
.Y(n_1308)
);

HB1xp67_ASAP7_75t_L g1309 ( 
.A(n_1267),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1201),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1281),
.Y(n_1311)
);

AO21x2_ASAP7_75t_L g1312 ( 
.A1(n_1277),
.A2(n_1224),
.B(n_1185),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1243),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1244),
.Y(n_1314)
);

HB1xp67_ASAP7_75t_L g1315 ( 
.A(n_1188),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1285),
.A2(n_1290),
.B1(n_1289),
.B2(n_1269),
.Y(n_1317)
);

OAI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1292),
.A2(n_1229),
.B(n_1285),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1273),
.A2(n_1275),
.B1(n_1287),
.B2(n_1278),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1186),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1235),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1279),
.B(n_1213),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1208),
.A2(n_1238),
.A3(n_1165),
.B(n_1242),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1250),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1155),
.A2(n_1161),
.B1(n_1209),
.B2(n_1208),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1215),
.A2(n_1169),
.B(n_1195),
.Y(n_1327)
);

AND2x4_ASAP7_75t_L g1328 ( 
.A(n_1199),
.B(n_1279),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1250),
.Y(n_1329)
);

O2A1O1Ixp33_ASAP7_75t_SL g1330 ( 
.A1(n_1173),
.A2(n_1200),
.B(n_1224),
.C(n_1181),
.Y(n_1330)
);

AO21x2_ASAP7_75t_L g1331 ( 
.A1(n_1185),
.A2(n_1262),
.B(n_1295),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1199),
.B(n_1279),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1273),
.B(n_1274),
.Y(n_1333)
);

OAI21x1_ASAP7_75t_L g1334 ( 
.A1(n_1156),
.A2(n_1176),
.B(n_1262),
.Y(n_1334)
);

INVx4_ASAP7_75t_L g1335 ( 
.A(n_1279),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1281),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1192),
.A2(n_1172),
.B(n_1276),
.Y(n_1338)
);

OAI21x1_ASAP7_75t_L g1339 ( 
.A1(n_1183),
.A2(n_1162),
.B(n_1175),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1300),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1274),
.B(n_1275),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1247),
.Y(n_1342)
);

AND2x4_ASAP7_75t_L g1343 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1227),
.A2(n_1231),
.B(n_1251),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_SL g1345 ( 
.A1(n_1251),
.A2(n_1253),
.B(n_1171),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1264),
.A2(n_1170),
.B(n_1248),
.Y(n_1346)
);

AOI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1181),
.A2(n_1286),
.B(n_1287),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1248),
.A2(n_1211),
.B(n_1246),
.Y(n_1348)
);

BUFx8_ASAP7_75t_L g1349 ( 
.A(n_1204),
.Y(n_1349)
);

OA21x2_ASAP7_75t_L g1350 ( 
.A1(n_1222),
.A2(n_1203),
.B(n_1180),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1178),
.B(n_1198),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1278),
.B(n_1286),
.Y(n_1352)
);

INVx6_ASAP7_75t_L g1353 ( 
.A(n_1174),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1258),
.A2(n_1253),
.B(n_1234),
.Y(n_1354)
);

INVx2_ASAP7_75t_SL g1355 ( 
.A(n_1174),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1159),
.A2(n_1299),
.B(n_1230),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1164),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1202),
.Y(n_1358)
);

OA21x2_ASAP7_75t_L g1359 ( 
.A1(n_1203),
.A2(n_1180),
.B(n_1179),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1179),
.A2(n_1193),
.B(n_1207),
.Y(n_1360)
);

OAI21x1_ASAP7_75t_L g1361 ( 
.A1(n_1193),
.A2(n_1207),
.B(n_1225),
.Y(n_1361)
);

OAI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1187),
.A2(n_1301),
.B(n_1228),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1212),
.A2(n_1301),
.B(n_1163),
.Y(n_1363)
);

OAI21x1_ASAP7_75t_L g1364 ( 
.A1(n_1166),
.A2(n_1160),
.B(n_1236),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1218),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1237),
.Y(n_1366)
);

OAI21xp5_ASAP7_75t_L g1367 ( 
.A1(n_1271),
.A2(n_1297),
.B(n_1221),
.Y(n_1367)
);

INVx2_ASAP7_75t_SL g1368 ( 
.A(n_1270),
.Y(n_1368)
);

INVx2_ASAP7_75t_SL g1369 ( 
.A(n_1282),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1239),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1272),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1167),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1184),
.B(n_1206),
.Y(n_1373)
);

OAI22xp5_ASAP7_75t_L g1374 ( 
.A1(n_1217),
.A2(n_1197),
.B1(n_1294),
.B2(n_1206),
.Y(n_1374)
);

OAI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1166),
.A2(n_1160),
.B(n_1236),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1205),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1216),
.A2(n_1168),
.B1(n_1190),
.B2(n_1295),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_1291),
.Y(n_1378)
);

AO32x2_ASAP7_75t_L g1379 ( 
.A1(n_1212),
.A2(n_1153),
.A3(n_1280),
.B1(n_1265),
.B2(n_1220),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1219),
.A2(n_1154),
.B(n_1263),
.Y(n_1380)
);

OAI21xp5_ASAP7_75t_L g1381 ( 
.A1(n_1219),
.A2(n_1190),
.B(n_1223),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1154),
.A2(n_1263),
.B(n_1245),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1223),
.B(n_1254),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1157),
.A2(n_1257),
.B(n_1296),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1245),
.A2(n_1256),
.B(n_1259),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1268),
.B(n_1302),
.Y(n_1386)
);

O2A1O1Ixp33_ASAP7_75t_SL g1387 ( 
.A1(n_1255),
.A2(n_1256),
.B(n_1249),
.C(n_1233),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1214),
.A2(n_1177),
.B(n_1288),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_L g1389 ( 
.A1(n_1191),
.A2(n_1153),
.B(n_1265),
.Y(n_1389)
);

INVx8_ASAP7_75t_L g1390 ( 
.A(n_1226),
.Y(n_1390)
);

AO21x2_ASAP7_75t_L g1391 ( 
.A1(n_1210),
.A2(n_1153),
.B(n_1265),
.Y(n_1391)
);

OAI22x1_ASAP7_75t_L g1392 ( 
.A1(n_1177),
.A2(n_1252),
.B1(n_1288),
.B2(n_1261),
.Y(n_1392)
);

AO31x2_ASAP7_75t_L g1393 ( 
.A1(n_1280),
.A2(n_1191),
.A3(n_1158),
.B(n_1232),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1158),
.B(n_1220),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1191),
.A2(n_1280),
.B(n_1158),
.Y(n_1395)
);

AO21x2_ASAP7_75t_L g1396 ( 
.A1(n_1232),
.A2(n_1277),
.B(n_1224),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1232),
.A2(n_1277),
.B(n_1276),
.Y(n_1397)
);

AOI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1189),
.A2(n_1285),
.B1(n_1290),
.B2(n_1289),
.Y(n_1398)
);

AOI21x1_ASAP7_75t_L g1399 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1240),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1401)
);

OAI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1289),
.A2(n_1292),
.B(n_1269),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1196),
.Y(n_1403)
);

BUFx2_ASAP7_75t_L g1404 ( 
.A(n_1182),
.Y(n_1404)
);

INVxp67_ASAP7_75t_SL g1405 ( 
.A(n_1182),
.Y(n_1405)
);

OAI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1155),
.A2(n_1289),
.B(n_1173),
.C(n_668),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1201),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1181),
.B(n_1299),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1410)
);

OA21x2_ASAP7_75t_L g1411 ( 
.A1(n_1277),
.A2(n_1276),
.B(n_1224),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1412)
);

CKINVDCx8_ASAP7_75t_R g1413 ( 
.A(n_1300),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1293),
.B(n_1303),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1277),
.A2(n_790),
.B(n_724),
.Y(n_1415)
);

INVx1_ASAP7_75t_SL g1416 ( 
.A(n_1267),
.Y(n_1416)
);

OA21x2_ASAP7_75t_L g1417 ( 
.A1(n_1277),
.A2(n_1276),
.B(n_1224),
.Y(n_1417)
);

AOI222xp33_ASAP7_75t_SL g1418 ( 
.A1(n_1289),
.A2(n_537),
.B1(n_483),
.B2(n_468),
.C1(n_443),
.C2(n_445),
.Y(n_1418)
);

INVx2_ASAP7_75t_L g1419 ( 
.A(n_1240),
.Y(n_1419)
);

AO21x2_ASAP7_75t_L g1420 ( 
.A1(n_1277),
.A2(n_1224),
.B(n_1185),
.Y(n_1420)
);

AO21x2_ASAP7_75t_L g1421 ( 
.A1(n_1277),
.A2(n_1224),
.B(n_1185),
.Y(n_1421)
);

BUFx12f_ASAP7_75t_L g1422 ( 
.A(n_1300),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1289),
.A2(n_1292),
.B(n_1269),
.Y(n_1423)
);

BUFx8_ASAP7_75t_L g1424 ( 
.A(n_1204),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1289),
.A2(n_1292),
.B(n_1269),
.Y(n_1425)
);

OR2x6_ASAP7_75t_SL g1426 ( 
.A(n_1269),
.B(n_1292),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1201),
.Y(n_1427)
);

HB1xp67_ASAP7_75t_L g1428 ( 
.A(n_1196),
.Y(n_1428)
);

OAI21x1_ASAP7_75t_L g1429 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1429)
);

INVx5_ASAP7_75t_L g1430 ( 
.A(n_1178),
.Y(n_1430)
);

NOR2x1_ASAP7_75t_R g1431 ( 
.A(n_1300),
.B(n_558),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1182),
.Y(n_1433)
);

NOR2xp67_ASAP7_75t_SL g1434 ( 
.A(n_1298),
.B(n_744),
.Y(n_1434)
);

NOR2xp67_ASAP7_75t_L g1435 ( 
.A(n_1188),
.B(n_877),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1201),
.Y(n_1436)
);

OAI211xp5_ASAP7_75t_L g1437 ( 
.A1(n_1289),
.A2(n_668),
.B(n_1285),
.C(n_1269),
.Y(n_1437)
);

INVx2_ASAP7_75t_SL g1438 ( 
.A(n_1241),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1285),
.A2(n_1290),
.B1(n_1289),
.B2(n_1269),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1266),
.A2(n_1283),
.B(n_1284),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1201),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1325),
.Y(n_1442)
);

O2A1O1Ixp33_ASAP7_75t_L g1443 ( 
.A1(n_1437),
.A2(n_1407),
.B(n_1425),
.C(n_1423),
.Y(n_1443)
);

O2A1O1Ixp5_ASAP7_75t_L g1444 ( 
.A1(n_1318),
.A2(n_1402),
.B(n_1407),
.C(n_1362),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1415),
.A2(n_1319),
.B(n_1431),
.Y(n_1446)
);

AND2x4_ASAP7_75t_L g1447 ( 
.A(n_1336),
.B(n_1343),
.Y(n_1447)
);

OR2x2_ASAP7_75t_L g1448 ( 
.A(n_1325),
.B(n_1329),
.Y(n_1448)
);

O2A1O1Ixp33_ASAP7_75t_L g1449 ( 
.A1(n_1316),
.A2(n_1401),
.B(n_1414),
.C(n_1412),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_L g1450 ( 
.A(n_1352),
.B(n_1347),
.Y(n_1450)
);

OAI22xp5_ASAP7_75t_L g1451 ( 
.A1(n_1317),
.A2(n_1439),
.B1(n_1398),
.B2(n_1426),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1329),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_L g1453 ( 
.A1(n_1374),
.A2(n_1330),
.B(n_1367),
.C(n_1344),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1400),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1390),
.Y(n_1455)
);

INVxp67_ASAP7_75t_L g1456 ( 
.A(n_1342),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1336),
.B(n_1343),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1426),
.A2(n_1326),
.B1(n_1377),
.B2(n_1376),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1373),
.A2(n_1416),
.B1(n_1403),
.B2(n_1428),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1383),
.B(n_1372),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_SL g1461 ( 
.A1(n_1381),
.A2(n_1335),
.B(n_1351),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1310),
.Y(n_1462)
);

AOI211xp5_ASAP7_75t_L g1463 ( 
.A1(n_1330),
.A2(n_1363),
.B(n_1384),
.C(n_1418),
.Y(n_1463)
);

AOI21xp5_ASAP7_75t_SL g1464 ( 
.A1(n_1335),
.A2(n_1351),
.B(n_1343),
.Y(n_1464)
);

BUFx6f_ASAP7_75t_L g1465 ( 
.A(n_1390),
.Y(n_1465)
);

NOR2xp67_ASAP7_75t_L g1466 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1466)
);

O2A1O1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1345),
.A2(n_1315),
.B(n_1307),
.C(n_1308),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1312),
.A2(n_1420),
.B(n_1421),
.C(n_1309),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1408),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1394),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_SL g1471 ( 
.A1(n_1321),
.A2(n_1353),
.B1(n_1340),
.B2(n_1413),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1427),
.Y(n_1472)
);

AND2x4_ASAP7_75t_L g1473 ( 
.A(n_1351),
.B(n_1328),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1383),
.B(n_1368),
.Y(n_1474)
);

OR2x2_ASAP7_75t_L g1475 ( 
.A(n_1306),
.B(n_1404),
.Y(n_1475)
);

OAI22xp5_ASAP7_75t_L g1476 ( 
.A1(n_1435),
.A2(n_1405),
.B1(n_1363),
.B2(n_1306),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1404),
.B(n_1433),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1386),
.B(n_1433),
.Y(n_1478)
);

A2O1A1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1338),
.A2(n_1346),
.B(n_1348),
.C(n_1361),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1357),
.B(n_1358),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1436),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1441),
.Y(n_1482)
);

AND2x2_ASAP7_75t_L g1483 ( 
.A(n_1365),
.B(n_1366),
.Y(n_1483)
);

AOI21xp5_ASAP7_75t_SL g1484 ( 
.A1(n_1335),
.A2(n_1332),
.B(n_1328),
.Y(n_1484)
);

AND2x2_ASAP7_75t_L g1485 ( 
.A(n_1370),
.B(n_1371),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1321),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1378),
.B(n_1380),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1342),
.B(n_1313),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_1340),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_SL g1490 ( 
.A1(n_1332),
.A2(n_1304),
.B(n_1438),
.Y(n_1490)
);

NOR2x1_ASAP7_75t_SL g1491 ( 
.A(n_1430),
.B(n_1331),
.Y(n_1491)
);

O2A1O1Ixp5_ASAP7_75t_L g1492 ( 
.A1(n_1409),
.A2(n_1388),
.B(n_1419),
.C(n_1399),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1422),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1380),
.B(n_1314),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1392),
.B(n_1322),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1392),
.B(n_1304),
.Y(n_1496)
);

AND2x4_ASAP7_75t_L g1497 ( 
.A(n_1430),
.B(n_1337),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1409),
.B(n_1382),
.Y(n_1498)
);

OAI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1353),
.A2(n_1413),
.B1(n_1355),
.B2(n_1438),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1430),
.B(n_1337),
.Y(n_1500)
);

A2O1A1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1346),
.A2(n_1361),
.B(n_1356),
.C(n_1375),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_L g1502 ( 
.A(n_1312),
.B(n_1420),
.Y(n_1502)
);

INVx5_ASAP7_75t_L g1503 ( 
.A(n_1430),
.Y(n_1503)
);

INVxp67_ASAP7_75t_L g1504 ( 
.A(n_1385),
.Y(n_1504)
);

AOI21x1_ASAP7_75t_SL g1505 ( 
.A1(n_1387),
.A2(n_1434),
.B(n_1353),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_L g1506 ( 
.A(n_1360),
.B(n_1359),
.Y(n_1506)
);

AOI221x1_ASAP7_75t_SL g1507 ( 
.A1(n_1411),
.A2(n_1417),
.B1(n_1353),
.B2(n_1331),
.C(n_1379),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1422),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_L g1509 ( 
.A(n_1360),
.B(n_1359),
.Y(n_1509)
);

AND2x4_ASAP7_75t_L g1510 ( 
.A(n_1430),
.B(n_1311),
.Y(n_1510)
);

OAI22xp5_ASAP7_75t_L g1511 ( 
.A1(n_1355),
.A2(n_1305),
.B1(n_1390),
.B2(n_1417),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1391),
.Y(n_1512)
);

OA22x2_ASAP7_75t_L g1513 ( 
.A1(n_1311),
.A2(n_1337),
.B1(n_1354),
.B2(n_1375),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1364),
.B(n_1350),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1364),
.B(n_1350),
.Y(n_1515)
);

OA21x2_ASAP7_75t_L g1516 ( 
.A1(n_1320),
.A2(n_1440),
.B(n_1432),
.Y(n_1516)
);

BUFx4_ASAP7_75t_R g1517 ( 
.A(n_1349),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_R g1518 ( 
.A(n_1349),
.B(n_1424),
.Y(n_1518)
);

OA21x2_ASAP7_75t_L g1519 ( 
.A1(n_1406),
.A2(n_1429),
.B(n_1410),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1311),
.B(n_1331),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1356),
.A2(n_1334),
.B(n_1395),
.C(n_1389),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1349),
.B(n_1424),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1411),
.B(n_1323),
.Y(n_1523)
);

OAI22xp5_ASAP7_75t_SL g1524 ( 
.A1(n_1397),
.A2(n_1324),
.B1(n_1379),
.B2(n_1396),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1334),
.A2(n_1395),
.B(n_1389),
.C(n_1339),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1393),
.B(n_1324),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1324),
.B(n_1397),
.Y(n_1527)
);

OAI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1324),
.A2(n_1379),
.B1(n_1393),
.B2(n_1327),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_R g1529 ( 
.A(n_1324),
.B(n_1393),
.Y(n_1529)
);

O2A1O1Ixp33_ASAP7_75t_L g1530 ( 
.A1(n_1437),
.A2(n_668),
.B(n_1407),
.C(n_1402),
.Y(n_1530)
);

O2A1O1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1437),
.A2(n_668),
.B(n_1407),
.C(n_1402),
.Y(n_1531)
);

OAI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1316),
.A2(n_1289),
.B1(n_1285),
.B2(n_1401),
.Y(n_1532)
);

CKINVDCx8_ASAP7_75t_R g1533 ( 
.A(n_1390),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1316),
.A2(n_1289),
.B1(n_1285),
.B2(n_1401),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1328),
.Y(n_1535)
);

O2A1O1Ixp33_ASAP7_75t_L g1536 ( 
.A1(n_1437),
.A2(n_668),
.B(n_1407),
.C(n_1402),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1316),
.A2(n_1289),
.B1(n_1285),
.B2(n_1401),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1333),
.B(n_1341),
.Y(n_1539)
);

AOI21xp5_ASAP7_75t_SL g1540 ( 
.A1(n_1407),
.A2(n_746),
.B(n_1208),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1520),
.B(n_1470),
.Y(n_1541)
);

INVxp67_ASAP7_75t_L g1542 ( 
.A(n_1477),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1494),
.Y(n_1543)
);

HB1xp67_ASAP7_75t_L g1544 ( 
.A(n_1456),
.Y(n_1544)
);

AOI211xp5_ASAP7_75t_L g1545 ( 
.A1(n_1451),
.A2(n_1534),
.B(n_1537),
.C(n_1532),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1454),
.Y(n_1546)
);

NAND2xp5_ASAP7_75t_L g1547 ( 
.A(n_1445),
.B(n_1538),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1486),
.Y(n_1548)
);

HB1xp67_ASAP7_75t_L g1549 ( 
.A(n_1456),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1539),
.B(n_1450),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1478),
.B(n_1460),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1448),
.Y(n_1552)
);

OR2x2_ASAP7_75t_L g1553 ( 
.A(n_1526),
.B(n_1502),
.Y(n_1553)
);

INVxp67_ASAP7_75t_SL g1554 ( 
.A(n_1487),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1523),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1449),
.B(n_1474),
.Y(n_1556)
);

OA21x2_ASAP7_75t_L g1557 ( 
.A1(n_1479),
.A2(n_1501),
.B(n_1521),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1495),
.B(n_1442),
.Y(n_1558)
);

AO21x2_ASAP7_75t_L g1559 ( 
.A1(n_1525),
.A2(n_1501),
.B(n_1529),
.Y(n_1559)
);

OR2x6_ASAP7_75t_L g1560 ( 
.A(n_1461),
.B(n_1464),
.Y(n_1560)
);

OR2x6_ASAP7_75t_L g1561 ( 
.A(n_1540),
.B(n_1468),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1488),
.B(n_1475),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_L g1563 ( 
.A(n_1452),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1443),
.B(n_1459),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1458),
.A2(n_1476),
.B1(n_1457),
.B2(n_1447),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1462),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1469),
.B(n_1472),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1489),
.B(n_1486),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1447),
.A2(n_1457),
.B1(n_1473),
.B2(n_1496),
.Y(n_1569)
);

OR2x6_ASAP7_75t_L g1570 ( 
.A(n_1446),
.B(n_1484),
.Y(n_1570)
);

NAND2xp5_ASAP7_75t_L g1571 ( 
.A(n_1483),
.B(n_1485),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1481),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1482),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1511),
.Y(n_1574)
);

NAND2xp5_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1536),
.Y(n_1575)
);

OR2x2_ASAP7_75t_L g1576 ( 
.A(n_1506),
.B(n_1509),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1527),
.A2(n_1515),
.B(n_1514),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1531),
.B(n_1480),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1453),
.B(n_1463),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1512),
.Y(n_1580)
);

OAI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1444),
.A2(n_1467),
.B(n_1492),
.Y(n_1581)
);

INVx3_ASAP7_75t_L g1582 ( 
.A(n_1497),
.Y(n_1582)
);

INVx2_ASAP7_75t_SL g1583 ( 
.A(n_1503),
.Y(n_1583)
);

NAND2x1p5_ASAP7_75t_L g1584 ( 
.A(n_1497),
.B(n_1510),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1513),
.B(n_1491),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1504),
.B(n_1500),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1504),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1528),
.B(n_1524),
.Y(n_1588)
);

NAND4xp25_ASAP7_75t_L g1589 ( 
.A(n_1466),
.B(n_1507),
.C(n_1499),
.D(n_1522),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1516),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1546),
.Y(n_1591)
);

INVx4_ASAP7_75t_L g1592 ( 
.A(n_1560),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1546),
.Y(n_1593)
);

OAI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1579),
.A2(n_1533),
.B1(n_1508),
.B2(n_1493),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1590),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1585),
.B(n_1519),
.Y(n_1596)
);

INVx2_ASAP7_75t_SL g1597 ( 
.A(n_1586),
.Y(n_1597)
);

OR2x2_ASAP7_75t_L g1598 ( 
.A(n_1576),
.B(n_1519),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1543),
.B(n_1554),
.Y(n_1599)
);

AOI22xp33_ASAP7_75t_L g1600 ( 
.A1(n_1575),
.A2(n_1471),
.B1(n_1518),
.B2(n_1473),
.Y(n_1600)
);

AOI221xp5_ASAP7_75t_L g1601 ( 
.A1(n_1545),
.A2(n_1518),
.B1(n_1508),
.B2(n_1493),
.C(n_1490),
.Y(n_1601)
);

BUFx2_ASAP7_75t_L g1602 ( 
.A(n_1586),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

OAI21xp5_ASAP7_75t_SL g1604 ( 
.A1(n_1564),
.A2(n_1565),
.B(n_1581),
.Y(n_1604)
);

HB1xp67_ASAP7_75t_L g1605 ( 
.A(n_1580),
.Y(n_1605)
);

AO22x1_ASAP7_75t_L g1606 ( 
.A1(n_1574),
.A2(n_1517),
.B1(n_1535),
.B2(n_1465),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1577),
.B(n_1535),
.Y(n_1607)
);

OR2x2_ASAP7_75t_L g1608 ( 
.A(n_1553),
.B(n_1455),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1551),
.B(n_1455),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1560),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1557),
.B(n_1465),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1557),
.B(n_1559),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1609),
.Y(n_1613)
);

INVx2_ASAP7_75t_L g1614 ( 
.A(n_1595),
.Y(n_1614)
);

INVxp67_ASAP7_75t_SL g1615 ( 
.A(n_1599),
.Y(n_1615)
);

OR2x2_ASAP7_75t_L g1616 ( 
.A(n_1598),
.B(n_1552),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1602),
.B(n_1596),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1603),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1603),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1598),
.B(n_1552),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_SL g1621 ( 
.A(n_1601),
.B(n_1556),
.Y(n_1621)
);

AO22x1_ASAP7_75t_L g1622 ( 
.A1(n_1612),
.A2(n_1548),
.B1(n_1568),
.B2(n_1550),
.Y(n_1622)
);

AND2x2_ASAP7_75t_SL g1623 ( 
.A(n_1612),
.B(n_1588),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1602),
.B(n_1555),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1599),
.B(n_1542),
.Y(n_1625)
);

AND2x4_ASAP7_75t_SL g1626 ( 
.A(n_1592),
.B(n_1560),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1609),
.B(n_1562),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1605),
.Y(n_1628)
);

OAI221xp5_ASAP7_75t_L g1629 ( 
.A1(n_1604),
.A2(n_1578),
.B1(n_1589),
.B2(n_1570),
.C(n_1561),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1602),
.B(n_1555),
.Y(n_1630)
);

AOI33xp33_ASAP7_75t_L g1631 ( 
.A1(n_1612),
.A2(n_1558),
.A3(n_1572),
.B1(n_1566),
.B2(n_1573),
.B3(n_1567),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1591),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1591),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1601),
.A2(n_1570),
.B1(n_1561),
.B2(n_1560),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1591),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1596),
.B(n_1541),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1604),
.A2(n_1547),
.B1(n_1588),
.B2(n_1544),
.C(n_1549),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1593),
.Y(n_1638)
);

BUFx10_ASAP7_75t_L g1639 ( 
.A(n_1593),
.Y(n_1639)
);

NOR2xp33_ASAP7_75t_SL g1640 ( 
.A(n_1592),
.B(n_1570),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1607),
.Y(n_1641)
);

NAND4xp75_ASAP7_75t_L g1642 ( 
.A(n_1612),
.B(n_1517),
.C(n_1557),
.D(n_1583),
.Y(n_1642)
);

AOI33xp33_ASAP7_75t_L g1643 ( 
.A1(n_1600),
.A2(n_1558),
.A3(n_1573),
.B1(n_1572),
.B2(n_1566),
.B3(n_1567),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1597),
.B(n_1586),
.Y(n_1644)
);

OAI211xp5_ASAP7_75t_SL g1645 ( 
.A1(n_1600),
.A2(n_1569),
.B(n_1571),
.C(n_1587),
.Y(n_1645)
);

OAI211xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1594),
.A2(n_1587),
.B(n_1563),
.C(n_1582),
.Y(n_1646)
);

NAND2xp5_ASAP7_75t_L g1647 ( 
.A(n_1615),
.B(n_1608),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1632),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1632),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1633),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1613),
.B(n_1608),
.Y(n_1651)
);

BUFx3_ASAP7_75t_L g1652 ( 
.A(n_1639),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1633),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1635),
.Y(n_1654)
);

INVxp67_ASAP7_75t_L g1655 ( 
.A(n_1621),
.Y(n_1655)
);

INVx1_ASAP7_75t_SL g1656 ( 
.A(n_1627),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1635),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1628),
.Y(n_1658)
);

AND2x4_ASAP7_75t_L g1659 ( 
.A(n_1644),
.B(n_1597),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1614),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1625),
.Y(n_1661)
);

AOI21xp33_ASAP7_75t_L g1662 ( 
.A1(n_1629),
.A2(n_1594),
.B(n_1561),
.Y(n_1662)
);

AND4x1_ASAP7_75t_L g1663 ( 
.A(n_1637),
.B(n_1611),
.C(n_1606),
.D(n_1505),
.Y(n_1663)
);

AND2x4_ASAP7_75t_L g1664 ( 
.A(n_1644),
.B(n_1597),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1643),
.B(n_1570),
.C(n_1561),
.Y(n_1665)
);

INVx2_ASAP7_75t_SL g1666 ( 
.A(n_1639),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1623),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1638),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1638),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1617),
.B(n_1596),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_SL g1671 ( 
.A1(n_1634),
.A2(n_1611),
.B(n_1584),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1623),
.A2(n_1570),
.B(n_1560),
.Y(n_1672)
);

INVx4_ASAP7_75t_L g1673 ( 
.A(n_1626),
.Y(n_1673)
);

AND2x6_ASAP7_75t_SL g1674 ( 
.A(n_1644),
.B(n_1548),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_SL g1675 ( 
.A1(n_1642),
.A2(n_1610),
.B(n_1561),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1667),
.B(n_1623),
.Y(n_1676)
);

OR2x2_ASAP7_75t_L g1677 ( 
.A(n_1647),
.B(n_1616),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1660),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1659),
.B(n_1624),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1656),
.B(n_1618),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1658),
.B(n_1620),
.Y(n_1681)
);

AND3x2_ASAP7_75t_L g1682 ( 
.A(n_1655),
.B(n_1640),
.C(n_1630),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1661),
.B(n_1618),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1648),
.B(n_1619),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1663),
.B(n_1622),
.C(n_1646),
.Y(n_1685)
);

NOR3xp33_ASAP7_75t_SL g1686 ( 
.A(n_1671),
.B(n_1642),
.C(n_1645),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1659),
.B(n_1624),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1660),
.Y(n_1688)
);

AND2x4_ASAP7_75t_SL g1689 ( 
.A(n_1673),
.B(n_1592),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1659),
.B(n_1630),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1649),
.Y(n_1691)
);

AND2x2_ASAP7_75t_L g1692 ( 
.A(n_1659),
.B(n_1636),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1664),
.B(n_1636),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1650),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1664),
.B(n_1644),
.Y(n_1695)
);

BUFx3_ASAP7_75t_L g1696 ( 
.A(n_1652),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1670),
.B(n_1641),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1653),
.B(n_1631),
.Y(n_1698)
);

OR2x6_ASAP7_75t_L g1699 ( 
.A(n_1675),
.B(n_1606),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1662),
.B(n_1622),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1653),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1654),
.B(n_1657),
.Y(n_1702)
);

CKINVDCx8_ASAP7_75t_R g1703 ( 
.A(n_1674),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1654),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1657),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1668),
.Y(n_1706)
);

AND3x2_ASAP7_75t_L g1707 ( 
.A(n_1675),
.B(n_1640),
.C(n_1611),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1668),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1706),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1698),
.B(n_1665),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1673),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1676),
.B(n_1673),
.Y(n_1712)
);

AOI21xp33_ASAP7_75t_SL g1713 ( 
.A1(n_1685),
.A2(n_1665),
.B(n_1606),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1698),
.B(n_1663),
.Y(n_1714)
);

NAND2x1p5_ASAP7_75t_L g1715 ( 
.A(n_1696),
.B(n_1673),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1692),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1681),
.B(n_1651),
.Y(n_1717)
);

HB1xp67_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1678),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1691),
.Y(n_1720)
);

AOI322xp5_ASAP7_75t_L g1721 ( 
.A1(n_1686),
.A2(n_1700),
.A3(n_1703),
.B1(n_1683),
.B2(n_1680),
.C1(n_1685),
.C2(n_1697),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1679),
.B(n_1687),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1679),
.B(n_1652),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1692),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1691),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1703),
.B(n_1674),
.Y(n_1726)
);

INVxp67_ASAP7_75t_L g1727 ( 
.A(n_1696),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1694),
.Y(n_1728)
);

HB1xp67_ASAP7_75t_L g1729 ( 
.A(n_1680),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1689),
.B(n_1652),
.Y(n_1730)
);

INVx1_ASAP7_75t_SL g1731 ( 
.A(n_1689),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1703),
.B(n_1669),
.Y(n_1732)
);

OR2x6_ASAP7_75t_L g1733 ( 
.A(n_1699),
.B(n_1672),
.Y(n_1733)
);

BUFx2_ASAP7_75t_L g1734 ( 
.A(n_1699),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1687),
.B(n_1666),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1694),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1701),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1690),
.B(n_1666),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1686),
.B(n_1669),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1677),
.B(n_1684),
.Y(n_1740)
);

OAI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1699),
.A2(n_1610),
.B1(n_1592),
.B2(n_1689),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1701),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1704),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1720),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1720),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1722),
.B(n_1699),
.Y(n_1746)
);

INVx1_ASAP7_75t_SL g1747 ( 
.A(n_1734),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1722),
.B(n_1699),
.Y(n_1748)
);

BUFx3_ASAP7_75t_L g1749 ( 
.A(n_1715),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1725),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1726),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1721),
.B(n_1696),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1730),
.B(n_1704),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1743),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1743),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1711),
.B(n_1690),
.Y(n_1756)
);

BUFx3_ASAP7_75t_L g1757 ( 
.A(n_1715),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1721),
.B(n_1693),
.Y(n_1758)
);

CKINVDCx16_ASAP7_75t_R g1759 ( 
.A(n_1734),
.Y(n_1759)
);

OAI22xp5_ASAP7_75t_L g1760 ( 
.A1(n_1714),
.A2(n_1693),
.B1(n_1677),
.B2(n_1697),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1739),
.A2(n_1682),
.B1(n_1707),
.B2(n_1592),
.Y(n_1761)
);

INVx2_ASAP7_75t_L g1762 ( 
.A(n_1719),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1715),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1727),
.B(n_1695),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1725),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1718),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1728),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1717),
.B(n_1702),
.Y(n_1768)
);

INVx1_ASAP7_75t_SL g1769 ( 
.A(n_1731),
.Y(n_1769)
);

OAI21xp33_ASAP7_75t_L g1770 ( 
.A1(n_1752),
.A2(n_1710),
.B(n_1713),
.Y(n_1770)
);

OAI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1758),
.A2(n_1713),
.B1(n_1710),
.B2(n_1733),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1751),
.A2(n_1732),
.B(n_1733),
.Y(n_1772)
);

AOI32xp33_ASAP7_75t_L g1773 ( 
.A1(n_1761),
.A2(n_1712),
.A3(n_1711),
.B1(n_1741),
.B2(n_1723),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1744),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_L g1775 ( 
.A(n_1759),
.B(n_1729),
.Y(n_1775)
);

OAI22xp5_ASAP7_75t_L g1776 ( 
.A1(n_1759),
.A2(n_1747),
.B1(n_1733),
.B2(n_1766),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1756),
.B(n_1712),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_L g1778 ( 
.A1(n_1747),
.A2(n_1733),
.B1(n_1709),
.B2(n_1724),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1744),
.Y(n_1779)
);

INVx3_ASAP7_75t_SL g1780 ( 
.A(n_1769),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1753),
.Y(n_1781)
);

OR2x2_ASAP7_75t_L g1782 ( 
.A(n_1769),
.B(n_1717),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1756),
.B(n_1746),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1749),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1749),
.Y(n_1785)
);

OAI31xp33_ASAP7_75t_L g1786 ( 
.A1(n_1760),
.A2(n_1730),
.A3(n_1723),
.B(n_1709),
.Y(n_1786)
);

NOR2x1p5_ASAP7_75t_L g1787 ( 
.A(n_1749),
.B(n_1716),
.Y(n_1787)
);

OAI21xp33_ASAP7_75t_L g1788 ( 
.A1(n_1764),
.A2(n_1716),
.B(n_1724),
.Y(n_1788)
);

AOI211xp5_ASAP7_75t_L g1789 ( 
.A1(n_1746),
.A2(n_1730),
.B(n_1740),
.C(n_1728),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1770),
.A2(n_1748),
.B1(n_1733),
.B2(n_1763),
.Y(n_1790)
);

INVxp33_ASAP7_75t_L g1791 ( 
.A(n_1782),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1781),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1780),
.B(n_1748),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1774),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1785),
.B(n_1753),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1784),
.B(n_1753),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_SL g1797 ( 
.A(n_1771),
.B(n_1763),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1779),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1777),
.B(n_1757),
.Y(n_1799)
);

INVx1_ASAP7_75t_SL g1800 ( 
.A(n_1783),
.Y(n_1800)
);

INVxp67_ASAP7_75t_L g1801 ( 
.A(n_1775),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1787),
.B(n_1757),
.Y(n_1802)
);

AOI21xp33_ASAP7_75t_L g1803 ( 
.A1(n_1791),
.A2(n_1771),
.B(n_1776),
.Y(n_1803)
);

AOI211xp5_ASAP7_75t_L g1804 ( 
.A1(n_1797),
.A2(n_1776),
.B(n_1772),
.C(n_1778),
.Y(n_1804)
);

OAI21xp5_ASAP7_75t_SL g1805 ( 
.A1(n_1791),
.A2(n_1786),
.B(n_1773),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1797),
.B(n_1763),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1792),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1801),
.A2(n_1778),
.B1(n_1772),
.B2(n_1789),
.C(n_1788),
.Y(n_1808)
);

O2A1O1Ixp33_ASAP7_75t_L g1809 ( 
.A1(n_1793),
.A2(n_1757),
.B(n_1767),
.C(n_1765),
.Y(n_1809)
);

AOI22xp5_ASAP7_75t_L g1810 ( 
.A1(n_1793),
.A2(n_1763),
.B1(n_1730),
.B2(n_1753),
.Y(n_1810)
);

A2O1A1Ixp33_ASAP7_75t_L g1811 ( 
.A1(n_1790),
.A2(n_1768),
.B(n_1767),
.C(n_1765),
.Y(n_1811)
);

AOI21xp33_ASAP7_75t_L g1812 ( 
.A1(n_1800),
.A2(n_1802),
.B(n_1799),
.Y(n_1812)
);

NOR5xp2_ASAP7_75t_L g1813 ( 
.A(n_1794),
.B(n_1745),
.C(n_1750),
.D(n_1755),
.E(n_1754),
.Y(n_1813)
);

OAI22xp33_ASAP7_75t_L g1814 ( 
.A1(n_1805),
.A2(n_1795),
.B1(n_1796),
.B2(n_1768),
.Y(n_1814)
);

AOI221xp5_ASAP7_75t_L g1815 ( 
.A1(n_1803),
.A2(n_1802),
.B1(n_1798),
.B2(n_1745),
.C(n_1755),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1804),
.B(n_1750),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1808),
.A2(n_1754),
.B(n_1762),
.Y(n_1817)
);

OAI311xp33_ASAP7_75t_L g1818 ( 
.A1(n_1810),
.A2(n_1740),
.A3(n_1742),
.B1(n_1736),
.C1(n_1737),
.Y(n_1818)
);

INVx2_ASAP7_75t_SL g1819 ( 
.A(n_1816),
.Y(n_1819)
);

NAND2x1_ASAP7_75t_SL g1820 ( 
.A(n_1818),
.B(n_1806),
.Y(n_1820)
);

AOI21xp5_ASAP7_75t_L g1821 ( 
.A1(n_1817),
.A2(n_1811),
.B(n_1812),
.Y(n_1821)
);

INVx1_ASAP7_75t_SL g1822 ( 
.A(n_1814),
.Y(n_1822)
);

HB1xp67_ASAP7_75t_L g1823 ( 
.A(n_1815),
.Y(n_1823)
);

INVx2_ASAP7_75t_L g1824 ( 
.A(n_1816),
.Y(n_1824)
);

AOI21xp33_ASAP7_75t_SL g1825 ( 
.A1(n_1819),
.A2(n_1809),
.B(n_1807),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1822),
.B(n_1735),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1820),
.Y(n_1827)
);

HB1xp67_ASAP7_75t_L g1828 ( 
.A(n_1822),
.Y(n_1828)
);

AOI22xp33_ASAP7_75t_R g1829 ( 
.A1(n_1823),
.A2(n_1813),
.B1(n_1762),
.B2(n_1719),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1826),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1828),
.Y(n_1831)
);

BUFx6f_ASAP7_75t_L g1832 ( 
.A(n_1827),
.Y(n_1832)
);

AND2x2_ASAP7_75t_L g1833 ( 
.A(n_1831),
.B(n_1824),
.Y(n_1833)
);

AOI322xp5_ASAP7_75t_L g1834 ( 
.A1(n_1833),
.A2(n_1831),
.A3(n_1830),
.B1(n_1832),
.B2(n_1829),
.C1(n_1821),
.C2(n_1825),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1834),
.B(n_1832),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1834),
.Y(n_1836)
);

OAI21x1_ASAP7_75t_L g1837 ( 
.A1(n_1835),
.A2(n_1832),
.B(n_1762),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1836),
.A2(n_1832),
.B(n_1719),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1838),
.A2(n_1742),
.B1(n_1737),
.B2(n_1736),
.Y(n_1839)
);

CKINVDCx20_ASAP7_75t_R g1840 ( 
.A(n_1839),
.Y(n_1840)
);

AOI21xp5_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1837),
.B(n_1738),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1738),
.B(n_1735),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1688),
.B1(n_1678),
.B2(n_1708),
.Y(n_1843)
);

AOI221xp5_ASAP7_75t_L g1844 ( 
.A1(n_1843),
.A2(n_1705),
.B1(n_1708),
.B2(n_1678),
.C(n_1688),
.Y(n_1844)
);

AOI211xp5_ASAP7_75t_L g1845 ( 
.A1(n_1844),
.A2(n_1705),
.B(n_1688),
.C(n_1702),
.Y(n_1845)
);


endmodule