module fake_jpeg_25030_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_6),
.B(n_2),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_42),
.Y(n_54)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx13_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_23),
.B(n_7),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_52),
.Y(n_78)
);

BUFx8_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_67),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_70),
.B(n_73),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_47),
.B1(n_43),
.B2(n_22),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_94),
.B1(n_69),
.B2(n_36),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_44),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_54),
.B(n_38),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_74),
.B(n_76),
.Y(n_112)
);

NAND2x2_ASAP7_75t_SL g75 ( 
.A(n_66),
.B(n_40),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_87),
.Y(n_129)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_81),
.Y(n_128)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_51),
.B(n_46),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_36),
.C(n_60),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_61),
.B(n_42),
.Y(n_81)
);

CKINVDCx12_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_53),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_34),
.B1(n_22),
.B2(n_30),
.Y(n_87)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_65),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_90),
.Y(n_133)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_56),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_38),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_92),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_55),
.A2(n_47),
.B1(n_22),
.B2(n_36),
.Y(n_94)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_32),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_99),
.C(n_20),
.Y(n_113)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_98),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_59),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_58),
.A2(n_34),
.B1(n_29),
.B2(n_30),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_26),
.Y(n_136)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_60),
.Y(n_105)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_105),
.Y(n_111)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_50),
.Y(n_106)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_46),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_107),
.B(n_110),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_75),
.A2(n_48),
.B1(n_25),
.B2(n_32),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_0),
.B(n_1),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_113),
.B(n_28),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_79),
.A2(n_47),
.B1(n_95),
.B2(n_78),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_117),
.A2(n_132),
.B1(n_135),
.B2(n_37),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_16),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_121),
.B(n_122),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_87),
.A2(n_0),
.B(n_1),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_124),
.B(n_130),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_40),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_126),
.B(n_136),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_104),
.B1(n_102),
.B2(n_82),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_86),
.A2(n_29),
.B1(n_25),
.B2(n_20),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_72),
.A2(n_48),
.B1(n_50),
.B2(n_45),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_94),
.A2(n_86),
.B1(n_97),
.B2(n_89),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_134),
.A2(n_82),
.B1(n_71),
.B2(n_93),
.Y(n_153)
);

O2A1O1Ixp33_ASAP7_75t_L g135 ( 
.A1(n_89),
.A2(n_37),
.B(n_41),
.C(n_19),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_137),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_L g140 ( 
.A1(n_121),
.A2(n_97),
.B1(n_88),
.B2(n_76),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_140),
.A2(n_151),
.B1(n_161),
.B2(n_167),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g141 ( 
.A1(n_136),
.A2(n_90),
.B1(n_104),
.B2(n_101),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g191 ( 
.A(n_141),
.B(n_166),
.Y(n_191)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_142),
.B(n_143),
.Y(n_184)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_125),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_133),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_145),
.B(n_155),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_100),
.B1(n_85),
.B2(n_80),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_146),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_118),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_147),
.Y(n_201)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_148),
.Y(n_178)
);

INVx3_ASAP7_75t_SL g149 ( 
.A(n_120),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_156),
.B1(n_158),
.B2(n_134),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_133),
.Y(n_155)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_157),
.A2(n_163),
.B(n_164),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_117),
.A2(n_37),
.B1(n_31),
.B2(n_27),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_125),
.Y(n_159)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_159),
.Y(n_181)
);

INVx13_ASAP7_75t_L g160 ( 
.A(n_125),
.Y(n_160)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_160),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_123),
.A2(n_93),
.B1(n_28),
.B2(n_33),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_109),
.B(n_112),
.Y(n_162)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_109),
.Y(n_163)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_115),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_147),
.B(n_128),
.Y(n_169)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_169),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_165),
.A2(n_152),
.B(n_154),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_171),
.A2(n_177),
.B(n_185),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_165),
.A2(n_132),
.B1(n_128),
.B2(n_122),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_150),
.B1(n_160),
.B2(n_143),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_154),
.B(n_107),
.Y(n_174)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_152),
.A2(n_129),
.B(n_110),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_175),
.A2(n_194),
.B(n_1),
.Y(n_204)
);

NAND2xp33_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_129),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_112),
.Y(n_180)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_139),
.A2(n_129),
.B(n_136),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_124),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_188),
.B(n_192),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_126),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_139),
.B(n_115),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_141),
.A2(n_135),
.B(n_113),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g195 ( 
.A(n_156),
.B(n_158),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_196),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_141),
.B(n_130),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_197),
.A2(n_27),
.B1(n_21),
.B2(n_24),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_142),
.B(n_127),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_198),
.B(n_199),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_164),
.B(n_135),
.Y(n_199)
);

O2A1O1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_119),
.B(n_131),
.C(n_37),
.Y(n_202)
);

OA22x2_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_167),
.B1(n_166),
.B2(n_137),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_148),
.C(n_144),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_203),
.B(n_229),
.C(n_195),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_204),
.B(n_175),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_167),
.B(n_149),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g256 ( 
.A1(n_205),
.A2(n_178),
.B(n_179),
.Y(n_256)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_206),
.A2(n_222),
.B(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_201),
.B(n_159),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_207),
.B(n_211),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_210),
.A2(n_200),
.B1(n_170),
.B2(n_187),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_119),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_35),
.Y(n_212)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_212),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_169),
.B(n_21),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_213),
.B(n_218),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_186),
.B(n_24),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_184),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_187),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_27),
.B1(n_21),
.B2(n_31),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_200),
.B1(n_202),
.B2(n_181),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_171),
.A2(n_1),
.B(n_2),
.Y(n_222)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_231),
.Y(n_243)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_172),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_225),
.A2(n_228),
.B1(n_230),
.B2(n_179),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_191),
.A2(n_2),
.B(n_3),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_197),
.A2(n_26),
.B1(n_24),
.B2(n_31),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_192),
.B(n_37),
.C(n_26),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_35),
.B1(n_28),
.B2(n_19),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_180),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_233),
.A2(n_235),
.B1(n_252),
.B2(n_230),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_234),
.B(n_242),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_170),
.B1(n_190),
.B2(n_194),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_210),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_236),
.A2(n_256),
.B(n_205),
.Y(n_259)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_227),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_240),
.B(n_246),
.Y(n_273)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_213),
.B(n_173),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_244),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_208),
.B(n_185),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_217),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_222),
.Y(n_246)
);

OAI22x1_ASAP7_75t_L g247 ( 
.A1(n_206),
.A2(n_191),
.B1(n_196),
.B2(n_176),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_247),
.A2(n_255),
.B1(n_221),
.B2(n_206),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_248),
.A2(n_254),
.B(n_226),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_209),
.B(n_174),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_203),
.B(n_190),
.C(n_178),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_229),
.C(n_216),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_181),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_205),
.Y(n_254)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_247),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_257),
.B(n_249),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_258),
.A2(n_266),
.B1(n_268),
.B2(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_259),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_208),
.C(n_217),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_261),
.B(n_265),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_263),
.B(n_276),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_251),
.B(n_216),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_228),
.B1(n_215),
.B2(n_212),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_271),
.C(n_275),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_252),
.A2(n_254),
.B1(n_240),
.B2(n_239),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_270),
.A2(n_206),
.B1(n_249),
.B2(n_255),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_215),
.C(n_220),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_243),
.A2(n_219),
.B(n_220),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_272),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_232),
.B(n_212),
.C(n_214),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_242),
.B(n_204),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_250),
.Y(n_279)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_281),
.B(n_285),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_256),
.B(n_249),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_282),
.A2(n_277),
.B(n_275),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_267),
.B(n_232),
.C(n_256),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_283),
.C(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_289),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_273),
.A2(n_238),
.B1(n_214),
.B2(n_237),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_294),
.Y(n_298)
);

AOI22xp33_ASAP7_75t_L g292 ( 
.A1(n_274),
.A2(n_241),
.B1(n_189),
.B2(n_183),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g305 ( 
.A(n_292),
.Y(n_305)
);

XNOR2x1_ASAP7_75t_L g293 ( 
.A(n_263),
.B(n_11),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_11),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_266),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_295),
.A2(n_284),
.B(n_293),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_261),
.C(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_296),
.B(n_300),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_278),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_287),
.B(n_260),
.C(n_265),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_291),
.B(n_276),
.C(n_33),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_306),
.Y(n_315)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_35),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_280),
.B(n_37),
.C(n_11),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_304),
.C(n_297),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_279),
.B(n_10),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_308),
.B(n_12),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_309),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_303),
.A2(n_288),
.B1(n_286),
.B2(n_282),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_298),
.B(n_294),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_312),
.B(n_316),
.Y(n_321)
);

HB1xp67_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g317 ( 
.A(n_299),
.B(n_278),
.Y(n_317)
);

OAI21x1_ASAP7_75t_SL g323 ( 
.A1(n_317),
.A2(n_305),
.B(n_307),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_318),
.B(n_7),
.C(n_14),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_302),
.A2(n_286),
.B1(n_4),
.B2(n_5),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_319),
.A2(n_311),
.B1(n_310),
.B2(n_6),
.Y(n_327)
);

OAI21x1_ASAP7_75t_L g320 ( 
.A1(n_314),
.A2(n_305),
.B(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_320),
.B(n_324),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_323),
.A2(n_315),
.B(n_319),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_327),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_318),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_331),
.C(n_324),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_322),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_327),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_329),
.B(n_325),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_10),
.B(n_13),
.Y(n_337)
);

AOI211xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_15),
.B(n_4),
.C(n_5),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_15),
.B(n_334),
.Y(n_340)
);


endmodule