module fake_aes_2256_n_700 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_700);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_700;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_12), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_69), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_23), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_61), .Y(n_82) );
INVx2_ASAP7_75t_L g83 ( .A(n_65), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_71), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_9), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_30), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_43), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_28), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_55), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_33), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_35), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_9), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_8), .Y(n_94) );
HB1xp67_ASAP7_75t_L g95 ( .A(n_12), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_18), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_15), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_15), .Y(n_98) );
INVx2_ASAP7_75t_L g99 ( .A(n_77), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_13), .Y(n_100) );
INVxp67_ASAP7_75t_SL g101 ( .A(n_60), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_51), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_49), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_29), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_74), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_70), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_5), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_19), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_26), .Y(n_109) );
BUFx3_ASAP7_75t_L g110 ( .A(n_0), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_50), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_27), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_45), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_57), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_78), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_31), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_68), .Y(n_117) );
CKINVDCx16_ASAP7_75t_R g118 ( .A(n_42), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_13), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_75), .Y(n_120) );
INVxp33_ASAP7_75t_SL g121 ( .A(n_53), .Y(n_121) );
INVxp67_ASAP7_75t_SL g122 ( .A(n_48), .Y(n_122) );
INVxp67_ASAP7_75t_L g123 ( .A(n_11), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_3), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_6), .Y(n_125) );
INVxp33_ASAP7_75t_SL g126 ( .A(n_40), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_110), .Y(n_127) );
AND2x2_ASAP7_75t_L g128 ( .A(n_98), .B(n_0), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
INVxp67_ASAP7_75t_L g130 ( .A(n_95), .Y(n_130) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_110), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_110), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_83), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_82), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_102), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_99), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_82), .Y(n_138) );
HB1xp67_ASAP7_75t_L g139 ( .A(n_123), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_94), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_86), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_99), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_89), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_94), .B(n_1), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_84), .B(n_1), .Y(n_148) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx3_ASAP7_75t_L g151 ( .A(n_106), .Y(n_151) );
BUFx3_ASAP7_75t_L g152 ( .A(n_106), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_106), .Y(n_153) );
HB1xp67_ASAP7_75t_L g154 ( .A(n_96), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_90), .Y(n_155) );
AND2x6_ASAP7_75t_L g156 ( .A(n_90), .B(n_36), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_91), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_91), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_92), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_84), .Y(n_160) );
AND2x2_ASAP7_75t_L g161 ( .A(n_102), .B(n_2), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_79), .B(n_2), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_108), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_103), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_103), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_105), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_108), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_105), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_131), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_129), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_133), .B(n_118), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_129), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_131), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_131), .Y(n_176) );
INVx3_ASAP7_75t_L g177 ( .A(n_162), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_131), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_131), .Y(n_179) );
BUFx6f_ASAP7_75t_L g180 ( .A(n_131), .Y(n_180) );
AND2x2_ASAP7_75t_L g181 ( .A(n_133), .B(n_118), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_134), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_130), .B(n_80), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_147), .Y(n_185) );
BUFx10_ASAP7_75t_L g186 ( .A(n_154), .Y(n_186) );
AND2x6_ASAP7_75t_L g187 ( .A(n_162), .B(n_114), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_135), .B(n_113), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g190 ( .A(n_136), .B(n_126), .Y(n_190) );
INVx2_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_134), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_135), .B(n_104), .Y(n_193) );
INVxp67_ASAP7_75t_L g194 ( .A(n_139), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_162), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_162), .Y(n_197) );
INVx2_ASAP7_75t_SL g198 ( .A(n_159), .Y(n_198) );
AND2x4_ASAP7_75t_SL g199 ( .A(n_161), .B(n_81), .Y(n_199) );
INVx2_ASAP7_75t_SL g200 ( .A(n_159), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_136), .B(n_125), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_137), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_128), .B(n_125), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_137), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_138), .B(n_121), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_134), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_134), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_128), .B(n_79), .Y(n_208) );
AND2x4_ASAP7_75t_L g209 ( .A(n_147), .B(n_119), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_147), .Y(n_210) );
INVx2_ASAP7_75t_SL g211 ( .A(n_159), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_156), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_161), .B(n_85), .Y(n_213) );
INVx1_ASAP7_75t_SL g214 ( .A(n_152), .Y(n_214) );
HB1xp67_ASAP7_75t_L g215 ( .A(n_138), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_140), .B(n_87), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_143), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_153), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_153), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_143), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_153), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_169), .B(n_119), .Y(n_222) );
INVx4_ASAP7_75t_SL g223 ( .A(n_156), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
BUFx2_ASAP7_75t_L g225 ( .A(n_152), .Y(n_225) );
BUFx6f_ASAP7_75t_L g226 ( .A(n_143), .Y(n_226) );
INVx4_ASAP7_75t_SL g227 ( .A(n_156), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_140), .B(n_124), .Y(n_228) );
AND2x4_ASAP7_75t_L g229 ( .A(n_142), .B(n_85), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_142), .B(n_111), .Y(n_230) );
OR2x2_ASAP7_75t_L g231 ( .A(n_169), .B(n_100), .Y(n_231) );
INVxp67_ASAP7_75t_L g232 ( .A(n_181), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_181), .B(n_100), .Y(n_233) );
NAND2x1p5_ASAP7_75t_L g234 ( .A(n_225), .B(n_107), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_215), .B(n_144), .Y(n_235) );
BUFx3_ASAP7_75t_L g236 ( .A(n_225), .Y(n_236) );
HB1xp67_ASAP7_75t_L g237 ( .A(n_194), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_205), .B(n_144), .Y(n_238) );
INVx3_ASAP7_75t_L g239 ( .A(n_177), .Y(n_239) );
BUFx4f_ASAP7_75t_SL g240 ( .A(n_186), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_222), .Y(n_241) );
INVx3_ASAP7_75t_L g242 ( .A(n_177), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_198), .Y(n_243) );
INVx2_ASAP7_75t_SL g244 ( .A(n_186), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_222), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_212), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_173), .Y(n_248) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_187), .Y(n_251) );
BUFx6f_ASAP7_75t_L g252 ( .A(n_212), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_229), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_229), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_229), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g256 ( .A(n_223), .B(n_159), .Y(n_256) );
A2O1A1Ixp33_ASAP7_75t_L g257 ( .A1(n_184), .A2(n_145), .B(n_167), .C(n_166), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_209), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g259 ( .A(n_223), .B(n_145), .Y(n_259) );
AND3x1_ASAP7_75t_L g260 ( .A(n_201), .B(n_107), .C(n_141), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_187), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_186), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_201), .B(n_146), .Y(n_263) );
BUFx8_ASAP7_75t_L g264 ( .A(n_213), .Y(n_264) );
BUFx2_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_200), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_214), .B(n_146), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_203), .B(n_150), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_213), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_209), .Y(n_270) );
HB1xp67_ASAP7_75t_L g271 ( .A(n_231), .Y(n_271) );
AND2x6_ASAP7_75t_L g272 ( .A(n_177), .B(n_109), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_228), .A2(n_120), .B1(n_167), .B2(n_166), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_188), .B(n_150), .Y(n_274) );
AOI22xp5_ASAP7_75t_L g275 ( .A1(n_187), .A2(n_165), .B1(n_163), .B2(n_155), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_199), .B(n_93), .Y(n_277) );
OR2x4_ASAP7_75t_L g278 ( .A(n_190), .B(n_155), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_203), .B(n_157), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_231), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_200), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_185), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_SL g283 ( .A1(n_230), .A2(n_151), .B(n_168), .C(n_164), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
INVx3_ASAP7_75t_L g285 ( .A(n_195), .Y(n_285) );
NOR2xp33_ASAP7_75t_R g286 ( .A(n_187), .B(n_156), .Y(n_286) );
CKINVDCx20_ASAP7_75t_R g287 ( .A(n_199), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_195), .Y(n_288) );
INVx2_ASAP7_75t_SL g289 ( .A(n_208), .Y(n_289) );
INVx5_ASAP7_75t_L g290 ( .A(n_187), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_193), .B(n_157), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_216), .B(n_158), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_183), .B(n_158), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_211), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_171), .Y(n_295) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_208), .A2(n_165), .B1(n_163), .B2(n_156), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_211), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_271), .Y(n_298) );
OR2x6_ASAP7_75t_L g299 ( .A(n_244), .B(n_195), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g300 ( .A(n_251), .B(n_197), .Y(n_300) );
INVx5_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_240), .Y(n_302) );
BUFx3_ASAP7_75t_L g303 ( .A(n_264), .Y(n_303) );
AOI22xp33_ASAP7_75t_L g304 ( .A1(n_280), .A2(n_197), .B1(n_156), .B2(n_152), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_261), .Y(n_305) );
CKINVDCx5p33_ASAP7_75t_R g306 ( .A(n_240), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_264), .Y(n_307) );
INVx3_ASAP7_75t_SL g308 ( .A(n_287), .Y(n_308) );
NAND2x1p5_ASAP7_75t_L g309 ( .A(n_251), .B(n_197), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_237), .B(n_171), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_271), .Y(n_311) );
O2A1O1Ixp33_ASAP7_75t_L g312 ( .A1(n_257), .A2(n_148), .B(n_221), .C(n_219), .Y(n_312) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_237), .B(n_262), .Y(n_313) );
CKINVDCx8_ASAP7_75t_R g314 ( .A(n_263), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_241), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_245), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_250), .Y(n_317) );
A2O1A1Ixp33_ASAP7_75t_L g318 ( .A1(n_257), .A2(n_174), .B(n_172), .C(n_202), .Y(n_318) );
BUFx6f_ASAP7_75t_L g319 ( .A(n_261), .Y(n_319) );
NAND3xp33_ASAP7_75t_L g320 ( .A(n_296), .B(n_174), .C(n_204), .Y(n_320) );
INVx1_ASAP7_75t_SL g321 ( .A(n_269), .Y(n_321) );
AOI22xp5_ASAP7_75t_L g322 ( .A1(n_232), .A2(n_156), .B1(n_97), .B2(n_221), .Y(n_322) );
NAND2x1_ASAP7_75t_SL g323 ( .A(n_273), .B(n_172), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_274), .A2(n_189), .B(n_219), .Y(n_324) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_236), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_239), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_263), .B(n_189), .Y(n_327) );
OAI22x1_ASAP7_75t_L g328 ( .A1(n_234), .A2(n_101), .B1(n_122), .B2(n_109), .Y(n_328) );
AOI22xp5_ASAP7_75t_L g329 ( .A1(n_232), .A2(n_156), .B1(n_204), .B2(n_218), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_253), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_254), .Y(n_331) );
CKINVDCx20_ASAP7_75t_R g332 ( .A(n_287), .Y(n_332) );
INVx4_ASAP7_75t_L g333 ( .A(n_261), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_255), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_263), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_258), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_270), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_248), .Y(n_338) );
INVx3_ASAP7_75t_L g339 ( .A(n_239), .Y(n_339) );
INVx4_ASAP7_75t_L g340 ( .A(n_290), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_248), .B(n_202), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_236), .Y(n_342) );
AOI22xp5_ASAP7_75t_L g343 ( .A1(n_260), .A2(n_218), .B1(n_223), .B2(n_227), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_276), .Y(n_344) );
OAI22xp33_ASAP7_75t_L g345 ( .A1(n_278), .A2(n_141), .B1(n_151), .B2(n_168), .Y(n_345) );
BUFx3_ASAP7_75t_L g346 ( .A(n_289), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_268), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_242), .Y(n_348) );
INVx3_ASAP7_75t_L g349 ( .A(n_242), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_305), .Y(n_350) );
OAI22xp5_ASAP7_75t_L g351 ( .A1(n_341), .A2(n_267), .B1(n_275), .B2(n_233), .Y(n_351) );
INVx3_ASAP7_75t_L g352 ( .A(n_333), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_338), .A2(n_233), .B1(n_277), .B2(n_279), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_298), .A2(n_279), .B1(n_272), .B2(n_234), .Y(n_354) );
AND2x4_ASAP7_75t_L g355 ( .A(n_327), .B(n_290), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_314), .A2(n_235), .B1(n_278), .B2(n_295), .Y(n_356) );
AOI22xp33_ASAP7_75t_SL g357 ( .A1(n_335), .A2(n_272), .B1(n_286), .B2(n_265), .Y(n_357) );
OAI22xp33_ASAP7_75t_L g358 ( .A1(n_308), .A2(n_293), .B1(n_291), .B2(n_292), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_305), .Y(n_359) );
BUFx12f_ASAP7_75t_L g360 ( .A(n_302), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_315), .Y(n_361) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_304), .A2(n_282), .B1(n_284), .B2(n_238), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_305), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_321), .B(n_285), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_310), .B(n_311), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_316), .Y(n_366) );
A2O1A1Ixp33_ASAP7_75t_L g367 ( .A1(n_312), .A2(n_285), .B(n_288), .C(n_283), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_317), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_347), .A2(n_272), .B1(n_288), .B2(n_286), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_305), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_319), .Y(n_372) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_325), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_330), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g375 ( .A1(n_308), .A2(n_290), .B1(n_246), .B2(n_249), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_319), .Y(n_376) );
AO31x2_ASAP7_75t_L g377 ( .A1(n_318), .A2(n_164), .A3(n_168), .B(n_127), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_319), .Y(n_378) );
INVx1_ASAP7_75t_SL g379 ( .A(n_325), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_304), .A2(n_290), .B1(n_294), .B2(n_281), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_345), .B(n_272), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_331), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_365), .Y(n_383) );
AOI22xp5_ASAP7_75t_L g384 ( .A1(n_358), .A2(n_332), .B1(n_313), .B2(n_307), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_346), .B1(n_345), .B2(n_342), .Y(n_385) );
AOI221xp5_ASAP7_75t_L g386 ( .A1(n_353), .A2(n_328), .B1(n_312), .B2(n_334), .C(n_337), .Y(n_386) );
INVx5_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_365), .B(n_342), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_360), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_351), .A2(n_329), .B1(n_299), .B2(n_318), .Y(n_390) );
AOI22xp33_ASAP7_75t_SL g391 ( .A1(n_381), .A2(n_332), .B1(n_303), .B2(n_306), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_379), .A2(n_299), .B1(n_343), .B2(n_322), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_373), .A2(n_272), .B1(n_299), .B2(n_344), .Y(n_393) );
OAI22xp33_ASAP7_75t_L g394 ( .A1(n_379), .A2(n_336), .B1(n_324), .B2(n_309), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_382), .Y(n_395) );
AOI22xp33_ASAP7_75t_L g396 ( .A1(n_362), .A2(n_348), .B1(n_349), .B2(n_339), .Y(n_396) );
OAI221xp5_ASAP7_75t_L g397 ( .A1(n_354), .A2(n_323), .B1(n_283), .B2(n_324), .C(n_320), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_357), .A2(n_300), .B1(n_309), .B2(n_301), .Y(n_398) );
CKINVDCx5p33_ASAP7_75t_R g399 ( .A(n_360), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g400 ( .A1(n_382), .A2(n_349), .B1(n_339), .B2(n_326), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g401 ( .A1(n_360), .A2(n_151), .B1(n_300), .B2(n_301), .Y(n_401) );
NOR2x1_ASAP7_75t_L g402 ( .A(n_364), .B(n_340), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_378), .Y(n_403) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_333), .B(n_340), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_369), .A2(n_301), .B1(n_151), .B2(n_281), .Y(n_405) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_382), .A2(n_297), .B1(n_266), .B2(n_243), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_364), .A2(n_301), .B1(n_141), .B2(n_111), .Y(n_407) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_361), .A2(n_141), .B1(n_132), .B2(n_127), .C(n_164), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_378), .Y(n_409) );
OAI22xp33_ASAP7_75t_L g410 ( .A1(n_361), .A2(n_112), .B1(n_114), .B2(n_115), .Y(n_410) );
OAI211xp5_ASAP7_75t_L g411 ( .A1(n_384), .A2(n_368), .B(n_366), .C(n_374), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_395), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_385), .B(n_112), .C(n_115), .D(n_116), .Y(n_413) );
NAND3xp33_ASAP7_75t_L g414 ( .A(n_386), .B(n_160), .C(n_143), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_383), .B(n_366), .Y(n_415) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_389), .A2(n_374), .B1(n_368), .B2(n_352), .Y(n_416) );
BUFx2_ASAP7_75t_L g417 ( .A(n_409), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_388), .B(n_377), .Y(n_418) );
OAI21xp33_ASAP7_75t_L g419 ( .A1(n_391), .A2(n_367), .B(n_116), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_395), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_388), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_387), .Y(n_422) );
AO21x2_ASAP7_75t_L g423 ( .A1(n_394), .A2(n_372), .B(n_350), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_408), .Y(n_424) );
OAI222xp33_ASAP7_75t_L g425 ( .A1(n_402), .A2(n_117), .B1(n_352), .B2(n_355), .C1(n_372), .C2(n_371), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_409), .Y(n_426) );
AOI221xp5_ASAP7_75t_SL g427 ( .A1(n_410), .A2(n_117), .B1(n_132), .B2(n_160), .C(n_149), .Y(n_427) );
OAI22xp5_ASAP7_75t_L g428 ( .A1(n_390), .A2(n_352), .B1(n_355), .B2(n_380), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g429 ( .A1(n_393), .A2(n_355), .B1(n_378), .B2(n_372), .Y(n_429) );
AOI21x1_ASAP7_75t_L g430 ( .A1(n_398), .A2(n_363), .B(n_376), .Y(n_430) );
INVx3_ASAP7_75t_L g431 ( .A(n_387), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_403), .Y(n_432) );
OA21x2_ASAP7_75t_L g433 ( .A1(n_397), .A2(n_350), .B(n_376), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_403), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_387), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_387), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_403), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g438 ( .A1(n_392), .A2(n_355), .B1(n_376), .B2(n_371), .Y(n_438) );
OA21x2_ASAP7_75t_L g439 ( .A1(n_396), .A2(n_350), .B(n_371), .Y(n_439) );
OR2x6_ASAP7_75t_L g440 ( .A(n_389), .B(n_359), .Y(n_440) );
AOI211xp5_ASAP7_75t_L g441 ( .A1(n_407), .A2(n_160), .B(n_143), .C(n_149), .Y(n_441) );
AOI33xp33_ASAP7_75t_L g442 ( .A1(n_401), .A2(n_179), .A3(n_191), .B1(n_192), .B2(n_196), .B3(n_206), .Y(n_442) );
AND2x4_ASAP7_75t_L g443 ( .A(n_387), .B(n_359), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_405), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_400), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_420), .Y(n_446) );
AND2x2_ASAP7_75t_SL g447 ( .A(n_417), .B(n_359), .Y(n_447) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_431), .B(n_363), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_418), .B(n_377), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_418), .B(n_377), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_412), .B(n_377), .Y(n_451) );
BUFx2_ASAP7_75t_L g452 ( .A(n_417), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_412), .Y(n_453) );
AND2x2_ASAP7_75t_L g454 ( .A(n_421), .B(n_377), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_422), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_422), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_426), .B(n_377), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_421), .B(n_149), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_420), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_432), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_432), .B(n_363), .Y(n_461) );
INVx1_ASAP7_75t_SL g462 ( .A(n_431), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_419), .A2(n_399), .B1(n_406), .B2(n_404), .C(n_160), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_424), .A2(n_399), .B1(n_160), .B2(n_149), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_426), .B(n_149), .Y(n_465) );
NAND3xp33_ASAP7_75t_L g466 ( .A(n_411), .B(n_149), .C(n_160), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_434), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_437), .Y(n_469) );
AND2x4_ASAP7_75t_SL g470 ( .A(n_431), .B(n_370), .Y(n_470) );
AND2x2_ASAP7_75t_SL g471 ( .A(n_438), .B(n_370), .Y(n_471) );
INVx5_ASAP7_75t_L g472 ( .A(n_440), .Y(n_472) );
INVx2_ASAP7_75t_SL g473 ( .A(n_436), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_415), .B(n_3), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_436), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_445), .A2(n_370), .B1(n_220), .B2(n_180), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_439), .Y(n_479) );
OAI33xp33_ASAP7_75t_L g480 ( .A1(n_413), .A2(n_4), .A3(n_5), .B1(n_6), .B2(n_7), .B3(n_8), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_439), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_440), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_443), .B(n_4), .Y(n_483) );
AND2x4_ASAP7_75t_SL g484 ( .A(n_440), .B(n_294), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_433), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
AOI211xp5_ASAP7_75t_SL g488 ( .A1(n_416), .A2(n_7), .B(n_10), .C(n_11), .Y(n_488) );
AND2x2_ASAP7_75t_SL g489 ( .A(n_433), .B(n_246), .Y(n_489) );
NOR3xp33_ASAP7_75t_L g490 ( .A(n_435), .B(n_196), .C(n_178), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_443), .B(n_67), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
OAI33xp33_ASAP7_75t_L g493 ( .A1(n_445), .A2(n_10), .A3(n_14), .B1(n_16), .B2(n_17), .B3(n_18), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_442), .B(n_175), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_443), .B(n_72), .Y(n_495) );
INVx2_ASAP7_75t_L g496 ( .A(n_453), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_469), .B(n_423), .Y(n_497) );
BUFx2_ASAP7_75t_L g498 ( .A(n_455), .Y(n_498) );
OAI221xp5_ASAP7_75t_L g499 ( .A1(n_475), .A2(n_440), .B1(n_427), .B2(n_428), .C(n_414), .Y(n_499) );
OR2x2_ASAP7_75t_L g500 ( .A(n_456), .B(n_444), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_453), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_483), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_477), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_454), .B(n_444), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_446), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_480), .B(n_425), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_483), .B(n_429), .Y(n_507) );
NAND2xp33_ASAP7_75t_L g508 ( .A(n_472), .B(n_441), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
NOR3xp33_ASAP7_75t_L g510 ( .A(n_493), .B(n_430), .C(n_217), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_454), .B(n_423), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_460), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_460), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_472), .B(n_430), .Y(n_514) );
AOI33xp33_ASAP7_75t_L g515 ( .A1(n_467), .A2(n_14), .A3(n_16), .B1(n_17), .B2(n_206), .B3(n_217), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_449), .B(n_450), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_449), .B(n_423), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_473), .B(n_207), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_467), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_472), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_450), .B(n_170), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_468), .Y(n_522) );
NOR3xp33_ASAP7_75t_L g523 ( .A(n_463), .B(n_192), .C(n_178), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_468), .B(n_451), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_473), .B(n_20), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_451), .B(n_170), .Y(n_526) );
AND4x1_ASAP7_75t_L g527 ( .A(n_488), .B(n_466), .C(n_448), .D(n_464), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_452), .B(n_21), .Y(n_528) );
NOR2x1_ASAP7_75t_L g529 ( .A(n_466), .B(n_207), .Y(n_529) );
INVxp33_ASAP7_75t_L g530 ( .A(n_452), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_462), .B(n_465), .Y(n_531) );
INVxp67_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_469), .Y(n_533) );
AND2x2_ASAP7_75t_L g534 ( .A(n_465), .B(n_22), .Y(n_534) );
NAND3xp33_ASAP7_75t_L g535 ( .A(n_458), .B(n_224), .C(n_176), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_474), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_447), .B(n_24), .Y(n_537) );
OR2x6_ASAP7_75t_L g538 ( .A(n_482), .B(n_175), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_457), .B(n_191), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_457), .B(n_179), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_458), .B(n_259), .C(n_256), .Y(n_542) );
INVx2_ASAP7_75t_L g543 ( .A(n_486), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_486), .Y(n_544) );
NAND4xp25_ASAP7_75t_L g545 ( .A(n_487), .B(n_256), .C(n_259), .D(n_247), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_461), .B(n_25), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_461), .B(n_32), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_447), .B(n_34), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_447), .B(n_37), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_461), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_461), .B(n_38), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_448), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_484), .B(n_39), .Y(n_554) );
AOI211x1_ASAP7_75t_L g555 ( .A1(n_527), .A2(n_492), .B(n_494), .C(n_481), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_503), .B(n_471), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_503), .B(n_492), .C(n_490), .Y(n_557) );
NAND2xp5_ASAP7_75t_SL g558 ( .A(n_505), .B(n_472), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_498), .B(n_476), .Y(n_559) );
NAND4xp25_ASAP7_75t_L g560 ( .A(n_506), .B(n_491), .C(n_495), .D(n_479), .Y(n_560) );
O2A1O1Ixp33_ASAP7_75t_SL g561 ( .A1(n_502), .A2(n_472), .B(n_476), .C(n_481), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_512), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_509), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_516), .B(n_479), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_524), .B(n_471), .Y(n_565) );
OAI22xp5_ASAP7_75t_SL g566 ( .A1(n_506), .A2(n_472), .B1(n_471), .B2(n_491), .Y(n_566) );
AOI21xp5_ASAP7_75t_SL g567 ( .A1(n_537), .A2(n_495), .B(n_491), .Y(n_567) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_507), .A2(n_495), .B1(n_491), .B2(n_489), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_509), .Y(n_569) );
NOR3xp33_ASAP7_75t_L g570 ( .A(n_515), .B(n_495), .C(n_485), .Y(n_570) );
OAI32xp33_ASAP7_75t_L g571 ( .A1(n_530), .A2(n_485), .A3(n_484), .B1(n_478), .B2(n_489), .Y(n_571) );
NAND4xp25_ASAP7_75t_L g572 ( .A(n_515), .B(n_247), .C(n_489), .D(n_470), .Y(n_572) );
OAI31xp33_ASAP7_75t_L g573 ( .A1(n_499), .A2(n_470), .A3(n_44), .B(n_46), .Y(n_573) );
NAND2xp5_ASAP7_75t_SL g574 ( .A(n_520), .B(n_529), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_504), .B(n_470), .Y(n_575) );
NAND4xp25_ASAP7_75t_SL g576 ( .A(n_548), .B(n_41), .C(n_47), .D(n_52), .Y(n_576) );
OAI31xp33_ASAP7_75t_L g577 ( .A1(n_549), .A2(n_54), .A3(n_56), .B(n_58), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_513), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_531), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_500), .B(n_182), .Y(n_580) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_530), .A2(n_182), .B1(n_226), .B2(n_224), .Y(n_581) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_514), .A2(n_59), .B(n_62), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_550), .B(n_64), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_496), .B(n_66), .Y(n_584) );
NAND2x1_ASAP7_75t_L g585 ( .A(n_520), .B(n_180), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_519), .B(n_180), .Y(n_586) );
NOR2xp67_ASAP7_75t_SL g587 ( .A(n_554), .B(n_252), .Y(n_587) );
INVxp67_ASAP7_75t_L g588 ( .A(n_552), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_496), .B(n_73), .Y(n_589) );
NOR2x1_ASAP7_75t_L g590 ( .A(n_508), .B(n_182), .Y(n_590) );
OAI221xp5_ASAP7_75t_SL g591 ( .A1(n_517), .A2(n_76), .B1(n_175), .B2(n_176), .C(n_180), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_522), .B(n_175), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_501), .B(n_175), .Y(n_593) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_510), .A2(n_176), .B1(n_180), .B2(n_182), .Y(n_594) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_508), .A2(n_176), .B1(n_182), .B2(n_220), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_532), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_532), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_533), .B(n_176), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_539), .B(n_220), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_536), .B(n_220), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_511), .B(n_224), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_553), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_553), .Y(n_603) );
OAI21xp5_ASAP7_75t_L g604 ( .A1(n_523), .A2(n_224), .B(n_226), .Y(n_604) );
INVxp67_ASAP7_75t_L g605 ( .A(n_497), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_602), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_562), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_605), .B(n_497), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_578), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g610 ( .A1(n_560), .A2(n_528), .B1(n_523), .B2(n_510), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_596), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_579), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_597), .B(n_544), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_564), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_559), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_603), .Y(n_616) );
OAI22xp5_ASAP7_75t_L g617 ( .A1(n_567), .A2(n_538), .B1(n_547), .B2(n_546), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_563), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_569), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_588), .Y(n_620) );
AOI311xp33_ASAP7_75t_L g621 ( .A1(n_566), .A2(n_521), .A3(n_542), .B(n_526), .C(n_497), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_565), .B(n_543), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_588), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_575), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_558), .Y(n_625) );
XOR2x2_ASAP7_75t_L g626 ( .A(n_555), .B(n_551), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_586), .Y(n_627) );
AND2x2_ASAP7_75t_L g628 ( .A(n_605), .B(n_543), .Y(n_628) );
NAND2xp33_ASAP7_75t_SL g629 ( .A(n_558), .B(n_525), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_592), .Y(n_630) );
OAI22xp5_ASAP7_75t_L g631 ( .A1(n_568), .A2(n_538), .B1(n_535), .B2(n_514), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_580), .Y(n_632) );
NOR2xp33_ASAP7_75t_SL g633 ( .A(n_590), .B(n_534), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
XOR2xp5_ASAP7_75t_L g635 ( .A(n_556), .B(n_541), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_593), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_568), .B(n_540), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_598), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_600), .Y(n_639) );
OAI21xp33_ASAP7_75t_SL g640 ( .A1(n_574), .A2(n_538), .B(n_545), .Y(n_640) );
INVxp67_ASAP7_75t_L g641 ( .A(n_557), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g642 ( .A1(n_573), .A2(n_542), .B1(n_518), .B2(n_226), .C(n_224), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_599), .Y(n_643) );
NOR2x1_ASAP7_75t_L g644 ( .A(n_572), .B(n_226), .Y(n_644) );
AOI22xp5_ASAP7_75t_L g645 ( .A1(n_570), .A2(n_226), .B1(n_223), .B2(n_227), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_570), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_574), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g648 ( .A1(n_561), .A2(n_576), .B(n_571), .C(n_591), .Y(n_648) );
INVxp67_ASAP7_75t_L g649 ( .A(n_587), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_585), .Y(n_650) );
AOI221xp5_ASAP7_75t_SL g651 ( .A1(n_594), .A2(n_246), .B1(n_249), .B2(n_252), .C(n_227), .Y(n_651) );
XNOR2xp5_ASAP7_75t_L g652 ( .A(n_595), .B(n_227), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_604), .B(n_246), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_583), .A2(n_249), .B1(n_252), .B2(n_581), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_561), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_584), .Y(n_656) );
INVx3_ASAP7_75t_L g657 ( .A(n_582), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_589), .Y(n_658) );
INVx1_ASAP7_75t_L g659 ( .A(n_583), .Y(n_659) );
NAND3xp33_ASAP7_75t_L g660 ( .A(n_594), .B(n_577), .C(n_581), .Y(n_660) );
AOI22xp33_ASAP7_75t_SL g661 ( .A1(n_566), .A2(n_249), .B1(n_252), .B2(n_503), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_596), .B(n_597), .Y(n_662) );
INVxp67_ASAP7_75t_L g663 ( .A(n_559), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_646), .A2(n_644), .B1(n_626), .B2(n_637), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_L g665 ( .A1(n_640), .A2(n_629), .B(n_648), .C(n_641), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_608), .Y(n_666) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_626), .A2(n_617), .B1(n_629), .B2(n_624), .Y(n_667) );
AOI32xp33_ASAP7_75t_L g668 ( .A1(n_621), .A2(n_612), .A3(n_661), .B1(n_655), .B2(n_625), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_L g669 ( .A1(n_642), .A2(n_657), .B(n_649), .C(n_631), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_662), .Y(n_670) );
NAND3xp33_ASAP7_75t_L g671 ( .A(n_647), .B(n_623), .C(n_620), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g672 ( .A1(n_637), .A2(n_659), .B1(n_635), .B2(n_657), .Y(n_672) );
NOR3xp33_ASAP7_75t_L g673 ( .A(n_642), .B(n_660), .C(n_661), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_662), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_610), .A2(n_663), .B1(n_635), .B2(n_614), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g676 ( .A1(n_633), .A2(n_645), .B1(n_615), .B2(n_623), .C(n_611), .Y(n_676) );
AO22x2_ASAP7_75t_L g677 ( .A1(n_607), .A2(n_609), .B1(n_650), .B2(n_616), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_668), .B(n_608), .Y(n_678) );
NOR3xp33_ASAP7_75t_L g679 ( .A(n_665), .B(n_654), .C(n_653), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_670), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_664), .B(n_673), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g682 ( .A1(n_667), .A2(n_675), .B1(n_672), .B2(n_674), .Y(n_682) );
AO22x2_ASAP7_75t_L g683 ( .A1(n_671), .A2(n_606), .B1(n_616), .B2(n_619), .Y(n_683) );
NAND2xp5_ASAP7_75t_SL g684 ( .A(n_669), .B(n_651), .Y(n_684) );
AOI211xp5_ASAP7_75t_L g685 ( .A1(n_676), .A2(n_627), .B(n_630), .C(n_643), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_681), .B(n_677), .Y(n_686) );
INVxp33_ASAP7_75t_SL g687 ( .A(n_682), .Y(n_687) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_678), .B(n_666), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_679), .B(n_677), .Y(n_689) );
XOR2xp5_ASAP7_75t_L g690 ( .A(n_684), .B(n_632), .Y(n_690) );
AOI221xp5_ASAP7_75t_L g691 ( .A1(n_687), .A2(n_683), .B1(n_685), .B2(n_680), .C(n_638), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_689), .B(n_613), .C(n_622), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_686), .A2(n_606), .B1(n_636), .B2(n_634), .C(n_656), .Y(n_693) );
AOI22xp5_ASAP7_75t_SL g694 ( .A1(n_691), .A2(n_690), .B1(n_688), .B2(n_652), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_693), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_695), .Y(n_696) );
OAI22x1_ASAP7_75t_L g697 ( .A1(n_694), .A2(n_692), .B1(n_658), .B2(n_634), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_696), .Y(n_698) );
OA22x2_ASAP7_75t_L g699 ( .A1(n_698), .A2(n_697), .B1(n_628), .B2(n_618), .Y(n_699) );
OAI21xp33_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_628), .B(n_639), .Y(n_700) );
endmodule