module real_jpeg_5775_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx8_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_42),
.B1(n_80),
.B2(n_83),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_1),
.A2(n_83),
.B1(n_158),
.B2(n_160),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_1),
.A2(n_83),
.B1(n_187),
.B2(n_189),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_1),
.A2(n_22),
.B1(n_83),
.B2(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_2),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_2),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_3),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_3),
.Y(n_114)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_3),
.Y(n_146)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_4),
.Y(n_61)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_5),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_5),
.Y(n_230)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_5),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_5),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_22),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_49),
.B1(n_86),
.B2(n_90),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_6),
.A2(n_49),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_6),
.A2(n_49),
.B1(n_260),
.B2(n_262),
.Y(n_259)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_9),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_21),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_10),
.B(n_40),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_10),
.A2(n_21),
.B1(n_172),
.B2(n_173),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_21),
.B1(n_91),
.B2(n_206),
.Y(n_205)
);

O2A1O1Ixp33_ASAP7_75t_L g219 ( 
.A1(n_10),
.A2(n_220),
.B(n_221),
.C(n_227),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_10),
.B(n_248),
.C(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_10),
.B(n_92),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_10),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_10),
.B(n_106),
.Y(n_293)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_11),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_11),
.Y(n_102)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_208),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_14),
.B(n_207),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_177),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_16),
.B(n_177),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_123),
.C(n_162),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_17),
.B(n_212),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_52),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_18),
.B(n_53),
.C(n_94),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B(n_24),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_21),
.B(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g221 ( 
.A1(n_21),
.A2(n_222),
.B(n_224),
.Y(n_221)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g132 ( 
.A(n_24),
.Y(n_132)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_27),
.B(n_48),
.Y(n_200)
);

NOR2x1_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_40),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_30),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_32),
.B(n_134),
.Y(n_133)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_40),
.B(n_197),
.Y(n_196)
);

AO22x1_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_44),
.B2(n_46),
.Y(n_40)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_41),
.Y(n_129)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_43),
.Y(n_128)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_43),
.Y(n_136)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_44),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_93),
.B1(n_94),
.B2(n_122),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_84),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_78),
.Y(n_55)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_56),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_69),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_64),
.Y(n_220)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_69),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B1(n_74),
.B2(n_76),
.Y(n_69)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_72),
.Y(n_98)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_73),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_73),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_76),
.Y(n_223)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_79),
.B(n_92),
.Y(n_164)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_84),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_85),
.B(n_92),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_85),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_115),
.B(n_116),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_96),
.B(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_96),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_96),
.B(n_186),
.Y(n_303)
);

NOR2x1_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_106),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_97)
);

AO22x1_ASAP7_75t_SL g106 ( 
.A1(n_99),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_106)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_101),
.Y(n_248)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx5_ASAP7_75t_L g226 ( 
.A(n_105),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_105),
.Y(n_239)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_106),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_106),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_106),
.B(n_236),
.Y(n_251)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_112),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_112),
.Y(n_262)
);

INVx8_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_114),
.Y(n_261)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_114),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_115),
.B(n_116),
.Y(n_234)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_123),
.A2(n_124),
.B1(n_162),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_137),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_125),
.B(n_137),
.Y(n_193)
);

AOI32xp33_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_129),
.A3(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

INVx6_ASAP7_75t_SL g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_134),
.Y(n_227)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_147),
.B(n_151),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_138),
.A2(n_176),
.B(n_182),
.Y(n_181)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_145),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_146),
.Y(n_175)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_148),
.B(n_157),
.Y(n_176)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_150),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_151),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_157),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_152),
.B(n_171),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_152),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_152),
.A2(n_171),
.B(n_229),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_152),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_155),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_161),
.Y(n_249)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_169),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_163),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_202),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_166),
.B(n_205),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_169),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_176),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_170),
.B(n_274),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_171),
.Y(n_256)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_176),
.B(n_258),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_192),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

AND2x2_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_184),
.B(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_185),
.B(n_235),
.Y(n_264)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_200),
.Y(n_195)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_240),
.B(n_316),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_211),
.B(n_214),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_231),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_215),
.B(n_312),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_218),
.A2(n_231),
.B1(n_232),
.B2(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_218),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_228),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_219),
.A2(n_228),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_219),
.Y(n_308)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_247),
.Y(n_246)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_228),
.Y(n_307)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_235),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_241),
.A2(n_310),
.B(n_315),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_242),
.A2(n_297),
.B(n_309),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_268),
.B(n_296),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_252),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_244),
.B(n_252),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_250),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_245),
.A2(n_246),
.B1(n_250),
.B2(n_271),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_303),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_263),
.Y(n_252)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_253),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_259),
.B(n_275),
.Y(n_274)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_265),
.B(n_266),
.C(n_299),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_279),
.B(n_295),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_272),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_272),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_278),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_280),
.A2(n_291),
.B(n_294),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_290),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g283 ( 
.A(n_284),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_292),
.B(n_293),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_300),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_306),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_302),
.B(n_304),
.C(n_306),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_314),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_314),
.Y(n_315)
);


endmodule