module fake_jpeg_26155_n_49 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_49);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_49;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

CKINVDCx14_ASAP7_75t_R g7 ( 
.A(n_5),
.Y(n_7)
);

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx5_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_2),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_17),
.Y(n_27)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_12),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_19),
.A2(n_21),
.B1(n_22),
.B2(n_14),
.Y(n_24)
);

CKINVDCx11_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_11),
.C(n_2),
.Y(n_26)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_26),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_8),
.B1(n_11),
.B2(n_7),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_25),
.A2(n_29),
.B1(n_24),
.B2(n_21),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_21),
.A2(n_17),
.B1(n_18),
.B2(n_22),
.Y(n_29)
);

FAx1_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_20),
.CI(n_15),
.CON(n_31),
.SN(n_31)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_32),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_33),
.A2(n_35),
.B1(n_31),
.B2(n_37),
.Y(n_42)
);

OA21x2_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_1),
.B(n_3),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_28),
.B1(n_4),
.B2(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_27),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_6),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_30),
.C(n_28),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_42),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_31),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_38),
.C(n_33),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_45),
.B(n_41),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_47),
.B(n_43),
.Y(n_48)
);

NOR3xp33_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_34),
.C(n_47),
.Y(n_49)
);


endmodule