module fake_jpeg_25377_n_216 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_SL g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_22),
.B(n_10),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_34),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_28),
.Y(n_43)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_31),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx6_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_30),
.C(n_27),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_17),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_26),
.A2(n_24),
.B1(n_15),
.B2(n_21),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_25),
.B1(n_23),
.B2(n_13),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_30),
.A2(n_15),
.B1(n_20),
.B2(n_21),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_40),
.A2(n_41),
.B1(n_25),
.B2(n_20),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_32),
.A2(n_15),
.B1(n_23),
.B2(n_21),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_18),
.B1(n_25),
.B2(n_20),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_23),
.B1(n_13),
.B2(n_12),
.Y(n_59)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_56),
.B1(n_13),
.B2(n_12),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_58),
.Y(n_68)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_54),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_34),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_28),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_61),
.Y(n_74)
);

INVxp67_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_16),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_59),
.A2(n_63),
.B1(n_12),
.B2(n_19),
.Y(n_73)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

NOR2x1_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_33),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_62),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_18),
.B1(n_33),
.B2(n_28),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_42),
.B(n_19),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_67),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_42),
.C(n_46),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_44),
.Y(n_66)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_72),
.B(n_65),
.C(n_59),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_73),
.A2(n_87),
.B1(n_56),
.B2(n_67),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_43),
.B(n_47),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_83),
.B(n_63),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_77),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_46),
.B1(n_19),
.B2(n_14),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_79),
.A2(n_84),
.B1(n_62),
.B2(n_60),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_82),
.B(n_17),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_55),
.A2(n_46),
.B1(n_14),
.B2(n_39),
.Y(n_84)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx13_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_65),
.A2(n_39),
.B1(n_45),
.B2(n_14),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_17),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_0),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_65),
.A2(n_11),
.B(n_9),
.C(n_8),
.Y(n_89)
);

A2O1A1O1Ixp25_ASAP7_75t_L g94 ( 
.A1(n_89),
.A2(n_52),
.B(n_58),
.C(n_64),
.D(n_11),
.Y(n_94)
);

CKINVDCx12_ASAP7_75t_R g90 ( 
.A(n_48),
.Y(n_90)
);

CKINVDCx12_ASAP7_75t_R g107 ( 
.A(n_90),
.Y(n_107)
);

BUFx5_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_93),
.B1(n_83),
.B2(n_81),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_94),
.A2(n_95),
.B(n_108),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_99),
.Y(n_117)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_70),
.Y(n_97)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_106),
.C(n_82),
.Y(n_127)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_71),
.B(n_61),
.Y(n_100)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_100),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_71),
.B(n_61),
.Y(n_102)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_102),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_17),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_0),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_109),
.A2(n_112),
.B1(n_113),
.B2(n_78),
.Y(n_119)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_80),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_7),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_111),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_2),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_2),
.Y(n_113)
);

NOR3xp33_ASAP7_75t_SL g114 ( 
.A(n_89),
.B(n_7),
.C(n_8),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_9),
.B(n_86),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_116),
.B(n_136),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_119),
.B(n_125),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_99),
.A2(n_81),
.B1(n_73),
.B2(n_87),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_132),
.B1(n_93),
.B2(n_97),
.Y(n_146)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_68),
.C(n_81),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_127),
.C(n_2),
.Y(n_153)
);

OA21x2_ASAP7_75t_L g123 ( 
.A1(n_100),
.A2(n_85),
.B(n_80),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_130),
.B(n_113),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_103),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_126),
.Y(n_139)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_102),
.A2(n_85),
.B(n_80),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_103),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_131),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_95),
.A2(n_70),
.B1(n_77),
.B2(n_76),
.Y(n_132)
);

AOI32xp33_ASAP7_75t_L g134 ( 
.A1(n_96),
.A2(n_86),
.A3(n_70),
.B1(n_76),
.B2(n_7),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_134),
.A2(n_104),
.B(n_114),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_107),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_137),
.B(n_91),
.Y(n_143)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_132),
.Y(n_138)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_141),
.A2(n_142),
.B1(n_146),
.B2(n_148),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_143),
.Y(n_161)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_145),
.A2(n_149),
.B1(n_115),
.B2(n_124),
.Y(n_170)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

INVx4_ASAP7_75t_SL g167 ( 
.A(n_147),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_94),
.B1(n_108),
.B2(n_101),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_109),
.B(n_112),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_101),
.B(n_110),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_150),
.A2(n_151),
.B1(n_152),
.B2(n_155),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_123),
.A2(n_101),
.B(n_106),
.Y(n_151)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_120),
.A2(n_128),
.A3(n_116),
.B1(n_122),
.B2(n_130),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_153),
.B(n_135),
.Y(n_160)
);

AOI21x1_ASAP7_75t_L g154 ( 
.A1(n_130),
.A2(n_2),
.B(n_3),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_154),
.B(n_133),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_120),
.A2(n_5),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_L g158 ( 
.A(n_152),
.B(n_135),
.Y(n_158)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_150),
.C(n_154),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_127),
.C(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_159),
.B(n_166),
.C(n_169),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_160),
.B(n_165),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_144),
.A2(n_129),
.B1(n_133),
.B2(n_136),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_162),
.A2(n_170),
.B1(n_148),
.B2(n_142),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_156),
.B(n_125),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_129),
.Y(n_166)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_155),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_151),
.B(n_125),
.C(n_118),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_171),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_139),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_172),
.B(n_174),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_140),
.Y(n_173)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_173),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_140),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_176),
.A2(n_157),
.B1(n_164),
.B2(n_138),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_177),
.A2(n_181),
.B1(n_147),
.B2(n_143),
.Y(n_191)
);

BUFx12_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_178),
.B(n_160),
.C(n_165),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_180),
.B(n_141),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_139),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_183),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g183 ( 
.A(n_175),
.B(n_169),
.C(n_159),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_177),
.A2(n_145),
.B1(n_167),
.B2(n_146),
.Y(n_186)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_186),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_188),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_179),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_178),
.B(n_4),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_184),
.B(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_196),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_190),
.A2(n_179),
.B(n_124),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_197),
.B(n_198),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_190),
.B(n_3),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_199),
.B(n_187),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_183),
.C(n_188),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_197),
.B(n_185),
.Y(n_202)
);

NOR2xp67_ASAP7_75t_SL g206 ( 
.A(n_203),
.B(n_204),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_195),
.A2(n_189),
.B1(n_178),
.B2(n_5),
.Y(n_204)
);

NOR2xp67_ASAP7_75t_L g207 ( 
.A(n_205),
.B(n_194),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_207),
.B(n_209),
.Y(n_210)
);

NOR3xp33_ASAP7_75t_SL g209 ( 
.A(n_203),
.B(n_192),
.C(n_4),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_208),
.B(n_200),
.C(n_201),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_211),
.B(n_206),
.Y(n_213)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_213),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_214),
.B(n_3),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_215),
.B(n_5),
.Y(n_216)
);


endmodule