module fake_jpeg_31572_n_219 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_219);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_219;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_2),
.B(n_8),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_33),
.B(n_35),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_17),
.B(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx11_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_17),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_45),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_0),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_18),
.B(n_1),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_48),
.Y(n_76)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_18),
.B(n_12),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_49),
.B(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_44),
.A2(n_28),
.B1(n_14),
.B2(n_21),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_53),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_47),
.A2(n_28),
.B1(n_14),
.B2(n_23),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_36),
.A2(n_28),
.B1(n_29),
.B2(n_27),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_56),
.A2(n_72),
.B1(n_73),
.B2(n_77),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_33),
.B(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_58),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_39),
.A2(n_23),
.B1(n_30),
.B2(n_20),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_39),
.A2(n_23),
.B1(n_30),
.B2(n_20),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_65),
.Y(n_102)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_36),
.A2(n_27),
.B1(n_19),
.B2(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_37),
.A2(n_16),
.B1(n_15),
.B2(n_24),
.Y(n_73)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_SL g104 ( 
.A(n_75),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_37),
.A2(n_24),
.B1(n_26),
.B2(n_3),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_39),
.A2(n_24),
.B1(n_26),
.B2(n_4),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_84),
.B1(n_91),
.B2(n_88),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_50),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_81),
.Y(n_107)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_51),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_82),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_26),
.B1(n_2),
.B2(n_4),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_85),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_42),
.B(n_1),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g88 ( 
.A1(n_49),
.A2(n_26),
.B1(n_2),
.B2(n_5),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g100 ( 
.A1(n_88),
.A2(n_34),
.B(n_10),
.C(n_11),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_34),
.B(n_1),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_90),
.B(n_70),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_34),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_93),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_78),
.Y(n_93)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_85),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_97),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_9),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_100),
.A2(n_101),
.B1(n_104),
.B2(n_92),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_69),
.A2(n_88),
.B1(n_67),
.B2(n_82),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_89),
.B(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_108),
.A2(n_67),
.B1(n_54),
.B2(n_78),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_61),
.B(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_70),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_113),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_54),
.B(n_75),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_104),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_58),
.B(n_65),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_68),
.B(n_63),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_120),
.A2(n_126),
.B1(n_128),
.B2(n_143),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_63),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_96),
.A2(n_74),
.B1(n_83),
.B2(n_66),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_112),
.A2(n_59),
.B1(n_62),
.B2(n_83),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_105),
.B(n_79),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_127),
.B(n_138),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_112),
.A2(n_62),
.B1(n_74),
.B2(n_79),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_136),
.B1(n_139),
.B2(n_124),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_100),
.A2(n_95),
.B(n_113),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_100),
.A2(n_93),
.B(n_117),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_114),
.B1(n_104),
.B2(n_102),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_118),
.Y(n_137)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_137),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_139),
.B(n_142),
.Y(n_148)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_111),
.A2(n_98),
.B(n_102),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_107),
.Y(n_153)
);

NOR3xp33_ASAP7_75t_SL g142 ( 
.A(n_114),
.B(n_116),
.C(n_94),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_116),
.A2(n_103),
.B1(n_114),
.B2(n_107),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_121),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_149),
.B(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_121),
.B(n_137),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_154),
.B(n_158),
.Y(n_176)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_129),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_159),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_142),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_157),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_123),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_132),
.B(n_133),
.Y(n_159)
);

AO22x1_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_142),
.B1(n_141),
.B2(n_128),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_160),
.A2(n_120),
.B(n_126),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_133),
.B(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_162),
.B(n_122),
.Y(n_172)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_151),
.Y(n_165)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_165),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_125),
.C(n_119),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_170),
.C(n_146),
.Y(n_189)
);

OR2x2_ASAP7_75t_L g167 ( 
.A(n_148),
.B(n_119),
.Y(n_167)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_175),
.B1(n_157),
.B2(n_153),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_138),
.C(n_129),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_172),
.B(n_173),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_150),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_145),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_174),
.B(n_145),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_131),
.B1(n_140),
.B2(n_122),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_178),
.A2(n_160),
.B1(n_152),
.B2(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_177),
.Y(n_180)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_180),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_171),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_184),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_176),
.B(n_158),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_186),
.B(n_190),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_147),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_189),
.B(n_166),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_167),
.B1(n_146),
.B2(n_168),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_147),
.C(n_170),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_167),
.B(n_177),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_198),
.B(n_185),
.Y(n_203)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_191),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_200),
.B(n_201),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_195),
.B(n_188),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_192),
.A2(n_186),
.B1(n_175),
.B2(n_187),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_195),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_196),
.A2(n_183),
.B1(n_168),
.B2(n_149),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_194),
.B(n_197),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_205),
.B(n_208),
.Y(n_213)
);

NAND3xp33_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_198),
.C(n_164),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_206),
.A2(n_169),
.B(n_181),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_209),
.B(n_169),
.Y(n_211)
);

OAI221xp5_ASAP7_75t_L g210 ( 
.A1(n_206),
.A2(n_181),
.B1(n_201),
.B2(n_144),
.C(n_155),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_210),
.A2(n_212),
.B1(n_161),
.B2(n_144),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_211),
.B(n_207),
.C(n_163),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_214),
.B(n_215),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_214),
.A2(n_213),
.B(n_151),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g218 ( 
.A1(n_216),
.A2(n_163),
.B(n_131),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_218),
.B(n_217),
.Y(n_219)
);


endmodule