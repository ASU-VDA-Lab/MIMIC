module real_aes_9099_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_537;
wire n_551;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_310;
wire n_504;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g462 ( .A1(n_0), .A2(n_142), .B(n_463), .C(n_466), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_1), .B(n_457), .Y(n_468) );
INVx1_ASAP7_75t_L g109 ( .A(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g180 ( .A(n_3), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_4), .B(n_143), .Y(n_540) );
OAI22xp5_ASAP7_75t_SL g120 ( .A1(n_5), .A2(n_121), .B1(n_122), .B2(n_428), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g428 ( .A(n_5), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g737 ( .A1(n_5), .A2(n_94), .B1(n_428), .B2(n_738), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_6), .A2(n_442), .B(n_489), .Y(n_488) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_7), .A2(n_149), .B(n_520), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g211 ( .A1(n_8), .A2(n_36), .B1(n_146), .B2(n_198), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_9), .B(n_149), .Y(n_166) );
AND2x6_ASAP7_75t_L g151 ( .A(n_10), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_11), .A2(n_151), .B(n_445), .C(n_513), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g110 ( .A(n_12), .B(n_38), .Y(n_110) );
INVx1_ASAP7_75t_L g133 ( .A(n_13), .Y(n_133) );
INVx1_ASAP7_75t_L g172 ( .A(n_14), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_15), .B(n_139), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g525 ( .A(n_16), .B(n_143), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g128 ( .A(n_17), .B(n_129), .Y(n_128) );
AO32x2_ASAP7_75t_L g209 ( .A1(n_18), .A2(n_149), .A3(n_150), .B1(n_169), .B2(n_210), .Y(n_209) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_19), .B(n_146), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_20), .B(n_129), .Y(n_182) );
AOI22xp33_ASAP7_75t_L g212 ( .A1(n_21), .A2(n_54), .B1(n_146), .B2(n_198), .Y(n_212) );
AOI22xp33_ASAP7_75t_SL g206 ( .A1(n_22), .A2(n_79), .B1(n_139), .B2(n_146), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_23), .B(n_146), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g444 ( .A1(n_24), .A2(n_150), .B(n_445), .C(n_447), .Y(n_444) );
A2O1A1Ixp33_ASAP7_75t_L g522 ( .A1(n_25), .A2(n_150), .B(n_445), .C(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_26), .Y(n_137) );
OAI22xp5_ASAP7_75t_L g115 ( .A1(n_27), .A2(n_95), .B1(n_116), .B2(n_117), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_27), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_28), .B(n_188), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_29), .A2(n_442), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_30), .B(n_188), .Y(n_225) );
INVx2_ASAP7_75t_L g141 ( .A(n_31), .Y(n_141) );
A2O1A1Ixp33_ASAP7_75t_L g476 ( .A1(n_32), .A2(n_477), .B(n_478), .C(n_482), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_33), .B(n_146), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_34), .B(n_188), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_35), .B(n_194), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_37), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_39), .B(n_441), .Y(n_440) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_40), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_41), .B(n_143), .Y(n_504) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_42), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_43), .B(n_442), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g501 ( .A1(n_44), .A2(n_477), .B(n_482), .C(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_45), .B(n_146), .Y(n_159) );
INVx1_ASAP7_75t_L g464 ( .A(n_46), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g101 ( .A1(n_47), .A2(n_102), .B1(n_114), .B2(n_725), .C(n_731), .Y(n_101) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_47), .A2(n_736), .B1(n_739), .B2(n_740), .Y(n_735) );
INVx1_ASAP7_75t_L g740 ( .A(n_47), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g204 ( .A1(n_48), .A2(n_88), .B1(n_198), .B2(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g503 ( .A(n_49), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_50), .B(n_146), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_51), .B(n_146), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_52), .B(n_442), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_53), .B(n_164), .Y(n_163) );
AOI22xp33_ASAP7_75t_SL g145 ( .A1(n_55), .A2(n_59), .B1(n_139), .B2(n_146), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_56), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_57), .B(n_146), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g245 ( .A(n_58), .B(n_146), .Y(n_245) );
INVx1_ASAP7_75t_L g152 ( .A(n_60), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_61), .B(n_442), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_62), .B(n_457), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g491 ( .A1(n_63), .A2(n_164), .B(n_175), .C(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_64), .B(n_146), .Y(n_181) );
INVx1_ASAP7_75t_L g132 ( .A(n_65), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_66), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g480 ( .A(n_67), .B(n_143), .Y(n_480) );
AO32x2_ASAP7_75t_L g202 ( .A1(n_68), .A2(n_149), .A3(n_150), .B1(n_203), .B2(n_207), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_69), .B(n_144), .Y(n_514) );
INVx1_ASAP7_75t_L g244 ( .A(n_70), .Y(n_244) );
INVx1_ASAP7_75t_L g220 ( .A(n_71), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g460 ( .A(n_72), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_73), .B(n_449), .Y(n_448) );
A2O1A1Ixp33_ASAP7_75t_L g537 ( .A1(n_74), .A2(n_445), .B(n_482), .C(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_75), .B(n_139), .Y(n_221) );
CKINVDCx16_ASAP7_75t_R g490 ( .A(n_76), .Y(n_490) );
INVx1_ASAP7_75t_L g113 ( .A(n_77), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g450 ( .A(n_78), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_80), .B(n_198), .Y(n_197) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_81), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_82), .B(n_139), .Y(n_224) );
INVx2_ASAP7_75t_L g130 ( .A(n_83), .Y(n_130) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_84), .Y(n_544) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_85), .B(n_136), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_86), .B(n_139), .Y(n_160) );
OR2x2_ASAP7_75t_L g106 ( .A(n_87), .B(n_107), .Y(n_106) );
OR2x2_ASAP7_75t_L g431 ( .A(n_87), .B(n_108), .Y(n_431) );
INVx2_ASAP7_75t_L g717 ( .A(n_87), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g138 ( .A1(n_89), .A2(n_100), .B1(n_139), .B2(n_140), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_90), .B(n_442), .Y(n_475) );
INVx1_ASAP7_75t_L g479 ( .A(n_91), .Y(n_479) );
INVxp67_ASAP7_75t_L g493 ( .A(n_92), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_93), .B(n_139), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_94), .Y(n_738) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_95), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_96), .B(n_113), .Y(n_112) );
INVx1_ASAP7_75t_L g510 ( .A(n_97), .Y(n_510) );
INVx1_ASAP7_75t_L g539 ( .A(n_98), .Y(n_539) );
AND2x2_ASAP7_75t_L g505 ( .A(n_99), .B(n_188), .Y(n_505) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
OA21x2_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_105), .B(n_111), .Y(n_103) );
NOR2xp33_ASAP7_75t_SL g728 ( .A(n_104), .B(n_112), .Y(n_728) );
INVx1_ASAP7_75t_L g749 ( .A(n_104), .Y(n_749) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx1_ASAP7_75t_SL g730 ( .A(n_106), .Y(n_730) );
INVx1_ASAP7_75t_SL g734 ( .A(n_106), .Y(n_734) );
INVx2_ASAP7_75t_L g745 ( .A(n_106), .Y(n_745) );
NOR2x2_ASAP7_75t_L g724 ( .A(n_107), .B(n_717), .Y(n_724) );
INVx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g716 ( .A(n_108), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x2_ASAP7_75t_L g747 ( .A(n_111), .B(n_748), .Y(n_747) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
OAI222xp33_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_118), .B1(n_718), .B2(n_719), .C1(n_722), .C2(n_723), .Y(n_114) );
INVx1_ASAP7_75t_L g718 ( .A(n_115), .Y(n_718) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI22xp5_ASAP7_75t_SL g119 ( .A1(n_120), .A2(n_429), .B1(n_432), .B2(n_714), .Y(n_119) );
INVx1_ASAP7_75t_L g721 ( .A(n_120), .Y(n_721) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
XNOR2xp5_ASAP7_75t_L g736 ( .A(n_122), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_SL g122 ( .A(n_123), .B(n_362), .Y(n_122) );
NOR5xp2_ASAP7_75t_L g123 ( .A(n_124), .B(n_275), .C(n_321), .D(n_334), .E(n_346), .Y(n_123) );
OAI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_183), .B(n_229), .C(n_256), .Y(n_124) );
INVx1_ASAP7_75t_SL g357 ( .A(n_125), .Y(n_357) );
OR2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_153), .Y(n_125) );
AND2x2_ASAP7_75t_L g281 ( .A(n_126), .B(n_154), .Y(n_281) );
AND2x2_ASAP7_75t_L g309 ( .A(n_126), .B(n_255), .Y(n_309) );
AND2x2_ASAP7_75t_L g317 ( .A(n_126), .B(n_260), .Y(n_317) );
INVx3_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g247 ( .A(n_127), .B(n_155), .Y(n_247) );
INVx2_ASAP7_75t_L g259 ( .A(n_127), .Y(n_259) );
AND2x2_ASAP7_75t_L g384 ( .A(n_127), .B(n_326), .Y(n_384) );
OR2x2_ASAP7_75t_L g386 ( .A(n_127), .B(n_387), .Y(n_386) );
AND2x4_ASAP7_75t_L g127 ( .A(n_128), .B(n_134), .Y(n_127) );
INVx1_ASAP7_75t_L g253 ( .A(n_128), .Y(n_253) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_129), .Y(n_149) );
INVx1_ASAP7_75t_L g169 ( .A(n_129), .Y(n_169) );
AND2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g188 ( .A(n_130), .B(n_131), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g131 ( .A(n_132), .B(n_133), .Y(n_131) );
NAND3xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_148), .C(n_150), .Y(n_134) );
AO21x1_ASAP7_75t_L g252 ( .A1(n_135), .A2(n_148), .B(n_253), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_138), .B1(n_142), .B2(n_145), .Y(n_135) );
INVx2_ASAP7_75t_L g199 ( .A(n_136), .Y(n_199) );
OAI22xp5_ASAP7_75t_SL g203 ( .A1(n_136), .A2(n_144), .B1(n_204), .B2(n_206), .Y(n_203) );
OAI22xp5_ASAP7_75t_L g210 ( .A1(n_136), .A2(n_142), .B1(n_211), .B2(n_212), .Y(n_210) );
INVx4_ASAP7_75t_L g465 ( .A(n_136), .Y(n_465) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx3_ASAP7_75t_L g144 ( .A(n_137), .Y(n_144) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_137), .Y(n_177) );
INVx1_ASAP7_75t_L g194 ( .A(n_137), .Y(n_194) );
AND2x2_ASAP7_75t_L g443 ( .A(n_137), .B(n_165), .Y(n_443) );
INVx1_ASAP7_75t_L g446 ( .A(n_137), .Y(n_446) );
INVx2_ASAP7_75t_L g173 ( .A(n_139), .Y(n_173) );
INVx3_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g147 ( .A(n_141), .Y(n_147) );
INVx1_ASAP7_75t_L g165 ( .A(n_141), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_142), .A2(n_162), .B(n_163), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g178 ( .A1(n_142), .A2(n_179), .B(n_180), .C(n_181), .Y(n_178) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_143), .A2(n_159), .B(n_160), .Y(n_158) );
O2A1O1Ixp5_ASAP7_75t_SL g218 ( .A1(n_143), .A2(n_219), .B(n_220), .C(n_221), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_143), .A2(n_241), .B(n_242), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g492 ( .A(n_143), .B(n_493), .Y(n_492) );
INVx5_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx3_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_146), .Y(n_541) );
BUFx6f_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g198 ( .A(n_147), .Y(n_198) );
BUFx3_ASAP7_75t_L g205 ( .A(n_147), .Y(n_205) );
AND2x6_ASAP7_75t_L g445 ( .A(n_147), .B(n_446), .Y(n_445) );
INVx3_ASAP7_75t_L g457 ( .A(n_148), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_148), .B(n_484), .Y(n_483) );
AO21x2_ASAP7_75t_L g508 ( .A1(n_148), .A2(n_509), .B(n_516), .Y(n_508) );
AO21x2_ASAP7_75t_L g535 ( .A1(n_148), .A2(n_536), .B(n_543), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g543 ( .A(n_148), .B(n_544), .Y(n_543) );
INVx4_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_149), .A2(n_157), .B(n_166), .Y(n_156) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_149), .Y(n_487) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_149), .A2(n_521), .B(n_522), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g239 ( .A1(n_150), .A2(n_240), .B(n_243), .Y(n_239) );
BUFx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI21xp5_ASAP7_75t_L g157 ( .A1(n_151), .A2(n_158), .B(n_161), .Y(n_157) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_151), .A2(n_171), .B(n_178), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g189 ( .A1(n_151), .A2(n_190), .B(n_195), .Y(n_189) );
OAI21xp5_ASAP7_75t_L g217 ( .A1(n_151), .A2(n_218), .B(n_222), .Y(n_217) );
AND2x4_ASAP7_75t_L g442 ( .A(n_151), .B(n_443), .Y(n_442) );
INVx4_ASAP7_75t_SL g467 ( .A(n_151), .Y(n_467) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_151), .B(n_443), .Y(n_511) );
INVx2_ASAP7_75t_SL g153 ( .A(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g297 ( .A(n_154), .B(n_269), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_154), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g411 ( .A(n_154), .B(n_251), .Y(n_411) );
AND2x2_ASAP7_75t_L g154 ( .A(n_155), .B(n_167), .Y(n_154) );
AND2x2_ASAP7_75t_L g254 ( .A(n_155), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g301 ( .A(n_155), .Y(n_301) );
AND2x2_ASAP7_75t_L g326 ( .A(n_155), .B(n_238), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_155), .B(n_359), .Y(n_396) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x2_ASAP7_75t_L g260 ( .A(n_156), .B(n_238), .Y(n_260) );
AND2x2_ASAP7_75t_L g274 ( .A(n_156), .B(n_237), .Y(n_274) );
AND2x2_ASAP7_75t_L g291 ( .A(n_156), .B(n_167), .Y(n_291) );
AND2x2_ASAP7_75t_L g348 ( .A(n_156), .B(n_349), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_156), .B(n_255), .Y(n_361) );
AND2x2_ASAP7_75t_L g413 ( .A(n_156), .B(n_338), .Y(n_413) );
INVx2_ASAP7_75t_L g179 ( .A(n_164), .Y(n_179) );
INVx1_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g236 ( .A(n_167), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g255 ( .A(n_167), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_167), .B(n_238), .Y(n_332) );
OA21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B(n_182), .Y(n_167) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_168), .A2(n_239), .B(n_246), .Y(n_238) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g516 ( .A(n_169), .B(n_517), .Y(n_516) );
O2A1O1Ixp33_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_173), .B(n_174), .C(n_175), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_173), .A2(n_514), .B(n_515), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_173), .A2(n_524), .B(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g538 ( .A1(n_175), .A2(n_539), .B(n_540), .C(n_541), .Y(n_538) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_176), .A2(n_223), .B(n_224), .Y(n_222) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g449 ( .A(n_177), .Y(n_449) );
O2A1O1Ixp5_ASAP7_75t_L g243 ( .A1(n_179), .A2(n_199), .B(n_244), .C(n_245), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_179), .A2(n_448), .B(n_450), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_213), .B(n_226), .Y(n_183) );
INVx1_ASAP7_75t_SL g345 ( .A(n_184), .Y(n_345) );
AND2x4_ASAP7_75t_L g184 ( .A(n_185), .B(n_201), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
AND2x2_ASAP7_75t_SL g233 ( .A(n_186), .B(n_234), .Y(n_233) );
INVx1_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g228 ( .A(n_187), .Y(n_228) );
INVx1_ASAP7_75t_L g265 ( .A(n_187), .Y(n_265) );
AND2x2_ASAP7_75t_L g286 ( .A(n_187), .B(n_208), .Y(n_286) );
AND2x2_ASAP7_75t_L g320 ( .A(n_187), .B(n_209), .Y(n_320) );
OR2x2_ASAP7_75t_L g339 ( .A(n_187), .B(n_215), .Y(n_339) );
HB1xp67_ASAP7_75t_L g353 ( .A(n_187), .Y(n_353) );
AND2x2_ASAP7_75t_L g366 ( .A(n_187), .B(n_367), .Y(n_366) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_189), .B(n_200), .Y(n_187) );
INVx2_ASAP7_75t_L g207 ( .A(n_188), .Y(n_207) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_188), .A2(n_217), .B(n_225), .Y(n_216) );
INVx1_ASAP7_75t_L g455 ( .A(n_188), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_188), .A2(n_475), .B(n_476), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_188), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
INVx1_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B(n_199), .Y(n_195) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_201), .A2(n_288), .B1(n_289), .B2(n_298), .Y(n_287) );
AND2x2_ASAP7_75t_L g371 ( .A(n_201), .B(n_372), .Y(n_371) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_208), .Y(n_201) );
INVx1_ASAP7_75t_L g232 ( .A(n_202), .Y(n_232) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
INVx1_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
AND2x2_ASAP7_75t_L g295 ( .A(n_202), .B(n_209), .Y(n_295) );
INVx2_ASAP7_75t_L g466 ( .A(n_205), .Y(n_466) );
HB1xp67_ASAP7_75t_L g481 ( .A(n_205), .Y(n_481) );
INVx1_ASAP7_75t_L g452 ( .A(n_207), .Y(n_452) );
OR2x2_ASAP7_75t_L g249 ( .A(n_208), .B(n_234), .Y(n_249) );
AND2x2_ASAP7_75t_L g279 ( .A(n_208), .B(n_280), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g367 ( .A(n_208), .B(n_368), .Y(n_367) );
INVx2_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g227 ( .A(n_209), .B(n_228), .Y(n_227) );
BUFx2_ASAP7_75t_L g336 ( .A(n_209), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_213), .B(n_352), .Y(n_351) );
BUFx2_ASAP7_75t_L g213 ( .A(n_214), .Y(n_213) );
AND2x2_ASAP7_75t_L g314 ( .A(n_214), .B(n_280), .Y(n_314) );
INVx2_ASAP7_75t_L g214 ( .A(n_215), .Y(n_214) );
AND2x2_ASAP7_75t_L g226 ( .A(n_215), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g285 ( .A(n_215), .Y(n_285) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g234 ( .A(n_216), .Y(n_234) );
OR2x2_ASAP7_75t_L g264 ( .A(n_216), .B(n_265), .Y(n_264) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_216), .Y(n_319) );
AOI32xp33_ASAP7_75t_L g356 ( .A1(n_226), .A2(n_286), .A3(n_357), .B1(n_358), .B2(n_360), .Y(n_356) );
AND2x2_ASAP7_75t_L g282 ( .A(n_227), .B(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_227), .B(n_381), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_227), .B(n_314), .Y(n_400) );
INVx1_ASAP7_75t_L g405 ( .A(n_227), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_235), .B1(n_248), .B2(n_250), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_231), .B(n_233), .Y(n_230) );
AND2x2_ASAP7_75t_L g335 ( .A(n_231), .B(n_336), .Y(n_335) );
HB1xp67_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_232), .B(n_234), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_233), .A2(n_257), .B1(n_261), .B2(n_271), .Y(n_256) );
AND2x2_ASAP7_75t_L g278 ( .A(n_233), .B(n_279), .Y(n_278) );
A2O1A1Ixp33_ASAP7_75t_L g329 ( .A1(n_233), .A2(n_247), .B(n_295), .C(n_330), .Y(n_329) );
OAI332xp33_ASAP7_75t_L g334 ( .A1(n_233), .A2(n_335), .A3(n_337), .B1(n_339), .B2(n_340), .B3(n_342), .C1(n_343), .C2(n_345), .Y(n_334) );
INVx2_ASAP7_75t_L g375 ( .A(n_233), .Y(n_375) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_234), .Y(n_293) );
INVx1_ASAP7_75t_L g368 ( .A(n_234), .Y(n_368) );
AND2x2_ASAP7_75t_L g422 ( .A(n_234), .B(n_286), .Y(n_422) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_247), .Y(n_235) );
AND2x2_ASAP7_75t_L g302 ( .A(n_237), .B(n_252), .Y(n_302) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g251 ( .A(n_238), .B(n_252), .Y(n_251) );
OR2x2_ASAP7_75t_L g350 ( .A(n_238), .B(n_252), .Y(n_350) );
INVx1_ASAP7_75t_L g359 ( .A(n_238), .Y(n_359) );
INVx1_ASAP7_75t_L g333 ( .A(n_247), .Y(n_333) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g417 ( .A(n_249), .B(n_269), .Y(n_417) );
INVx1_ASAP7_75t_SL g328 ( .A(n_250), .Y(n_328) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
AND2x2_ASAP7_75t_L g355 ( .A(n_251), .B(n_313), .Y(n_355) );
INVx1_ASAP7_75t_L g374 ( .A(n_251), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g376 ( .A(n_251), .B(n_341), .Y(n_376) );
INVx1_ASAP7_75t_L g273 ( .A(n_252), .Y(n_273) );
AND2x2_ASAP7_75t_L g277 ( .A(n_254), .B(n_258), .Y(n_277) );
AND2x2_ASAP7_75t_L g344 ( .A(n_254), .B(n_302), .Y(n_344) );
INVx2_ASAP7_75t_L g387 ( .A(n_254), .Y(n_387) );
INVx2_ASAP7_75t_L g270 ( .A(n_255), .Y(n_270) );
AND2x2_ASAP7_75t_L g272 ( .A(n_255), .B(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
INVx1_ASAP7_75t_L g288 ( .A(n_258), .Y(n_288) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
NOR2xp33_ASAP7_75t_L g338 ( .A(n_259), .B(n_332), .Y(n_338) );
OR2x2_ASAP7_75t_L g402 ( .A(n_259), .B(n_361), .Y(n_402) );
INVx1_ASAP7_75t_L g426 ( .A(n_259), .Y(n_426) );
INVx1_ASAP7_75t_L g382 ( .A(n_260), .Y(n_382) );
AND2x2_ASAP7_75t_L g427 ( .A(n_260), .B(n_270), .Y(n_427) );
INVx1_ASAP7_75t_L g261 ( .A(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_266), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_264), .A2(n_290), .B1(n_292), .B2(n_296), .Y(n_289) );
INVx1_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OAI322xp33_ASAP7_75t_SL g373 ( .A1(n_267), .A2(n_374), .A3(n_375), .B1(n_376), .B2(n_377), .C1(n_380), .C2(n_382), .Y(n_373) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_270), .Y(n_267) );
AND2x2_ASAP7_75t_L g370 ( .A(n_268), .B(n_286), .Y(n_370) );
OR2x2_ASAP7_75t_L g404 ( .A(n_268), .B(n_405), .Y(n_404) );
OR2x2_ASAP7_75t_L g407 ( .A(n_268), .B(n_339), .Y(n_407) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g352 ( .A(n_269), .B(n_353), .Y(n_352) );
OR2x2_ASAP7_75t_L g408 ( .A(n_269), .B(n_339), .Y(n_408) );
INVx3_ASAP7_75t_L g341 ( .A(n_270), .Y(n_341) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g397 ( .A(n_272), .Y(n_397) );
AOI222xp33_ASAP7_75t_L g276 ( .A1(n_274), .A2(n_277), .B1(n_278), .B2(n_281), .C1(n_282), .C2(n_284), .Y(n_276) );
INVx1_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
NAND3xp33_ASAP7_75t_SL g275 ( .A(n_276), .B(n_287), .C(n_304), .Y(n_275) );
AND2x2_ASAP7_75t_L g392 ( .A(n_279), .B(n_293), .Y(n_392) );
BUFx2_ASAP7_75t_L g283 ( .A(n_280), .Y(n_283) );
INVx1_ASAP7_75t_L g324 ( .A(n_280), .Y(n_324) );
AOI221xp5_ASAP7_75t_L g369 ( .A1(n_281), .A2(n_317), .B1(n_370), .B2(n_371), .C(n_373), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_283), .B(n_366), .Y(n_365) );
AND2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_286), .Y(n_310) );
AND2x2_ASAP7_75t_L g323 ( .A(n_286), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_291), .B(n_302), .Y(n_303) );
OR2x2_ASAP7_75t_L g292 ( .A(n_293), .B(n_294), .Y(n_292) );
OAI21xp33_ASAP7_75t_L g298 ( .A1(n_293), .A2(n_299), .B(n_303), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_293), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_SL g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g390 ( .A(n_295), .B(n_372), .Y(n_390) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g313 ( .A(n_301), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_302), .B(n_313), .Y(n_312) );
INVx2_ASAP7_75t_L g419 ( .A(n_302), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g304 ( .A1(n_305), .A2(n_310), .B1(n_311), .B2(n_314), .C(n_315), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_SL g394 ( .A(n_306), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g306 ( .A(n_307), .B(n_308), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g415 ( .A(n_314), .B(n_320), .Y(n_415) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
OAI31xp33_ASAP7_75t_SL g383 ( .A1(n_318), .A2(n_357), .A3(n_384), .B(n_385), .Y(n_383) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
INVx1_ASAP7_75t_L g372 ( .A(n_319), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g423 ( .A(n_320), .B(n_324), .Y(n_423) );
OAI221xp5_ASAP7_75t_SL g321 ( .A1(n_322), .A2(n_325), .B1(n_327), .B2(n_328), .C(n_329), .Y(n_321) );
INVx1_ASAP7_75t_L g327 ( .A(n_323), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_326), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_332), .B(n_333), .Y(n_331) );
INVx1_ASAP7_75t_L g342 ( .A(n_335), .Y(n_342) );
INVx2_ASAP7_75t_L g378 ( .A(n_336), .Y(n_378) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g364 ( .A(n_341), .B(n_350), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g414 ( .A1(n_341), .A2(n_358), .B(n_415), .C(n_416), .Y(n_414) );
OAI221xp5_ASAP7_75t_SL g346 ( .A1(n_342), .A2(n_347), .B1(n_351), .B2(n_354), .C(n_356), .Y(n_346) );
INVx1_ASAP7_75t_SL g343 ( .A(n_344), .Y(n_343) );
A2O1A1Ixp33_ASAP7_75t_L g409 ( .A1(n_345), .A2(n_410), .B(n_412), .C(n_414), .Y(n_409) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_348), .A2(n_399), .B1(n_401), .B2(n_403), .C(n_406), .Y(n_398) );
INVx1_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
NOR4xp25_ASAP7_75t_L g362 ( .A(n_363), .B(n_388), .C(n_409), .D(n_420), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_365), .B(n_369), .C(n_383), .Y(n_363) );
INVx1_ASAP7_75t_SL g418 ( .A(n_370), .Y(n_418) );
OR2x2_ASAP7_75t_L g377 ( .A(n_378), .B(n_379), .Y(n_377) );
INVx1_ASAP7_75t_SL g381 ( .A(n_379), .Y(n_381) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
OAI22xp5_ASAP7_75t_L g406 ( .A1(n_386), .A2(n_395), .B1(n_407), .B2(n_408), .Y(n_406) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_389), .A2(n_391), .B(n_393), .C(n_398), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI31xp33_ASAP7_75t_L g420 ( .A1(n_391), .A2(n_421), .A3(n_423), .B(n_424), .Y(n_420) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVxp67_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_397), .Y(n_395) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_SL g412 ( .A(n_413), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B(n_419), .Y(n_416) );
INVx1_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_427), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_431), .A2(n_433), .B1(n_716), .B2(n_721), .Y(n_720) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_434), .B(n_650), .Y(n_433) );
NOR5xp2_ASAP7_75t_L g434 ( .A(n_435), .B(n_581), .C(n_610), .D(n_630), .E(n_637), .Y(n_434) );
OAI211xp5_ASAP7_75t_SL g435 ( .A1(n_436), .A2(n_469), .B(n_526), .C(n_568), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g652 ( .A1(n_437), .A2(n_653), .B1(n_655), .B2(n_656), .Y(n_652) );
AND2x2_ASAP7_75t_L g437 ( .A(n_438), .B(n_456), .Y(n_437) );
HB1xp67_ASAP7_75t_L g529 ( .A(n_438), .Y(n_529) );
AND2x4_ASAP7_75t_L g561 ( .A(n_438), .B(n_562), .Y(n_561) );
INVx5_ASAP7_75t_L g579 ( .A(n_438), .Y(n_579) );
AND2x2_ASAP7_75t_L g588 ( .A(n_438), .B(n_580), .Y(n_588) );
AND2x2_ASAP7_75t_L g600 ( .A(n_438), .B(n_473), .Y(n_600) );
AND2x2_ASAP7_75t_L g696 ( .A(n_438), .B(n_564), .Y(n_696) );
OR2x6_ASAP7_75t_L g438 ( .A(n_439), .B(n_453), .Y(n_438) );
AOI21xp5_ASAP7_75t_SL g439 ( .A1(n_440), .A2(n_444), .B(n_452), .Y(n_439) );
BUFx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx5_ASAP7_75t_L g461 ( .A(n_445), .Y(n_461) );
INVx2_ASAP7_75t_L g451 ( .A(n_449), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g478 ( .A1(n_451), .A2(n_479), .B(n_480), .C(n_481), .Y(n_478) );
O2A1O1Ixp33_ASAP7_75t_L g502 ( .A1(n_451), .A2(n_481), .B(n_503), .C(n_504), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
INVx2_ASAP7_75t_L g562 ( .A(n_456), .Y(n_562) );
AND2x2_ASAP7_75t_L g580 ( .A(n_456), .B(n_535), .Y(n_580) );
AND2x2_ASAP7_75t_L g599 ( .A(n_456), .B(n_534), .Y(n_599) );
AND2x2_ASAP7_75t_L g639 ( .A(n_456), .B(n_579), .Y(n_639) );
OA21x2_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_468), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_SL g459 ( .A1(n_460), .A2(n_461), .B(n_462), .C(n_467), .Y(n_459) );
INVx2_ASAP7_75t_L g477 ( .A(n_461), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_L g489 ( .A1(n_461), .A2(n_467), .B(n_490), .C(n_491), .Y(n_489) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_465), .Y(n_463) );
INVx1_ASAP7_75t_L g482 ( .A(n_467), .Y(n_482) );
INVxp67_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_495), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI322xp5_ASAP7_75t_L g698 ( .A1(n_472), .A2(n_506), .A3(n_553), .B1(n_561), .B2(n_615), .C1(n_699), .C2(n_702), .Y(n_698) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_485), .Y(n_472) );
INVx5_ASAP7_75t_L g531 ( .A(n_473), .Y(n_531) );
AND2x2_ASAP7_75t_L g547 ( .A(n_473), .B(n_533), .Y(n_547) );
BUFx2_ASAP7_75t_L g625 ( .A(n_473), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_473), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g702 ( .A(n_473), .B(n_609), .Y(n_702) );
OR2x6_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_485), .B(n_497), .Y(n_556) );
INVx1_ASAP7_75t_L g583 ( .A(n_485), .Y(n_583) );
AND2x2_ASAP7_75t_L g596 ( .A(n_485), .B(n_518), .Y(n_596) );
AND2x2_ASAP7_75t_L g697 ( .A(n_485), .B(n_615), .Y(n_697) );
INVx3_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g551 ( .A(n_486), .B(n_497), .Y(n_551) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_486), .Y(n_559) );
OR2x2_ASAP7_75t_L g566 ( .A(n_486), .B(n_518), .Y(n_566) );
AND2x2_ASAP7_75t_L g576 ( .A(n_486), .B(n_577), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_486), .B(n_508), .Y(n_605) );
INVxp67_ASAP7_75t_L g629 ( .A(n_486), .Y(n_629) );
AND2x2_ASAP7_75t_L g636 ( .A(n_486), .B(n_506), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_486), .B(n_518), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_486), .B(n_507), .Y(n_662) );
OA21x2_ASAP7_75t_L g486 ( .A1(n_487), .A2(n_488), .B(n_494), .Y(n_486) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_497), .B(n_519), .Y(n_606) );
OR2x2_ASAP7_75t_L g628 ( .A(n_497), .B(n_507), .Y(n_628) );
AND2x2_ASAP7_75t_L g641 ( .A(n_497), .B(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_497), .B(n_596), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g651 ( .A1(n_497), .A2(n_652), .B(n_657), .C(n_666), .Y(n_651) );
AND2x2_ASAP7_75t_L g712 ( .A(n_497), .B(n_518), .Y(n_712) );
INVx5_ASAP7_75t_SL g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g565 ( .A(n_498), .B(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_498), .B(n_571), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_498), .B(n_560), .Y(n_572) );
HB1xp67_ASAP7_75t_L g574 ( .A(n_498), .Y(n_574) );
OR2x2_ASAP7_75t_L g585 ( .A(n_498), .B(n_507), .Y(n_585) );
AND2x2_ASAP7_75t_SL g590 ( .A(n_498), .B(n_576), .Y(n_590) );
AND2x2_ASAP7_75t_L g615 ( .A(n_498), .B(n_507), .Y(n_615) );
AND2x2_ASAP7_75t_L g635 ( .A(n_498), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g673 ( .A(n_498), .B(n_506), .Y(n_673) );
OR2x2_ASAP7_75t_L g676 ( .A(n_498), .B(n_662), .Y(n_676) );
OR2x6_ASAP7_75t_L g498 ( .A(n_499), .B(n_505), .Y(n_498) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_518), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_507), .A2(n_620), .B(n_623), .C(n_629), .Y(n_619) );
INVx5_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_508), .B(n_518), .Y(n_550) );
AND2x2_ASAP7_75t_L g554 ( .A(n_508), .B(n_519), .Y(n_554) );
OR2x2_ASAP7_75t_L g560 ( .A(n_508), .B(n_518), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_511), .B(n_512), .Y(n_509) );
INVx1_ASAP7_75t_SL g577 ( .A(n_518), .Y(n_577) );
OR2x2_ASAP7_75t_L g705 ( .A(n_518), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_545), .B(n_548), .C(n_557), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
AOI31xp33_ASAP7_75t_L g630 ( .A1(n_528), .A2(n_631), .A3(n_633), .B(n_634), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_529), .B(n_530), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_529), .B(n_547), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_530), .B(n_561), .Y(n_567) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_531), .B(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g587 ( .A(n_531), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g592 ( .A(n_531), .B(n_562), .Y(n_592) );
AND2x2_ASAP7_75t_L g602 ( .A(n_531), .B(n_561), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_531), .B(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g622 ( .A(n_531), .B(n_579), .Y(n_622) );
AND2x2_ASAP7_75t_L g627 ( .A(n_531), .B(n_599), .Y(n_627) );
OR2x2_ASAP7_75t_L g646 ( .A(n_531), .B(n_533), .Y(n_646) );
OR2x2_ASAP7_75t_L g648 ( .A(n_531), .B(n_649), .Y(n_648) );
HB1xp67_ASAP7_75t_L g695 ( .A(n_531), .Y(n_695) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x2_ASAP7_75t_L g595 ( .A(n_533), .B(n_562), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_533), .B(n_579), .Y(n_618) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx2_ASAP7_75t_L g564 ( .A(n_535), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_542), .Y(n_536) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g655 ( .A(n_547), .B(n_579), .Y(n_655) );
AOI322xp5_ASAP7_75t_L g657 ( .A1(n_547), .A2(n_561), .A3(n_599), .B1(n_658), .B2(n_659), .C1(n_660), .C2(n_663), .Y(n_657) );
INVx1_ASAP7_75t_L g665 ( .A(n_547), .Y(n_665) );
NAND2xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_552), .Y(n_548) );
INVx1_ASAP7_75t_SL g659 ( .A(n_549), .Y(n_659) );
OR2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
OR2x2_ASAP7_75t_L g611 ( .A(n_550), .B(n_556), .Y(n_611) );
INVx1_ASAP7_75t_L g642 ( .A(n_550), .Y(n_642) );
INVx2_ASAP7_75t_SL g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OAI32xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .A3(n_563), .B1(n_565), .B2(n_567), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
AOI21xp33_ASAP7_75t_SL g597 ( .A1(n_560), .A2(n_575), .B(n_598), .Y(n_597) );
INVx1_ASAP7_75t_SL g612 ( .A(n_561), .Y(n_612) );
AND2x4_ASAP7_75t_L g609 ( .A(n_562), .B(n_579), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_562), .B(n_645), .Y(n_644) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_563), .A2(n_590), .A3(n_609), .B1(n_642), .B2(n_675), .C1(n_677), .C2(n_678), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g703 ( .A1(n_563), .A2(n_640), .B1(n_704), .B2(n_705), .C(n_707), .Y(n_703) );
AND2x2_ASAP7_75t_L g591 ( .A(n_564), .B(n_592), .Y(n_591) );
INVx1_ASAP7_75t_SL g571 ( .A(n_566), .Y(n_571) );
OR2x2_ASAP7_75t_L g643 ( .A(n_566), .B(n_628), .Y(n_643) );
OAI31xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_572), .A3(n_573), .B(n_578), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_569), .A2(n_602), .B1(n_603), .B2(n_607), .Y(n_601) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g614 ( .A(n_571), .B(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_573), .A2(n_614), .B1(n_667), .B2(n_670), .Y(n_666) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g656 ( .A(n_576), .B(n_625), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_576), .B(n_615), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_577), .B(n_683), .Y(n_682) );
OR2x2_ASAP7_75t_L g690 ( .A(n_577), .B(n_628), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_578), .A2(n_673), .B1(n_686), .B2(n_689), .Y(n_685) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
INVx2_ASAP7_75t_L g594 ( .A(n_579), .Y(n_594) );
AND2x2_ASAP7_75t_L g677 ( .A(n_579), .B(n_599), .Y(n_677) );
OR2x2_ASAP7_75t_L g679 ( .A(n_579), .B(n_646), .Y(n_679) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_579), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_580), .B(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_580), .B(n_625), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_586), .B(n_589), .C(n_601), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_SL g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_593), .B2(n_596), .C(n_597), .Y(n_589) );
INVxp67_ASAP7_75t_L g701 ( .A(n_592), .Y(n_701) );
INVx1_ASAP7_75t_L g668 ( .A(n_593), .Y(n_668) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g632 ( .A(n_594), .B(n_599), .Y(n_632) );
INVx1_ASAP7_75t_L g649 ( .A(n_595), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_595), .B(n_622), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g664 ( .A(n_599), .Y(n_664) );
AND2x2_ASAP7_75t_L g670 ( .A(n_599), .B(n_625), .Y(n_670) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_SL g658 ( .A(n_606), .Y(n_658) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_609), .B(n_645), .Y(n_669) );
OAI221xp5_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_612), .B1(n_613), .B2(n_616), .C(n_619), .Y(n_610) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g706 ( .A(n_615), .Y(n_706) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OR2x2_ASAP7_75t_L g624 ( .A(n_618), .B(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_622), .B(n_681), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_626), .B(n_628), .Y(n_623) );
OAI211xp5_ASAP7_75t_SL g671 ( .A1(n_626), .A2(n_672), .B(n_674), .C(n_680), .Y(n_671) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g683 ( .A(n_628), .Y(n_683) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
OAI222xp33_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_640), .B1(n_643), .B2(n_644), .C1(n_647), .C2(n_648), .Y(n_637) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
INVx1_ASAP7_75t_L g713 ( .A(n_644), .Y(n_713) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_645), .B(n_688), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_645), .A2(n_692), .B1(n_694), .B2(n_697), .Y(n_691) );
INVx2_ASAP7_75t_SL g645 ( .A(n_646), .Y(n_645) );
NOR4xp25_ASAP7_75t_L g650 ( .A(n_651), .B(n_671), .C(n_684), .D(n_703), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_653), .B(n_683), .Y(n_693) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g660 ( .A(n_658), .B(n_661), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_661), .B(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g661 ( .A(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_664), .B(n_665), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g667 ( .A(n_668), .B(n_669), .Y(n_667) );
INVx1_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g684 ( .A(n_685), .B(n_691), .C(n_698), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx2_ASAP7_75t_L g700 ( .A(n_696), .Y(n_700) );
NOR2xp33_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
OAI21xp5_ASAP7_75t_SL g707 ( .A1(n_708), .A2(n_710), .B(n_713), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
NAND2xp33_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
AOI21xp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_741), .B(n_746), .Y(n_731) );
INVxp33_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_735), .Y(n_733) );
INVx1_ASAP7_75t_L g739 ( .A(n_736), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
endmodule