module fake_jpeg_23264_n_25 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_25);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_25;

wire n_13;
wire n_21;
wire n_23;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_24;
wire n_17;
wire n_12;
wire n_15;

INVx3_ASAP7_75t_SL g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_10),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_SL g15 ( 
.A1(n_11),
.A2(n_0),
.B1(n_3),
.B2(n_6),
.Y(n_15)
);

OAI21xp5_ASAP7_75t_SL g16 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_17),
.C(n_18),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_13),
.B(n_2),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_2),
.B(n_3),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_12),
.B1(n_15),
.B2(n_13),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_19),
.B(n_12),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_18),
.A2(n_12),
.B1(n_5),
.B2(n_7),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g23 ( 
.A(n_21),
.B(n_4),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_22),
.B(n_23),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_24),
.A2(n_20),
.B(n_9),
.Y(n_25)
);


endmodule