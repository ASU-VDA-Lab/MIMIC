module real_aes_5122_n_234 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_234);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_234;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_461;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_856;
wire n_594;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_578;
wire n_372;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_656;
wire n_532;
wire n_316;
wire n_755;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_246;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_269;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_854;
wire n_403;
wire n_877;
wire n_424;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_0), .A2(n_56), .B1(n_426), .B2(n_432), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_1), .A2(n_211), .B1(n_386), .B2(n_387), .Y(n_603) );
AO22x2_ASAP7_75t_L g585 ( .A1(n_2), .A2(n_586), .B1(n_605), .B2(n_606), .Y(n_585) );
INVxp67_ASAP7_75t_SL g605 ( .A(n_2), .Y(n_605) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_3), .Y(n_635) );
AND2x4_ASAP7_75t_L g645 ( .A(n_3), .B(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g651 ( .A(n_3), .B(n_228), .Y(n_651) );
INVx1_ASAP7_75t_L g411 ( .A(n_4), .Y(n_411) );
AO22x1_ASAP7_75t_L g655 ( .A1(n_4), .A2(n_6), .B1(n_656), .B2(n_657), .Y(n_655) );
INVx1_ASAP7_75t_L g473 ( .A(n_5), .Y(n_473) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_7), .A2(n_169), .B1(n_642), .B2(n_662), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_8), .A2(n_180), .B1(n_328), .B2(n_432), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_9), .A2(n_83), .B1(n_386), .B2(n_387), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_10), .A2(n_204), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_11), .A2(n_15), .B1(n_380), .B2(n_381), .Y(n_602) );
AOI22xp5_ASAP7_75t_L g420 ( .A1(n_12), .A2(n_18), .B1(n_421), .B2(n_422), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_13), .A2(n_190), .B1(n_397), .B2(n_421), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_14), .A2(n_66), .B1(n_333), .B2(n_394), .Y(n_393) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_16), .A2(n_102), .B1(n_321), .B2(n_327), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g458 ( .A1(n_17), .A2(n_28), .B1(n_459), .B2(n_461), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_19), .A2(n_24), .B1(n_368), .B2(n_476), .Y(n_475) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_20), .A2(n_133), .B1(n_383), .B2(n_384), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_21), .A2(n_69), .B1(n_350), .B2(n_427), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_22), .A2(n_110), .B1(n_380), .B2(n_381), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_23), .A2(n_116), .B1(n_378), .B2(n_387), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g689 ( .A1(n_25), .A2(n_104), .B1(n_652), .B2(n_690), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_26), .A2(n_105), .B1(n_514), .B2(n_862), .Y(n_861) );
CKINVDCx20_ASAP7_75t_R g484 ( .A(n_27), .Y(n_484) );
AOI221xp5_ASAP7_75t_L g404 ( .A1(n_29), .A2(n_34), .B1(n_405), .B2(n_406), .C(n_409), .Y(n_404) );
INVx1_ASAP7_75t_L g544 ( .A(n_30), .Y(n_544) );
INVx1_ASAP7_75t_L g489 ( .A(n_31), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g501 ( .A1(n_32), .A2(n_93), .B1(n_244), .B2(n_269), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_33), .A2(n_146), .B1(n_383), .B2(n_384), .Y(n_621) );
XNOR2x1_ASAP7_75t_L g536 ( .A(n_35), .B(n_537), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_36), .A2(n_154), .B1(n_332), .B2(n_339), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_37), .A2(n_406), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g518 ( .A(n_38), .Y(n_518) );
INVx1_ASAP7_75t_L g265 ( .A(n_39), .Y(n_265) );
INVxp67_ASAP7_75t_L g305 ( .A(n_39), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_39), .B(n_176), .Y(n_314) );
AOI22xp33_ASAP7_75t_L g391 ( .A1(n_40), .A2(n_135), .B1(n_350), .B2(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_41), .A2(n_71), .B1(n_285), .B2(n_402), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_42), .A2(n_111), .B1(n_365), .B2(n_380), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_43), .A2(n_112), .B1(n_343), .B2(n_345), .Y(n_342) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_44), .A2(n_90), .B1(n_426), .B2(n_427), .Y(n_425) );
XNOR2x1_ASAP7_75t_L g239 ( .A(n_45), .B(n_240), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_46), .B(n_249), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_47), .A2(n_77), .B1(n_853), .B2(n_854), .Y(n_852) );
AOI21xp33_ASAP7_75t_SL g588 ( .A1(n_48), .A2(n_476), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g579 ( .A(n_49), .Y(n_579) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_50), .A2(n_220), .B1(n_368), .B2(n_369), .Y(n_367) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_51), .A2(n_195), .B1(n_366), .B2(n_368), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_52), .A2(n_149), .B1(n_402), .B2(n_865), .Y(n_864) );
BUFx2_ASAP7_75t_L g595 ( .A(n_53), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_54), .A2(n_89), .B1(n_380), .B2(n_381), .Y(n_379) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_55), .A2(n_141), .B1(n_650), .B2(n_657), .Y(n_660) );
INVx1_ASAP7_75t_L g410 ( .A(n_57), .Y(n_410) );
INVx2_ASAP7_75t_L g633 ( .A(n_58), .Y(n_633) );
INVx1_ASAP7_75t_L g644 ( .A(n_59), .Y(n_644) );
AND2x4_ASAP7_75t_L g648 ( .A(n_59), .B(n_633), .Y(n_648) );
INVx1_ASAP7_75t_SL g688 ( .A(n_59), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_60), .A2(n_207), .B1(n_402), .B2(n_476), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_61), .A2(n_132), .B1(n_402), .B2(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_62), .B(n_444), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_63), .A2(n_156), .B1(n_656), .B2(n_680), .Y(n_725) );
AOI22xp33_ASAP7_75t_L g860 ( .A1(n_64), .A2(n_143), .B1(n_437), .B2(n_567), .Y(n_860) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_65), .A2(n_202), .B1(n_366), .B2(n_369), .Y(n_477) );
AOI22xp33_ASAP7_75t_SL g431 ( .A1(n_67), .A2(n_215), .B1(n_328), .B2(n_432), .Y(n_431) );
BUFx6f_ASAP7_75t_L g249 ( .A(n_68), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_70), .A2(n_178), .B1(n_383), .B2(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g559 ( .A(n_72), .Y(n_559) );
INVx1_ASAP7_75t_L g575 ( .A(n_73), .Y(n_575) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_74), .A2(n_166), .B1(n_463), .B2(n_464), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_75), .A2(n_230), .B1(n_381), .B2(n_386), .Y(n_620) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_76), .A2(n_516), .B(n_517), .Y(n_515) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_78), .A2(n_136), .B1(n_642), .B2(n_647), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_79), .A2(n_159), .B1(n_346), .B2(n_856), .Y(n_855) );
AOI22xp5_ASAP7_75t_L g614 ( .A1(n_80), .A2(n_81), .B1(n_369), .B2(n_377), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_82), .A2(n_189), .B1(n_269), .B2(n_441), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_84), .A2(n_130), .B1(n_285), .B2(n_511), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_85), .A2(n_148), .B1(n_656), .B2(n_657), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g669 ( .A1(n_86), .A2(n_167), .B1(n_650), .B2(n_657), .Y(n_669) );
INVx1_ASAP7_75t_L g253 ( .A(n_87), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_87), .B(n_175), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_88), .A2(n_129), .B1(n_328), .B2(n_399), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g676 ( .A1(n_91), .A2(n_140), .B1(n_642), .B2(n_677), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g364 ( .A1(n_92), .A2(n_186), .B1(n_365), .B2(n_366), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_94), .A2(n_97), .B1(n_642), .B2(n_662), .Y(n_667) );
XNOR2x1_ASAP7_75t_L g610 ( .A(n_95), .B(n_611), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_96), .A2(n_158), .B1(n_448), .B2(n_450), .Y(n_447) );
INVx1_ASAP7_75t_L g417 ( .A(n_98), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_99), .A2(n_181), .B1(n_328), .B2(n_430), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_100), .A2(n_179), .B1(n_677), .B2(n_723), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_101), .A2(n_229), .B1(n_377), .B2(n_378), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_103), .A2(n_117), .B1(n_243), .B2(n_268), .Y(n_242) );
XNOR2x1_ASAP7_75t_L g455 ( .A(n_104), .B(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g306 ( .A(n_106), .Y(n_306) );
INVx1_ASAP7_75t_L g590 ( .A(n_107), .Y(n_590) );
INVx1_ASAP7_75t_L g466 ( .A(n_108), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g661 ( .A1(n_109), .A2(n_219), .B1(n_642), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g573 ( .A1(n_113), .A2(n_216), .B1(n_386), .B2(n_387), .Y(n_573) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_114), .A2(n_371), .B(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_115), .A2(n_205), .B1(n_383), .B2(n_384), .Y(n_569) );
INVx1_ASAP7_75t_L g546 ( .A(n_118), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_119), .A2(n_163), .B1(n_494), .B2(n_495), .Y(n_493) );
INVx1_ASAP7_75t_L g618 ( .A(n_120), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_121), .A2(n_227), .B1(n_377), .B2(n_378), .Y(n_480) );
AOI22xp33_ASAP7_75t_SL g599 ( .A1(n_122), .A2(n_203), .B1(n_369), .B2(n_468), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_123), .A2(n_124), .B1(n_285), .B2(n_500), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_125), .A2(n_126), .B1(n_350), .B2(n_552), .Y(n_551) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_127), .A2(n_153), .B1(n_541), .B2(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_128), .A2(n_218), .B1(n_662), .B2(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_131), .B(n_592), .Y(n_613) );
AOI22xp33_ASAP7_75t_L g348 ( .A1(n_134), .A2(n_161), .B1(n_349), .B2(n_352), .Y(n_348) );
INVx1_ASAP7_75t_L g359 ( .A(n_137), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g649 ( .A1(n_137), .A2(n_183), .B1(n_650), .B2(n_652), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_138), .A2(n_191), .B1(n_340), .B2(n_463), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_139), .B(n_491), .Y(n_866) );
XOR2xp5_ASAP7_75t_L g507 ( .A(n_142), .B(n_508), .Y(n_507) );
AOI22xp33_ASAP7_75t_L g278 ( .A1(n_144), .A2(n_164), .B1(n_279), .B2(n_283), .Y(n_278) );
AOI22xp5_ASAP7_75t_L g497 ( .A1(n_145), .A2(n_209), .B1(n_333), .B2(n_432), .Y(n_497) );
AO221x2_ASAP7_75t_L g654 ( .A1(n_147), .A2(n_200), .B1(n_642), .B2(n_647), .C(n_655), .Y(n_654) );
OA22x2_ASAP7_75t_L g247 ( .A1(n_150), .A2(n_176), .B1(n_248), .B2(n_249), .Y(n_247) );
INVx1_ASAP7_75t_L g275 ( .A(n_150), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g288 ( .A1(n_151), .A2(n_289), .B(n_295), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_152), .A2(n_232), .B1(n_328), .B2(n_494), .Y(n_555) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_155), .A2(n_196), .B1(n_343), .B2(n_397), .Y(n_396) );
XOR2x2_ASAP7_75t_L g847 ( .A(n_156), .B(n_848), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_156), .A2(n_873), .B1(n_875), .B2(n_879), .Y(n_872) );
INVx1_ASAP7_75t_L g318 ( .A(n_157), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_160), .A2(n_223), .B1(n_650), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_162), .A2(n_197), .B1(n_280), .B2(n_297), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_165), .A2(n_222), .B1(n_350), .B2(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_168), .A2(n_174), .B1(n_377), .B2(n_378), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_170), .B(n_522), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_171), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_L g580 ( .A(n_172), .Y(n_580) );
BUFx2_ASAP7_75t_L g597 ( .A(n_173), .Y(n_597) );
INVx1_ASAP7_75t_L g267 ( .A(n_175), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_175), .B(n_273), .Y(n_317) );
OAI21xp33_ASAP7_75t_L g276 ( .A1(n_176), .A2(n_192), .B(n_277), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_177), .A2(n_201), .B1(n_383), .B2(n_384), .Y(n_604) );
INVx1_ASAP7_75t_L g542 ( .A(n_182), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_184), .A2(n_217), .B1(n_377), .B2(n_378), .Y(n_376) );
AOI221x1_ASAP7_75t_SL g486 ( .A1(n_185), .A2(n_188), .B1(n_437), .B2(n_487), .C(n_488), .Y(n_486) );
INVx1_ASAP7_75t_L g439 ( .A(n_187), .Y(n_439) );
INVx1_ASAP7_75t_L g255 ( .A(n_192), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_192), .B(n_221), .Y(n_315) );
AOI21xp33_ASAP7_75t_L g436 ( .A1(n_193), .A2(n_437), .B(n_438), .Y(n_436) );
OAI22xp5_ASAP7_75t_L g875 ( .A1(n_194), .A2(n_876), .B1(n_877), .B2(n_878), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_194), .Y(n_876) );
AOI221xp5_ASAP7_75t_L g556 ( .A1(n_198), .A2(n_225), .B1(n_405), .B2(n_557), .C(n_558), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_199), .A2(n_408), .B(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g373 ( .A(n_206), .Y(n_373) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_208), .A2(n_224), .B1(n_343), .B2(n_397), .Y(n_503) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_210), .A2(n_371), .B(n_372), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_212), .A2(n_214), .B1(n_322), .B2(n_429), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g591 ( .A1(n_213), .A2(n_592), .B(n_593), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_221), .B(n_260), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_226), .B(n_297), .Y(n_548) );
INVx1_ASAP7_75t_L g646 ( .A(n_228), .Y(n_646) );
HB1xp67_ASAP7_75t_L g882 ( .A(n_228), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_231), .A2(n_233), .B1(n_397), .B2(n_421), .Y(n_554) );
O2A1O1Ixp33_ASAP7_75t_SL g234 ( .A1(n_235), .A2(n_532), .B(n_627), .C(n_636), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_235), .A2(n_532), .B(n_628), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_237), .B1(n_412), .B2(n_531), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
XNOR2xp5_ASAP7_75t_L g237 ( .A(n_238), .B(n_356), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
OR2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_319), .Y(n_240) );
NAND3xp33_ASAP7_75t_L g241 ( .A(n_242), .B(n_278), .C(n_288), .Y(n_241) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
INVx1_ASAP7_75t_L g576 ( .A(n_244), .Y(n_576) );
BUFx8_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
BUFx3_ASAP7_75t_L g405 ( .A(n_245), .Y(n_405) );
INVx2_ASAP7_75t_L g442 ( .A(n_245), .Y(n_442) );
BUFx6f_ASAP7_75t_L g468 ( .A(n_245), .Y(n_468) );
AND2x4_ASAP7_75t_L g245 ( .A(n_246), .B(n_256), .Y(n_245) );
AND2x4_ASAP7_75t_L g281 ( .A(n_246), .B(n_282), .Y(n_281) );
AND2x4_ASAP7_75t_L g365 ( .A(n_246), .B(n_282), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_246), .B(n_256), .Y(n_371) );
AND2x2_ASAP7_75t_L g246 ( .A(n_247), .B(n_250), .Y(n_246) );
AND2x2_ASAP7_75t_L g287 ( .A(n_247), .B(n_251), .Y(n_287) );
AND2x2_ASAP7_75t_L g303 ( .A(n_247), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g336 ( .A(n_247), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_248), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp33_ASAP7_75t_L g252 ( .A(n_249), .B(n_253), .Y(n_252) );
INVx3_ASAP7_75t_L g260 ( .A(n_249), .Y(n_260) );
NAND2xp33_ASAP7_75t_L g266 ( .A(n_249), .B(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g277 ( .A(n_249), .Y(n_277) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_249), .Y(n_301) );
AND2x4_ASAP7_75t_L g335 ( .A(n_250), .B(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_253), .B(n_275), .Y(n_274) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_255), .A2(n_277), .B(n_305), .Y(n_304) );
AND2x4_ASAP7_75t_L g270 ( .A(n_256), .B(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g294 ( .A(n_256), .B(n_287), .Y(n_294) );
AND2x2_ASAP7_75t_L g347 ( .A(n_256), .B(n_335), .Y(n_347) );
AND2x4_ASAP7_75t_L g369 ( .A(n_256), .B(n_271), .Y(n_369) );
AND2x4_ASAP7_75t_L g384 ( .A(n_256), .B(n_335), .Y(n_384) );
AND2x2_ASAP7_75t_L g408 ( .A(n_256), .B(n_287), .Y(n_408) );
AND2x4_ASAP7_75t_L g256 ( .A(n_257), .B(n_262), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g282 ( .A(n_258), .B(n_262), .Y(n_282) );
AND2x2_ASAP7_75t_L g299 ( .A(n_258), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g325 ( .A(n_258), .B(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g337 ( .A(n_258), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_261), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_260), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g273 ( .A(n_260), .Y(n_273) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_261), .B(n_272), .C(n_317), .Y(n_316) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g326 ( .A(n_263), .Y(n_326) );
AND2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_266), .Y(n_263) );
BUFx3_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx6f_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_270), .Y(n_402) );
AND2x4_ASAP7_75t_L g329 ( .A(n_271), .B(n_330), .Y(n_329) );
AND2x4_ASAP7_75t_L g355 ( .A(n_271), .B(n_337), .Y(n_355) );
AND2x4_ASAP7_75t_L g378 ( .A(n_271), .B(n_330), .Y(n_378) );
AND2x4_ASAP7_75t_L g387 ( .A(n_271), .B(n_337), .Y(n_387) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_276), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
BUFx2_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
BUFx6f_ASAP7_75t_L g437 ( .A(n_281), .Y(n_437) );
BUFx3_ASAP7_75t_L g476 ( .A(n_281), .Y(n_476) );
INVx1_ASAP7_75t_L g512 ( .A(n_281), .Y(n_512) );
AND2x2_ASAP7_75t_L g286 ( .A(n_282), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g344 ( .A(n_282), .B(n_335), .Y(n_344) );
AND2x4_ASAP7_75t_L g366 ( .A(n_282), .B(n_287), .Y(n_366) );
AND2x4_ASAP7_75t_L g383 ( .A(n_282), .B(n_335), .Y(n_383) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx3_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx2_ASAP7_75t_L g452 ( .A(n_286), .Y(n_452) );
BUFx6f_ASAP7_75t_L g541 ( .A(n_286), .Y(n_541) );
AND2x4_ASAP7_75t_L g323 ( .A(n_287), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g351 ( .A(n_287), .B(n_337), .Y(n_351) );
AND2x4_ASAP7_75t_L g380 ( .A(n_287), .B(n_337), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_287), .B(n_330), .Y(n_381) );
AND2x2_ASAP7_75t_L g460 ( .A(n_287), .B(n_337), .Y(n_460) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g487 ( .A(n_292), .Y(n_487) );
INVx2_ASAP7_75t_L g557 ( .A(n_292), .Y(n_557) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx2_ASAP7_75t_L g363 ( .A(n_293), .Y(n_363) );
INVx2_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx3_ASAP7_75t_L g446 ( .A(n_294), .Y(n_446) );
BUFx3_ASAP7_75t_L g592 ( .A(n_294), .Y(n_592) );
OAI22xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_306), .B1(n_307), .B2(n_318), .Y(n_295) );
INVx2_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
INVx5_ASAP7_75t_L g449 ( .A(n_298), .Y(n_449) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
AND2x2_ASAP7_75t_L g368 ( .A(n_299), .B(n_303), .Y(n_368) );
AND2x4_ASAP7_75t_L g520 ( .A(n_299), .B(n_303), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g312 ( .A(n_301), .Y(n_312) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
INVx4_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR2xp33_ASAP7_75t_L g409 ( .A(n_309), .B(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_309), .B(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_309), .B(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g589 ( .A(n_309), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx4_ASAP7_75t_L g374 ( .A(n_310), .Y(n_374) );
INVx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_311), .Y(n_472) );
AO21x2_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_313), .B(n_316), .Y(n_311) );
HB1xp67_ASAP7_75t_L g634 ( .A(n_313), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
NAND4xp25_ASAP7_75t_SL g319 ( .A(n_320), .B(n_331), .C(n_342), .D(n_348), .Y(n_319) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_323), .Y(n_392) );
BUFx3_ASAP7_75t_L g430 ( .A(n_323), .Y(n_430) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_323), .Y(n_461) );
BUFx12f_ASAP7_75t_L g494 ( .A(n_323), .Y(n_494) );
AND2x4_ASAP7_75t_L g377 ( .A(n_324), .B(n_335), .Y(n_377) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_L g330 ( .A(n_325), .Y(n_330) );
INVx1_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
BUFx3_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
BUFx12f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx6_ASAP7_75t_L g496 ( .A(n_329), .Y(n_496) );
AND2x4_ASAP7_75t_L g341 ( .A(n_330), .B(n_335), .Y(n_341) );
BUFx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_334), .Y(n_426) );
BUFx12f_ASAP7_75t_L g463 ( .A(n_334), .Y(n_463) );
AND2x4_ASAP7_75t_L g334 ( .A(n_335), .B(n_337), .Y(n_334) );
AND2x4_ASAP7_75t_L g386 ( .A(n_335), .B(n_337), .Y(n_386) );
BUFx3_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_341), .Y(n_399) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_341), .Y(n_432) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_344), .Y(n_421) );
INVx3_ASAP7_75t_L g858 ( .A(n_344), .Y(n_858) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx5_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_347), .Y(n_397) );
INVx1_ASAP7_75t_L g424 ( .A(n_347), .Y(n_424) );
BUFx3_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx6f_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx8_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
BUFx2_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
INVx4_ASAP7_75t_L g394 ( .A(n_354), .Y(n_394) );
INVx4_ASAP7_75t_L g427 ( .A(n_354), .Y(n_427) );
INVx1_ASAP7_75t_L g464 ( .A(n_354), .Y(n_464) );
INVx2_ASAP7_75t_L g505 ( .A(n_354), .Y(n_505) );
INVx2_ASAP7_75t_L g552 ( .A(n_354), .Y(n_552) );
INVx1_ASAP7_75t_L g854 ( .A(n_354), .Y(n_854) );
INVx8_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
XNOR2x1_ASAP7_75t_L g357 ( .A(n_358), .B(n_388), .Y(n_357) );
XNOR2x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
OR2x2_ASAP7_75t_L g360 ( .A(n_361), .B(n_375), .Y(n_360) );
NAND4xp25_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .C(n_367), .D(n_370), .Y(n_361) );
BUFx3_ASAP7_75t_L g516 ( .A(n_363), .Y(n_516) );
INVx2_ASAP7_75t_L g598 ( .A(n_366), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx4_ASAP7_75t_L g561 ( .A(n_374), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_374), .B(n_618), .Y(n_617) );
NAND4xp25_ASAP7_75t_L g375 ( .A(n_376), .B(n_379), .C(n_382), .D(n_385), .Y(n_375) );
XNOR2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_411), .Y(n_388) );
NAND4xp75_ASAP7_75t_L g389 ( .A(n_390), .B(n_395), .C(n_400), .D(n_404), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_398), .Y(n_395) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_403), .Y(n_400) );
INVx3_ASAP7_75t_L g543 ( .A(n_402), .Y(n_543) );
INVx2_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g531 ( .A(n_412), .Y(n_531) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_481), .B1(n_529), .B2(n_530), .Y(n_412) );
INVx1_ASAP7_75t_L g529 ( .A(n_413), .Y(n_529) );
XNOR2xp5_ASAP7_75t_L g413 ( .A(n_414), .B(n_453), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_416), .Y(n_415) );
XNOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
NOR2x1_ASAP7_75t_L g418 ( .A(n_419), .B(n_433), .Y(n_418) );
NAND4xp25_ASAP7_75t_L g419 ( .A(n_420), .B(n_425), .C(n_428), .D(n_431), .Y(n_419) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
NAND3xp33_ASAP7_75t_L g433 ( .A(n_434), .B(n_443), .C(n_447), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_440), .Y(n_435) );
INVx4_ASAP7_75t_L g547 ( .A(n_437), .Y(n_547) );
INVx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx2_ASAP7_75t_L g514 ( .A(n_442), .Y(n_514) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g500 ( .A(n_449), .Y(n_500) );
INVx3_ASAP7_75t_L g567 ( .A(n_449), .Y(n_567) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g865 ( .A(n_451), .Y(n_865) );
BUFx6f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND4xp75_ASAP7_75t_L g456 ( .A(n_457), .B(n_465), .C(n_474), .D(n_478), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_462), .Y(n_457) );
BUFx6f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
BUFx12f_ASAP7_75t_L g853 ( .A(n_463), .Y(n_853) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_467), .B(n_469), .Y(n_465) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_471), .B(n_473), .Y(n_470) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_SL g491 ( .A(n_472), .Y(n_491) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
AND2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_477), .Y(n_474) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g530 ( .A(n_481), .Y(n_530) );
XNOR2x1_ASAP7_75t_L g481 ( .A(n_482), .B(n_506), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
XOR2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
NAND4xp75_ASAP7_75t_L g485 ( .A(n_486), .B(n_492), .C(n_498), .D(n_502), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_489), .B(n_490), .Y(n_488) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
AND2x2_ASAP7_75t_L g492 ( .A(n_493), .B(n_497), .Y(n_492) );
INVx5_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_501), .Y(n_498) );
AND2x2_ASAP7_75t_L g502 ( .A(n_503), .B(n_504), .Y(n_502) );
INVx1_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2x1_ASAP7_75t_SL g508 ( .A(n_509), .B(n_524), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_510), .B(n_513), .C(n_515), .Y(n_509) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
OAI21xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_519), .B(n_521), .Y(n_517) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_519), .A2(n_594), .B1(n_596), .B2(n_598), .Y(n_593) );
INVx4_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx1_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
NAND4xp25_ASAP7_75t_SL g524 ( .A(n_525), .B(n_526), .C(n_527), .D(n_528), .Y(n_524) );
XNOR2x1_ASAP7_75t_L g532 ( .A(n_533), .B(n_581), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
XNOR2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_562), .Y(n_535) );
NAND4xp75_ASAP7_75t_L g537 ( .A(n_538), .B(n_549), .C(n_553), .D(n_556), .Y(n_537) );
NOR2xp67_ASAP7_75t_L g538 ( .A(n_539), .B(n_545), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_540), .A2(n_542), .B1(n_543), .B2(n_544), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_547), .B(n_548), .Y(n_545) );
AND2x2_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
XOR2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_580), .Y(n_562) );
NOR4xp75_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .C(n_571), .D(n_574), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_SL g571 ( .A(n_572), .B(n_573), .Y(n_571) );
OAI21x1_ASAP7_75t_SL g574 ( .A1(n_575), .A2(n_576), .B(n_577), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_607), .B1(n_624), .B2(n_625), .Y(n_581) );
INVx1_ASAP7_75t_L g624 ( .A(n_582), .Y(n_624) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g606 ( .A(n_586), .Y(n_606) );
NOR2x1_ASAP7_75t_L g586 ( .A(n_587), .B(n_600), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .C(n_599), .Y(n_587) );
INVx2_ASAP7_75t_L g863 ( .A(n_592), .Y(n_863) );
CKINVDCx16_ASAP7_75t_R g594 ( .A(n_595), .Y(n_594) );
CKINVDCx9p33_ASAP7_75t_R g596 ( .A(n_597), .Y(n_596) );
NAND4xp25_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .C(n_603), .D(n_604), .Y(n_600) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
HB1xp67_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_609), .Y(n_626) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_619), .Y(n_611) );
NAND4xp25_ASAP7_75t_L g612 ( .A(n_613), .B(n_614), .C(n_615), .D(n_616), .Y(n_612) );
NAND4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .C(n_622), .D(n_623), .Y(n_619) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
BUFx3_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
HB1xp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
NAND3xp33_ASAP7_75t_L g630 ( .A(n_631), .B(n_634), .C(n_635), .Y(n_630) );
AND2x2_ASAP7_75t_L g869 ( .A(n_631), .B(n_870), .Y(n_869) );
AND2x2_ASAP7_75t_L g874 ( .A(n_631), .B(n_871), .Y(n_874) );
AOI21xp5_ASAP7_75t_L g883 ( .A1(n_631), .A2(n_635), .B(n_688), .Y(n_883) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AO21x1_ASAP7_75t_L g880 ( .A1(n_632), .A2(n_881), .B(n_883), .Y(n_880) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g643 ( .A(n_633), .B(n_644), .Y(n_643) );
AND3x4_ASAP7_75t_L g687 ( .A(n_633), .B(n_645), .C(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g870 ( .A(n_634), .B(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_635), .Y(n_871) );
OAI221xp5_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_843), .B1(n_845), .B2(n_867), .C(n_872), .Y(n_636) );
AOI221x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_720), .B1(n_721), .B2(n_726), .C(n_765), .Y(n_637) );
OAI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_658), .B(n_671), .C(n_715), .Y(n_638) );
INVx1_ASAP7_75t_L g737 ( .A(n_639), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_653), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g704 ( .A(n_640), .B(n_684), .Y(n_704) );
CKINVDCx6p67_ASAP7_75t_R g707 ( .A(n_640), .Y(n_707) );
AND2x2_ASAP7_75t_L g714 ( .A(n_640), .B(n_710), .Y(n_714) );
AND2x2_ASAP7_75t_L g729 ( .A(n_640), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g759 ( .A(n_640), .B(n_750), .Y(n_759) );
AND2x2_ASAP7_75t_L g787 ( .A(n_640), .B(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g793 ( .A(n_640), .B(n_708), .Y(n_793) );
AND2x2_ASAP7_75t_L g811 ( .A(n_640), .B(n_717), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_640), .B(n_654), .Y(n_825) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_649), .Y(n_640) );
INVx3_ASAP7_75t_L g724 ( .A(n_642), .Y(n_724) );
AND2x4_ASAP7_75t_L g642 ( .A(n_643), .B(n_645), .Y(n_642) );
AND2x2_ASAP7_75t_L g650 ( .A(n_643), .B(n_651), .Y(n_650) );
AND2x4_ASAP7_75t_L g656 ( .A(n_643), .B(n_651), .Y(n_656) );
AND2x2_ASAP7_75t_L g690 ( .A(n_643), .B(n_651), .Y(n_690) );
AND2x4_ASAP7_75t_L g647 ( .A(n_645), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g662 ( .A(n_645), .B(n_648), .Y(n_662) );
AND2x2_ASAP7_75t_L g652 ( .A(n_648), .B(n_651), .Y(n_652) );
AND2x2_ASAP7_75t_L g657 ( .A(n_648), .B(n_651), .Y(n_657) );
AND2x4_ASAP7_75t_L g680 ( .A(n_648), .B(n_651), .Y(n_680) );
AND2x2_ASAP7_75t_L g750 ( .A(n_653), .B(n_685), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_653), .B(n_707), .Y(n_820) );
NOR3xp33_ASAP7_75t_L g841 ( .A(n_653), .B(n_659), .C(n_721), .Y(n_841) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g708 ( .A(n_654), .B(n_685), .Y(n_708) );
AND2x2_ASAP7_75t_L g710 ( .A(n_654), .B(n_684), .Y(n_710) );
OR2x2_ASAP7_75t_L g718 ( .A(n_654), .B(n_685), .Y(n_718) );
AND2x2_ASAP7_75t_L g757 ( .A(n_654), .B(n_707), .Y(n_757) );
OAI221xp5_ASAP7_75t_L g770 ( .A1(n_654), .A2(n_658), .B1(n_771), .B2(n_773), .C(n_774), .Y(n_770) );
BUFx2_ASAP7_75t_L g844 ( .A(n_656), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_663), .Y(n_658) );
INVx2_ASAP7_75t_L g692 ( .A(n_659), .Y(n_692) );
NOR2xp33_ASAP7_75t_L g695 ( .A(n_659), .B(n_668), .Y(n_695) );
INVx3_ASAP7_75t_L g709 ( .A(n_659), .Y(n_709) );
INVx2_ASAP7_75t_L g733 ( .A(n_659), .Y(n_733) );
AND2x2_ASAP7_75t_L g744 ( .A(n_659), .B(n_707), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g781 ( .A(n_659), .B(n_751), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_659), .B(n_674), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_659), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_SL g678 ( .A(n_662), .Y(n_678) );
A2O1A1Ixp33_ASAP7_75t_L g715 ( .A1(n_663), .A2(n_714), .B(n_716), .C(n_719), .Y(n_715) );
AND2x2_ASAP7_75t_L g663 ( .A(n_664), .B(n_668), .Y(n_663) );
INVx2_ASAP7_75t_L g681 ( .A(n_664), .Y(n_681) );
AND2x2_ASAP7_75t_L g702 ( .A(n_664), .B(n_674), .Y(n_702) );
OR2x2_ASAP7_75t_L g747 ( .A(n_664), .B(n_701), .Y(n_747) );
INVxp67_ASAP7_75t_L g777 ( .A(n_664), .Y(n_777) );
OR2x2_ASAP7_75t_L g779 ( .A(n_664), .B(n_668), .Y(n_779) );
INVx2_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OR2x2_ASAP7_75t_L g734 ( .A(n_665), .B(n_668), .Y(n_734) );
AND2x2_ASAP7_75t_L g796 ( .A(n_665), .B(n_675), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_666), .B(n_667), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_668), .B(n_692), .Y(n_691) );
INVx4_ASAP7_75t_L g701 ( .A(n_668), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_668), .B(n_692), .Y(n_753) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AOI211xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_682), .B(n_693), .C(n_711), .Y(n_671) );
O2A1O1Ixp33_ASAP7_75t_L g758 ( .A1(n_672), .A2(n_759), .B(n_760), .C(n_761), .Y(n_758) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_673), .B(n_769), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_681), .Y(n_673) );
INVx2_ASAP7_75t_L g736 ( .A(n_674), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_674), .B(n_743), .Y(n_742) );
AND2x2_ASAP7_75t_L g754 ( .A(n_674), .B(n_713), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_674), .B(n_734), .Y(n_764) );
OR2x2_ASAP7_75t_L g802 ( .A(n_674), .B(n_777), .Y(n_802) );
INVx4_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g719 ( .A(n_675), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_675), .B(n_740), .Y(n_739) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_675), .B(n_747), .Y(n_746) );
NOR3xp33_ASAP7_75t_SL g752 ( .A(n_675), .B(n_749), .C(n_753), .Y(n_752) );
AND2x2_ASAP7_75t_L g812 ( .A(n_675), .B(n_813), .Y(n_812) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
INVx3_ASAP7_75t_SL g727 ( .A(n_681), .Y(n_727) );
INVxp67_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_684), .B(n_691), .Y(n_683) );
AOI211xp5_ASAP7_75t_L g774 ( .A1(n_684), .A2(n_695), .B(n_775), .C(n_781), .Y(n_774) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
NOR2xp33_ASAP7_75t_L g760 ( .A(n_692), .B(n_703), .Y(n_760) );
AND2x2_ASAP7_75t_L g827 ( .A(n_692), .B(n_757), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_692), .B(n_699), .Y(n_840) );
A2O1A1Ixp33_ASAP7_75t_SL g693 ( .A1(n_694), .A2(n_696), .B(n_703), .C(n_705), .Y(n_693) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_694), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
AOI32xp33_ASAP7_75t_L g705 ( .A1(n_695), .A2(n_702), .A3(n_706), .B1(n_709), .B2(n_710), .Y(n_705) );
INVx1_ASAP7_75t_L g807 ( .A(n_696), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_697), .B(n_702), .Y(n_696) );
HB1xp67_ASAP7_75t_L g768 ( .A(n_697), .Y(n_768) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g803 ( .A(n_698), .Y(n_803) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_699), .Y(n_795) );
INVx1_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx1_ASAP7_75t_L g740 ( .A(n_700), .Y(n_740) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx2_ASAP7_75t_L g713 ( .A(n_701), .Y(n_713) );
INVx1_ASAP7_75t_L g791 ( .A(n_702), .Y(n_791) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g778 ( .A(n_704), .B(n_709), .Y(n_778) );
INVx1_ASAP7_75t_L g762 ( .A(n_706), .Y(n_762) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
AND2x2_ASAP7_75t_L g716 ( .A(n_707), .B(n_717), .Y(n_716) );
AOI322xp5_ASAP7_75t_L g745 ( .A1(n_707), .A2(n_727), .A3(n_746), .B1(n_748), .B2(n_752), .C1(n_754), .C2(n_755), .Y(n_745) );
AND2x2_ASAP7_75t_L g772 ( .A(n_707), .B(n_710), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_707), .B(n_750), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_707), .B(n_730), .Y(n_809) );
AND2x2_ASAP7_75t_L g730 ( .A(n_708), .B(n_709), .Y(n_730) );
INVx1_ASAP7_75t_L g780 ( .A(n_708), .Y(n_780) );
INVx3_ASAP7_75t_L g788 ( .A(n_709), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_709), .B(n_772), .Y(n_815) );
AND2x2_ASAP7_75t_L g743 ( .A(n_710), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g751 ( .A(n_710), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_710), .B(n_787), .Y(n_801) );
INVxp67_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_713), .B(n_714), .Y(n_712) );
INVx1_ASAP7_75t_L g741 ( .A(n_714), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_714), .B(n_790), .Y(n_789) );
AND2x2_ASAP7_75t_L g786 ( .A(n_717), .B(n_787), .Y(n_786) );
AND2x2_ASAP7_75t_L g817 ( .A(n_717), .B(n_744), .Y(n_817) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_720), .B(n_736), .Y(n_783) );
CKINVDCx5p33_ASAP7_75t_R g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_722), .B(n_725), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B(n_731), .C(n_758), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_727), .A2(n_773), .B1(n_823), .B2(n_826), .Y(n_822) );
INVx1_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
O2A1O1Ixp33_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_735), .B(n_737), .C(n_738), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_734), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g755 ( .A(n_733), .B(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_733), .B(n_759), .Y(n_769) );
AND2x2_ASAP7_75t_L g830 ( .A(n_733), .B(n_813), .Y(n_830) );
OAI21xp33_ASAP7_75t_L g808 ( .A1(n_734), .A2(n_809), .B(n_810), .Y(n_808) );
INVx1_ASAP7_75t_L g842 ( .A(n_734), .Y(n_842) );
AOI221xp5_ASAP7_75t_SL g818 ( .A1(n_736), .A2(n_813), .B1(n_819), .B2(n_822), .C(n_828), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_737), .B(n_830), .Y(n_829) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_739), .A2(n_741), .B(n_742), .C(n_745), .Y(n_738) );
INVx2_ASAP7_75t_L g773 ( .A(n_740), .Y(n_773) );
A2O1A1Ixp33_ASAP7_75t_SL g819 ( .A1(n_741), .A2(n_816), .B(n_820), .C(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g813 ( .A(n_747), .Y(n_813) );
AND2x2_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g790 ( .A(n_753), .Y(n_790) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g835 ( .A(n_759), .Y(n_835) );
NOR2xp33_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
NAND5xp2_ASAP7_75t_L g765 ( .A(n_766), .B(n_804), .C(n_818), .D(n_831), .E(n_833), .Y(n_765) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_770), .B(n_782), .C(n_784), .Y(n_766) );
NOR2xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_769), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g834 ( .A(n_771), .B(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
AOI222xp33_ASAP7_75t_L g833 ( .A1(n_772), .A2(n_834), .B1(n_836), .B2(n_838), .C1(n_841), .C2(n_842), .Y(n_833) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_773), .B(n_786), .Y(n_785) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_776), .A2(n_778), .B1(n_779), .B2(n_780), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g799 ( .A(n_779), .Y(n_799) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
A2O1A1Ixp33_ASAP7_75t_L g784 ( .A1(n_785), .A2(n_789), .B(n_791), .C(n_792), .Y(n_784) );
NOR2x1_ASAP7_75t_L g797 ( .A(n_788), .B(n_798), .Y(n_797) );
AND2x2_ASAP7_75t_L g805 ( .A(n_788), .B(n_806), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g837 ( .A(n_788), .B(n_799), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g838 ( .A(n_791), .B(n_839), .Y(n_838) );
AOI221xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_797), .B2(n_799), .C(n_800), .Y(n_792) );
AND2x2_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx1_ASAP7_75t_L g806 ( .A(n_798), .Y(n_806) );
NOR3xp33_ASAP7_75t_L g800 ( .A(n_801), .B(n_802), .C(n_803), .Y(n_800) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_802), .A2(n_815), .B(n_816), .Y(n_814) );
AOI211xp5_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B(n_808), .C(n_814), .Y(n_804) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_812), .Y(n_810) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVxp33_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g843 ( .A(n_844), .Y(n_843) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g877 ( .A(n_848), .Y(n_877) );
NOR2x1_ASAP7_75t_L g848 ( .A(n_849), .B(n_859), .Y(n_848) );
NAND4xp25_ASAP7_75t_SL g849 ( .A(n_850), .B(n_851), .C(n_852), .D(n_855), .Y(n_849) );
BUFx4f_ASAP7_75t_L g856 ( .A(n_857), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
NAND4xp25_ASAP7_75t_L g859 ( .A(n_860), .B(n_861), .C(n_864), .D(n_866), .Y(n_859) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
HB1xp67_ASAP7_75t_L g868 ( .A(n_869), .Y(n_868) );
BUFx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g878 ( .A(n_877), .Y(n_878) );
BUFx2_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_882), .Y(n_881) );
endmodule