module fake_jpeg_3512_n_435 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_435);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_435;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_17),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_3),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_11),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_6),
.Y(n_52)
);

BUFx6f_ASAP7_75t_SL g53 ( 
.A(n_13),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g165 ( 
.A(n_54),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_14),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_55),
.B(n_73),
.Y(n_119)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_57),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_58),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_59),
.Y(n_174)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_60),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_32),
.B(n_14),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_61),
.A2(n_62),
.B(n_68),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_0),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_63),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_19),
.B(n_21),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_66),
.B(n_86),
.Y(n_150)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_67),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_19),
.B(n_0),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_24),
.Y(n_69)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_72),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_13),
.Y(n_73)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_74),
.Y(n_143)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_75),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_76),
.Y(n_146)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_43),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_18),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_80),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_81),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_82),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx10_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx5_ASAP7_75t_SL g183 ( 
.A(n_84),
.Y(n_183)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_38),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_85),
.A2(n_35),
.B1(n_39),
.B2(n_49),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_87),
.Y(n_136)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_37),
.Y(n_88)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_22),
.B(n_13),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_90),
.B(n_95),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_31),
.Y(n_91)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_91),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_31),
.Y(n_92)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_92),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_31),
.Y(n_93)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_93),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_30),
.Y(n_94)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_22),
.B(n_1),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

BUFx24_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_97),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_98),
.B(n_105),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_24),
.B(n_4),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_99),
.B(n_35),
.Y(n_131)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_12),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_101),
.B(n_102),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_20),
.B(n_12),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g103 ( 
.A(n_33),
.Y(n_103)
);

NAND2x1_ASAP7_75t_SL g152 ( 
.A(n_103),
.B(n_109),
.Y(n_152)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_23),
.B(n_4),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_106),
.Y(n_188)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_42),
.Y(n_108)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_108),
.Y(n_172)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g110 ( 
.A(n_29),
.Y(n_110)
);

INVx6_ASAP7_75t_SL g178 ( 
.A(n_110),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_23),
.B(n_4),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_112),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_34),
.B(n_5),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_38),
.Y(n_113)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_113),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_44),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_114),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_118),
.B(n_176),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_62),
.A2(n_53),
.B1(n_45),
.B2(n_52),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g247 ( 
.A1(n_120),
.A2(n_142),
.B1(n_149),
.B2(n_153),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_99),
.A2(n_41),
.B1(n_46),
.B2(n_45),
.Y(n_123)
);

AOI22x1_ASAP7_75t_L g251 ( 
.A1(n_123),
.A2(n_158),
.B1(n_166),
.B2(n_118),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_85),
.A2(n_53),
.B1(n_34),
.B2(n_49),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_126),
.A2(n_148),
.B1(n_171),
.B2(n_175),
.Y(n_226)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_127),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_131),
.B(n_133),
.Y(n_193)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_68),
.B(n_39),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_61),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_141),
.B(n_143),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_88),
.A2(n_52),
.B1(n_37),
.B2(n_46),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_94),
.B(n_46),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_144),
.B(n_152),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_78),
.A2(n_52),
.B1(n_40),
.B2(n_7),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_65),
.A2(n_52),
.B1(n_33),
.B2(n_40),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_114),
.A2(n_74),
.B1(n_82),
.B2(n_81),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_83),
.A2(n_29),
.B1(n_6),
.B2(n_7),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_57),
.A2(n_29),
.B1(n_7),
.B2(n_8),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_58),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_167)
);

OA22x2_ASAP7_75t_L g248 ( 
.A1(n_167),
.A2(n_149),
.B1(n_148),
.B2(n_142),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_59),
.A2(n_5),
.B1(n_10),
.B2(n_11),
.Y(n_171)
);

A2O1A1Ixp33_ASAP7_75t_L g173 ( 
.A1(n_84),
.A2(n_104),
.B(n_110),
.C(n_11),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_149),
.B(n_142),
.C(n_171),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_89),
.A2(n_5),
.B1(n_10),
.B2(n_12),
.Y(n_175)
);

NAND2x1_ASAP7_75t_L g176 ( 
.A(n_77),
.B(n_10),
.Y(n_176)
);

NAND2x1_ASAP7_75t_L g177 ( 
.A(n_91),
.B(n_93),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_177),
.B(n_180),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_92),
.A2(n_72),
.B1(n_76),
.B2(n_84),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_182),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_L g186 ( 
.A1(n_85),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_85),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_85),
.A2(n_86),
.B1(n_81),
.B2(n_82),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_115),
.Y(n_190)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_190),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_173),
.A2(n_120),
.B(n_176),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_191),
.A2(n_213),
.B(n_247),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g192 ( 
.A(n_116),
.B(n_119),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_192),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_194),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_165),
.A2(n_170),
.B1(n_136),
.B2(n_156),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_195),
.Y(n_254)
);

AO22x1_ASAP7_75t_SL g196 ( 
.A1(n_159),
.A2(n_189),
.B1(n_187),
.B2(n_186),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g283 ( 
.A1(n_196),
.A2(n_210),
.B(n_234),
.Y(n_283)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_140),
.Y(n_197)
);

INVxp67_ASAP7_75t_SL g288 ( 
.A(n_197),
.Y(n_288)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_165),
.A2(n_170),
.B1(n_127),
.B2(n_125),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_198),
.A2(n_200),
.B1(n_207),
.B2(n_215),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_155),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_199),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_118),
.A2(n_166),
.B1(n_126),
.B2(n_159),
.Y(n_200)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g271 ( 
.A(n_201),
.Y(n_271)
);

INVx11_ASAP7_75t_L g202 ( 
.A(n_132),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_151),
.B(n_134),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_203),
.B(n_246),
.C(n_250),
.Y(n_284)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_145),
.Y(n_204)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_204),
.Y(n_253)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_138),
.Y(n_205)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_205),
.Y(n_264)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_206),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g207 ( 
.A1(n_172),
.A2(n_137),
.B1(n_181),
.B2(n_162),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_150),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_208),
.B(n_211),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_169),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_209),
.B(n_217),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_135),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_148),
.A2(n_153),
.B1(n_144),
.B2(n_133),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_212),
.A2(n_219),
.B1(n_242),
.B2(n_244),
.Y(n_266)
);

A2O1A1Ixp33_ASAP7_75t_L g213 ( 
.A1(n_179),
.A2(n_178),
.B(n_152),
.C(n_188),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_213),
.A2(n_234),
.B(n_193),
.C(n_210),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_121),
.B(n_184),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_214),
.B(n_223),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_125),
.A2(n_135),
.B1(n_129),
.B2(n_130),
.Y(n_215)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_132),
.Y(n_216)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_216),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_177),
.B(n_117),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_167),
.A2(n_122),
.B1(n_124),
.B2(n_128),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_220),
.B(n_222),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_143),
.B(n_130),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_139),
.B(n_157),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_225),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_147),
.B(n_154),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_168),
.B(n_160),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_227),
.B(n_230),
.Y(n_287)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

INVx8_ASAP7_75t_L g229 ( 
.A(n_155),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_146),
.B(n_164),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_183),
.B(n_164),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_233),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_146),
.B(n_174),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_232),
.B(n_245),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_174),
.B(n_180),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_155),
.Y(n_236)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_236),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_141),
.B(n_156),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_237),
.B(n_238),
.Y(n_269)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_178),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_239),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_141),
.B(n_156),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_240),
.B(n_238),
.Y(n_290)
);

INVx5_ASAP7_75t_L g241 ( 
.A(n_138),
.Y(n_241)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_241),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_126),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_123),
.A2(n_53),
.B1(n_98),
.B2(n_141),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_243),
.A2(n_251),
.B1(n_217),
.B2(n_234),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_126),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_115),
.B(n_116),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g293 ( 
.A1(n_248),
.A2(n_249),
.B1(n_247),
.B2(n_205),
.Y(n_293)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_186),
.A2(n_189),
.B1(n_187),
.B2(n_126),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_115),
.B(n_116),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_252),
.B(n_274),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_SL g256 ( 
.A(n_192),
.B(n_203),
.C(n_221),
.Y(n_256)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_256),
.B(n_239),
.C(n_241),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_191),
.A2(n_221),
.B1(n_196),
.B2(n_251),
.Y(n_262)
);

A2O1A1Ixp33_ASAP7_75t_SL g297 ( 
.A1(n_262),
.A2(n_272),
.B(n_273),
.C(n_280),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_202),
.B1(n_218),
.B2(n_235),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_221),
.A2(n_196),
.B1(n_251),
.B2(n_192),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_246),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_275),
.A2(n_273),
.B(n_262),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_279),
.B(n_280),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_242),
.A2(n_244),
.B1(n_226),
.B2(n_230),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_232),
.A2(n_247),
.B1(n_248),
.B2(n_227),
.Y(n_281)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_281),
.A2(n_293),
.B(n_229),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_286),
.B(n_290),
.Y(n_298)
);

OAI32xp33_ASAP7_75t_L g289 ( 
.A1(n_250),
.A2(n_248),
.A3(n_247),
.B1(n_219),
.B2(n_190),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_289),
.B(n_206),
.Y(n_296)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_292),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_266),
.A2(n_248),
.B1(n_199),
.B2(n_236),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_295),
.A2(n_296),
.B1(n_313),
.B2(n_266),
.Y(n_329)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_255),
.Y(n_299)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_299),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_276),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_300),
.B(n_307),
.Y(n_334)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_253),
.Y(n_302)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_302),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_253),
.Y(n_304)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_304),
.Y(n_344)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_275),
.B(n_235),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_305),
.A2(n_318),
.B(n_254),
.Y(n_336)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_285),
.Y(n_306)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_306),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_228),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_287),
.B(n_201),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_308),
.B(n_309),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_252),
.B(n_238),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_272),
.B(n_216),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_310),
.B(n_314),
.Y(n_350)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_268),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_311),
.B(n_315),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_312),
.A2(n_286),
.B1(n_292),
.B2(n_254),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_263),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_277),
.B(n_284),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_316),
.B(n_319),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_257),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_317),
.Y(n_342)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_283),
.B(n_256),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_259),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_320),
.A2(n_321),
.B1(n_324),
.B2(n_325),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_288),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_261),
.B(n_263),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g330 ( 
.A1(n_322),
.A2(n_326),
.B(n_274),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_323),
.A2(n_269),
.B(n_291),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_265),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_259),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_258),
.B(n_281),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_305),
.A2(n_283),
.B(n_289),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g365 ( 
.A1(n_328),
.A2(n_336),
.B(n_345),
.Y(n_365)
);

OAI22xp33_ASAP7_75t_L g360 ( 
.A1(n_329),
.A2(n_297),
.B1(n_309),
.B2(n_315),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_330),
.B(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_332),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_314),
.A2(n_293),
.B1(n_283),
.B2(n_282),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_339),
.B1(n_310),
.B2(n_294),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_313),
.A2(n_293),
.B1(n_260),
.B2(n_284),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_337),
.A2(n_346),
.B1(n_347),
.B2(n_313),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_L g338 ( 
.A1(n_297),
.A2(n_323),
.B(n_326),
.C(n_322),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_296),
.A2(n_293),
.B1(n_278),
.B2(n_265),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_313),
.A2(n_278),
.B1(n_291),
.B2(n_271),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_295),
.A2(n_264),
.B1(n_257),
.B2(n_271),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g348 ( 
.A1(n_305),
.A2(n_264),
.B(n_267),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_348),
.B(n_301),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_367),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_334),
.B(n_307),
.Y(n_355)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_355),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_334),
.B(n_308),
.Y(n_356)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_356),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_357),
.A2(n_360),
.B1(n_362),
.B2(n_364),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_300),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_358),
.B(n_366),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_359),
.A2(n_350),
.B1(n_335),
.B2(n_331),
.Y(n_372)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_341),
.B(n_318),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_361),
.B(n_363),
.Y(n_376)
);

OAI22x1_ASAP7_75t_SL g362 ( 
.A1(n_329),
.A2(n_297),
.B1(n_318),
.B2(n_301),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_303),
.C(n_294),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_328),
.A2(n_297),
.B1(n_298),
.B2(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_327),
.B(n_299),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_340),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_371),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_343),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_369),
.Y(n_380)
);

OAI22x1_ASAP7_75t_SL g370 ( 
.A1(n_328),
.A2(n_297),
.B1(n_298),
.B2(n_304),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_370),
.A2(n_338),
.B1(n_345),
.B2(n_342),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_343),
.B(n_302),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_374),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_336),
.B(n_348),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_373),
.B(n_385),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g374 ( 
.A1(n_359),
.A2(n_350),
.B1(n_337),
.B2(n_331),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_357),
.A2(n_346),
.B1(n_347),
.B2(n_348),
.Y(n_378)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_378),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_354),
.A2(n_339),
.B1(n_333),
.B2(n_332),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_379),
.B(n_359),
.Y(n_399)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_383),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_354),
.A2(n_335),
.B1(n_342),
.B2(n_330),
.Y(n_385)
);

AO22x2_ASAP7_75t_L g387 ( 
.A1(n_364),
.A2(n_344),
.B1(n_349),
.B2(n_351),
.Y(n_387)
);

FAx1_ASAP7_75t_L g389 ( 
.A(n_387),
.B(n_370),
.CI(n_362),
.CON(n_389),
.SN(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_376),
.B(n_361),
.C(n_363),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g403 ( 
.A(n_390),
.B(n_394),
.C(n_396),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_377),
.B(n_366),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_391),
.B(n_393),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_381),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_376),
.B(n_361),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_363),
.C(n_364),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_311),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_397),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_385),
.B(n_365),
.C(n_370),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_362),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g409 ( 
.A1(n_399),
.A2(n_378),
.B(n_379),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_395),
.A2(n_383),
.B(n_375),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_401),
.A2(n_398),
.B1(n_389),
.B2(n_380),
.Y(n_412)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_392),
.Y(n_402)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

AO221x1_ASAP7_75t_L g405 ( 
.A1(n_389),
.A2(n_375),
.B1(n_377),
.B2(n_358),
.C(n_380),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_405),
.B(n_406),
.Y(n_411)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_388),
.Y(n_407)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_407),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_409),
.B(n_352),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_408),
.A2(n_388),
.B1(n_392),
.B2(n_400),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_410),
.B(n_412),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_404),
.B(n_386),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_414),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_401),
.A2(n_400),
.B1(n_352),
.B2(n_369),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_417),
.B(n_404),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_415),
.B(n_403),
.C(n_402),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_419),
.B(n_422),
.Y(n_426)
);

XOR2x2_ASAP7_75t_L g420 ( 
.A(n_410),
.B(n_406),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_420),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_417),
.B(n_403),
.Y(n_422)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_423),
.A2(n_408),
.B(n_419),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g425 ( 
.A1(n_421),
.A2(n_411),
.B(n_413),
.Y(n_425)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_425),
.Y(n_429)
);

OAI21x1_ASAP7_75t_L g428 ( 
.A1(n_427),
.A2(n_426),
.B(n_418),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_424),
.Y(n_430)
);

AOI321xp33_ASAP7_75t_L g431 ( 
.A1(n_430),
.A2(n_429),
.A3(n_416),
.B1(n_415),
.B2(n_409),
.C(n_316),
.Y(n_431)
);

OAI211xp5_ASAP7_75t_L g432 ( 
.A1(n_431),
.A2(n_371),
.B(n_384),
.C(n_381),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g433 ( 
.A1(n_432),
.A2(n_372),
.B(n_384),
.Y(n_433)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_433),
.A2(n_382),
.B1(n_407),
.B2(n_356),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_434),
.B(n_420),
.Y(n_435)
);


endmodule