module fake_jpeg_2279_n_564 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_564);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_564;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx2_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx8_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_4),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_56),
.Y(n_150)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_57),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_27),
.B(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_59),
.B(n_66),
.Y(n_128)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g156 ( 
.A(n_62),
.Y(n_156)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_63),
.Y(n_113)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_64),
.Y(n_123)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_27),
.A2(n_1),
.B(n_2),
.Y(n_66)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_67),
.Y(n_125)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_46),
.Y(n_68)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_68),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_19),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_70),
.Y(n_124)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx11_ASAP7_75t_L g157 ( 
.A(n_72),
.Y(n_157)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_73),
.Y(n_137)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

INVx2_ASAP7_75t_SL g121 ( 
.A(n_76),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_77),
.B(n_88),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_22),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_78),
.Y(n_153)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_22),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_79),
.Y(n_154)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx3_ASAP7_75t_SL g172 ( 
.A(n_80),
.Y(n_172)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_81),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g82 ( 
.A(n_39),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_85),
.Y(n_155)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_86),
.Y(n_142)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_87),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_18),
.B(n_1),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_89),
.Y(n_175)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_45),
.Y(n_90)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_90),
.Y(n_159)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_92),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_17),
.Y(n_93)
);

NAND2xp33_ASAP7_75t_SL g168 ( 
.A(n_93),
.B(n_37),
.Y(n_168)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_94),
.Y(n_176)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_48),
.Y(n_95)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_43),
.Y(n_96)
);

INVx4_ASAP7_75t_L g147 ( 
.A(n_96),
.Y(n_147)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

BUFx10_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_43),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_98),
.B(n_100),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_99),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_51),
.B(n_2),
.Y(n_100)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_25),
.Y(n_101)
);

BUFx10_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_25),
.Y(n_102)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_102),
.Y(n_149)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_104),
.Y(n_164)
);

INVx11_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_105),
.Y(n_173)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_25),
.Y(n_106)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_106),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_17),
.Y(n_107)
);

CKINVDCx6p67_ASAP7_75t_R g115 ( 
.A(n_107),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_18),
.B(n_3),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_108),
.B(n_6),
.Y(n_132)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_17),
.Y(n_109)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_109),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_3),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_110),
.B(n_112),
.Y(n_178)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_52),
.Y(n_111)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_111),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_31),
.Y(n_112)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_97),
.Y(n_118)
);

INVx5_ASAP7_75t_L g239 ( 
.A(n_118),
.Y(n_239)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_104),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_122),
.A2(n_58),
.B1(n_85),
.B2(n_75),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_132),
.B(n_152),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_67),
.A2(n_54),
.B1(n_31),
.B2(n_29),
.Y(n_134)
);

AO22x1_ASAP7_75t_L g224 ( 
.A1(n_134),
.A2(n_50),
.B1(n_69),
.B2(n_106),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_79),
.A2(n_54),
.B1(n_29),
.B2(n_34),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_141),
.A2(n_162),
.B1(n_37),
.B2(n_105),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_63),
.B(n_33),
.C(n_53),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_144),
.B(n_171),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_61),
.B(n_36),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_145),
.B(n_53),
.Y(n_210)
);

AND2x2_ASAP7_75t_SL g146 ( 
.A(n_71),
.B(n_37),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_146),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_76),
.B(n_33),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_82),
.B(n_36),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_161),
.B(n_166),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_97),
.A2(n_37),
.B1(n_50),
.B2(n_29),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_84),
.B(n_20),
.Y(n_166)
);

INVx1_ASAP7_75t_SL g219 ( 
.A(n_168),
.Y(n_219)
);

NAND2x1_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_54),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_174),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_101),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_177),
.Y(n_245)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_179),
.Y(n_186)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_72),
.Y(n_182)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_91),
.Y(n_183)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_183),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_184),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_131),
.B(n_178),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_187),
.B(n_209),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_189),
.A2(n_147),
.B1(n_151),
.B2(n_148),
.Y(n_269)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_190),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_117),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_192),
.Y(n_254)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_116),
.Y(n_193)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_193),
.Y(n_260)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_60),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g277 ( 
.A(n_195),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_56),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_196),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_128),
.A2(n_78),
.B1(n_102),
.B2(n_99),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_197),
.A2(n_224),
.B1(n_148),
.B2(n_130),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_199),
.A2(n_226),
.B1(n_219),
.B2(n_149),
.Y(n_262)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_200),
.Y(n_265)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g304 ( 
.A(n_201),
.Y(n_304)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_137),
.Y(n_203)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_203),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_115),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_204),
.B(n_212),
.Y(n_285)
);

BUFx12_ASAP7_75t_L g205 ( 
.A(n_115),
.Y(n_205)
);

BUFx2_ASAP7_75t_SL g267 ( 
.A(n_205),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_115),
.Y(n_206)
);

INVx5_ASAP7_75t_L g259 ( 
.A(n_206),
.Y(n_259)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_207),
.Y(n_292)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_170),
.Y(n_208)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_208),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_131),
.B(n_49),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_210),
.B(n_230),
.Y(n_273)
);

AO22x2_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_80),
.B1(n_62),
.B2(n_28),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_211),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_178),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_177),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_213),
.B(n_217),
.Y(n_299)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_175),
.Y(n_215)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_216),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_128),
.B(n_24),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_248),
.Y(n_275)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_119),
.Y(n_220)
);

BUFx2_ASAP7_75t_SL g294 ( 
.A(n_220),
.Y(n_294)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_165),
.Y(n_221)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_221),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_20),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_222),
.B(n_225),
.Y(n_305)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_163),
.B(n_23),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_130),
.Y(n_227)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_227),
.Y(n_289)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_129),
.Y(n_228)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_228),
.Y(n_293)
);

O2A1O1Ixp33_ASAP7_75t_L g229 ( 
.A1(n_122),
.A2(n_32),
.B(n_24),
.C(n_28),
.Y(n_229)
);

O2A1O1Ixp33_ASAP7_75t_L g291 ( 
.A1(n_229),
.A2(n_127),
.B(n_47),
.C(n_30),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_124),
.B(n_23),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_121),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_231),
.Y(n_290)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_133),
.Y(n_232)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_150),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_233),
.B(n_236),
.Y(n_283)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_121),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_138),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_143),
.B(n_49),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_135),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_237),
.Y(n_272)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_136),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

AOI32xp33_ASAP7_75t_L g240 ( 
.A1(n_159),
.A2(n_32),
.A3(n_28),
.B1(n_24),
.B2(n_50),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_240),
.B(n_242),
.Y(n_298)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_142),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_160),
.B(n_32),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_126),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_243),
.B(n_249),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_150),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_244),
.B(n_247),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_169),
.A2(n_42),
.B(n_35),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_162),
.C(n_172),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_42),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_113),
.B(n_42),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_173),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_120),
.B(n_42),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_250),
.Y(n_263)
);

AO22x1_ASAP7_75t_L g251 ( 
.A1(n_157),
.A2(n_35),
.B1(n_34),
.B2(n_47),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_251),
.B(n_211),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_252),
.B(n_276),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_219),
.A2(n_158),
.B1(n_125),
.B2(n_154),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_258),
.A2(n_227),
.B1(n_192),
.B2(n_223),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_262),
.A2(n_268),
.B1(n_279),
.B2(n_282),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_188),
.B(n_114),
.C(n_139),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_264),
.B(n_271),
.C(n_274),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_269),
.A2(n_288),
.B1(n_206),
.B2(n_252),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_188),
.B(n_172),
.C(n_156),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_202),
.B(n_156),
.C(n_154),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_125),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_278),
.B(n_300),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_199),
.A2(n_153),
.B1(n_180),
.B2(n_35),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_218),
.A2(n_153),
.B1(n_34),
.B2(n_140),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_195),
.B(n_140),
.C(n_127),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_284),
.B(n_301),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_197),
.A2(n_140),
.B1(n_47),
.B2(n_127),
.Y(n_288)
);

O2A1O1Ixp33_ASAP7_75t_L g354 ( 
.A1(n_291),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_196),
.A2(n_47),
.B1(n_30),
.B2(n_21),
.Y(n_295)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_295),
.A2(n_307),
.B1(n_198),
.B2(n_239),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_246),
.B(n_30),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_194),
.B(n_21),
.C(n_7),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_221),
.A2(n_21),
.B1(n_7),
.B2(n_8),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_266),
.B(n_186),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g364 ( 
.A(n_309),
.B(n_335),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g380 ( 
.A1(n_310),
.A2(n_353),
.B1(n_304),
.B2(n_270),
.Y(n_380)
);

BUFx4f_ASAP7_75t_SL g311 ( 
.A(n_254),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g385 ( 
.A(n_311),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_302),
.A2(n_211),
.B1(n_224),
.B2(n_229),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_312),
.A2(n_282),
.B1(n_277),
.B2(n_288),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_290),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_313),
.B(n_314),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

INVx2_ASAP7_75t_SL g315 ( 
.A(n_281),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_315),
.Y(n_392)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_317),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_261),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_318),
.B(n_324),
.Y(n_384)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_297),
.Y(n_319)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_319),
.Y(n_365)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_320),
.Y(n_382)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_260),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g393 ( 
.A(n_321),
.Y(n_393)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_283),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

INVxp67_ASAP7_75t_L g377 ( 
.A(n_325),
.Y(n_377)
);

INVx13_ASAP7_75t_L g326 ( 
.A(n_267),
.Y(n_326)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_326),
.Y(n_359)
);

OAI22xp33_ASAP7_75t_SL g369 ( 
.A1(n_328),
.A2(n_334),
.B1(n_339),
.B2(n_354),
.Y(n_369)
);

OAI21xp33_ASAP7_75t_L g329 ( 
.A1(n_275),
.A2(n_211),
.B(n_243),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g376 ( 
.A(n_329),
.Y(n_376)
);

BUFx4f_ASAP7_75t_SL g330 ( 
.A(n_281),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g395 ( 
.A(n_330),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_276),
.A2(n_245),
.B(n_190),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_331),
.A2(n_332),
.B(n_352),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_298),
.A2(n_245),
.B(n_235),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_251),
.B1(n_200),
.B2(n_193),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_333),
.A2(n_337),
.B1(n_346),
.B2(n_259),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_261),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_300),
.A2(n_232),
.B1(n_228),
.B2(n_185),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_291),
.A2(n_249),
.B(n_237),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_338),
.A2(n_306),
.B(n_272),
.Y(n_387)
);

AOI22x1_ASAP7_75t_SL g339 ( 
.A1(n_275),
.A2(n_214),
.B1(n_241),
.B2(n_185),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_306),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_340),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_278),
.B(n_207),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_341),
.B(n_351),
.Y(n_356)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_260),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_342),
.B(n_344),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_285),
.B(n_214),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_343),
.B(n_345),
.Y(n_368)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_265),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_263),
.B(n_239),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_268),
.A2(n_201),
.B1(n_205),
.B2(n_8),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_296),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_347),
.B(n_350),
.Y(n_373)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_265),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_348),
.B(n_349),
.Y(n_381)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_308),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_296),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_264),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_277),
.A2(n_205),
.B(n_7),
.Y(n_352)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_253),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_274),
.B(n_6),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_355),
.B(n_259),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_316),
.B(n_271),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_362),
.C(n_367),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_361),
.B(n_379),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_322),
.C(n_323),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g418 ( 
.A1(n_363),
.A2(n_370),
.B1(n_380),
.B2(n_386),
.Y(n_418)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_322),
.A2(n_279),
.B1(n_256),
.B2(n_273),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_366),
.A2(n_372),
.B1(n_375),
.B2(n_390),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_284),
.Y(n_367)
);

MAJx2_ASAP7_75t_L g371 ( 
.A(n_322),
.B(n_305),
.C(n_256),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_318),
.C(n_350),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_327),
.A2(n_287),
.B1(n_257),
.B2(n_303),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_327),
.A2(n_286),
.B1(n_304),
.B2(n_289),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_341),
.B(n_355),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_312),
.A2(n_270),
.B1(n_289),
.B2(n_292),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_387),
.Y(n_407)
);

AOI32xp33_ASAP7_75t_L g388 ( 
.A1(n_314),
.A2(n_253),
.A3(n_272),
.B1(n_255),
.B2(n_280),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_388),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g389 ( 
.A1(n_310),
.A2(n_292),
.B1(n_306),
.B2(n_280),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_389),
.A2(n_338),
.B1(n_334),
.B2(n_346),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_333),
.A2(n_293),
.B1(n_255),
.B2(n_301),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_SL g391 ( 
.A(n_309),
.B(n_293),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_391),
.B(n_394),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_331),
.B(n_343),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_398),
.B1(n_415),
.B2(n_390),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_363),
.A2(n_336),
.B1(n_337),
.B2(n_332),
.Y(n_398)
);

OA21x2_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_345),
.B(n_354),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_399),
.B(n_373),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_336),
.B(n_352),
.Y(n_402)
);

AOI21xp33_ASAP7_75t_L g455 ( 
.A1(n_402),
.A2(n_408),
.B(n_412),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_336),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_410),
.Y(n_447)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_358),
.Y(n_404)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_404),
.Y(n_450)
);

OAI21x1_ASAP7_75t_R g405 ( 
.A1(n_387),
.A2(n_330),
.B(n_339),
.Y(n_405)
);

AOI21xp5_ASAP7_75t_L g457 ( 
.A1(n_405),
.A2(n_414),
.B(n_424),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_313),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_406),
.A2(n_413),
.B1(n_425),
.B2(n_428),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_376),
.A2(n_347),
.B(n_335),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_320),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_368),
.Y(n_448)
);

OAI21xp5_ASAP7_75t_L g412 ( 
.A1(n_383),
.A2(n_317),
.B(n_319),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_384),
.B(n_348),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_383),
.A2(n_315),
.B(n_326),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_356),
.A2(n_315),
.B1(n_325),
.B2(n_342),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_356),
.B(n_344),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_417),
.C(n_419),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_367),
.B(n_321),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_371),
.B(n_326),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_373),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_420),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_379),
.B(n_330),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_422),
.B(n_426),
.C(n_427),
.Y(n_434)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_358),
.Y(n_423)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_423),
.Y(n_431)
);

AOI211xp5_ASAP7_75t_SL g424 ( 
.A1(n_369),
.A2(n_330),
.B(n_311),
.C(n_325),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_372),
.A2(n_311),
.B1(n_9),
.B2(n_10),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_361),
.B(n_311),
.C(n_10),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_366),
.B(n_6),
.C(n_10),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_389),
.A2(n_15),
.B1(n_12),
.B2(n_13),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_365),
.Y(n_429)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_429),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_396),
.B(n_368),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_403),
.Y(n_461)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_396),
.B(n_374),
.C(n_365),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_435),
.B(n_417),
.C(n_410),
.Y(n_464)
);

OAI21xp5_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_399),
.B(n_414),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_437),
.A2(n_453),
.B1(n_454),
.B2(n_456),
.Y(n_468)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_400),
.Y(n_439)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_415),
.Y(n_440)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_440),
.Y(n_478)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_416),
.Y(n_442)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_442),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_421),
.A2(n_386),
.B1(n_374),
.B2(n_375),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_443),
.A2(n_449),
.B1(n_397),
.B2(n_399),
.Y(n_466)
);

CKINVDCx16_ASAP7_75t_R g444 ( 
.A(n_412),
.Y(n_444)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_444),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_364),
.Y(n_445)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_364),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_446),
.B(n_452),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_448),
.B(n_359),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_378),
.B1(n_382),
.B2(n_395),
.Y(n_449)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_425),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_451),
.Y(n_469)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_401),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g453 ( 
.A1(n_409),
.A2(n_391),
.B1(n_382),
.B2(n_393),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_408),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g456 ( 
.A1(n_398),
.A2(n_393),
.B1(n_392),
.B2(n_377),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_426),
.B(n_393),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g471 ( 
.A(n_458),
.B(n_459),
.Y(n_471)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_418),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g487 ( 
.A(n_461),
.B(n_480),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_437),
.A2(n_407),
.B1(n_405),
.B2(n_424),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_462),
.A2(n_457),
.B1(n_465),
.B2(n_469),
.Y(n_500)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_436),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_463),
.B(n_473),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_467),
.C(n_470),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g499 ( 
.A1(n_465),
.A2(n_457),
.B(n_456),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_466),
.A2(n_459),
.B1(n_440),
.B2(n_454),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_447),
.B(n_435),
.C(n_430),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_447),
.B(n_411),
.C(n_419),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_432),
.B(n_407),
.C(n_405),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_472),
.B(n_458),
.C(n_439),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_SL g473 ( 
.A(n_433),
.B(n_427),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_432),
.B(n_428),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_481),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g475 ( 
.A(n_446),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_475),
.B(n_452),
.Y(n_492)
);

INVx13_ASAP7_75t_L g476 ( 
.A(n_445),
.Y(n_476)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_476),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_479),
.B(n_442),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_448),
.B(n_392),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_455),
.B(n_392),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_485),
.A2(n_468),
.B1(n_462),
.B2(n_469),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_486),
.B(n_494),
.Y(n_506)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_477),
.Y(n_491)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_491),
.Y(n_522)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_492),
.Y(n_507)
);

CKINVDCx14_ASAP7_75t_R g493 ( 
.A(n_482),
.Y(n_493)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_493),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_467),
.B(n_449),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_434),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_495),
.B(n_497),
.C(n_503),
.Y(n_515)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_482),
.Y(n_496)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_496),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_461),
.B(n_434),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_471),
.Y(n_498)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_498),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g516 ( 
.A1(n_499),
.A2(n_504),
.B(n_476),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_466),
.B1(n_460),
.B2(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_471),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_501),
.B(n_484),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_460),
.A2(n_443),
.B(n_451),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_464),
.B(n_450),
.C(n_438),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_505),
.B(n_480),
.C(n_472),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_L g532 ( 
.A1(n_509),
.A2(n_511),
.B1(n_519),
.B2(n_489),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_510),
.A2(n_518),
.B1(n_509),
.B2(n_513),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_504),
.A2(n_478),
.B1(n_484),
.B2(n_483),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_512),
.A2(n_490),
.B1(n_502),
.B2(n_503),
.Y(n_523)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_505),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_514),
.B(n_516),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_518),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_500),
.Y(n_518)
);

AOI22xp5_ASAP7_75t_L g519 ( 
.A1(n_499),
.A2(n_481),
.B1(n_441),
.B2(n_470),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g520 ( 
.A(n_488),
.B(n_479),
.C(n_438),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_520),
.B(n_497),
.C(n_487),
.Y(n_527)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_523),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_525),
.A2(n_530),
.B1(n_535),
.B2(n_516),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_SL g526 ( 
.A1(n_514),
.A2(n_488),
.B(n_494),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_526),
.B(n_527),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_495),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_528),
.B(n_531),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_508),
.A2(n_489),
.B1(n_487),
.B2(n_431),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_507),
.B(n_431),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_532),
.B(n_524),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_515),
.B(n_486),
.C(n_377),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_533),
.B(n_534),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_517),
.B(n_385),
.C(n_12),
.Y(n_534)
);

AOI22xp5_ASAP7_75t_L g535 ( 
.A1(n_510),
.A2(n_385),
.B1(n_13),
.B2(n_14),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g537 ( 
.A(n_530),
.B(n_519),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_537),
.B(n_542),
.Y(n_548)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_541),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_525),
.A2(n_521),
.B1(n_511),
.B2(n_522),
.Y(n_542)
);

NOR2x1_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_520),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g549 ( 
.A(n_543),
.B(n_506),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_527),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_544),
.B(n_545),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_543),
.B(n_528),
.Y(n_546)
);

NAND3xp33_ASAP7_75t_L g555 ( 
.A(n_546),
.B(n_549),
.C(n_506),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g547 ( 
.A1(n_536),
.A2(n_538),
.B(n_544),
.Y(n_547)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_547),
.A2(n_535),
.B(n_545),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g550 ( 
.A(n_537),
.B(n_534),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g553 ( 
.A(n_550),
.B(n_540),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_553),
.B(n_554),
.Y(n_557)
);

OAI21xp33_ASAP7_75t_L g554 ( 
.A1(n_551),
.A2(n_539),
.B(n_541),
.Y(n_554)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_555),
.Y(n_558)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_558),
.A2(n_552),
.B(n_551),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_559),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g560 ( 
.A1(n_557),
.A2(n_556),
.B(n_548),
.Y(n_560)
);

AO21x1_ASAP7_75t_L g562 ( 
.A1(n_561),
.A2(n_560),
.B(n_385),
.Y(n_562)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_10),
.C(n_14),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_563),
.B(n_15),
.Y(n_564)
);


endmodule