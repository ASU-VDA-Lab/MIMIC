module fake_jpeg_26336_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx16f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_4),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_38),
.Y(n_51)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_20),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_42),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_21),
.Y(n_42)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_21),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_17),
.Y(n_59)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_32),
.Y(n_47)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g88 ( 
.A(n_54),
.Y(n_88)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_59),
.B(n_60),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

AO22x2_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_22),
.B1(n_33),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_61),
.A2(n_38),
.B1(n_37),
.B2(n_45),
.Y(n_97)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_34),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_63),
.B(n_48),
.Y(n_78)
);

OAI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_43),
.A2(n_44),
.B1(n_40),
.B2(n_46),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_66),
.A2(n_44),
.B1(n_47),
.B2(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_68),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_61),
.A2(n_35),
.B1(n_25),
.B2(n_46),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_70),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_44),
.B1(n_43),
.B2(n_46),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_75),
.B1(n_80),
.B2(n_53),
.Y(n_109)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_72),
.B(n_76),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_48),
.Y(n_73)
);

A2O1A1Ixp33_ASAP7_75t_L g106 ( 
.A1(n_73),
.A2(n_83),
.B(n_95),
.C(n_42),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_78),
.B(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_79),
.B(n_81),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_61),
.A2(n_45),
.B1(n_42),
.B2(n_25),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_39),
.Y(n_82)
);

NOR2xp67_ASAP7_75t_R g83 ( 
.A(n_64),
.B(n_59),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_50),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_85),
.Y(n_113)
);

INVx5_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g87 ( 
.A(n_67),
.B(n_48),
.Y(n_87)
);

NAND2xp33_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_19),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_65),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_49),
.Y(n_90)
);

HB1xp67_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_92),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_48),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_18),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_94),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_22),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_97),
.A2(n_55),
.B1(n_58),
.B2(n_62),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_83),
.A2(n_57),
.B1(n_54),
.B2(n_52),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_98),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_99),
.A2(n_117),
.B1(n_126),
.B2(n_88),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_93),
.Y(n_103)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_103),
.Y(n_132)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_104),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_125),
.B(n_115),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_121),
.B1(n_88),
.B2(n_95),
.Y(n_135)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_77),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_111),
.B(n_112),
.Y(n_148)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_114),
.B(n_73),
.C(n_87),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_85),
.A2(n_35),
.B1(n_27),
.B2(n_23),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_116),
.A2(n_27),
.B1(n_120),
.B2(n_105),
.Y(n_152)
);

AO22x1_ASAP7_75t_SL g117 ( 
.A1(n_81),
.A2(n_28),
.B1(n_34),
.B2(n_33),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_30),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_124),
.Y(n_130)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_82),
.B1(n_68),
.B2(n_72),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_122),
.A2(n_95),
.B(n_73),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_86),
.B(n_30),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_37),
.B1(n_31),
.B2(n_26),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_96),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_128),
.B(n_24),
.Y(n_184)
);

INVx13_ASAP7_75t_L g129 ( 
.A(n_104),
.Y(n_129)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_131),
.A2(n_150),
.B(n_151),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_101),
.B(n_90),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_133),
.B(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_113),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_135),
.A2(n_136),
.B1(n_142),
.B2(n_140),
.Y(n_159)
);

AO22x2_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_88),
.B1(n_74),
.B2(n_92),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_136),
.A2(n_142),
.B1(n_108),
.B2(n_127),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_99),
.Y(n_157)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_139),
.B(n_141),
.Y(n_170)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_105),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_74),
.B1(n_94),
.B2(n_34),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_30),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_144),
.B(n_145),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_122),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_34),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_146),
.B(n_147),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_112),
.B(n_100),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_17),
.B(n_23),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_152),
.A2(n_0),
.B(n_1),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_118),
.A2(n_33),
.B1(n_28),
.B2(n_19),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_117),
.B1(n_31),
.B2(n_26),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_33),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_154),
.Y(n_172)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_158),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_157),
.A2(n_161),
.B(n_174),
.Y(n_205)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_148),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_159),
.A2(n_168),
.B1(n_180),
.B2(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_163),
.Y(n_202)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_115),
.B(n_111),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_114),
.C(n_107),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_162),
.B(n_183),
.Y(n_190)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_132),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_165),
.B(n_173),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_136),
.Y(n_166)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_140),
.A2(n_108),
.B(n_107),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_167),
.A2(n_186),
.B(n_149),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_137),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_169),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_117),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_137),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_176),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_141),
.A2(n_117),
.B1(n_126),
.B2(n_19),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_130),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_178),
.B(n_139),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_24),
.B1(n_18),
.B2(n_31),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_24),
.A3(n_18),
.B1(n_26),
.B2(n_3),
.Y(n_181)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_181),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_131),
.B(n_24),
.C(n_18),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_162),
.Y(n_213)
);

FAx1_ASAP7_75t_SL g185 ( 
.A(n_153),
.B(n_10),
.CI(n_15),
.CON(n_185),
.SN(n_185)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_152),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_0),
.Y(n_187)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_187),
.Y(n_206)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_182),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_194),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_173),
.B1(n_161),
.B2(n_166),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_191),
.A2(n_197),
.B1(n_129),
.B2(n_0),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_193),
.B(n_208),
.Y(n_244)
);

INVx13_ASAP7_75t_L g194 ( 
.A(n_182),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_165),
.A2(n_187),
.B(n_175),
.Y(n_195)
);

NOR3xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_183),
.C(n_179),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_169),
.Y(n_196)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_135),
.B1(n_142),
.B2(n_134),
.Y(n_197)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_198),
.A2(n_180),
.B1(n_135),
.B2(n_185),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g203 ( 
.A1(n_167),
.A2(n_135),
.B(n_1),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_209),
.B(n_160),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_207),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_137),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_172),
.B(n_149),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_211),
.Y(n_228)
);

INVx13_ASAP7_75t_L g211 ( 
.A(n_170),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_212),
.B(n_216),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_129),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_156),
.B(n_143),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_214),
.B(n_219),
.Y(n_234)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_168),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_217),
.B(n_218),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_186),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_178),
.B(n_143),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_220),
.A2(n_221),
.B1(n_243),
.B2(n_245),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_179),
.B(n_158),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_222),
.A2(n_232),
.B(n_233),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_241),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_188),
.B(n_184),
.Y(n_224)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_224),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_181),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_226),
.B(n_230),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_201),
.A2(n_185),
.B(n_0),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_229),
.A2(n_239),
.B(n_5),
.Y(n_263)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_202),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_191),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_207),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_235),
.B(n_211),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_139),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_236),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_209),
.A2(n_11),
.B(n_2),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_240),
.B(n_190),
.C(n_213),
.Y(n_250)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_192),
.Y(n_258)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_197),
.B(n_2),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_232),
.A2(n_201),
.B1(n_218),
.B2(n_199),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_246),
.A2(n_227),
.B1(n_229),
.B2(n_239),
.Y(n_274)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_244),
.Y(n_269)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_225),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_251),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_190),
.C(n_205),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_257),
.C(n_262),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_255),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_233),
.A2(n_216),
.B1(n_199),
.B2(n_192),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_254),
.B(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_228),
.B(n_206),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_237),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_224),
.B(n_206),
.C(n_198),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_263),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_237),
.A2(n_200),
.B1(n_204),
.B2(n_196),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_259),
.B(n_245),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_204),
.C(n_200),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_189),
.C(n_196),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_265),
.B(n_227),
.C(n_231),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_270),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_222),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_221),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_SL g293 ( 
.A(n_273),
.B(n_275),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_274),
.A2(n_278),
.B1(n_220),
.B2(n_194),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_SL g275 ( 
.A(n_257),
.B(n_226),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_277),
.B(n_6),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_238),
.B1(n_231),
.B2(n_242),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_262),
.B(n_238),
.C(n_243),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_279),
.B(n_247),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_253),
.B(n_236),
.Y(n_280)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_280),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_245),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_282),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_260),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_8),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_284),
.A2(n_249),
.B(n_251),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_299),
.C(n_296),
.Y(n_301)
);

AOI22x1_ASAP7_75t_R g286 ( 
.A1(n_275),
.A2(n_246),
.B1(n_263),
.B2(n_256),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_294),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_261),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_289),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_296),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_271),
.A2(n_220),
.B(n_8),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_267),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_297),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_283),
.A2(n_220),
.B(n_8),
.Y(n_296)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_281),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_300),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_268),
.B(n_9),
.Y(n_300)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_301),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_276),
.C(n_269),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_302),
.B(n_304),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_292),
.B(n_270),
.C(n_273),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_293),
.B(n_281),
.C(n_10),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_307),
.B(n_311),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_293),
.B(n_9),
.C(n_10),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_287),
.C(n_299),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_312),
.B(n_313),
.C(n_298),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_9),
.C(n_11),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_314),
.B(n_303),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_12),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_317),
.B(n_318),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_308),
.B(n_309),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_305),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_319),
.B(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_305),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_306),
.A2(n_12),
.B(n_13),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_321),
.B(n_310),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_323),
.A2(n_329),
.B(n_14),
.Y(n_330)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_324),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_328),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g328 ( 
.A1(n_322),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_315),
.A2(n_16),
.B(n_13),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_330),
.B(n_317),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_L g334 ( 
.A1(n_333),
.A2(n_326),
.B(n_314),
.C(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_331),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_325),
.B(n_328),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_318),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_16),
.Y(n_339)
);


endmodule