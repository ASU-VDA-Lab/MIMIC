module real_jpeg_19528_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_321, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;
input n_321;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_0),
.A2(n_47),
.B1(n_49),
.B2(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_68),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_0),
.A2(n_32),
.B1(n_33),
.B2(n_68),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_26),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_1),
.A2(n_36),
.B1(n_63),
.B2(n_64),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_1),
.A2(n_36),
.B1(n_47),
.B2(n_49),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_2),
.A2(n_47),
.B1(n_49),
.B2(n_160),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_2),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_2),
.A2(n_63),
.B1(n_64),
.B2(n_160),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_2),
.A2(n_32),
.B1(n_33),
.B2(n_160),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_2),
.A2(n_26),
.B1(n_35),
.B2(n_160),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_3),
.A2(n_47),
.B1(n_49),
.B2(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_3),
.A2(n_26),
.B1(n_35),
.B2(n_52),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_3),
.A2(n_52),
.B1(n_63),
.B2(n_64),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_4),
.A2(n_26),
.B1(n_35),
.B2(n_131),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_4),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_4),
.A2(n_63),
.B1(n_64),
.B2(n_131),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_47),
.B1(n_49),
.B2(n_131),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_131),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g145 ( 
.A1(n_5),
.A2(n_49),
.B(n_59),
.C(n_146),
.D(n_147),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_5),
.B(n_49),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_5),
.B(n_46),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_5),
.Y(n_182)
);

OAI21xp33_ASAP7_75t_L g184 ( 
.A1(n_5),
.A2(n_82),
.B(n_165),
.Y(n_184)
);

A2O1A1O1Ixp25_ASAP7_75t_L g197 ( 
.A1(n_5),
.A2(n_32),
.B(n_43),
.C(n_198),
.D(n_199),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_5),
.B(n_32),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_133),
.Y(n_223)
);

AOI21xp33_ASAP7_75t_L g241 ( 
.A1(n_5),
.A2(n_31),
.B(n_33),
.Y(n_241)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_5),
.A2(n_26),
.B1(n_35),
.B2(n_182),
.Y(n_257)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_7),
.Y(n_83)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_7),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_7),
.B(n_166),
.Y(n_165)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_9),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_11),
.A2(n_26),
.B1(n_35),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_11),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_11),
.A2(n_47),
.B1(n_49),
.B2(n_92),
.Y(n_148)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_92),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g200 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_92),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_12),
.A2(n_26),
.B1(n_35),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_12),
.A2(n_32),
.B1(n_33),
.B2(n_38),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_12),
.A2(n_38),
.B1(n_47),
.B2(n_49),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_12),
.A2(n_38),
.B1(n_63),
.B2(n_64),
.Y(n_222)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_15),
.A2(n_32),
.B1(n_33),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_15),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_15),
.A2(n_47),
.B1(n_49),
.B2(n_55),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_15),
.A2(n_55),
.B1(n_63),
.B2(n_64),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_108),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_107),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_94),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_21),
.B(n_94),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.C(n_78),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_22),
.A2(n_70),
.B1(n_71),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_22),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_39),
.B2(n_40),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_23),
.A2(n_24),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_24),
.B(n_56),
.C(n_69),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_37),
.Y(n_24)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_30),
.B1(n_37),
.B2(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_25),
.A2(n_130),
.B(n_132),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_25),
.A2(n_30),
.B1(n_130),
.B2(n_266),
.Y(n_286)
);

A2O1A1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_28),
.Y(n_29)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g240 ( 
.A1(n_26),
.A2(n_28),
.B(n_182),
.C(n_241),
.Y(n_240)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_30),
.A2(n_34),
.B(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_30),
.Y(n_133)
);

OAI21xp33_ASAP7_75t_L g265 ( 
.A1(n_30),
.A2(n_90),
.B(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

O2A1O1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_44),
.B(n_45),
.C(n_46),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_44),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_56),
.B1(n_57),
.B2(n_69),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_41),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_50),
.B1(n_53),
.B2(n_54),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_42),
.A2(n_53),
.B1(n_54),
.B2(n_103),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_42),
.A2(n_53),
.B1(n_217),
.B2(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_42),
.A2(n_254),
.B(n_269),
.Y(n_268)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_43),
.A2(n_46),
.B1(n_51),
.B2(n_73),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_43),
.A2(n_46),
.B1(n_73),
.B2(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_43),
.B(n_219),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_44),
.B(n_49),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_45),
.A2(n_47),
.B1(n_205),
.B2(n_206),
.Y(n_204)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_60),
.B(n_61),
.C(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_60),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_53),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_53),
.A2(n_217),
.B(n_218),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_53),
.A2(n_218),
.B(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_56),
.A2(n_57),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_66),
.B(n_67),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_58),
.A2(n_66),
.B1(n_76),
.B2(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_58),
.A2(n_66),
.B1(n_87),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_58),
.A2(n_66),
.B1(n_159),
.B2(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_58),
.A2(n_196),
.B(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_58),
.A2(n_66),
.B1(n_125),
.B2(n_251),
.Y(n_274)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_62),
.B1(n_75),
.B2(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_59),
.B(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_60),
.A2(n_63),
.B1(n_64),
.B2(n_65),
.Y(n_62)
);

CKINVDCx9p33_ASAP7_75t_R g65 ( 
.A(n_60),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_60),
.B(n_64),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_61),
.A2(n_63),
.B1(n_151),
.B2(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_62),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g64 ( 
.A(n_63),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_64),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_66),
.B(n_148),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_66),
.A2(n_159),
.B(n_161),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_66),
.B(n_182),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_66),
.A2(n_161),
.B(n_251),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_72),
.B(n_74),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_78),
.B(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_88),
.B(n_89),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_79),
.A2(n_80),
.B1(n_112),
.B2(n_114),
.Y(n_111)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_86),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_81),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_113),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_81),
.A2(n_86),
.B1(n_88),
.B2(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_84),
.B(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_82),
.A2(n_85),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_82),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_82),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_82),
.A2(n_84),
.B1(n_208),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_82),
.A2(n_84),
.B1(n_222),
.B2(n_244),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_82),
.A2(n_121),
.B1(n_122),
.B2(n_244),
.Y(n_273)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_83),
.A2(n_171),
.B(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_84),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_84),
.B(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_86),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_93),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_93),
.A2(n_257),
.B(n_258),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_106),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_105),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g108 ( 
.A1(n_109),
.A2(n_137),
.B(n_319),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_134),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_110),
.B(n_134),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_115),
.C(n_117),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_111),
.A2(n_115),
.B1(n_116),
.B2(n_306),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_111),
.Y(n_306)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_112),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_117),
.A2(n_118),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_126),
.C(n_128),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_119),
.B(n_298),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_124),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_120),
.B(n_124),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_122),
.A2(n_180),
.B(n_208),
.Y(n_207)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_126),
.A2(n_128),
.B1(n_129),
.B2(n_299),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_126),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_127),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_132),
.Y(n_258)
);

AOI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_294),
.A3(n_307),
.B1(n_313),
.B2(n_318),
.C(n_321),
.Y(n_137)
);

NOR3xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_260),
.C(n_290),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_234),
.B(n_259),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_211),
.B(n_233),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_190),
.B(n_210),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_167),
.B(n_189),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_153),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_144),
.B(n_153),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_145),
.A2(n_149),
.B1(n_150),
.B2(n_176),
.Y(n_175)
);

CKINVDCx14_ASAP7_75t_R g176 ( 
.A(n_145),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_147),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_148),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_155),
.B(n_158),
.C(n_163),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_164),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_166),
.B(n_172),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_168),
.A2(n_177),
.B(n_188),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_175),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_175),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_172),
.B1(n_173),
.B2(n_174),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_183),
.B(n_187),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_181),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_179),
.B(n_181),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_185),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_192),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_191),
.B(n_192),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_193),
.A2(n_194),
.B1(n_203),
.B2(n_209),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_197),
.B1(n_201),
.B2(n_202),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_195),
.Y(n_202)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_197),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_202),
.C(n_209),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_198),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_199),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_200),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_203),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_207),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_207),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_212),
.B(n_213),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_227),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_229),
.C(n_231),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_220),
.B2(n_226),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_215),
.B(n_223),
.C(n_224),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_220),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_221),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_221),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_223),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_229),
.B1(n_231),
.B2(n_232),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_228),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_229),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_236),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_235),
.B(n_236),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_248),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_238),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_238),
.B(n_247),
.C(n_248),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B1(n_242),
.B2(n_243),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_239),
.B(n_243),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g247 ( 
.A(n_245),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_256),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_250),
.A2(n_252),
.B1(n_253),
.B2(n_255),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_250),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_255),
.C(n_256),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g314 ( 
.A1(n_261),
.A2(n_315),
.B(n_316),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_276),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_262),
.B(n_276),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_272),
.C(n_275),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_263),
.B(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_271),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_265),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_270),
.C(n_271),
.Y(n_288)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_272),
.B(n_275),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_273),
.B(n_274),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_288),
.B2(n_289),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_280),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_279),
.B(n_280),
.C(n_289),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_285),
.C(n_287),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_285),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_283),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_288),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_291),
.B(n_292),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_303),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_295),
.B(n_303),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_300),
.C(n_302),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_296),
.A2(n_297),
.B1(n_300),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_300),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_302),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_308),
.A2(n_314),
.B(n_317),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_309),
.B(n_310),
.Y(n_317)
);


endmodule