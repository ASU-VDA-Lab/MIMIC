module fake_jpeg_1809_n_680 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_680);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_680;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_574;
wire n_542;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_615;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_650;
wire n_328;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_1),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_18),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_14),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_9),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_4),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_61),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_9),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_62),
.B(n_73),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_63),
.Y(n_192)
);

NAND2x1_ASAP7_75t_SL g64 ( 
.A(n_29),
.B(n_9),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_64),
.B(n_0),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_28),
.Y(n_66)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_66),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_67),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_69),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_70),
.Y(n_216)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_72),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_74),
.Y(n_184)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_75),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_76),
.Y(n_202)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_56),
.Y(n_77)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_77),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_25),
.Y(n_78)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

INVx3_ASAP7_75t_SL g161 ( 
.A(n_79),
.Y(n_161)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_80),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_53),
.Y(n_81)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_81),
.Y(n_183)
);

BUFx24_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g155 ( 
.A(n_82),
.Y(n_155)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_28),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_50),
.B(n_10),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_84),
.B(n_91),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_85),
.A2(n_92),
.B1(n_54),
.B2(n_32),
.Y(n_167)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_25),
.Y(n_88)
);

INVx6_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_89),
.Y(n_162)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_31),
.Y(n_90)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_24),
.B(n_7),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_55),
.A2(n_10),
.B1(n_15),
.B2(n_13),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_19),
.Y(n_94)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_19),
.Y(n_95)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_95),
.Y(n_137)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_19),
.Y(n_96)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_97),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_98),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_99),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_30),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_100),
.B(n_45),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_27),
.Y(n_101)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_101),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_24),
.B(n_17),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_102),
.B(n_113),
.Y(n_164)
);

BUFx8_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_29),
.Y(n_104)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_35),
.Y(n_105)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_41),
.Y(n_106)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_106),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_27),
.Y(n_107)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_107),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_108),
.Y(n_150)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_109),
.Y(n_177)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_110),
.Y(n_170)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx6_ASAP7_75t_L g220 ( 
.A(n_112),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_42),
.B(n_17),
.Y(n_113)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_56),
.Y(n_116)
);

INVx8_ASAP7_75t_L g188 ( 
.A(n_116),
.Y(n_188)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_37),
.Y(n_117)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_117),
.Y(n_203)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_35),
.Y(n_118)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_118),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_119),
.Y(n_178)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_20),
.Y(n_120)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_120),
.Y(n_204)
);

INVx4_ASAP7_75t_SL g121 ( 
.A(n_39),
.Y(n_121)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_121),
.Y(n_194)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_20),
.Y(n_122)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_122),
.Y(n_205)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_30),
.Y(n_123)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_123),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_39),
.Y(n_124)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_124),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_39),
.Y(n_125)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_125),
.Y(n_213)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_60),
.Y(n_126)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_20),
.Y(n_127)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_20),
.Y(n_128)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_34),
.Y(n_129)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_129),
.Y(n_214)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_34),
.Y(n_130)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_34),
.Y(n_131)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_39),
.Y(n_132)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_45),
.B1(n_58),
.B2(n_57),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_133),
.A2(n_151),
.B1(n_169),
.B2(n_51),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_103),
.B(n_59),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_136),
.B(n_149),
.Y(n_285)
);

BUFx4f_ASAP7_75t_L g140 ( 
.A(n_103),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_140),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_121),
.A2(n_20),
.B1(n_58),
.B2(n_57),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_148),
.A2(n_154),
.B1(n_167),
.B2(n_186),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_66),
.B(n_59),
.Y(n_149)
);

OAI22xp33_ASAP7_75t_L g151 ( 
.A1(n_65),
.A2(n_69),
.B1(n_125),
.B2(n_124),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_123),
.A2(n_58),
.B1(n_57),
.B2(n_45),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_68),
.A2(n_58),
.B1(n_57),
.B2(n_45),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_64),
.B(n_32),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_171),
.B(n_191),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_181),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_116),
.B(n_44),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_182),
.B(n_187),
.Y(n_262)
);

OR2x4_ASAP7_75t_L g185 ( 
.A(n_82),
.B(n_42),
.Y(n_185)
);

NAND2x1_ASAP7_75t_SL g272 ( 
.A(n_185),
.B(n_208),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_130),
.A2(n_43),
.B1(n_33),
.B2(n_22),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_116),
.B(n_44),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_111),
.B(n_52),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_189),
.B(n_224),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_95),
.B(n_21),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_96),
.B(n_21),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_221),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_131),
.A2(n_43),
.B1(n_33),
.B2(n_22),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_201),
.A2(n_207),
.B1(n_211),
.B2(n_128),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_75),
.A2(n_106),
.B1(n_114),
.B2(n_110),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_97),
.A2(n_43),
.B1(n_33),
.B2(n_22),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_126),
.Y(n_215)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_63),
.B(n_52),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_72),
.Y(n_223)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_223),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_67),
.B(n_47),
.Y(n_224)
);

INVx11_ASAP7_75t_L g226 ( 
.A(n_144),
.Y(n_226)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_226),
.Y(n_349)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_227),
.Y(n_332)
);

AO22x2_ASAP7_75t_L g228 ( 
.A1(n_169),
.A2(n_82),
.B1(n_92),
.B2(n_54),
.Y(n_228)
);

OA22x2_ASAP7_75t_L g348 ( 
.A1(n_228),
.A2(n_233),
.B1(n_237),
.B2(n_292),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_79),
.Y(n_229)
);

CKINVDCx14_ASAP7_75t_R g318 ( 
.A(n_229),
.Y(n_318)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_140),
.A2(n_40),
.B1(n_38),
.B2(n_47),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_231),
.A2(n_234),
.B1(n_258),
.B2(n_265),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_194),
.A2(n_40),
.B1(n_38),
.B2(n_26),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_204),
.Y(n_235)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_235),
.Y(n_328)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_205),
.Y(n_236)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_236),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_153),
.A2(n_81),
.B1(n_119),
.B2(n_115),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_237),
.A2(n_168),
.B(n_202),
.Y(n_356)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_135),
.Y(n_238)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_238),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_161),
.Y(n_240)
);

INVxp33_ASAP7_75t_L g315 ( 
.A(n_240),
.Y(n_315)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_241),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_154),
.A2(n_76),
.B1(n_112),
.B2(n_107),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_242),
.A2(n_279),
.B1(n_293),
.B2(n_300),
.Y(n_320)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_135),
.Y(n_243)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_244),
.Y(n_341)
);

INVx4_ASAP7_75t_SL g245 ( 
.A(n_190),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_245),
.B(n_250),
.Y(n_306)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_170),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_246),
.Y(n_358)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_180),
.Y(n_247)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_174),
.Y(n_248)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_248),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_143),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_155),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_251),
.Y(n_338)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_222),
.Y(n_253)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_253),
.Y(n_351)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_178),
.Y(n_254)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_254),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_160),
.B(n_51),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_255),
.B(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_166),
.B(n_36),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_176),
.B(n_36),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_257),
.B(n_271),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_139),
.A2(n_40),
.B1(n_26),
.B2(n_54),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_155),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_259),
.B(n_263),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g261 ( 
.A(n_137),
.B(n_141),
.Y(n_261)
);

OAI21xp33_ASAP7_75t_L g354 ( 
.A1(n_261),
.A2(n_280),
.B(n_283),
.Y(n_354)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_156),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_264),
.Y(n_363)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_164),
.A2(n_70),
.B1(n_93),
.B2(n_217),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_143),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_267),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_158),
.B(n_138),
.C(n_162),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_268),
.B(n_179),
.C(n_150),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_142),
.B(n_74),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g361 ( 
.A(n_269),
.B(n_302),
.Y(n_361)
);

HB1xp67_ASAP7_75t_L g270 ( 
.A(n_163),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_270),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_147),
.B(n_0),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_133),
.A2(n_101),
.B1(n_99),
.B2(n_88),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_273),
.A2(n_276),
.B1(n_292),
.B2(n_211),
.Y(n_305)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_183),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_274),
.Y(n_312)
);

AOI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_275),
.A2(n_278),
.B1(n_290),
.B2(n_175),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_151),
.A2(n_127),
.B1(n_78),
.B2(n_43),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

OR2x2_ASAP7_75t_L g319 ( 
.A(n_277),
.B(n_284),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_209),
.A2(n_17),
.B1(n_15),
.B2(n_13),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_148),
.A2(n_12),
.B1(n_11),
.B2(n_2),
.Y(n_279)
);

A2O1A1Ixp33_ASAP7_75t_L g280 ( 
.A1(n_157),
.A2(n_12),
.B(n_11),
.C(n_2),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_165),
.B(n_0),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_281),
.B(n_304),
.Y(n_314)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_161),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_282),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_177),
.B(n_0),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_203),
.Y(n_284)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_286),
.Y(n_330)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_200),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_287),
.B(n_294),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_145),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_288),
.B(n_299),
.Y(n_310)
);

NAND2x1_ASAP7_75t_L g289 ( 
.A(n_196),
.B(n_0),
.Y(n_289)
);

OR2x2_ASAP7_75t_L g345 ( 
.A(n_289),
.B(n_291),
.Y(n_345)
);

INVx11_ASAP7_75t_L g290 ( 
.A(n_155),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_216),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_134),
.A2(n_11),
.B1(n_12),
.B2(n_3),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_186),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_146),
.Y(n_294)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_146),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_295),
.B(n_297),
.Y(n_365)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_188),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_296),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx6_ASAP7_75t_L g298 ( 
.A(n_134),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_298),
.Y(n_326)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_145),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_201),
.A2(n_6),
.B1(n_1),
.B2(n_5),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_188),
.B(n_5),
.Y(n_302)
);

INVx6_ASAP7_75t_L g303 ( 
.A(n_152),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_303),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_193),
.B(n_5),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_305),
.A2(n_329),
.B1(n_337),
.B2(n_344),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_307),
.B(n_322),
.C(n_327),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_L g311 ( 
.A1(n_260),
.A2(n_184),
.B1(n_202),
.B2(n_172),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_311),
.A2(n_360),
.B1(n_364),
.B2(n_291),
.Y(n_400)
);

NOR2x1_ASAP7_75t_R g313 ( 
.A(n_272),
.B(n_301),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_313),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_268),
.B(n_239),
.C(n_252),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_225),
.B(n_150),
.C(n_219),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_233),
.A2(n_220),
.B1(n_218),
.B2(n_212),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_271),
.B(n_281),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_336),
.B(n_353),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_273),
.A2(n_220),
.B1(n_218),
.B2(n_212),
.Y(n_337)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_339),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_242),
.A2(n_179),
.B1(n_207),
.B2(n_152),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_342),
.A2(n_266),
.B(n_296),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_228),
.A2(n_159),
.B1(n_206),
.B2(n_172),
.Y(n_344)
);

AND2x2_ASAP7_75t_SL g347 ( 
.A(n_283),
.B(n_184),
.Y(n_347)
);

CKINVDCx14_ASAP7_75t_R g384 ( 
.A(n_347),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_348),
.A2(n_359),
.B1(n_286),
.B2(n_251),
.Y(n_409)
);

OA21x2_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_193),
.B(n_206),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_350),
.A2(n_261),
.B(n_266),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_285),
.B(n_159),
.Y(n_353)
);

CKINVDCx14_ASAP7_75t_R g398 ( 
.A(n_356),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_255),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_357),
.B(n_229),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_228),
.A2(n_168),
.B1(n_5),
.B2(n_6),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g360 ( 
.A1(n_256),
.A2(n_6),
.B1(n_257),
.B2(n_228),
.Y(n_360)
);

OA22x2_ASAP7_75t_L g362 ( 
.A1(n_228),
.A2(n_6),
.B1(n_289),
.B2(n_284),
.Y(n_362)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_280),
.A2(n_283),
.B1(n_272),
.B2(n_262),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_367),
.B(n_380),
.Y(n_423)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_330),
.Y(n_369)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_305),
.A2(n_290),
.B1(n_227),
.B2(n_247),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_370),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_309),
.B(n_229),
.Y(n_371)
);

MAJx2_ASAP7_75t_L g417 ( 
.A(n_371),
.B(n_347),
.C(n_361),
.Y(n_417)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_341),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_373),
.B(n_375),
.Y(n_416)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_374),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_358),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_320),
.A2(n_299),
.B1(n_303),
.B2(n_298),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_376),
.A2(n_391),
.B1(n_397),
.B2(n_400),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_312),
.Y(n_377)
);

CKINVDCx14_ASAP7_75t_R g418 ( 
.A(n_377),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_297),
.C(n_261),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_378),
.B(n_411),
.C(n_318),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_306),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_241),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_382),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_312),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_383),
.A2(n_395),
.B(n_408),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_309),
.B(n_244),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_385),
.B(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_386),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_238),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g456 ( 
.A(n_387),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_314),
.B(n_232),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_320),
.A2(n_232),
.B1(n_248),
.B2(n_246),
.Y(n_391)
);

OA21x2_ASAP7_75t_R g392 ( 
.A1(n_331),
.A2(n_235),
.B(n_236),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_392),
.B(n_402),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_314),
.B(n_243),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_393),
.B(n_396),
.Y(n_430)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_316),
.Y(n_394)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_394),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g395 ( 
.A1(n_345),
.A2(n_254),
.B(n_287),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_331),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_348),
.A2(n_264),
.B1(n_277),
.B2(n_230),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_405),
.Y(n_438)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_323),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_348),
.A2(n_362),
.B1(n_364),
.B2(n_345),
.Y(n_403)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_403),
.A2(n_407),
.B1(n_319),
.B2(n_324),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_330),
.Y(n_404)
);

INVxp33_ASAP7_75t_SL g455 ( 
.A(n_404),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_306),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g407 ( 
.A1(n_348),
.A2(n_362),
.B1(n_345),
.B2(n_342),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_L g408 ( 
.A1(n_354),
.A2(n_274),
.B(n_253),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g431 ( 
.A1(n_409),
.A2(n_388),
.B1(n_344),
.B2(n_350),
.Y(n_431)
);

INVx5_ASAP7_75t_SL g410 ( 
.A(n_330),
.Y(n_410)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_410),
.B(n_349),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_307),
.B(n_230),
.C(n_245),
.Y(n_411)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_332),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_317),
.Y(n_444)
);

CKINVDCx16_ASAP7_75t_R g413 ( 
.A(n_319),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_413),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_414),
.A2(n_356),
.B(n_350),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_335),
.A2(n_240),
.B(n_294),
.Y(n_415)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_415),
.A2(n_383),
.B(n_414),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_417),
.B(n_424),
.Y(n_477)
);

OAI22x1_ASAP7_75t_SL g419 ( 
.A1(n_406),
.A2(n_348),
.B1(n_362),
.B2(n_359),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_419),
.A2(n_431),
.B1(n_435),
.B2(n_441),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_420),
.B(n_432),
.Y(n_485)
);

AND2x2_ASAP7_75t_SL g422 ( 
.A(n_403),
.B(n_407),
.Y(n_422)
);

CKINVDCx16_ASAP7_75t_R g492 ( 
.A(n_422),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_368),
.B(n_327),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_313),
.C(n_353),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_378),
.B(n_347),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_434),
.B(n_445),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_409),
.A2(n_362),
.B1(n_347),
.B2(n_329),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g483 ( 
.A1(n_439),
.A2(n_448),
.B(n_452),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_406),
.A2(n_350),
.B1(n_337),
.B2(n_319),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_442),
.A2(n_446),
.B1(n_450),
.B2(n_408),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_444),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_371),
.B(n_321),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_388),
.A2(n_310),
.B1(n_326),
.B2(n_355),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_375),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_447),
.B(n_373),
.Y(n_468)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_398),
.A2(n_326),
.B1(n_355),
.B2(n_324),
.Y(n_450)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_451),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_390),
.A2(n_321),
.B(n_365),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_411),
.B(n_323),
.C(n_363),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_453),
.B(n_434),
.Y(n_486)
);

AO22x1_ASAP7_75t_SL g454 ( 
.A1(n_397),
.A2(n_363),
.B1(n_352),
.B2(n_325),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_454),
.B(n_391),
.Y(n_457)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_457),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_445),
.B(n_424),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_459),
.B(n_486),
.C(n_417),
.Y(n_513)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_416),
.Y(n_460)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_460),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_396),
.Y(n_461)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_461),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_448),
.A2(n_415),
.B(n_398),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_SL g511 ( 
.A1(n_463),
.A2(n_471),
.B(n_474),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_430),
.B(n_374),
.Y(n_464)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_464),
.Y(n_508)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_416),
.Y(n_465)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_465),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_456),
.B(n_379),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_480),
.Y(n_501)
);

INVxp67_ASAP7_75t_SL g519 ( 
.A(n_468),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_436),
.B(n_372),
.Y(n_469)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_469),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_392),
.B1(n_384),
.B2(n_400),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g496 ( 
.A1(n_470),
.A2(n_472),
.B1(n_482),
.B2(n_484),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_437),
.A2(n_399),
.B(n_395),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_442),
.A2(n_384),
.B1(n_379),
.B2(n_381),
.Y(n_472)
);

BUFx2_ASAP7_75t_L g473 ( 
.A(n_429),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_473),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_441),
.A2(n_405),
.B1(n_380),
.B2(n_413),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_436),
.B(n_385),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_476),
.B(n_478),
.Y(n_512)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_449),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_440),
.B(n_389),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_479),
.B(n_481),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_440),
.B(n_387),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_418),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_433),
.A2(n_380),
.B1(n_405),
.B2(n_393),
.Y(n_484)
);

AOI22xp33_ASAP7_75t_L g487 ( 
.A1(n_439),
.A2(n_367),
.B1(n_386),
.B2(n_394),
.Y(n_487)
);

OAI22x1_ASAP7_75t_L g505 ( 
.A1(n_487),
.A2(n_489),
.B1(n_423),
.B2(n_438),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g488 ( 
.A(n_429),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_488),
.Y(n_499)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_428),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_490),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_419),
.A2(n_376),
.B1(n_402),
.B2(n_382),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g517 ( 
.A1(n_491),
.A2(n_433),
.B1(n_426),
.B2(n_422),
.Y(n_517)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_426),
.Y(n_493)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_493),
.A2(n_494),
.B(n_452),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_453),
.B(n_366),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_420),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_495),
.B(n_500),
.Y(n_539)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_486),
.B(n_432),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g504 ( 
.A1(n_483),
.A2(n_437),
.B(n_423),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_SL g536 ( 
.A1(n_504),
.A2(n_514),
.B(n_529),
.Y(n_536)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_505),
.Y(n_551)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_485),
.B(n_417),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_506),
.B(n_513),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g507 ( 
.A1(n_475),
.A2(n_450),
.B(n_454),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_507),
.B(n_489),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_475),
.A2(n_435),
.B1(n_446),
.B2(n_443),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g538 ( 
.A1(n_509),
.A2(n_518),
.B1(n_530),
.B2(n_491),
.Y(n_538)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_483),
.A2(n_438),
.B(n_425),
.Y(n_514)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_515),
.Y(n_554)
);

AOI22xp5_ASAP7_75t_L g544 ( 
.A1(n_517),
.A2(n_522),
.B1(n_492),
.B2(n_465),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_470),
.A2(n_443),
.B1(n_422),
.B2(n_427),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g520 ( 
.A(n_485),
.B(n_427),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_520),
.B(n_478),
.Y(n_561)
);

OAI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_474),
.A2(n_422),
.B1(n_425),
.B2(n_421),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_458),
.B(n_365),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_523),
.B(n_524),
.C(n_526),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_458),
.B(n_447),
.C(n_454),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_468),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_525),
.B(n_527),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_477),
.B(n_454),
.C(n_444),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_469),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g529 ( 
.A1(n_471),
.A2(n_451),
.B(n_455),
.Y(n_529)
);

AOI22xp5_ASAP7_75t_L g530 ( 
.A1(n_484),
.A2(n_451),
.B1(n_410),
.B2(n_401),
.Y(n_530)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_529),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_531),
.B(n_550),
.Y(n_574)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_521),
.Y(n_532)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_532),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_500),
.B(n_477),
.C(n_460),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_534),
.B(n_545),
.C(n_547),
.Y(n_578)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_535),
.Y(n_573)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_521),
.Y(n_537)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_537),
.Y(n_571)
);

AOI22xp5_ASAP7_75t_L g567 ( 
.A1(n_538),
.A2(n_496),
.B1(n_517),
.B2(n_535),
.Y(n_567)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_540),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_505),
.B(n_504),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_541),
.A2(n_536),
.B(n_511),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_519),
.B(n_464),
.Y(n_543)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_543),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_SL g565 ( 
.A1(n_544),
.A2(n_509),
.B1(n_530),
.B2(n_498),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_495),
.B(n_472),
.C(n_493),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_512),
.Y(n_546)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_546),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_513),
.B(n_463),
.C(n_467),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_506),
.B(n_467),
.C(n_461),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_549),
.B(n_562),
.C(n_503),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_510),
.B(n_476),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_510),
.B(n_479),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_553),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_508),
.B(n_481),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g555 ( 
.A(n_528),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_555),
.B(n_502),
.Y(n_577)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_516),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_556),
.B(n_557),
.Y(n_564)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_516),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_508),
.B(n_490),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_560),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g559 ( 
.A(n_523),
.B(n_462),
.Y(n_559)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_559),
.B(n_561),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_497),
.B(n_457),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_520),
.B(n_482),
.C(n_462),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_501),
.B(n_473),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g589 ( 
.A(n_563),
.B(n_473),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_SL g610 ( 
.A1(n_565),
.A2(n_573),
.B1(n_571),
.B2(n_570),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_499),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_566),
.B(n_583),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_567),
.A2(n_585),
.B1(n_546),
.B2(n_553),
.Y(n_606)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_539),
.B(n_524),
.Y(n_572)
);

XOR2xp5_ASAP7_75t_L g599 ( 
.A(n_572),
.B(n_575),
.Y(n_599)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_539),
.B(n_526),
.Y(n_575)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_577),
.Y(n_598)
);

XOR2x2_ASAP7_75t_L g594 ( 
.A(n_579),
.B(n_587),
.Y(n_594)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_514),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g602 ( 
.A(n_580),
.B(n_536),
.Y(n_602)
);

FAx1_ASAP7_75t_SL g581 ( 
.A(n_549),
.B(n_503),
.CI(n_522),
.CON(n_581),
.SN(n_581)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_581),
.B(n_559),
.Y(n_596)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_532),
.A2(n_537),
.B1(n_556),
.B2(n_557),
.Y(n_585)
);

OAI21xp5_ASAP7_75t_SL g587 ( 
.A1(n_541),
.A2(n_507),
.B(n_518),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g588 ( 
.A(n_533),
.B(n_507),
.C(n_498),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_588),
.B(n_590),
.Y(n_597)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_589),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g590 ( 
.A(n_533),
.B(n_412),
.C(n_340),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g591 ( 
.A1(n_567),
.A2(n_544),
.B1(n_551),
.B2(n_540),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_591),
.A2(n_606),
.B1(n_568),
.B2(n_589),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_590),
.B(n_534),
.C(n_545),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_592),
.B(n_595),
.Y(n_614)
);

MAJIxp5_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_548),
.C(n_562),
.Y(n_595)
);

MAJx2_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_602),
.C(n_315),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_588),
.B(n_578),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_600),
.B(n_564),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_572),
.B(n_548),
.C(n_561),
.Y(n_601)
);

MAJIxp5_ASAP7_75t_L g615 ( 
.A(n_601),
.B(n_604),
.C(n_574),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_578),
.B(n_580),
.C(n_575),
.Y(n_604)
);

XOR2xp5_ASAP7_75t_L g605 ( 
.A(n_569),
.B(n_531),
.Y(n_605)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_605),
.B(n_607),
.Y(n_619)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_569),
.B(n_579),
.Y(n_607)
);

NOR2xp33_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_542),
.Y(n_608)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_608),
.Y(n_616)
);

XOR2xp5_ASAP7_75t_L g609 ( 
.A(n_587),
.B(n_543),
.Y(n_609)
);

XOR2xp5_ASAP7_75t_L g628 ( 
.A(n_609),
.B(n_369),
.Y(n_628)
);

OAI22xp5_ASAP7_75t_SL g631 ( 
.A1(n_610),
.A2(n_404),
.B1(n_340),
.B2(n_317),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_576),
.B(n_563),
.Y(n_611)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_611),
.Y(n_617)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_573),
.A2(n_560),
.B1(n_552),
.B2(n_550),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_612),
.B(n_613),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_586),
.B(n_565),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_615),
.B(n_620),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_594),
.A2(n_574),
.B(n_585),
.Y(n_618)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_618),
.B(n_621),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g621 ( 
.A1(n_609),
.A2(n_582),
.B(n_581),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_SL g622 ( 
.A1(n_598),
.A2(n_582),
.B1(n_558),
.B2(n_581),
.Y(n_622)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_622),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g646 ( 
.A1(n_623),
.A2(n_603),
.B1(n_607),
.B2(n_605),
.Y(n_646)
);

INVx6_ASAP7_75t_L g624 ( 
.A(n_593),
.Y(n_624)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_624),
.B(n_631),
.Y(n_635)
);

OAI21xp5_ASAP7_75t_L g625 ( 
.A1(n_610),
.A2(n_568),
.B(n_377),
.Y(n_625)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_625),
.A2(n_594),
.B(n_596),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_598),
.B(n_488),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_626),
.B(n_630),
.Y(n_641)
);

XOR2xp5_ASAP7_75t_L g639 ( 
.A(n_628),
.B(n_629),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g630 ( 
.A(n_595),
.B(n_404),
.C(n_332),
.Y(n_630)
);

MAJIxp5_ASAP7_75t_L g632 ( 
.A(n_597),
.B(n_338),
.C(n_351),
.Y(n_632)
);

HB1xp67_ASAP7_75t_L g633 ( 
.A(n_632),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g636 ( 
.A(n_614),
.B(n_604),
.C(n_592),
.Y(n_636)
);

NOR2xp67_ASAP7_75t_SL g651 ( 
.A(n_636),
.B(n_637),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_615),
.B(n_602),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_624),
.B(n_616),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_638),
.B(n_645),
.Y(n_656)
);

AOI21x1_ASAP7_75t_L g655 ( 
.A1(n_642),
.A2(n_625),
.B(n_629),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g644 ( 
.A(n_617),
.B(n_601),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_644),
.B(n_619),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g645 ( 
.A(n_627),
.B(n_591),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_646),
.B(n_647),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_619),
.B(n_599),
.C(n_603),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_627),
.B(n_599),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_648),
.B(n_308),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_636),
.B(n_630),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_649),
.B(n_650),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_SL g650 ( 
.A(n_634),
.B(n_637),
.Y(n_650)
);

OAI21xp5_ASAP7_75t_SL g652 ( 
.A1(n_640),
.A2(n_618),
.B(n_621),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_652),
.A2(n_657),
.B(n_659),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g663 ( 
.A1(n_653),
.A2(n_654),
.B(n_655),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_641),
.B(n_632),
.Y(n_654)
);

OAI21xp5_ASAP7_75t_SL g657 ( 
.A1(n_642),
.A2(n_623),
.B(n_628),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_633),
.B(n_631),
.C(n_346),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_660),
.B(n_639),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_656),
.A2(n_635),
.B(n_647),
.C(n_646),
.Y(n_662)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_662),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_664),
.B(n_325),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g665 ( 
.A1(n_651),
.A2(n_658),
.B(n_643),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_SL g670 ( 
.A1(n_665),
.A2(n_667),
.B(n_668),
.Y(n_670)
);

OAI21xp5_ASAP7_75t_SL g667 ( 
.A1(n_655),
.A2(n_643),
.B(n_639),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_SL g668 ( 
.A1(n_659),
.A2(n_410),
.B(n_352),
.Y(n_668)
);

HB1xp67_ASAP7_75t_L g669 ( 
.A(n_666),
.Y(n_669)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_669),
.B(n_671),
.C(n_673),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g673 ( 
.A(n_663),
.B(n_351),
.C(n_338),
.Y(n_673)
);

A2O1A1O1Ixp25_ASAP7_75t_L g674 ( 
.A1(n_672),
.A2(n_661),
.B(n_334),
.C(n_328),
.D(n_343),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g677 ( 
.A1(n_674),
.A2(n_676),
.B(n_349),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g676 ( 
.A1(n_670),
.A2(n_328),
.B(n_334),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g678 ( 
.A(n_677),
.B(n_675),
.C(n_266),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_678),
.B(n_343),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_679),
.A2(n_282),
.B(n_226),
.Y(n_680)
);


endmodule