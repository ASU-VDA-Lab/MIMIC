module fake_jpeg_11974_n_351 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_351);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_10),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g110 ( 
.A(n_43),
.Y(n_110)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_22),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g89 ( 
.A(n_44),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_18),
.B(n_42),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_27),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_22),
.Y(n_49)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_68),
.Y(n_87)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_55),
.Y(n_88)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_18),
.B(n_8),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_57),
.B(n_42),
.Y(n_71)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_60),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_61),
.Y(n_83)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_62),
.Y(n_117)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_64),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_69),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_36),
.Y(n_70)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_71),
.B(n_78),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_19),
.B1(n_34),
.B2(n_40),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_112),
.B1(n_34),
.B2(n_38),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_43),
.B(n_30),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_74),
.A2(n_106),
.B(n_28),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_70),
.A2(n_41),
.B1(n_37),
.B2(n_25),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_77),
.A2(n_82),
.B1(n_96),
.B2(n_38),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_23),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_81),
.B(n_85),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_41),
.B1(n_37),
.B2(n_25),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_67),
.B(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_45),
.B(n_21),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_91),
.B(n_92),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_95),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_39),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_53),
.A2(n_41),
.B1(n_37),
.B2(n_25),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_39),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_99),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_35),
.Y(n_99)
);

NAND2x1_ASAP7_75t_L g101 ( 
.A(n_56),
.B(n_40),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_31),
.C(n_32),
.Y(n_124)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_60),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_103),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_61),
.B(n_35),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_104),
.B(n_109),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_65),
.B(n_30),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_30),
.Y(n_131)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_45),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_47),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_45),
.A2(n_34),
.B1(n_40),
.B2(n_26),
.Y(n_112)
);

INVx11_ASAP7_75t_L g115 ( 
.A(n_51),
.Y(n_115)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

HB1xp67_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_122),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_123),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_124),
.B(n_131),
.Y(n_168)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_125),
.Y(n_188)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_126),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_129),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_130),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_105),
.A2(n_23),
.B1(n_32),
.B2(n_24),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_132),
.A2(n_138),
.B(n_156),
.Y(n_177)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_118),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_135),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_31),
.B1(n_24),
.B2(n_30),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g181 ( 
.A(n_137),
.B(n_117),
.Y(n_181)
);

NAND2xp33_ASAP7_75t_SL g138 ( 
.A(n_78),
.B(n_30),
.Y(n_138)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_84),
.B1(n_80),
.B2(n_83),
.Y(n_174)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_141),
.B(n_147),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_73),
.A2(n_26),
.B1(n_28),
.B2(n_10),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_151),
.B1(n_86),
.B2(n_113),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_28),
.A3(n_8),
.B1(n_11),
.B2(n_16),
.Y(n_145)
);

AOI32xp33_ASAP7_75t_L g191 ( 
.A1(n_145),
.A2(n_98),
.A3(n_88),
.B1(n_13),
.B2(n_4),
.Y(n_191)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_89),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_146),
.Y(n_165)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_100),
.Y(n_147)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_76),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_148),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g149 ( 
.A(n_101),
.B(n_0),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_0),
.Y(n_163)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_150),
.B(n_153),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_112),
.A2(n_28),
.B1(n_11),
.B2(n_12),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_110),
.B(n_7),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_152),
.B(n_155),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_13),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_110),
.B(n_7),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_74),
.B(n_0),
.Y(n_156)
);

BUFx4f_ASAP7_75t_SL g157 ( 
.A(n_103),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_157),
.Y(n_195)
);

O2A1O1Ixp33_ASAP7_75t_SL g160 ( 
.A1(n_144),
.A2(n_111),
.B(n_76),
.C(n_79),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g216 ( 
.A1(n_160),
.A2(n_170),
.B(n_176),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_163),
.B(n_164),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_114),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_166),
.B(n_178),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_127),
.B(n_121),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_167),
.B(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_140),
.A2(n_132),
.B1(n_133),
.B2(n_124),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_114),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_84),
.B1(n_80),
.B2(n_83),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_173),
.A2(n_175),
.B1(n_190),
.B2(n_191),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_174),
.B(n_160),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_156),
.A2(n_72),
.B1(n_113),
.B2(n_86),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_72),
.B1(n_117),
.B2(n_79),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_149),
.B(n_131),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_142),
.B(n_157),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_196),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_145),
.A2(n_111),
.B1(n_98),
.B2(n_88),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g212 ( 
.A1(n_184),
.A2(n_187),
.B1(n_142),
.B2(n_157),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_131),
.A2(n_98),
.B1(n_88),
.B2(n_28),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_0),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_126),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_134),
.A2(n_148),
.B1(n_119),
.B2(n_135),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_146),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_197),
.B(n_213),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_168),
.B(n_122),
.C(n_153),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_198),
.B(n_181),
.C(n_168),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_158),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_199),
.B(n_201),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_158),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_139),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_206),
.Y(n_248)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_193),
.Y(n_204)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_204),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_214),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_1),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_207),
.A2(n_215),
.B(n_230),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_163),
.B(n_1),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_211),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_212),
.A2(n_181),
.B1(n_164),
.B2(n_195),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_192),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_165),
.B(n_6),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g215 ( 
.A1(n_178),
.A2(n_177),
.B(n_161),
.C(n_183),
.D(n_168),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_217),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_159),
.B(n_12),
.Y(n_220)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_220),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g221 ( 
.A1(n_161),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_221),
.A2(n_223),
.B1(n_174),
.B2(n_184),
.Y(n_232)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_171),
.Y(n_222)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_222),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_2),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_169),
.Y(n_225)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_186),
.B(n_14),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_226),
.B(n_228),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_3),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_227),
.B(n_209),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_179),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_177),
.B(n_14),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_232),
.A2(n_256),
.B(n_214),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_233),
.A2(n_216),
.B1(n_223),
.B2(n_215),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_242),
.C(n_243),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_216),
.A2(n_173),
.B1(n_191),
.B2(n_160),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_241),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_176),
.B1(n_182),
.B2(n_194),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_190),
.C(n_159),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_203),
.B(n_185),
.C(n_182),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_185),
.A3(n_169),
.B1(n_195),
.B2(n_188),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_216),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_198),
.B(n_188),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_202),
.C(n_205),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_200),
.B(n_16),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_200),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_207),
.A2(n_3),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_218),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_247),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_258),
.B(n_265),
.Y(n_294)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_237),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_260),
.B(n_264),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_263),
.A2(n_234),
.B1(n_256),
.B2(n_233),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_269),
.C(n_275),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_208),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_267),
.B(n_273),
.Y(n_292)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_245),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_268),
.B(n_271),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_218),
.C(n_228),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_270),
.B(n_272),
.Y(n_286)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_251),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_244),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_241),
.A2(n_242),
.B(n_249),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_274),
.A2(n_248),
.B(n_239),
.Y(n_282)
);

OAI22x1_ASAP7_75t_R g276 ( 
.A1(n_234),
.A2(n_219),
.B1(n_223),
.B2(n_227),
.Y(n_276)
);

NOR2x1_ASAP7_75t_R g285 ( 
.A(n_276),
.B(n_275),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_219),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_235),
.C(n_227),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_218),
.Y(n_278)
);

INVxp33_ASAP7_75t_SL g295 ( 
.A(n_278),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_226),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_279),
.A2(n_250),
.B1(n_217),
.B2(n_210),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_261),
.A2(n_232),
.B1(n_240),
.B2(n_252),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_280),
.A2(n_287),
.B1(n_290),
.B2(n_293),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_288),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_261),
.A2(n_235),
.B1(n_231),
.B2(n_257),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_262),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g293 ( 
.A1(n_276),
.A2(n_204),
.B1(n_231),
.B2(n_254),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_264),
.A2(n_221),
.B(n_211),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_296),
.B(n_293),
.Y(n_298)
);

AOI211xp5_ASAP7_75t_SL g297 ( 
.A1(n_276),
.A2(n_211),
.B(n_225),
.C(n_206),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_297),
.B(n_278),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_310),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_281),
.B(n_262),
.C(n_269),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_306),
.C(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_301),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_277),
.B1(n_274),
.B2(n_266),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_302),
.A2(n_308),
.B1(n_290),
.B2(n_295),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_294),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_281),
.B(n_265),
.C(n_259),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_307),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_270),
.B1(n_260),
.B2(n_268),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_289),
.Y(n_309)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_309),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_271),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_286),
.B(n_272),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_311),
.B(n_312),
.Y(n_318)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_284),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_303),
.A2(n_282),
.B(n_300),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_319),
.Y(n_327)
);

BUFx24_ASAP7_75t_SL g314 ( 
.A(n_304),
.Y(n_314)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_314),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_283),
.CI(n_285),
.CON(n_317),
.SN(n_317)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_302),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_286),
.Y(n_321)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_321),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_306),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_299),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_319),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_330),
.Y(n_335)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_315),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g337 ( 
.A(n_331),
.Y(n_337)
);

OAI22xp33_ASAP7_75t_L g332 ( 
.A1(n_316),
.A2(n_299),
.B1(n_301),
.B2(n_303),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_332),
.B(n_320),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_324),
.A2(n_296),
.B1(n_283),
.B2(n_297),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_333),
.B(n_332),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_334),
.B(n_336),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_323),
.C(n_318),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_338),
.A2(n_339),
.B(n_340),
.Y(n_344)
);

NOR2x1_ASAP7_75t_L g339 ( 
.A(n_325),
.B(n_322),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g341 ( 
.A1(n_335),
.A2(n_320),
.B(n_326),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_341),
.B(n_342),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_337),
.A2(n_317),
.B(n_331),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_339),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_346),
.B(n_344),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_348),
.B(n_337),
.CI(n_317),
.CON(n_349),
.SN(n_349)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_349),
.Y(n_351)
);


endmodule