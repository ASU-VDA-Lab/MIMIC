module fake_jpeg_19184_n_317 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_317);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_317;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_11;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_12;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_8),
.Y(n_15)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_27),
.Y(n_45)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_26),
.B(n_34),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_12),
.B(n_10),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_35),
.B(n_23),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_36),
.B(n_31),
.Y(n_61)
);

OR2x2_ASAP7_75t_SL g46 ( 
.A(n_27),
.B(n_22),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_33),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_49),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_50),
.B(n_46),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_41),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_60),
.Y(n_63)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_52),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_57),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_55),
.Y(n_73)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_58),
.B(n_59),
.Y(n_78)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_36),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_62),
.B(n_69),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_46),
.B1(n_43),
.B2(n_45),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_36),
.B1(n_43),
.B2(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_46),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_65),
.B(n_38),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_51),
.A2(n_41),
.B1(n_34),
.B2(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_40),
.B1(n_55),
.B2(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_53),
.B(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_75),
.B(n_54),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_57),
.A2(n_43),
.B(n_41),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_87),
.B1(n_69),
.B2(n_55),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_58),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_78),
.Y(n_108)
);

XOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_69),
.B(n_43),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_24),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_71),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_82),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_67),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_92),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_63),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_66),
.B(n_59),
.Y(n_86)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_43),
.C(n_39),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_24),
.C(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_91),
.B(n_93),
.Y(n_99)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_66),
.B(n_56),
.Y(n_94)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_48),
.Y(n_95)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_95),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_75),
.B(n_15),
.Y(n_97)
);

NOR2x1_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_84),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_64),
.B1(n_65),
.B2(n_63),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_107),
.B1(n_115),
.B2(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_97),
.Y(n_129)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_92),
.Y(n_103)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_118),
.B1(n_95),
.B2(n_85),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_86),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_92),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_80),
.A2(n_63),
.B1(n_78),
.B2(n_76),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_108),
.A2(n_13),
.B(n_21),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_116),
.C(n_121),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_110),
.B(n_112),
.Y(n_136)
);

OAI32xp33_ASAP7_75t_L g111 ( 
.A1(n_90),
.A2(n_73),
.A3(n_16),
.B1(n_20),
.B2(n_67),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_77),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_90),
.B(n_26),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_80),
.A2(n_38),
.B1(n_34),
.B2(n_39),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_70),
.C(n_73),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_81),
.B(n_26),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_96),
.A2(n_73),
.B1(n_74),
.B2(n_25),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_119),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_70),
.C(n_60),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_122),
.A2(n_85),
.B1(n_93),
.B2(n_94),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_154),
.B1(n_82),
.B2(n_74),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_102),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_126),
.B(n_128),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_127),
.B(n_140),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_129),
.B(n_133),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_130),
.A2(n_74),
.B1(n_37),
.B2(n_29),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_32),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_98),
.B(n_83),
.C(n_95),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_132),
.B(n_138),
.C(n_144),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_108),
.B(n_91),
.Y(n_133)
);

CKINVDCx12_ASAP7_75t_R g134 ( 
.A(n_120),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_150),
.Y(n_160)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_119),
.Y(n_135)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_83),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_12),
.B(n_22),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_91),
.C(n_70),
.Y(n_138)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_148),
.Y(n_180)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_79),
.B1(n_88),
.B2(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_142),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_107),
.B(n_112),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_143),
.B(n_54),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_109),
.B(n_117),
.C(n_114),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_88),
.Y(n_145)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_103),
.Y(n_146)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_17),
.Y(n_168)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_60),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_52),
.C(n_48),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_71),
.C(n_52),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_105),
.B(n_68),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_101),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_151),
.B(n_153),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_152),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_99),
.B(n_77),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_118),
.B(n_100),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_155),
.B(n_16),
.Y(n_182)
);

NOR2x1_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_18),
.Y(n_159)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_159),
.Y(n_188)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_162),
.B(n_165),
.Y(n_193)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_164),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_123),
.B(n_52),
.C(n_71),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_167),
.Y(n_190)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_168),
.Y(n_187)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_141),
.Y(n_170)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_170),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_123),
.B(n_31),
.C(n_32),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_171),
.B(n_149),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_172),
.A2(n_137),
.B1(n_139),
.B2(n_140),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_173),
.A2(n_124),
.B1(n_138),
.B2(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_154),
.A2(n_14),
.B1(n_18),
.B2(n_74),
.Y(n_174)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_174),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_179),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_29),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_184),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_127),
.B(n_128),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_16),
.B1(n_22),
.B2(n_15),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_47),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_136),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_194),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_169),
.B(n_147),
.Y(n_192)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g194 ( 
.A(n_184),
.B(n_132),
.CI(n_137),
.CON(n_194),
.SN(n_194)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_206),
.B1(n_173),
.B2(n_170),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_175),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_197),
.B(n_202),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_198),
.A2(n_161),
.B1(n_180),
.B2(n_179),
.Y(n_212)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_183),
.Y(n_199)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_199),
.Y(n_230)
);

XOR2x2_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_144),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_200),
.A2(n_167),
.B1(n_160),
.B2(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_176),
.A2(n_136),
.B1(n_37),
.B2(n_22),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_201),
.A2(n_209),
.B1(n_13),
.B2(n_19),
.Y(n_232)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_170),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_185),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g215 ( 
.A(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_14),
.B1(n_18),
.B2(n_16),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_77),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_208),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_SL g208 ( 
.A(n_159),
.B(n_10),
.C(n_9),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_156),
.A2(n_37),
.B1(n_16),
.B2(n_14),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_212),
.B(n_229),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_163),
.C(n_166),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_220),
.C(n_221),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_193),
.B(n_163),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_214),
.B(n_217),
.Y(n_248)
);

FAx1_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_178),
.CI(n_162),
.CON(n_219),
.SN(n_219)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_161),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_196),
.B(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_196),
.B(n_190),
.C(n_165),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_229),
.C(n_231),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_223),
.A2(n_225),
.B1(n_232),
.B2(n_208),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_188),
.A2(n_168),
.B1(n_158),
.B2(n_18),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_14),
.B1(n_1),
.B2(n_2),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_226),
.B(n_210),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_187),
.B(n_47),
.Y(n_227)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_21),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_194),
.B(n_31),
.C(n_23),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_194),
.B(n_13),
.C(n_19),
.Y(n_231)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_195),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_235),
.A2(n_245),
.B(n_17),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_233),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_239),
.A2(n_226),
.B1(n_232),
.B2(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_218),
.B(n_209),
.Y(n_240)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_240),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_212),
.A2(n_186),
.B1(n_202),
.B2(n_189),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_241),
.A2(n_220),
.B1(n_213),
.B2(n_2),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_204),
.Y(n_242)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_216),
.Y(n_244)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_244),
.Y(n_259)
);

BUFx12f_ASAP7_75t_SL g245 ( 
.A(n_231),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g246 ( 
.A1(n_215),
.A2(n_186),
.B(n_204),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_246),
.A2(n_249),
.B1(n_252),
.B2(n_219),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_222),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_250),
.A2(n_21),
.B(n_19),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_217),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_261),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_257),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_214),
.B(n_219),
.Y(n_260)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_260),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_234),
.B(n_221),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_264),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_243),
.B(n_248),
.C(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_263),
.B(n_267),
.C(n_10),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_251),
.A2(n_7),
.B(n_10),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_235),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_266),
.B(n_8),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_243),
.B(n_17),
.C(n_1),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_244),
.Y(n_268)
);

AOI21xp33_ASAP7_75t_L g292 ( 
.A1(n_268),
.A2(n_1),
.B(n_2),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_237),
.C(n_246),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_271),
.C(n_267),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_246),
.C(n_247),
.Y(n_271)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_272),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_266),
.A2(n_238),
.B(n_241),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_274),
.A2(n_281),
.B(n_0),
.Y(n_288)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_275),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_257),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_0),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_0),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_8),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_262),
.C(n_260),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_293),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_255),
.B1(n_254),
.B2(n_258),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_285),
.B(n_286),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_264),
.C(n_1),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_288),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_290),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_275),
.B(n_278),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_291),
.B(n_3),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_294),
.B(n_281),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_278),
.B(n_2),
.C(n_3),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_276),
.Y(n_294)
);

NOR2xp67_ASAP7_75t_SL g295 ( 
.A(n_284),
.B(n_273),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_304),
.B(n_4),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_298),
.B(n_299),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_282),
.A2(n_283),
.B(n_294),
.Y(n_299)
);

NOR2x1_ASAP7_75t_L g301 ( 
.A(n_293),
.B(n_280),
.Y(n_301)
);

OR2x2_ASAP7_75t_L g309 ( 
.A(n_301),
.B(n_4),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_4),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g304 ( 
.A1(n_290),
.A2(n_3),
.B(n_4),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_300),
.B(n_6),
.Y(n_306)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_308),
.A3(n_300),
.B1(n_303),
.B2(n_6),
.C1(n_4),
.C2(n_5),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_297),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_305),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_296),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_310),
.B1(n_5),
.B2(n_6),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_5),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_316),
.A2(n_5),
.B(n_306),
.Y(n_317)
);


endmodule