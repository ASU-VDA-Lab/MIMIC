module fake_jpeg_7639_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_37),
.Y(n_54)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_22),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_27),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_41),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_22),
.B(n_15),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_43),
.Y(n_63)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_53),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g46 ( 
.A(n_36),
.Y(n_46)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_49),
.Y(n_86)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_38),
.B(n_31),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_25),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_50),
.A2(n_21),
.B(n_28),
.Y(n_90)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_51),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_39),
.Y(n_52)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_37),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_18),
.B1(n_35),
.B2(n_33),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_60),
.B1(n_21),
.B2(n_28),
.Y(n_89)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_24),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_20),
.B1(n_33),
.B2(n_32),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_62),
.Y(n_88)
);

INVx1_ASAP7_75t_SL g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_64),
.B(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_31),
.Y(n_65)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_50),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_44),
.B1(n_59),
.B2(n_51),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_69),
.A2(n_78),
.B1(n_45),
.B2(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_71),
.B(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_63),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_46),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_59),
.A2(n_25),
.B1(n_32),
.B2(n_20),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_42),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_79),
.B(n_90),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_47),
.A2(n_26),
.B1(n_19),
.B2(n_30),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_81),
.A2(n_23),
.B1(n_26),
.B2(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_29),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_67),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_84),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_18),
.B1(n_32),
.B2(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_87),
.A2(n_89),
.B1(n_91),
.B2(n_19),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_21),
.B1(n_30),
.B2(n_17),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_SL g125 ( 
.A(n_94),
.B(n_103),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g95 ( 
.A(n_84),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_99),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_96),
.B(n_100),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_98),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_82),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_83),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_73),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_106),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_50),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_76),
.B(n_54),
.C(n_58),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_113),
.C(n_117),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_54),
.Y(n_106)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_108),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_86),
.B(n_58),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_109),
.B(n_90),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_72),
.B(n_75),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_66),
.B(n_57),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

AND2x6_ASAP7_75t_L g117 ( 
.A(n_86),
.B(n_0),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_97),
.A2(n_80),
.B1(n_45),
.B2(n_88),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_121),
.A2(n_132),
.B1(n_140),
.B2(n_95),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g122 ( 
.A(n_97),
.B(n_66),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_SL g157 ( 
.A(n_122),
.B(n_96),
.C(n_61),
.Y(n_157)
);

AO21x2_ASAP7_75t_L g123 ( 
.A1(n_113),
.A2(n_74),
.B(n_75),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_123),
.A2(n_128),
.B1(n_142),
.B2(n_107),
.Y(n_145)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_113),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_130),
.B(n_136),
.Y(n_151)
);

OAI22xp33_ASAP7_75t_L g128 ( 
.A1(n_101),
.A2(n_85),
.B1(n_82),
.B2(n_77),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_103),
.A2(n_46),
.B1(n_81),
.B2(n_70),
.Y(n_132)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_137),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_109),
.B(n_23),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_138),
.Y(n_170)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_94),
.A2(n_61),
.B1(n_29),
.B2(n_34),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_61),
.B1(n_29),
.B2(n_34),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_143),
.Y(n_163)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_108),
.Y(n_144)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_145),
.A2(n_153),
.B1(n_169),
.B2(n_130),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_126),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_147),
.B(n_149),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_125),
.B(n_102),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_167),
.C(n_119),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_131),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_144),
.A2(n_117),
.B1(n_111),
.B2(n_109),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_128),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_118),
.A2(n_107),
.B1(n_116),
.B2(n_110),
.Y(n_155)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_155),
.Y(n_174)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_159),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_157),
.A2(n_158),
.B(n_165),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_118),
.A2(n_96),
.B1(n_92),
.B2(n_99),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_122),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_123),
.A2(n_99),
.B1(n_115),
.B2(n_92),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g193 ( 
.A1(n_160),
.A2(n_124),
.B(n_141),
.Y(n_193)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_123),
.B(n_1),
.C(n_3),
.D(n_4),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_161),
.B(n_142),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_120),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_168),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_133),
.A2(n_29),
.B1(n_34),
.B2(n_114),
.Y(n_164)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_164),
.Y(n_179)
);

AOI32xp33_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_95),
.A3(n_27),
.B1(n_114),
.B2(n_5),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_123),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_124),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_27),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_120),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_139),
.A2(n_114),
.B1(n_95),
.B2(n_27),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_140),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_167),
.B(n_119),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_176),
.B(n_183),
.C(n_194),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_136),
.B(n_127),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_177),
.A2(n_191),
.B(n_193),
.Y(n_206)
);

FAx1_ASAP7_75t_SL g213 ( 
.A(n_178),
.B(n_4),
.CI(n_6),
.CON(n_213),
.SN(n_213)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_147),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_143),
.C(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_184),
.B(n_188),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_132),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_7),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_186),
.A2(n_192),
.B1(n_159),
.B2(n_156),
.Y(n_197)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_158),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_146),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_189),
.B(n_195),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_171),
.B1(n_149),
.B2(n_172),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_157),
.B1(n_134),
.B2(n_163),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_151),
.B(n_138),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_145),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_196),
.B(n_8),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_197),
.B(n_192),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_212),
.B1(n_217),
.B2(n_179),
.Y(n_230)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_173),
.Y(n_199)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_199),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_152),
.C(n_129),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_204),
.C(n_210),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_202),
.B(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_129),
.Y(n_203)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_191),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_175),
.Y(n_207)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

INVx13_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_137),
.C(n_170),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_1),
.C(n_3),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_211),
.B(n_215),
.C(n_178),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_195),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_214),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_181),
.B(n_6),
.Y(n_214)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_221),
.B(n_213),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_198),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_175),
.C(n_194),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_223),
.B(n_213),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_181),
.C(n_193),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_224),
.B(n_226),
.C(n_233),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_190),
.C(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_230),
.Y(n_245)
);

AOI21xp33_ASAP7_75t_L g231 ( 
.A1(n_206),
.A2(n_188),
.B(n_174),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_231),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_200),
.B(n_8),
.C(n_9),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_9),
.Y(n_234)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_234),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_234),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_238),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_208),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_240),
.A2(n_242),
.B(n_225),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_222),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_200),
.C(n_210),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_219),
.C(n_226),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_228),
.A2(n_206),
.B1(n_212),
.B2(n_211),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_246),
.B(n_233),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_248),
.C(n_256),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_239),
.A2(n_238),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_253),
.B(n_237),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_245),
.A2(n_224),
.B1(n_229),
.B2(n_221),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_236),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_225),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_252),
.B(n_255),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_235),
.A2(n_220),
.B(n_229),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_215),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_247),
.B(n_244),
.C(n_236),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_260),
.C(n_254),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_259),
.B(n_10),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_251),
.B(n_248),
.C(n_256),
.Y(n_260)
);

NOR2xp67_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_241),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_10),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_263),
.B(n_10),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_265),
.B(n_269),
.Y(n_272)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_261),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_268),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_11),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_270),
.A2(n_262),
.B(n_12),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_271),
.B(n_11),
.C(n_13),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_275),
.B(n_276),
.C(n_274),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_257),
.C(n_267),
.Y(n_276)
);

AOI33xp33_ASAP7_75t_L g278 ( 
.A1(n_277),
.A2(n_13),
.A3(n_14),
.B1(n_15),
.B2(n_273),
.B3(n_262),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_13),
.Y(n_279)
);


endmodule