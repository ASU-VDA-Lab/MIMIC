module real_aes_7496_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_182;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_217;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_420;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g107 ( .A(n_0), .Y(n_107) );
A2O1A1Ixp33_ASAP7_75t_L g455 ( .A1(n_1), .A2(n_144), .B(n_156), .C(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g263 ( .A(n_2), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_3), .A2(n_171), .B(n_495), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_4), .B(n_167), .Y(n_500) );
AOI21xp33_ASAP7_75t_L g170 ( .A1(n_5), .A2(n_171), .B(n_172), .Y(n_170) );
AND2x6_ASAP7_75t_L g144 ( .A(n_6), .B(n_145), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_7), .A2(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g105 ( .A(n_8), .Y(n_105) );
NOR2xp33_ASAP7_75t_L g124 ( .A(n_8), .B(n_39), .Y(n_124) );
INVx1_ASAP7_75t_L g471 ( .A(n_9), .Y(n_471) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_10), .B(n_177), .Y(n_459) );
INVx1_ASAP7_75t_L g179 ( .A(n_11), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_12), .B(n_231), .Y(n_230) );
INVx1_ASAP7_75t_L g141 ( .A(n_13), .Y(n_141) );
INVx1_ASAP7_75t_L g245 ( .A(n_14), .Y(n_245) );
A2O1A1Ixp33_ASAP7_75t_L g479 ( .A1(n_15), .A2(n_180), .B(n_246), .C(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_16), .B(n_167), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_17), .B(n_190), .Y(n_217) );
NAND2xp5_ASAP7_75t_SL g199 ( .A(n_18), .B(n_171), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_19), .B(n_513), .Y(n_512) );
A2O1A1Ixp33_ASAP7_75t_L g487 ( .A1(n_20), .A2(n_147), .B(n_231), .C(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_21), .B(n_167), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_22), .B(n_177), .Y(n_534) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_23), .A2(n_243), .B(n_244), .C(n_246), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_24), .B(n_177), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g530 ( .A(n_25), .Y(n_530) );
INVx1_ASAP7_75t_L g520 ( .A(n_26), .Y(n_520) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_27), .Y(n_152) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_28), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_29), .B(n_177), .Y(n_264) );
INVx1_ASAP7_75t_L g509 ( .A(n_30), .Y(n_509) );
INVx1_ASAP7_75t_L g155 ( .A(n_31), .Y(n_155) );
INVx2_ASAP7_75t_L g149 ( .A(n_32), .Y(n_149) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_33), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g497 ( .A1(n_34), .A2(n_181), .B(n_231), .C(n_498), .Y(n_497) );
INVxp67_ASAP7_75t_L g510 ( .A(n_35), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g200 ( .A1(n_36), .A2(n_144), .B(n_156), .C(n_201), .Y(n_200) );
CKINVDCx14_ASAP7_75t_R g496 ( .A(n_37), .Y(n_496) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_38), .A2(n_156), .B(n_519), .C(n_523), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_39), .B(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g153 ( .A(n_40), .Y(n_153) );
A2O1A1Ixp33_ASAP7_75t_L g469 ( .A1(n_41), .A2(n_176), .B(n_206), .C(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_42), .B(n_177), .Y(n_216) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_43), .Y(n_525) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_44), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_45), .Y(n_125) );
INVx1_ASAP7_75t_L g486 ( .A(n_46), .Y(n_486) );
CKINVDCx16_ASAP7_75t_R g159 ( .A(n_47), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_48), .B(n_171), .Y(n_233) );
AOI222xp33_ASAP7_75t_SL g126 ( .A1(n_49), .A2(n_58), .B1(n_127), .B2(n_713), .C1(n_714), .C2(n_718), .Y(n_126) );
AOI22xp5_ASAP7_75t_L g146 ( .A1(n_50), .A2(n_147), .B1(n_150), .B2(n_156), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_51), .Y(n_210) );
CKINVDCx16_ASAP7_75t_R g260 ( .A(n_52), .Y(n_260) );
A2O1A1Ixp33_ASAP7_75t_L g175 ( .A1(n_53), .A2(n_176), .B(n_178), .C(n_181), .Y(n_175) );
CKINVDCx14_ASAP7_75t_R g468 ( .A(n_54), .Y(n_468) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_55), .Y(n_220) );
INVx1_ASAP7_75t_L g173 ( .A(n_56), .Y(n_173) );
INVx1_ASAP7_75t_L g145 ( .A(n_57), .Y(n_145) );
CKINVDCx20_ASAP7_75t_R g713 ( .A(n_58), .Y(n_713) );
INVx1_ASAP7_75t_L g140 ( .A(n_59), .Y(n_140) );
INVx1_ASAP7_75t_SL g499 ( .A(n_60), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_61), .Y(n_117) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_62), .B(n_167), .Y(n_490) );
OAI22xp5_ASAP7_75t_SL g723 ( .A1(n_63), .A2(n_445), .B1(n_715), .B2(n_724), .Y(n_723) );
CKINVDCx20_ASAP7_75t_R g724 ( .A(n_63), .Y(n_724) );
INVx1_ASAP7_75t_L g533 ( .A(n_64), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_SL g189 ( .A1(n_65), .A2(n_181), .B(n_190), .C(n_191), .Y(n_189) );
INVxp67_ASAP7_75t_L g192 ( .A(n_66), .Y(n_192) );
INVx1_ASAP7_75t_L g110 ( .A(n_67), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_68), .A2(n_171), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g537 ( .A(n_69), .Y(n_537) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_70), .Y(n_164) );
AOI21xp5_ASAP7_75t_L g476 ( .A1(n_71), .A2(n_171), .B(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g213 ( .A(n_72), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_73), .A2(n_239), .B(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g478 ( .A(n_74), .Y(n_478) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_75), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g214 ( .A1(n_76), .A2(n_144), .B(n_156), .C(n_215), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_77), .A2(n_171), .B(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g481 ( .A(n_78), .Y(n_481) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_79), .B(n_203), .Y(n_202) );
INVx2_ASAP7_75t_L g138 ( .A(n_80), .Y(n_138) );
INVx1_ASAP7_75t_L g457 ( .A(n_81), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_82), .B(n_190), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_83), .A2(n_144), .B(n_156), .C(n_262), .Y(n_261) );
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_84), .B(n_107), .C(n_108), .Y(n_106) );
OR2x2_ASAP7_75t_L g121 ( .A(n_84), .B(n_122), .Y(n_121) );
INVx2_ASAP7_75t_L g444 ( .A(n_84), .Y(n_444) );
OR2x2_ASAP7_75t_L g712 ( .A(n_84), .B(n_123), .Y(n_712) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_85), .A2(n_156), .B(n_532), .C(n_535), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_86), .B(n_184), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g267 ( .A(n_87), .Y(n_267) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_88), .A2(n_144), .B(n_156), .C(n_228), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_89), .Y(n_235) );
INVx1_ASAP7_75t_L g188 ( .A(n_90), .Y(n_188) );
CKINVDCx16_ASAP7_75t_R g241 ( .A(n_91), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_92), .B(n_203), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_93), .B(n_169), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_94), .B(n_169), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_95), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_96), .A2(n_171), .B(n_187), .Y(n_186) );
INVx2_ASAP7_75t_L g489 ( .A(n_97), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g99 ( .A1(n_98), .A2(n_100), .B1(n_111), .B2(n_727), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g100 ( .A(n_101), .Y(n_100) );
INVx5_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
CKINVDCx9p33_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
BUFx4f_ASAP7_75t_SL g727 ( .A(n_103), .Y(n_727) );
OR2x4_ASAP7_75t_L g103 ( .A(n_104), .B(n_106), .Y(n_103) );
AND2x2_ASAP7_75t_L g123 ( .A(n_107), .B(n_124), .Y(n_123) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_126), .B1(n_721), .B2(n_722), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_118), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_SL g721 ( .A(n_115), .Y(n_721) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g722 ( .A1(n_118), .A2(n_723), .B(n_725), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g118 ( .A(n_119), .B(n_125), .Y(n_118) );
INVx1_ASAP7_75t_SL g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_SL g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g726 ( .A(n_121), .Y(n_726) );
NOR2x2_ASAP7_75t_L g720 ( .A(n_122), .B(n_444), .Y(n_720) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g443 ( .A(n_123), .B(n_444), .Y(n_443) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_441), .B1(n_445), .B2(n_712), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
OAI22xp5_ASAP7_75t_SL g714 ( .A1(n_129), .A2(n_441), .B1(n_715), .B2(n_716), .Y(n_714) );
AND3x1_ASAP7_75t_L g129 ( .A(n_130), .B(n_366), .C(n_415), .Y(n_129) );
NOR3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_273), .C(n_311), .Y(n_130) );
OAI222xp33_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_194), .B1(n_248), .B2(n_254), .C1(n_268), .C2(n_271), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_133), .B(n_165), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g340 ( .A(n_133), .B(n_341), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_133), .B(n_316), .Y(n_407) );
BUFx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OR2x2_ASAP7_75t_L g284 ( .A(n_134), .B(n_185), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_134), .B(n_166), .Y(n_292) );
AND2x2_ASAP7_75t_L g327 ( .A(n_134), .B(n_304), .Y(n_327) );
OR2x2_ASAP7_75t_L g351 ( .A(n_134), .B(n_166), .Y(n_351) );
OR2x2_ASAP7_75t_L g359 ( .A(n_134), .B(n_258), .Y(n_359) );
AND2x2_ASAP7_75t_L g362 ( .A(n_134), .B(n_185), .Y(n_362) );
INVx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
OR2x2_ASAP7_75t_L g256 ( .A(n_135), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g270 ( .A(n_135), .B(n_185), .Y(n_270) );
AND2x2_ASAP7_75t_L g320 ( .A(n_135), .B(n_258), .Y(n_320) );
AND2x2_ASAP7_75t_L g333 ( .A(n_135), .B(n_166), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_135), .B(n_419), .Y(n_440) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_142), .B(n_163), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g163 ( .A(n_136), .B(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g208 ( .A(n_136), .Y(n_208) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_136), .A2(n_259), .B(n_266), .Y(n_258) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_137), .Y(n_169) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_138), .B(n_139), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
OAI22xp33_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_146), .B1(n_159), .B2(n_160), .Y(n_142) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_143), .A2(n_173), .B(n_174), .C(n_175), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g187 ( .A1(n_143), .A2(n_174), .B(n_188), .C(n_189), .Y(n_187) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_143), .A2(n_174), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g467 ( .A1(n_143), .A2(n_174), .B(n_468), .C(n_469), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_SL g477 ( .A1(n_143), .A2(n_174), .B(n_478), .C(n_479), .Y(n_477) );
O2A1O1Ixp33_ASAP7_75t_SL g485 ( .A1(n_143), .A2(n_174), .B(n_486), .C(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g495 ( .A1(n_143), .A2(n_174), .B(n_496), .C(n_497), .Y(n_495) );
O2A1O1Ixp33_ASAP7_75t_SL g505 ( .A1(n_143), .A2(n_174), .B(n_506), .C(n_507), .Y(n_505) );
INVx1_ASAP7_75t_L g535 ( .A(n_143), .Y(n_535) );
INVx4_ASAP7_75t_SL g143 ( .A(n_144), .Y(n_143) );
NAND2x1p5_ASAP7_75t_L g160 ( .A(n_144), .B(n_161), .Y(n_160) );
AND2x4_ASAP7_75t_L g171 ( .A(n_144), .B(n_161), .Y(n_171) );
BUFx3_ASAP7_75t_L g523 ( .A(n_144), .Y(n_523) );
INVx2_ASAP7_75t_L g265 ( .A(n_147), .Y(n_265) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g157 ( .A(n_149), .Y(n_157) );
INVx1_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
OAI22xp5_ASAP7_75t_SL g150 ( .A1(n_151), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_150) );
INVx2_ASAP7_75t_L g154 ( .A(n_151), .Y(n_154) );
INVx4_ASAP7_75t_L g243 ( .A(n_151), .Y(n_243) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g158 ( .A(n_152), .Y(n_158) );
AND2x2_ASAP7_75t_L g161 ( .A(n_152), .B(n_162), .Y(n_161) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_152), .Y(n_177) );
INVx3_ASAP7_75t_L g180 ( .A(n_152), .Y(n_180) );
INVx1_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx2_ASAP7_75t_L g458 ( .A(n_154), .Y(n_458) );
INVx5_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_158), .Y(n_156) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_157), .Y(n_182) );
BUFx3_ASAP7_75t_L g207 ( .A(n_157), .Y(n_207) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_160), .A2(n_213), .B(n_214), .Y(n_212) );
OAI21xp5_ASAP7_75t_L g259 ( .A1(n_160), .A2(n_260), .B(n_261), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_160), .A2(n_454), .B(n_455), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_160), .A2(n_184), .B(n_517), .C(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_160), .A2(n_530), .B(n_531), .Y(n_529) );
INVx1_ASAP7_75t_L g511 ( .A(n_162), .Y(n_511) );
O2A1O1Ixp33_ASAP7_75t_L g358 ( .A1(n_165), .A2(n_359), .B(n_360), .C(n_363), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_165), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_165), .B(n_303), .Y(n_425) );
AND2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_185), .Y(n_165) );
AND2x2_ASAP7_75t_SL g269 ( .A(n_166), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g283 ( .A(n_166), .Y(n_283) );
AND2x2_ASAP7_75t_L g310 ( .A(n_166), .B(n_304), .Y(n_310) );
INVx1_ASAP7_75t_SL g318 ( .A(n_166), .Y(n_318) );
AND2x2_ASAP7_75t_L g341 ( .A(n_166), .B(n_342), .Y(n_341) );
BUFx2_ASAP7_75t_L g419 ( .A(n_166), .Y(n_419) );
OA21x2_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_183), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g209 ( .A(n_168), .B(n_210), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_168), .B(n_461), .Y(n_460) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_168), .B(n_525), .Y(n_524) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_168), .A2(n_529), .B(n_536), .Y(n_528) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_169), .A2(n_186), .B(n_193), .Y(n_185) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_169), .Y(n_475) );
BUFx2_ASAP7_75t_L g239 ( .A(n_171), .Y(n_239) );
INVx2_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx4_ASAP7_75t_L g231 ( .A(n_177), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_179), .B(n_180), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_180), .B(n_192), .Y(n_191) );
INVx5_ASAP7_75t_L g203 ( .A(n_180), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_180), .B(n_471), .Y(n_470) );
INVx3_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
HB1xp67_ASAP7_75t_L g232 ( .A(n_182), .Y(n_232) );
INVx1_ASAP7_75t_L g221 ( .A(n_184), .Y(n_221) );
INVx2_ASAP7_75t_L g225 ( .A(n_184), .Y(n_225) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_184), .A2(n_238), .B(n_247), .Y(n_237) );
OA21x2_ASAP7_75t_L g465 ( .A1(n_184), .A2(n_466), .B(n_472), .Y(n_465) );
BUFx2_ASAP7_75t_L g255 ( .A(n_185), .Y(n_255) );
INVx1_ASAP7_75t_L g317 ( .A(n_185), .Y(n_317) );
INVx3_ASAP7_75t_L g342 ( .A(n_185), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_194), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_222), .Y(n_194) );
INVx1_ASAP7_75t_L g338 ( .A(n_195), .Y(n_338) );
OAI32xp33_ASAP7_75t_L g344 ( .A1(n_195), .A2(n_283), .A3(n_345), .B1(n_346), .B2(n_347), .Y(n_344) );
OAI22xp5_ASAP7_75t_L g348 ( .A1(n_195), .A2(n_349), .B1(n_352), .B2(n_357), .Y(n_348) );
INVx4_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
AND2x2_ASAP7_75t_L g286 ( .A(n_196), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g364 ( .A(n_196), .B(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g434 ( .A(n_196), .B(n_380), .Y(n_434) );
AND2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_211), .Y(n_196) );
AND2x2_ASAP7_75t_L g249 ( .A(n_197), .B(n_250), .Y(n_249) );
INVx2_ASAP7_75t_L g279 ( .A(n_197), .Y(n_279) );
INVx1_ASAP7_75t_L g298 ( .A(n_197), .Y(n_298) );
OR2x2_ASAP7_75t_L g306 ( .A(n_197), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g313 ( .A(n_197), .B(n_287), .Y(n_313) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_197), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g334 ( .A(n_197), .B(n_252), .Y(n_334) );
INVx3_ASAP7_75t_L g356 ( .A(n_197), .Y(n_356) );
AND2x2_ASAP7_75t_L g381 ( .A(n_197), .B(n_253), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g429 ( .A(n_197), .B(n_346), .Y(n_429) );
OR2x6_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
AOI21xp5_ASAP7_75t_SL g198 ( .A1(n_199), .A2(n_200), .B(n_208), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_202), .A2(n_204), .B(n_205), .Y(n_201) );
O2A1O1Ixp33_ASAP7_75t_L g262 ( .A1(n_203), .A2(n_263), .B(n_264), .C(n_265), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g508 ( .A1(n_203), .A2(n_243), .B1(n_509), .B2(n_510), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_203), .A2(n_520), .B(n_521), .C(n_522), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_205), .A2(n_216), .B(n_217), .Y(n_215) );
O2A1O1Ixp5_ASAP7_75t_L g456 ( .A1(n_205), .A2(n_457), .B(n_458), .C(n_459), .Y(n_456) );
O2A1O1Ixp33_ASAP7_75t_L g532 ( .A1(n_205), .A2(n_458), .B(n_533), .C(n_534), .Y(n_532) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx1_ASAP7_75t_L g246 ( .A(n_207), .Y(n_246) );
INVx1_ASAP7_75t_L g218 ( .A(n_208), .Y(n_218) );
INVx2_ASAP7_75t_L g253 ( .A(n_211), .Y(n_253) );
AND2x2_ASAP7_75t_L g385 ( .A(n_211), .B(n_223), .Y(n_385) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_211) );
INVx1_ASAP7_75t_L g503 ( .A(n_218), .Y(n_503) );
AO21x2_ASAP7_75t_L g555 ( .A1(n_218), .A2(n_556), .B(n_557), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g219 ( .A(n_220), .B(n_221), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_221), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g266 ( .A(n_221), .B(n_267), .Y(n_266) );
AO21x2_ASAP7_75t_L g452 ( .A1(n_221), .A2(n_453), .B(n_460), .Y(n_452) );
INVx2_ASAP7_75t_L g427 ( .A(n_222), .Y(n_427) );
OR2x2_ASAP7_75t_L g222 ( .A(n_223), .B(n_236), .Y(n_222) );
INVx1_ASAP7_75t_L g272 ( .A(n_223), .Y(n_272) );
AND2x2_ASAP7_75t_L g299 ( .A(n_223), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_223), .B(n_253), .Y(n_307) );
AND2x2_ASAP7_75t_L g365 ( .A(n_223), .B(n_288), .Y(n_365) );
INVx2_ASAP7_75t_L g223 ( .A(n_224), .Y(n_223) );
INVx1_ASAP7_75t_L g251 ( .A(n_224), .Y(n_251) );
AND2x2_ASAP7_75t_L g278 ( .A(n_224), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g287 ( .A(n_224), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_224), .B(n_253), .Y(n_353) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_234), .Y(n_224) );
INVx1_ASAP7_75t_L g513 ( .A(n_225), .Y(n_513) );
NOR2xp33_ASAP7_75t_L g536 ( .A(n_225), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_233), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g228 ( .A1(n_229), .A2(n_230), .B(n_232), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_231), .B(n_499), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_236), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_236), .B(n_253), .Y(n_346) );
AND2x2_ASAP7_75t_L g355 ( .A(n_236), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g380 ( .A(n_236), .Y(n_380) );
INVx2_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g252 ( .A(n_237), .B(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g288 ( .A(n_237), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_243), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_243), .B(n_481), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_243), .B(n_489), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_248), .A2(n_258), .B1(n_417), .B2(n_420), .Y(n_416) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
OAI21xp5_ASAP7_75t_SL g439 ( .A1(n_250), .A2(n_361), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g373 ( .A(n_251), .B(n_356), .Y(n_373) );
INVx1_ASAP7_75t_L g398 ( .A(n_251), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_252), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g325 ( .A(n_252), .B(n_278), .Y(n_325) );
INVx2_ASAP7_75t_L g281 ( .A(n_253), .Y(n_281) );
INVx1_ASAP7_75t_L g331 ( .A(n_253), .Y(n_331) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_254), .A2(n_406), .B1(n_423), .B2(n_426), .C(n_428), .Y(n_422) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
INVx1_ASAP7_75t_L g293 ( .A(n_255), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_255), .B(n_304), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g314 ( .A(n_256), .B(n_315), .Y(n_314) );
OR2x2_ASAP7_75t_L g347 ( .A(n_256), .B(n_293), .Y(n_347) );
INVx3_ASAP7_75t_SL g388 ( .A(n_256), .Y(n_388) );
AND2x2_ASAP7_75t_L g332 ( .A(n_257), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g361 ( .A(n_257), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_257), .B(n_270), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_257), .B(n_316), .Y(n_402) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g304 ( .A(n_258), .Y(n_304) );
OAI322xp33_ASAP7_75t_L g399 ( .A1(n_258), .A2(n_330), .A3(n_352), .B1(n_400), .B2(n_402), .C1(n_403), .C2(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
AOI21xp33_ASAP7_75t_L g423 ( .A1(n_269), .A2(n_272), .B(n_424), .Y(n_423) );
NOR2xp33_ASAP7_75t_SL g349 ( .A(n_270), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g371 ( .A(n_270), .B(n_283), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_270), .B(n_310), .Y(n_386) );
INVxp67_ASAP7_75t_L g337 ( .A(n_272), .Y(n_337) );
AOI211xp5_ASAP7_75t_L g343 ( .A1(n_272), .A2(n_344), .B(n_348), .C(n_358), .Y(n_343) );
OAI221xp5_ASAP7_75t_SL g273 ( .A1(n_274), .A2(n_282), .B1(n_285), .B2(n_289), .C(n_294), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AND2x2_ASAP7_75t_L g297 ( .A(n_281), .B(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g414 ( .A(n_281), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_282), .A2(n_431), .B1(n_436), .B2(n_437), .C(n_439), .Y(n_430) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_283), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_SL g330 ( .A(n_283), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_283), .B(n_361), .Y(n_368) );
AND2x2_ASAP7_75t_L g410 ( .A(n_283), .B(n_388), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g308 ( .A(n_284), .B(n_309), .Y(n_308) );
OAI22xp33_ASAP7_75t_L g405 ( .A1(n_284), .A2(n_296), .B1(n_406), .B2(n_407), .Y(n_405) );
OR2x2_ASAP7_75t_L g436 ( .A(n_284), .B(n_304), .Y(n_436) );
CKINVDCx16_ASAP7_75t_R g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g413 ( .A(n_287), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_287), .B(n_381), .Y(n_438) );
INVxp67_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
NOR2xp33_ASAP7_75t_SL g290 ( .A(n_291), .B(n_293), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
OR2x2_ASAP7_75t_L g302 ( .A(n_292), .B(n_303), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g294 ( .A1(n_295), .A2(n_301), .B1(n_305), .B2(n_308), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_L g369 ( .A(n_297), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_297), .B(n_337), .Y(n_404) );
AOI322xp5_ASAP7_75t_L g328 ( .A1(n_299), .A2(n_329), .A3(n_331), .B1(n_332), .B2(n_334), .C1(n_335), .C2(n_339), .Y(n_328) );
INVxp67_ASAP7_75t_L g322 ( .A(n_300), .Y(n_322) );
INVx1_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_302), .A2(n_307), .B1(n_324), .B2(n_326), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_303), .B(n_316), .Y(n_403) );
INVx1_ASAP7_75t_SL g303 ( .A(n_304), .Y(n_303) );
NOR2xp33_ASAP7_75t_L g412 ( .A(n_304), .B(n_342), .Y(n_412) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_304), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OR2x2_ASAP7_75t_L g400 ( .A(n_306), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
NAND3xp33_ASAP7_75t_SL g311 ( .A(n_312), .B(n_328), .C(n_343), .Y(n_311) );
AOI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_314), .B1(n_319), .B2(n_321), .C(n_323), .Y(n_312) );
AND2x2_ASAP7_75t_L g319 ( .A(n_315), .B(n_320), .Y(n_319) );
INVx3_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g329 ( .A(n_320), .B(n_330), .Y(n_329) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_322), .Y(n_401) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_327), .B(n_341), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_330), .B(n_388), .Y(n_394) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_331), .B(n_391), .Y(n_390) );
INVx1_ASAP7_75t_SL g406 ( .A(n_334), .Y(n_406) );
AND2x2_ASAP7_75t_L g421 ( .A(n_334), .B(n_398), .Y(n_421) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AOI211xp5_ASAP7_75t_L g415 ( .A1(n_345), .A2(n_416), .B(n_422), .C(n_430), .Y(n_415) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
OR2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_354), .Y(n_352) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
AND2x2_ASAP7_75t_L g384 ( .A(n_355), .B(n_385), .Y(n_384) );
NAND2x1_ASAP7_75t_SL g426 ( .A(n_356), .B(n_427), .Y(n_426) );
CKINVDCx16_ASAP7_75t_R g396 ( .A(n_359), .Y(n_396) );
INVx1_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g391 ( .A(n_365), .Y(n_391) );
AND2x2_ASAP7_75t_L g395 ( .A(n_365), .B(n_381), .Y(n_395) );
NOR5xp2_ASAP7_75t_L g366 ( .A(n_367), .B(n_382), .C(n_399), .D(n_405), .E(n_408), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B1(n_370), .B2(n_372), .C(n_374), .Y(n_367) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_371), .B(n_429), .Y(n_428) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_377), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_381), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
AND2x2_ASAP7_75t_L g397 ( .A(n_381), .B(n_398), .Y(n_397) );
OAI221xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_386), .B1(n_387), .B2(n_389), .C(n_392), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_395), .B1(n_396), .B2(n_397), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx1_ASAP7_75t_L g435 ( .A(n_395), .Y(n_435) );
AOI211xp5_ASAP7_75t_SL g408 ( .A1(n_409), .A2(n_411), .B(n_413), .C(n_414), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_433), .B(n_435), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
CKINVDCx14_ASAP7_75t_R g437 ( .A(n_438), .Y(n_437) );
INVx2_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g715 ( .A(n_445), .Y(n_715) );
OR2x2_ASAP7_75t_SL g445 ( .A(n_446), .B(n_667), .Y(n_445) );
NAND5xp2_ASAP7_75t_L g446 ( .A(n_447), .B(n_579), .C(n_617), .D(n_638), .E(n_655), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_448), .B(n_551), .C(n_572), .Y(n_447) );
OAI221xp5_ASAP7_75t_SL g448 ( .A1(n_449), .A2(n_491), .B1(n_514), .B2(n_538), .C(n_542), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_462), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_451), .B(n_540), .Y(n_559) );
OR2x2_ASAP7_75t_L g586 ( .A(n_451), .B(n_474), .Y(n_586) );
AND2x2_ASAP7_75t_L g600 ( .A(n_451), .B(n_474), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_451), .B(n_465), .Y(n_614) );
AND2x2_ASAP7_75t_L g652 ( .A(n_451), .B(n_616), .Y(n_652) );
AND2x2_ASAP7_75t_L g681 ( .A(n_451), .B(n_591), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_451), .B(n_563), .Y(n_698) );
INVx4_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g578 ( .A(n_452), .B(n_473), .Y(n_578) );
BUFx3_ASAP7_75t_L g603 ( .A(n_452), .Y(n_603) );
AND2x2_ASAP7_75t_L g632 ( .A(n_452), .B(n_474), .Y(n_632) );
AND3x2_ASAP7_75t_L g645 ( .A(n_452), .B(n_646), .C(n_647), .Y(n_645) );
INVx1_ASAP7_75t_L g568 ( .A(n_462), .Y(n_568) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
AOI32xp33_ASAP7_75t_L g623 ( .A1(n_463), .A2(n_575), .A3(n_624), .B1(n_627), .B2(n_628), .Y(n_623) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g550 ( .A(n_464), .B(n_473), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_464), .B(n_578), .Y(n_621) );
AND2x2_ASAP7_75t_L g628 ( .A(n_464), .B(n_600), .Y(n_628) );
OR2x2_ASAP7_75t_L g634 ( .A(n_464), .B(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g659 ( .A(n_464), .B(n_589), .Y(n_659) );
OR2x2_ASAP7_75t_L g677 ( .A(n_464), .B(n_502), .Y(n_677) );
BUFx3_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
AND2x2_ASAP7_75t_L g541 ( .A(n_465), .B(n_483), .Y(n_541) );
INVx2_ASAP7_75t_L g563 ( .A(n_465), .Y(n_563) );
OR2x2_ASAP7_75t_L g585 ( .A(n_465), .B(n_483), .Y(n_585) );
AND2x2_ASAP7_75t_L g590 ( .A(n_465), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_465), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g646 ( .A(n_465), .B(n_540), .Y(n_646) );
INVx1_ASAP7_75t_SL g697 ( .A(n_473), .Y(n_697) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_483), .Y(n_473) );
INVx1_ASAP7_75t_SL g540 ( .A(n_474), .Y(n_540) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_474), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_474), .B(n_626), .Y(n_625) );
NAND3xp33_ASAP7_75t_L g692 ( .A(n_474), .B(n_563), .C(n_681), .Y(n_692) );
OA21x2_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B(n_482), .Y(n_474) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_475), .A2(n_484), .B(n_490), .Y(n_483) );
OA21x2_ASAP7_75t_L g493 ( .A1(n_475), .A2(n_494), .B(n_500), .Y(n_493) );
INVx2_ASAP7_75t_L g591 ( .A(n_483), .Y(n_591) );
HB1xp67_ASAP7_75t_L g605 ( .A(n_483), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
INVx1_ASAP7_75t_L g627 ( .A(n_492), .Y(n_627) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g545 ( .A(n_493), .B(n_527), .Y(n_545) );
INVx2_ASAP7_75t_L g562 ( .A(n_493), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_493), .B(n_528), .Y(n_567) );
AND2x2_ASAP7_75t_L g582 ( .A(n_493), .B(n_515), .Y(n_582) );
AND2x2_ASAP7_75t_L g594 ( .A(n_493), .B(n_566), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_501), .B(n_610), .Y(n_609) );
NAND2x1p5_ASAP7_75t_L g666 ( .A(n_501), .B(n_567), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_501), .B(n_686), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_501), .B(n_561), .Y(n_689) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g526 ( .A(n_502), .B(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_502), .B(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g571 ( .A(n_502), .B(n_515), .Y(n_571) );
AND2x2_ASAP7_75t_L g597 ( .A(n_502), .B(n_527), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_502), .B(n_637), .Y(n_636) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_504), .B(n_512), .Y(n_502) );
INVx1_ASAP7_75t_L g556 ( .A(n_504), .Y(n_556) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_508), .B(n_511), .Y(n_507) );
INVx2_ASAP7_75t_L g522 ( .A(n_511), .Y(n_522) );
INVx1_ASAP7_75t_L g557 ( .A(n_512), .Y(n_557) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_526), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_515), .B(n_548), .Y(n_547) );
AND2x4_ASAP7_75t_L g561 ( .A(n_515), .B(n_562), .Y(n_561) );
INVx3_ASAP7_75t_SL g566 ( .A(n_515), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_515), .B(n_553), .Y(n_619) );
OR2x2_ASAP7_75t_L g629 ( .A(n_515), .B(n_555), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_515), .B(n_597), .Y(n_657) );
OR2x2_ASAP7_75t_L g687 ( .A(n_515), .B(n_527), .Y(n_687) );
AND2x2_ASAP7_75t_L g691 ( .A(n_515), .B(n_528), .Y(n_691) );
NAND2xp5_ASAP7_75t_SL g704 ( .A(n_515), .B(n_567), .Y(n_704) );
AND2x2_ASAP7_75t_L g711 ( .A(n_515), .B(n_593), .Y(n_711) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_524), .Y(n_515) );
INVx1_ASAP7_75t_SL g654 ( .A(n_526), .Y(n_654) );
AND2x2_ASAP7_75t_L g593 ( .A(n_527), .B(n_555), .Y(n_593) );
AND2x2_ASAP7_75t_L g607 ( .A(n_527), .B(n_562), .Y(n_607) );
AND2x2_ASAP7_75t_L g610 ( .A(n_527), .B(n_566), .Y(n_610) );
INVx1_ASAP7_75t_L g637 ( .A(n_527), .Y(n_637) );
INVx2_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
BUFx2_ASAP7_75t_L g549 ( .A(n_528), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_541), .Y(n_538) );
A2O1A1Ixp33_ASAP7_75t_L g708 ( .A1(n_539), .A2(n_585), .B(n_709), .C(n_710), .Y(n_708) );
HB1xp67_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g615 ( .A(n_540), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_541), .B(n_558), .Y(n_573) );
AND2x2_ASAP7_75t_L g599 ( .A(n_541), .B(n_600), .Y(n_599) );
OAI21xp5_ASAP7_75t_SL g542 ( .A1(n_543), .A2(n_546), .B(n_550), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g643 ( .A(n_544), .B(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g570 ( .A(n_545), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_545), .B(n_566), .Y(n_611) );
AND2x2_ASAP7_75t_L g702 ( .A(n_545), .B(n_553), .Y(n_702) );
INVxp67_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g575 ( .A(n_549), .B(n_562), .Y(n_575) );
OR2x2_ASAP7_75t_L g576 ( .A(n_549), .B(n_560), .Y(n_576) );
OAI322xp33_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_559), .A3(n_560), .B1(n_563), .B2(n_564), .C1(n_568), .C2(n_569), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_558), .Y(n_552) );
AND2x2_ASAP7_75t_L g663 ( .A(n_553), .B(n_575), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_553), .B(n_627), .Y(n_709) );
INVx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AND2x2_ASAP7_75t_L g606 ( .A(n_555), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
OR2x2_ASAP7_75t_L g672 ( .A(n_559), .B(n_585), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_560), .B(n_654), .Y(n_653) );
INVx3_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_561), .B(n_593), .Y(n_650) );
AND2x2_ASAP7_75t_L g596 ( .A(n_562), .B(n_566), .Y(n_596) );
AND2x2_ASAP7_75t_L g604 ( .A(n_563), .B(n_605), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g701 ( .A1(n_563), .A2(n_642), .B(n_702), .C(n_703), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g674 ( .A1(n_564), .A2(n_577), .B(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_566), .B(n_593), .Y(n_633) );
AND2x2_ASAP7_75t_L g639 ( .A(n_566), .B(n_607), .Y(n_639) );
AND2x2_ASAP7_75t_L g673 ( .A(n_566), .B(n_575), .Y(n_673) );
NOR2xp33_ASAP7_75t_L g581 ( .A(n_567), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_SL g683 ( .A(n_567), .Y(n_683) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g598 ( .A1(n_571), .A2(n_599), .B1(n_601), .B2(n_606), .Y(n_598) );
OAI22xp5_ASAP7_75t_SL g572 ( .A1(n_573), .A2(n_574), .B1(n_576), .B2(n_577), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g608 ( .A1(n_573), .A2(n_609), .B1(n_611), .B2(n_612), .Y(n_608) );
INVxp67_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_SL g577 ( .A(n_578), .Y(n_577) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_578), .A2(n_680), .B1(n_682), .B2(n_684), .C(n_688), .Y(n_679) );
AOI211xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_583), .B(n_587), .C(n_608), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
OR2x2_ASAP7_75t_L g649 ( .A(n_585), .B(n_602), .Y(n_649) );
INVx1_ASAP7_75t_L g700 ( .A(n_585), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g587 ( .A1(n_586), .A2(n_588), .B1(n_592), .B2(n_595), .C(n_598), .Y(n_587) );
INVx2_ASAP7_75t_SL g642 ( .A(n_586), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g707 ( .A(n_589), .Y(n_707) );
AND2x2_ASAP7_75t_L g631 ( .A(n_590), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g616 ( .A(n_591), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
INVx1_ASAP7_75t_L g678 ( .A(n_594), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
AND2x2_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
NOR2xp33_ASAP7_75t_L g703 ( .A(n_602), .B(n_704), .Y(n_703) );
CKINVDCx16_ASAP7_75t_R g602 ( .A(n_603), .Y(n_602) );
INVxp67_ASAP7_75t_L g647 ( .A(n_605), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g617 ( .A1(n_606), .A2(n_618), .B(n_620), .C(n_622), .Y(n_617) );
INVx1_ASAP7_75t_L g695 ( .A(n_609), .Y(n_695) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g670 ( .A(n_613), .B(n_671), .Y(n_670) );
AND2x2_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
INVx2_ASAP7_75t_L g626 ( .A(n_616), .Y(n_626) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
OAI222xp33_ASAP7_75t_L g622 ( .A1(n_623), .A2(n_629), .B1(n_630), .B2(n_633), .C1(n_634), .C2(n_636), .Y(n_622) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_SL g662 ( .A(n_626), .Y(n_662) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_629), .B(n_683), .Y(n_682) );
NAND2xp33_ASAP7_75t_SL g660 ( .A(n_630), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_SL g635 ( .A(n_632), .Y(n_635) );
AND2x2_ASAP7_75t_L g699 ( .A(n_632), .B(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g665 ( .A(n_635), .B(n_662), .Y(n_665) );
INVx1_ASAP7_75t_L g694 ( .A(n_636), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_643), .C(n_648), .Y(n_638) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_642), .B(n_662), .Y(n_661) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_645), .A2(n_673), .A3(n_678), .B1(n_694), .B2(n_695), .C1(n_696), .C2(n_699), .Y(n_693) );
AND2x2_ASAP7_75t_L g680 ( .A(n_646), .B(n_681), .Y(n_680) );
OAI22xp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_650), .B1(n_651), .B2(n_653), .Y(n_648) );
INVxp33_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g655 ( .A1(n_656), .A2(n_658), .B1(n_660), .B2(n_663), .C(n_664), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
NAND5xp2_ASAP7_75t_L g667 ( .A(n_668), .B(n_679), .C(n_693), .D(n_701), .E(n_705), .Y(n_667) );
AOI21xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_673), .B(n_674), .Y(n_668) );
INVxp67_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVxp33_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_678), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_681), .A2(n_706), .B(n_707), .C(n_708), .Y(n_705) );
AOI31xp33_ASAP7_75t_L g688 ( .A1(n_683), .A2(n_689), .A3(n_690), .B(n_692), .Y(n_688) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_698), .Y(n_696) );
INVx1_ASAP7_75t_L g706 ( .A(n_704), .Y(n_706) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_712), .Y(n_717) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
endmodule