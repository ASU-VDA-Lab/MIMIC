module real_aes_16568_n_312 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_19, n_40, n_239, n_100, n_54, n_112, n_35, n_42, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_73, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_292, n_116, n_94, n_289, n_280, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_93, n_182, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_183, n_266, n_205, n_177, n_22, n_140, n_219, n_180, n_212, n_210, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_312);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_19;
input n_40;
input n_239;
input n_100;
input n_54;
input n_112;
input n_35;
input n_42;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_73;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_93;
input n_182;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_183;
input n_266;
input n_205;
input n_177;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_312;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_1328;
wire n_571;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1250;
wire n_1284;
wire n_1095;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1666;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_328;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_1338;
wire n_981;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1671;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_1226;
wire n_525;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1257;
wire n_1082;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1352;
wire n_1280;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g896 ( .A(n_0), .Y(n_896) );
AO22x1_ASAP7_75t_L g922 ( .A1(n_0), .A2(n_205), .B1(n_596), .B2(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g327 ( .A(n_1), .Y(n_327) );
NOR2xp33_ASAP7_75t_L g363 ( .A(n_1), .B(n_337), .Y(n_363) );
AND2x2_ASAP7_75t_L g580 ( .A(n_1), .B(n_223), .Y(n_580) );
AND2x2_ASAP7_75t_L g598 ( .A(n_1), .B(n_484), .Y(n_598) );
INVx1_ASAP7_75t_L g905 ( .A(n_2), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_2), .A2(n_116), .B1(n_500), .B2(n_921), .Y(n_920) );
AOI22xp33_ASAP7_75t_SL g1202 ( .A1(n_3), .A2(n_277), .B1(n_844), .B2(n_1158), .Y(n_1202) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_3), .A2(n_5), .B1(n_601), .B2(n_608), .C(n_1217), .Y(n_1216) );
AOI22xp33_ASAP7_75t_SL g540 ( .A1(n_4), .A2(n_37), .B1(n_541), .B2(n_545), .Y(n_540) );
INVxp67_ASAP7_75t_SL g636 ( .A(n_4), .Y(n_636) );
AOI22xp33_ASAP7_75t_SL g1208 ( .A1(n_5), .A2(n_9), .B1(n_557), .B2(n_839), .Y(n_1208) );
AOI22xp33_ASAP7_75t_SL g1157 ( .A1(n_6), .A2(n_274), .B1(n_826), .B2(n_1158), .Y(n_1157) );
AOI221xp5_ASAP7_75t_L g1174 ( .A1(n_6), .A2(n_228), .B1(n_1087), .B2(n_1175), .C(n_1176), .Y(n_1174) );
INVx1_ASAP7_75t_L g1301 ( .A(n_7), .Y(n_1301) );
XOR2x2_ASAP7_75t_L g345 ( .A(n_8), .B(n_346), .Y(n_345) );
A2O1A1Ixp33_ASAP7_75t_L g1225 ( .A1(n_9), .A2(n_874), .B(n_1226), .C(n_1231), .Y(n_1225) );
OAI22xp5_ASAP7_75t_L g1366 ( .A1(n_10), .A2(n_195), .B1(n_821), .B2(n_1367), .Y(n_1366) );
AOI22xp33_ASAP7_75t_SL g835 ( .A1(n_11), .A2(n_198), .B1(n_836), .B2(n_837), .Y(n_835) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_11), .Y(n_872) );
INVxp67_ASAP7_75t_SL g1238 ( .A(n_12), .Y(n_1238) );
AND4x1_ASAP7_75t_L g1275 ( .A(n_12), .B(n_1240), .C(n_1243), .D(n_1260), .Y(n_1275) );
AOI22xp33_ASAP7_75t_L g1656 ( .A1(n_13), .A2(n_289), .B1(n_935), .B2(n_1133), .Y(n_1656) );
INVx1_ASAP7_75t_L g1674 ( .A(n_13), .Y(n_1674) );
INVx2_ASAP7_75t_L g398 ( .A(n_14), .Y(n_398) );
OAI22xp5_ASAP7_75t_SL g1079 ( .A1(n_15), .A2(n_252), .B1(n_973), .B2(n_1080), .Y(n_1079) );
OAI221xp5_ASAP7_75t_L g1093 ( .A1(n_15), .A2(n_252), .B1(n_626), .B2(n_628), .C(n_1094), .Y(n_1093) );
XNOR2x1_ASAP7_75t_L g1057 ( .A(n_16), .B(n_1058), .Y(n_1057) );
AOI22xp5_ASAP7_75t_L g1394 ( .A1(n_16), .A2(n_18), .B1(n_1378), .B2(n_1385), .Y(n_1394) );
INVx1_ASAP7_75t_L g1349 ( .A(n_17), .Y(n_1349) );
INVx1_ASAP7_75t_L g1347 ( .A(n_19), .Y(n_1347) );
AOI22xp33_ASAP7_75t_L g1358 ( .A1(n_19), .A2(n_60), .B1(n_859), .B2(n_1359), .Y(n_1358) );
OAI22xp5_ASAP7_75t_L g1242 ( .A1(n_20), .A2(n_145), .B1(n_585), .B2(n_589), .Y(n_1242) );
OAI211xp5_ASAP7_75t_L g1244 ( .A1(n_20), .A2(n_1034), .B(n_1245), .C(n_1248), .Y(n_1244) );
AOI22xp33_ASAP7_75t_L g1252 ( .A1(n_21), .A2(n_81), .B1(n_923), .B2(n_993), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1269 ( .A1(n_21), .A2(n_29), .B1(n_550), .B2(n_1268), .Y(n_1269) );
HB1xp67_ASAP7_75t_L g322 ( .A(n_22), .Y(n_322) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_22), .B(n_320), .Y(n_1379) );
INVx1_ASAP7_75t_L g1092 ( .A(n_23), .Y(n_1092) );
AOI22xp33_ASAP7_75t_L g1447 ( .A1(n_24), .A2(n_172), .B1(n_1378), .B2(n_1434), .Y(n_1447) );
CKINVDCx5p33_ASAP7_75t_R g810 ( .A(n_25), .Y(n_810) );
INVx1_ASAP7_75t_L g1007 ( .A(n_26), .Y(n_1007) );
OAI211xp5_ASAP7_75t_L g1016 ( .A1(n_26), .A2(n_863), .B(n_1017), .C(n_1024), .Y(n_1016) );
INVxp67_ASAP7_75t_L g1149 ( .A(n_27), .Y(n_1149) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_28), .Y(n_1241) );
AOI221xp5_ASAP7_75t_L g1258 ( .A1(n_29), .A2(n_295), .B1(n_646), .B2(n_921), .C(n_1259), .Y(n_1258) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_30), .A2(n_42), .B1(n_551), .B2(n_721), .Y(n_783) );
INVx1_ASAP7_75t_L g796 ( .A(n_30), .Y(n_796) );
INVx1_ASAP7_75t_L g693 ( .A(n_31), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g657 ( .A1(n_32), .A2(n_40), .B1(n_658), .B2(n_659), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_32), .A2(n_143), .B1(n_720), .B2(n_722), .Y(n_719) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_33), .A2(n_89), .B1(n_1155), .B2(n_1204), .Y(n_1203) );
AOI221xp5_ASAP7_75t_L g1227 ( .A1(n_33), .A2(n_177), .B1(n_1104), .B2(n_1176), .C(n_1228), .Y(n_1227) );
AOI221xp5_ASAP7_75t_L g1030 ( .A1(n_34), .A2(n_270), .B1(n_641), .B2(n_921), .C(n_1031), .Y(n_1030) );
INVxp67_ASAP7_75t_SL g1041 ( .A(n_34), .Y(n_1041) );
INVx1_ASAP7_75t_L g1013 ( .A(n_35), .Y(n_1013) );
OAI22xp5_ASAP7_75t_L g1032 ( .A1(n_35), .A2(n_189), .B1(n_1033), .B2(n_1034), .Y(n_1032) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_36), .A2(n_303), .B1(n_454), .B2(n_773), .C(n_774), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g794 ( .A1(n_36), .A2(n_109), .B1(n_787), .B2(n_788), .C(n_795), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_37), .A2(n_94), .B1(n_601), .B2(n_603), .C(n_607), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_38), .A2(n_251), .B1(n_829), .B2(n_833), .Y(n_832) );
INVx1_ASAP7_75t_L g865 ( .A(n_38), .Y(n_865) );
INVx1_ASAP7_75t_L g1659 ( .A(n_39), .Y(n_1659) );
AOI22xp33_ASAP7_75t_SL g706 ( .A1(n_40), .A2(n_152), .B1(n_707), .B2(n_709), .Y(n_706) );
INVx1_ASAP7_75t_L g1658 ( .A(n_41), .Y(n_1658) );
INVx1_ASAP7_75t_L g790 ( .A(n_42), .Y(n_790) );
INVxp67_ASAP7_75t_SL g1029 ( .A(n_43), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_43), .A2(n_125), .B1(n_1053), .B2(n_1054), .Y(n_1052) );
AOI22xp5_ASAP7_75t_L g1432 ( .A1(n_44), .A2(n_190), .B1(n_1385), .B2(n_1388), .Y(n_1432) );
AOI22xp5_ASAP7_75t_L g1403 ( .A1(n_45), .A2(n_292), .B1(n_1378), .B2(n_1382), .Y(n_1403) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_46), .Y(n_334) );
INVx1_ASAP7_75t_L g1246 ( .A(n_47), .Y(n_1246) );
OAI22xp33_ASAP7_75t_L g1262 ( .A1(n_47), .A2(n_96), .B1(n_559), .B2(n_1263), .Y(n_1262) );
AOI21xp33_ASAP7_75t_L g1614 ( .A1(n_48), .A2(n_788), .B(n_1104), .Y(n_1614) );
AOI221xp5_ASAP7_75t_L g1631 ( .A1(n_48), .A2(n_235), .B1(n_1155), .B2(n_1632), .C(n_1633), .Y(n_1631) );
AOI22xp5_ASAP7_75t_L g1433 ( .A1(n_49), .A2(n_276), .B1(n_1378), .B2(n_1434), .Y(n_1433) );
INVx1_ASAP7_75t_L g819 ( .A(n_50), .Y(n_819) );
AOI22xp5_ASAP7_75t_L g1384 ( .A1(n_51), .A2(n_118), .B1(n_1385), .B2(n_1388), .Y(n_1384) );
OAI222xp33_ASAP7_75t_L g1589 ( .A1(n_52), .A2(n_66), .B1(n_72), .B2(n_821), .C1(n_1590), .C2(n_1592), .Y(n_1589) );
INVx1_ASAP7_75t_L g1091 ( .A(n_53), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g546 ( .A1(n_54), .A2(n_230), .B1(n_547), .B2(n_550), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_54), .A2(n_127), .B1(n_610), .B2(n_612), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_55), .Y(n_1211) );
INVx1_ASAP7_75t_L g369 ( .A(n_56), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_57), .A2(n_141), .B1(n_833), .B2(n_1154), .Y(n_1161) );
AOI21xp33_ASAP7_75t_L g1184 ( .A1(n_57), .A2(n_646), .B(n_1185), .Y(n_1184) );
CKINVDCx5p33_ASAP7_75t_R g1598 ( .A(n_58), .Y(n_1598) );
AOI221xp5_ASAP7_75t_L g1249 ( .A1(n_59), .A2(n_294), .B1(n_856), .B2(n_1185), .C(n_1250), .Y(n_1249) );
AOI22xp33_ASAP7_75t_SL g1270 ( .A1(n_59), .A2(n_265), .B1(n_720), .B2(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1337 ( .A(n_60), .Y(n_1337) );
INVx1_ASAP7_75t_L g1199 ( .A(n_61), .Y(n_1199) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_62), .A2(n_291), .B1(n_662), .B2(n_664), .C(n_666), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g712 ( .A1(n_62), .A2(n_259), .B1(n_713), .B2(n_715), .C(n_718), .Y(n_712) );
AOI22xp33_ASAP7_75t_SL g825 ( .A1(n_63), .A2(n_155), .B1(n_713), .B2(n_826), .Y(n_825) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_63), .Y(n_871) );
OAI211xp5_ASAP7_75t_SL g763 ( .A1(n_64), .A2(n_731), .B(n_738), .C(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g799 ( .A(n_64), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_65), .A2(n_222), .B1(n_443), .B2(n_447), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_65), .A2(n_222), .B1(n_488), .B2(n_490), .Y(n_487) );
CKINVDCx5p33_ASAP7_75t_R g1164 ( .A(n_67), .Y(n_1164) );
OAI21xp5_ASAP7_75t_SL g1190 ( .A1(n_68), .A2(n_585), .B(n_1191), .Y(n_1190) );
AOI22xp33_ASAP7_75t_L g1293 ( .A1(n_69), .A2(n_209), .B1(n_545), .B2(n_836), .Y(n_1293) );
AOI22xp33_ASAP7_75t_SL g1321 ( .A1(n_69), .A2(n_257), .B1(n_993), .B2(n_1133), .Y(n_1321) );
INVxp67_ASAP7_75t_SL g699 ( .A(n_70), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_70), .A2(n_299), .B1(n_724), .B2(n_727), .Y(n_723) );
AOI22xp33_ASAP7_75t_SL g1160 ( .A1(n_71), .A2(n_228), .B1(n_557), .B2(n_837), .Y(n_1160) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_71), .A2(n_274), .B1(n_980), .B2(n_993), .Y(n_1183) );
OAI22xp5_ASAP7_75t_L g1620 ( .A1(n_72), .A2(n_305), .B1(n_1314), .B2(n_1621), .Y(n_1620) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_73), .A2(n_94), .B1(n_545), .B2(n_555), .Y(n_554) );
INVxp67_ASAP7_75t_SL g639 ( .A(n_73), .Y(n_639) );
OR2x2_ASAP7_75t_L g1011 ( .A(n_74), .B(n_575), .Y(n_1011) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_75), .A2(n_187), .B1(n_628), .B2(n_1026), .C(n_1027), .Y(n_1025) );
OAI322xp33_ASAP7_75t_L g1039 ( .A1(n_75), .A2(n_429), .A3(n_566), .B1(n_1040), .B2(n_1043), .C1(n_1044), .C2(n_1047), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1121 ( .A1(n_76), .A2(n_181), .B1(n_722), .B2(n_829), .Y(n_1121) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_76), .A2(n_86), .B1(n_613), .B2(n_1133), .Y(n_1132) );
AOI22xp33_ASAP7_75t_SL g1292 ( .A1(n_77), .A2(n_202), .B1(n_709), .B2(n_1290), .Y(n_1292) );
INVx1_ASAP7_75t_L g1316 ( .A(n_77), .Y(n_1316) );
INVx1_ASAP7_75t_L g1061 ( .A(n_78), .Y(n_1061) );
AOI22xp33_ASAP7_75t_SL g1069 ( .A1(n_79), .A2(n_254), .B1(n_963), .B2(n_1070), .Y(n_1069) );
AOI221xp5_ASAP7_75t_L g1086 ( .A1(n_79), .A2(n_88), .B1(n_855), .B2(n_1023), .C(n_1087), .Y(n_1086) );
INVx1_ASAP7_75t_L g880 ( .A(n_80), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g1267 ( .A1(n_81), .A2(n_295), .B1(n_550), .B2(n_1268), .Y(n_1267) );
AOI22xp5_ASAP7_75t_L g1410 ( .A1(n_82), .A2(n_304), .B1(n_1385), .B2(n_1388), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g971 ( .A1(n_83), .A2(n_243), .B1(n_541), .B2(n_963), .Y(n_971) );
AOI221xp5_ASAP7_75t_L g978 ( .A1(n_83), .A2(n_238), .B1(n_602), .B2(n_608), .C(n_788), .Y(n_978) );
AOI22xp33_ASAP7_75t_L g1615 ( .A1(n_84), .A2(n_139), .B1(n_613), .B2(n_1137), .Y(n_1615) );
INVx1_ASAP7_75t_L g1626 ( .A(n_84), .Y(n_1626) );
INVx1_ASAP7_75t_L g1063 ( .A(n_85), .Y(n_1063) );
AOI22xp33_ASAP7_75t_SL g1124 ( .A1(n_86), .A2(n_256), .B1(n_722), .B2(n_829), .Y(n_1124) );
INVx1_ASAP7_75t_L g961 ( .A(n_87), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g979 ( .A1(n_87), .A2(n_263), .B1(n_613), .B2(n_980), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_88), .A2(n_170), .B1(n_713), .B2(n_1053), .Y(n_1078) );
AOI22xp33_ASAP7_75t_SL g1219 ( .A1(n_89), .A2(n_124), .B1(n_612), .B2(n_1133), .Y(n_1219) );
INVx1_ASAP7_75t_L g365 ( .A(n_90), .Y(n_365) );
INVx1_ASAP7_75t_L g1346 ( .A(n_91), .Y(n_1346) );
AOI221xp5_ASAP7_75t_L g1354 ( .A1(n_91), .A2(n_203), .B1(n_641), .B2(n_646), .C(n_1175), .Y(n_1354) );
CKINVDCx5p33_ASAP7_75t_R g1117 ( .A(n_92), .Y(n_1117) );
CKINVDCx5p33_ASAP7_75t_R g1172 ( .A(n_93), .Y(n_1172) );
AOI22xp5_ASAP7_75t_SL g1411 ( .A1(n_95), .A2(n_200), .B1(n_1378), .B2(n_1382), .Y(n_1411) );
INVx1_ASAP7_75t_L g1247 ( .A(n_96), .Y(n_1247) );
INVx1_ASAP7_75t_L g1028 ( .A(n_97), .Y(n_1028) );
CKINVDCx5p33_ASAP7_75t_R g1167 ( .A(n_98), .Y(n_1167) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_98), .A2(n_114), .B1(n_1188), .B2(n_1189), .Y(n_1187) );
INVx1_ASAP7_75t_L g391 ( .A(n_99), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g1665 ( .A1(n_100), .A2(n_788), .B(n_1666), .Y(n_1665) );
INVx1_ASAP7_75t_L g1673 ( .A(n_100), .Y(n_1673) );
INVx1_ASAP7_75t_L g950 ( .A(n_101), .Y(n_950) );
OAI221xp5_ASAP7_75t_L g1253 ( .A1(n_102), .A2(n_240), .B1(n_624), .B2(n_875), .C(n_1254), .Y(n_1253) );
INVx1_ASAP7_75t_L g1274 ( .A(n_102), .Y(n_1274) );
INVx1_ASAP7_75t_L g320 ( .A(n_103), .Y(n_320) );
AOI221xp5_ASAP7_75t_L g1653 ( .A1(n_104), .A2(n_224), .B1(n_608), .B2(n_787), .C(n_1654), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1675 ( .A1(n_104), .A2(n_156), .B1(n_541), .B2(n_572), .Y(n_1675) );
INVx1_ASAP7_75t_L g1112 ( .A(n_105), .Y(n_1112) );
INVx1_ASAP7_75t_L g1111 ( .A(n_106), .Y(n_1111) );
AOI221xp5_ASAP7_75t_L g1119 ( .A1(n_107), .A2(n_255), .B1(n_839), .B2(n_1053), .C(n_1120), .Y(n_1119) );
AOI221xp5_ASAP7_75t_L g1131 ( .A1(n_107), .A2(n_207), .B1(n_602), .B2(n_604), .C(n_1087), .Y(n_1131) );
AOI22xp33_ASAP7_75t_L g828 ( .A1(n_108), .A2(n_162), .B1(n_829), .B2(n_830), .Y(n_828) );
INVx1_ASAP7_75t_L g869 ( .A(n_108), .Y(n_869) );
INVx1_ASAP7_75t_L g779 ( .A(n_109), .Y(n_779) );
OAI22xp33_ASAP7_75t_L g1333 ( .A1(n_110), .A2(n_267), .B1(n_559), .B2(n_1263), .Y(n_1333) );
INVx1_ASAP7_75t_L g1361 ( .A(n_110), .Y(n_1361) );
AOI22xp5_ASAP7_75t_L g1407 ( .A1(n_111), .A2(n_285), .B1(n_1382), .B2(n_1388), .Y(n_1407) );
OAI222xp33_ASAP7_75t_L g910 ( .A1(n_112), .A2(n_290), .B1(n_734), .B2(n_736), .C1(n_911), .C2(n_914), .Y(n_910) );
INVx1_ASAP7_75t_L g926 ( .A(n_112), .Y(n_926) );
INVx1_ASAP7_75t_L g531 ( .A(n_113), .Y(n_531) );
OAI221xp5_ASAP7_75t_L g623 ( .A1(n_113), .A2(n_115), .B1(n_624), .B2(n_628), .C(n_632), .Y(n_623) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_114), .Y(n_1166) );
INVx1_ASAP7_75t_L g522 ( .A(n_115), .Y(n_522) );
INVx1_ASAP7_75t_L g901 ( .A(n_116), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g968 ( .A(n_117), .Y(n_968) );
OAI22xp33_ASAP7_75t_L g741 ( .A1(n_119), .A2(n_148), .B1(n_742), .B2(n_745), .Y(n_741) );
INVxp67_ASAP7_75t_SL g750 ( .A(n_119), .Y(n_750) );
INVx1_ASAP7_75t_L g1338 ( .A(n_120), .Y(n_1338) );
AOI221xp5_ASAP7_75t_L g1357 ( .A1(n_120), .A2(n_248), .B1(n_607), .B2(n_641), .C(n_1228), .Y(n_1357) );
INVx1_ASAP7_75t_L g957 ( .A(n_121), .Y(n_957) );
AOI21xp33_ASAP7_75t_L g991 ( .A1(n_121), .A2(n_646), .B(n_788), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g951 ( .A1(n_122), .A2(n_147), .B1(n_589), .B2(n_952), .Y(n_951) );
OAI211xp5_ASAP7_75t_L g976 ( .A1(n_122), .A2(n_594), .B(n_977), .C(n_983), .Y(n_976) );
INVx1_ASAP7_75t_L g814 ( .A(n_123), .Y(n_814) );
OAI222xp33_ASAP7_75t_L g862 ( .A1(n_123), .A2(n_184), .B1(n_863), .B2(n_864), .C1(n_870), .C2(n_875), .Y(n_862) );
AOI22xp33_ASAP7_75t_L g1206 ( .A1(n_124), .A2(n_177), .B1(n_1155), .B2(n_1207), .Y(n_1206) );
AOI221xp5_ASAP7_75t_L g1022 ( .A1(n_125), .A2(n_197), .B1(n_608), .B2(n_921), .C(n_1023), .Y(n_1022) );
OAI22xp33_ASAP7_75t_L g762 ( .A1(n_126), .A2(n_310), .B1(n_742), .B2(n_745), .Y(n_762) );
INVxp33_ASAP7_75t_SL g803 ( .A(n_126), .Y(n_803) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_127), .A2(n_154), .B1(n_547), .B2(n_550), .Y(n_552) );
INVx1_ASAP7_75t_L g1283 ( .A(n_128), .Y(n_1283) );
OAI221xp5_ASAP7_75t_L g1313 ( .A1(n_128), .A2(n_129), .B1(n_876), .B2(n_1314), .C(n_1315), .Y(n_1313) );
INVx1_ASAP7_75t_L g1284 ( .A(n_129), .Y(n_1284) );
CKINVDCx5p33_ASAP7_75t_R g765 ( .A(n_130), .Y(n_765) );
OA21x2_ASAP7_75t_L g1059 ( .A1(n_131), .A2(n_575), .B(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g769 ( .A(n_132), .Y(n_769) );
AOI221xp5_ASAP7_75t_L g786 ( .A1(n_132), .A2(n_219), .B1(n_787), .B2(n_788), .C(n_789), .Y(n_786) );
AOI221xp5_ASAP7_75t_L g677 ( .A1(n_133), .A2(n_143), .B1(n_659), .B2(n_678), .C(n_680), .Y(n_677) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_133), .A2(n_291), .B1(n_541), .B2(n_545), .C(n_711), .Y(n_710) );
XNOR2xp5_ASAP7_75t_L g1647 ( .A(n_134), .B(n_1648), .Y(n_1647) );
OAI22xp33_ASAP7_75t_L g558 ( .A1(n_135), .A2(n_250), .B1(n_559), .B2(n_566), .Y(n_558) );
INVx1_ASAP7_75t_L g620 ( .A(n_135), .Y(n_620) );
INVx1_ASAP7_75t_L g845 ( .A(n_136), .Y(n_845) );
OAI22xp33_ASAP7_75t_L g467 ( .A1(n_137), .A2(n_144), .B1(n_468), .B2(n_471), .Y(n_467) );
OAI22xp33_ASAP7_75t_L g479 ( .A1(n_137), .A2(n_144), .B1(n_480), .B2(n_481), .Y(n_479) );
OAI221xp5_ASAP7_75t_L g1660 ( .A1(n_138), .A2(n_300), .B1(n_876), .B2(n_1314), .C(n_1661), .Y(n_1660) );
OAI22xp33_ASAP7_75t_L g1680 ( .A1(n_138), .A2(n_300), .B1(n_524), .B2(n_973), .Y(n_1680) );
INVxp67_ASAP7_75t_SL g1634 ( .A(n_139), .Y(n_1634) );
AO22x1_ASAP7_75t_L g1153 ( .A1(n_140), .A2(n_175), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_140), .B(n_1181), .Y(n_1180) );
AOI22xp33_ASAP7_75t_SL g1177 ( .A1(n_141), .A2(n_175), .B1(n_610), .B2(n_1178), .Y(n_1177) );
INVx1_ASAP7_75t_L g457 ( .A(n_142), .Y(n_457) );
INVx1_ASAP7_75t_L g379 ( .A(n_146), .Y(n_379) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_148), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g584 ( .A1(n_149), .A2(n_167), .B1(n_585), .B2(n_589), .Y(n_584) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_149), .A2(n_594), .B(n_599), .C(n_615), .Y(n_593) );
INVx1_ASAP7_75t_L g898 ( .A(n_150), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_150), .A2(n_231), .B1(n_923), .B2(n_935), .Y(n_934) );
INVx1_ASAP7_75t_L g1444 ( .A(n_151), .Y(n_1444) );
INVx1_ASAP7_75t_L g681 ( .A(n_152), .Y(n_681) );
AOI22xp5_ASAP7_75t_SL g1377 ( .A1(n_153), .A2(n_161), .B1(n_1378), .B2(n_1382), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_154), .A2(n_230), .B1(n_641), .B2(n_642), .C(n_646), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g850 ( .A1(n_155), .A2(n_198), .B1(n_851), .B2(n_854), .C(n_856), .Y(n_850) );
AOI22xp33_ASAP7_75t_SL g1667 ( .A1(n_156), .A2(n_275), .B1(n_596), .B2(n_610), .Y(n_1667) );
OAI211xp5_ASAP7_75t_L g1651 ( .A1(n_157), .A2(n_594), .B(n_1652), .C(n_1657), .Y(n_1651) );
OAI22xp5_ASAP7_75t_L g1683 ( .A1(n_157), .A2(n_293), .B1(n_589), .B2(n_952), .Y(n_1683) );
AOI22xp33_ASAP7_75t_SL g1289 ( .A1(n_158), .A2(n_260), .B1(n_709), .B2(n_1290), .Y(n_1289) );
AOI22xp33_ASAP7_75t_L g1308 ( .A1(n_158), .A2(n_202), .B1(n_613), .B2(n_1309), .Y(n_1308) );
INVx1_ASAP7_75t_L g1613 ( .A(n_159), .Y(n_1613) );
AOI221x1_ASAP7_75t_SL g1624 ( .A1(n_159), .A2(n_232), .B1(n_1155), .B2(n_1207), .C(n_1625), .Y(n_1624) );
INVx1_ASAP7_75t_L g1068 ( .A(n_160), .Y(n_1068) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_160), .A2(n_201), .B1(n_604), .B2(n_1101), .C(n_1104), .Y(n_1100) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_162), .A2(n_251), .B1(n_858), .B2(n_859), .Y(n_857) );
AOI21xp33_ASAP7_75t_L g1618 ( .A1(n_163), .A2(n_855), .B(n_1087), .Y(n_1618) );
INVx1_ASAP7_75t_L g1635 ( .A(n_163), .Y(n_1635) );
AOI221xp5_ASAP7_75t_L g1122 ( .A1(n_164), .A2(n_207), .B1(n_713), .B2(n_1053), .C(n_1123), .Y(n_1122) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_164), .A2(n_255), .B1(n_613), .B2(n_1137), .Y(n_1136) );
INVx2_ASAP7_75t_L g1381 ( .A(n_165), .Y(n_1381) );
AND2x2_ASAP7_75t_L g1383 ( .A(n_165), .B(n_264), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1389 ( .A(n_165), .B(n_1387), .Y(n_1389) );
CKINVDCx5p33_ASAP7_75t_R g1038 ( .A(n_166), .Y(n_1038) );
INVx1_ASAP7_75t_L g986 ( .A(n_168), .Y(n_986) );
AOI22xp5_ASAP7_75t_SL g1392 ( .A1(n_169), .A2(n_226), .B1(n_1388), .B2(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1099 ( .A(n_170), .Y(n_1099) );
OAI22xp5_ASAP7_75t_L g1212 ( .A1(n_171), .A2(n_253), .B1(n_585), .B2(n_821), .Y(n_1212) );
OAI211xp5_ASAP7_75t_L g1214 ( .A1(n_171), .A2(n_1034), .B(n_1215), .C(n_1220), .Y(n_1214) );
CKINVDCx5p33_ASAP7_75t_R g1171 ( .A(n_173), .Y(n_1171) );
XOR2x2_ASAP7_75t_L g517 ( .A(n_174), .B(n_518), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g1399 ( .A1(n_174), .A2(n_282), .B1(n_1378), .B2(n_1393), .Y(n_1399) );
AOI22xp5_ASAP7_75t_L g1402 ( .A1(n_176), .A2(n_229), .B1(n_1385), .B2(n_1388), .Y(n_1402) );
INVx1_ASAP7_75t_L g942 ( .A(n_178), .Y(n_942) );
INVx1_ASAP7_75t_L g842 ( .A(n_179), .Y(n_842) );
AOI22xp33_ASAP7_75t_SL g962 ( .A1(n_180), .A2(n_238), .B1(n_541), .B2(n_963), .Y(n_962) );
AOI22xp33_ASAP7_75t_SL g992 ( .A1(n_180), .A2(n_243), .B1(n_610), .B2(n_993), .Y(n_992) );
AOI221xp5_ASAP7_75t_L g1138 ( .A1(n_181), .A2(n_256), .B1(n_604), .B2(n_646), .C(n_787), .Y(n_1138) );
INVx1_ASAP7_75t_L g1342 ( .A(n_182), .Y(n_1342) );
INVx1_ASAP7_75t_L g1077 ( .A(n_183), .Y(n_1077) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_183), .A2(n_242), .B1(n_935), .B2(n_1089), .Y(n_1088) );
INVx1_ASAP7_75t_L g816 ( .A(n_184), .Y(n_816) );
OAI211xp5_ASAP7_75t_L g451 ( .A1(n_185), .A2(n_427), .B(n_452), .C(n_456), .Y(n_451) );
INVx1_ASAP7_75t_L g506 ( .A(n_185), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g1408 ( .A1(n_186), .A2(n_246), .B1(n_1378), .B2(n_1385), .Y(n_1408) );
INVx1_ASAP7_75t_L g1006 ( .A(n_187), .Y(n_1006) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_188), .Y(n_900) );
INVx1_ASAP7_75t_L g1009 ( .A(n_189), .Y(n_1009) );
CKINVDCx5p33_ASAP7_75t_R g1662 ( .A(n_191), .Y(n_1662) );
OAI22xp5_ASAP7_75t_L g1302 ( .A1(n_192), .A2(n_308), .B1(n_566), .B2(n_1303), .Y(n_1302) );
INVx1_ASAP7_75t_L g1311 ( .A(n_192), .Y(n_1311) );
INVx1_ASAP7_75t_L g1055 ( .A(n_193), .Y(n_1055) );
INVx2_ASAP7_75t_L g397 ( .A(n_194), .Y(n_397) );
INVx1_ASAP7_75t_L g436 ( .A(n_194), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_194), .B(n_398), .Y(n_565) );
OAI211xp5_ASAP7_75t_L g1355 ( .A1(n_195), .A2(n_594), .B(n_1356), .C(n_1360), .Y(n_1355) );
INVx1_ASAP7_75t_L g908 ( .A(n_196), .Y(n_908) );
NAND2xp33_ASAP7_75t_SL g936 ( .A(n_196), .B(n_500), .Y(n_936) );
INVx1_ASAP7_75t_L g1045 ( .A(n_197), .Y(n_1045) );
INVx1_ASAP7_75t_L g390 ( .A(n_199), .Y(n_390) );
INVx1_ASAP7_75t_L g1587 ( .A(n_200), .Y(n_1587) );
AOI22xp33_ASAP7_75t_L g1640 ( .A1(n_200), .A2(n_1641), .B1(n_1646), .B2(n_1685), .Y(n_1640) );
INVx1_ASAP7_75t_L g1076 ( .A(n_201), .Y(n_1076) );
INVx1_ASAP7_75t_L g1343 ( .A(n_203), .Y(n_1343) );
INVx1_ASAP7_75t_L g1021 ( .A(n_204), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g909 ( .A1(n_205), .A2(n_711), .B(n_721), .Y(n_909) );
INVx1_ASAP7_75t_L g938 ( .A(n_206), .Y(n_938) );
BUFx3_ASAP7_75t_L g403 ( .A(n_208), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g1307 ( .A1(n_209), .A2(n_216), .B1(n_602), .B2(n_608), .C(n_788), .Y(n_1307) );
INVx1_ASAP7_75t_L g1129 ( .A(n_210), .Y(n_1129) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_211), .Y(n_766) );
OAI22xp5_ASAP7_75t_L g1330 ( .A1(n_212), .A2(n_217), .B1(n_524), .B2(n_1331), .Y(n_1330) );
OAI221xp5_ASAP7_75t_L g1352 ( .A1(n_212), .A2(n_217), .B1(n_624), .B2(n_875), .C(n_1353), .Y(n_1352) );
AOI22xp5_ASAP7_75t_L g1398 ( .A1(n_213), .A2(n_244), .B1(n_1385), .B2(n_1388), .Y(n_1398) );
OAI22xp5_ASAP7_75t_SL g1600 ( .A1(n_214), .A2(n_247), .B1(n_576), .B2(n_588), .Y(n_1600) );
CKINVDCx5p33_ASAP7_75t_R g1608 ( .A(n_214), .Y(n_1608) );
INVx1_ASAP7_75t_L g891 ( .A(n_215), .Y(n_891) );
NOR2xp33_ASAP7_75t_L g893 ( .A(n_215), .B(n_742), .Y(n_893) );
AOI22xp33_ASAP7_75t_SL g1288 ( .A1(n_216), .A2(n_257), .B1(n_545), .B2(n_826), .Y(n_1288) );
AOI22xp5_ASAP7_75t_L g1326 ( .A1(n_218), .A2(n_1327), .B1(n_1328), .B2(n_1368), .Y(n_1326) );
INVx1_ASAP7_75t_L g1368 ( .A(n_218), .Y(n_1368) );
AOI21xp33_ASAP7_75t_L g782 ( .A1(n_219), .A2(n_717), .B(n_718), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_220), .B(n_1279), .Y(n_1278) );
AOI22xp5_ASAP7_75t_L g1297 ( .A1(n_220), .A2(n_1298), .B1(n_1299), .B2(n_1322), .Y(n_1297) );
INVx1_ASAP7_75t_L g1324 ( .A(n_220), .Y(n_1324) );
OAI22xp33_ASAP7_75t_L g1209 ( .A1(n_221), .A2(n_237), .B1(n_559), .B2(n_566), .Y(n_1209) );
INVx1_ASAP7_75t_L g1221 ( .A(n_221), .Y(n_1221) );
BUFx3_ASAP7_75t_L g337 ( .A(n_223), .Y(n_337) );
INVx1_ASAP7_75t_L g484 ( .A(n_223), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g1679 ( .A1(n_224), .A2(n_275), .B1(n_541), .B2(n_713), .Y(n_1679) );
XNOR2x1_ASAP7_75t_L g1108 ( .A(n_225), .B(n_1109), .Y(n_1108) );
CKINVDCx5p33_ASAP7_75t_R g771 ( .A(n_227), .Y(n_771) );
INVx1_ASAP7_75t_L g906 ( .A(n_231), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g1619 ( .A1(n_232), .A2(n_235), .B1(n_613), .B2(n_1137), .Y(n_1619) );
INVx1_ASAP7_75t_L g1128 ( .A(n_233), .Y(n_1128) );
CKINVDCx5p33_ASAP7_75t_R g1296 ( .A(n_234), .Y(n_1296) );
INVx1_ASAP7_75t_L g1200 ( .A(n_236), .Y(n_1200) );
INVx1_ASAP7_75t_L g1222 ( .A(n_237), .Y(n_1222) );
INVx1_ASAP7_75t_L g1018 ( .A(n_239), .Y(n_1018) );
INVx1_ASAP7_75t_L g1273 ( .A(n_240), .Y(n_1273) );
INVx1_ASAP7_75t_L g984 ( .A(n_241), .Y(n_984) );
NAND2xp33_ASAP7_75t_SL g1071 ( .A(n_242), .B(n_830), .Y(n_1071) );
INVx1_ASAP7_75t_L g753 ( .A(n_245), .Y(n_753) );
XNOR2x2_ASAP7_75t_L g1194 ( .A(n_246), .B(n_1195), .Y(n_1194) );
INVx1_ASAP7_75t_L g1604 ( .A(n_247), .Y(n_1604) );
INVx1_ASAP7_75t_L g1350 ( .A(n_248), .Y(n_1350) );
INVx1_ASAP7_75t_L g405 ( .A(n_249), .Y(n_405) );
INVx1_ASAP7_75t_L g412 ( .A(n_249), .Y(n_412) );
INVx1_ASAP7_75t_L g616 ( .A(n_250), .Y(n_616) );
INVx1_ASAP7_75t_L g1096 ( .A(n_254), .Y(n_1096) );
INVx1_ASAP7_75t_L g1617 ( .A(n_258), .Y(n_1617) );
INVx1_ASAP7_75t_L g682 ( .A(n_259), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g1318 ( .A1(n_260), .A2(n_646), .B(n_1319), .Y(n_1318) );
CKINVDCx5p33_ASAP7_75t_R g890 ( .A(n_261), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g1115 ( .A(n_262), .Y(n_1115) );
INVx1_ASAP7_75t_L g970 ( .A(n_263), .Y(n_970) );
AND2x2_ASAP7_75t_L g1380 ( .A(n_264), .B(n_1381), .Y(n_1380) );
INVx1_ASAP7_75t_L g1387 ( .A(n_264), .Y(n_1387) );
INVxp67_ASAP7_75t_SL g1257 ( .A(n_265), .Y(n_1257) );
INVx1_ASAP7_75t_L g463 ( .A(n_266), .Y(n_463) );
OAI211xp5_ASAP7_75t_L g496 ( .A1(n_266), .A2(n_356), .B(n_497), .C(n_502), .Y(n_496) );
INVx1_ASAP7_75t_L g1362 ( .A(n_267), .Y(n_1362) );
XNOR2xp5_ASAP7_75t_L g754 ( .A(n_268), .B(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g350 ( .A(n_269), .Y(n_350) );
INVxp67_ASAP7_75t_SL g1050 ( .A(n_270), .Y(n_1050) );
INVxp67_ASAP7_75t_SL g1286 ( .A(n_271), .Y(n_1286) );
OAI211xp5_ASAP7_75t_L g1305 ( .A1(n_271), .A2(n_594), .B(n_1306), .C(n_1310), .Y(n_1305) );
INVx1_ASAP7_75t_L g1446 ( .A(n_272), .Y(n_1446) );
CKINVDCx16_ASAP7_75t_R g912 ( .A(n_273), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_277), .B(n_1230), .Y(n_1229) );
OAI21xp33_ASAP7_75t_L g840 ( .A1(n_278), .A2(n_585), .B(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g757 ( .A(n_279), .Y(n_757) );
OAI21xp5_ASAP7_75t_SL g1141 ( .A1(n_280), .A2(n_952), .B(n_1142), .Y(n_1141) );
INVx1_ASAP7_75t_L g777 ( .A(n_281), .Y(n_777) );
INVx1_ASAP7_75t_L g378 ( .A(n_283), .Y(n_378) );
INVx1_ASAP7_75t_L g354 ( .A(n_284), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g1193 ( .A(n_286), .Y(n_1193) );
INVxp67_ASAP7_75t_SL g1255 ( .A(n_287), .Y(n_1255) );
AOI22xp33_ASAP7_75t_SL g1265 ( .A1(n_287), .A2(n_294), .B1(n_557), .B2(n_1266), .Y(n_1265) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_288), .Y(n_333) );
INVx1_ASAP7_75t_L g1678 ( .A(n_289), .Y(n_1678) );
NOR2xp33_ASAP7_75t_R g928 ( .A(n_290), .B(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g886 ( .A(n_292), .Y(n_886) );
INVxp67_ASAP7_75t_SL g697 ( .A(n_296), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g733 ( .A1(n_296), .A2(n_298), .B1(n_734), .B2(n_736), .C(n_738), .Y(n_733) );
INVx1_ASAP7_75t_L g1682 ( .A(n_297), .Y(n_1682) );
OAI221xp5_ASAP7_75t_L g668 ( .A1(n_298), .A2(n_299), .B1(n_669), .B2(n_674), .C(n_675), .Y(n_668) );
INVx2_ASAP7_75t_L g362 ( .A(n_301), .Y(n_362) );
INVx1_ASAP7_75t_L g387 ( .A(n_301), .Y(n_387) );
INVx1_ASAP7_75t_L g435 ( .A(n_301), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g583 ( .A(n_302), .Y(n_583) );
INVx1_ASAP7_75t_L g791 ( .A(n_303), .Y(n_791) );
INVx1_ASAP7_75t_L g1599 ( .A(n_305), .Y(n_1599) );
CKINVDCx5p33_ASAP7_75t_R g1365 ( .A(n_306), .Y(n_1365) );
OAI22xp33_ASAP7_75t_SL g972 ( .A1(n_307), .A2(n_311), .B1(n_524), .B2(n_973), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g987 ( .A1(n_307), .A2(n_311), .B1(n_624), .B2(n_876), .C(n_988), .Y(n_987) );
INVx1_ASAP7_75t_L g1312 ( .A(n_308), .Y(n_1312) );
XNOR2xp5_ASAP7_75t_L g947 ( .A(n_309), .B(n_948), .Y(n_947) );
INVxp67_ASAP7_75t_SL g760 ( .A(n_310), .Y(n_760) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_338), .B(n_1370), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
BUFx4f_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
INVx3_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_323), .Y(n_316) );
NOR2xp33_ASAP7_75t_L g1639 ( .A(n_317), .B(n_326), .Y(n_1639) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
NOR2xp33_ASAP7_75t_L g1645 ( .A(n_319), .B(n_322), .Y(n_1645) );
INVx1_ASAP7_75t_L g1688 ( .A(n_319), .Y(n_1688) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NOR2xp33_ASAP7_75t_L g1690 ( .A(n_322), .B(n_1688), .Y(n_1690) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_325), .B(n_328), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
AND2x4_ASAP7_75t_L g513 ( .A(n_326), .B(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x4_ASAP7_75t_L g388 ( .A(n_327), .B(n_337), .Y(n_388) );
AND2x4_ASAP7_75t_L g647 ( .A(n_327), .B(n_336), .Y(n_647) );
INVx1_ASAP7_75t_L g480 ( .A(n_328), .Y(n_480) );
AND2x4_ASAP7_75t_SL g1638 ( .A(n_328), .B(n_1639), .Y(n_1638) );
INVx3_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x6_ASAP7_75t_L g329 ( .A(n_330), .B(n_335), .Y(n_329) );
OR2x6_ASAP7_75t_L g489 ( .A(n_330), .B(n_483), .Y(n_489) );
INVxp67_ASAP7_75t_L g1230 ( .A(n_330), .Y(n_1230) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx3_ASAP7_75t_L g368 ( .A(n_331), .Y(n_368) );
BUFx4f_ASAP7_75t_L g635 ( .A(n_331), .Y(n_635) );
INVx3_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
OR2x2_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g353 ( .A(n_333), .Y(n_353) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_333), .B(n_334), .Y(n_358) );
INVx2_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
AND2x2_ASAP7_75t_L g485 ( .A(n_333), .B(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g501 ( .A(n_333), .B(n_334), .Y(n_501) );
INVx1_ASAP7_75t_L g511 ( .A(n_333), .Y(n_511) );
OR2x2_ASAP7_75t_L g352 ( .A(n_334), .B(n_353), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_334), .B(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g486 ( .A(n_334), .Y(n_486) );
BUFx2_ASAP7_75t_L g505 ( .A(n_334), .Y(n_505) );
INVx1_ASAP7_75t_L g582 ( .A(n_334), .Y(n_582) );
AND2x2_ASAP7_75t_L g597 ( .A(n_334), .B(n_376), .Y(n_597) );
INVxp67_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g499 ( .A(n_336), .Y(n_499) );
INVx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx2_ASAP7_75t_L g495 ( .A(n_337), .Y(n_495) );
AND2x4_ASAP7_75t_L g509 ( .A(n_337), .B(n_510), .Y(n_509) );
OAI22xp5_ASAP7_75t_L g338 ( .A1(n_339), .A2(n_340), .B1(n_998), .B2(n_1369), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B1(n_806), .B2(n_997), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_344), .B1(n_650), .B2(n_805), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OA22x2_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_516), .B1(n_517), .B2(n_649), .Y(n_344) );
INVx1_ASAP7_75t_L g649 ( .A(n_345), .Y(n_649) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_441), .C(n_478), .Y(n_346) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_348), .B(n_392), .Y(n_347) );
OAI33xp33_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_359), .A3(n_364), .B1(n_377), .B2(n_380), .B3(n_389), .Y(n_348) );
OAI22xp5_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_351), .B1(n_354), .B2(n_355), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_350), .A2(n_378), .B1(n_415), .B2(n_420), .Y(n_414) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_351), .A2(n_370), .B1(n_390), .B2(n_391), .Y(n_389) );
BUFx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g663 ( .A(n_352), .Y(n_663) );
BUFx2_ASAP7_75t_L g868 ( .A(n_352), .Y(n_868) );
INVx1_ASAP7_75t_L g933 ( .A(n_352), .Y(n_933) );
AND2x2_ASAP7_75t_L g581 ( .A(n_353), .B(n_582), .Y(n_581) );
HB1xp67_ASAP7_75t_L g1610 ( .A(n_353), .Y(n_1610) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_354), .A2(n_379), .B1(n_425), .B2(n_427), .Y(n_424) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp33_ASAP7_75t_L g377 ( .A1(n_356), .A2(n_366), .B1(n_378), .B2(n_379), .Y(n_377) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx4f_ASAP7_75t_L g665 ( .A(n_357), .Y(n_665) );
OR2x6_ASAP7_75t_L g675 ( .A(n_357), .B(n_676), .Y(n_675) );
INVx4_ASAP7_75t_L g990 ( .A(n_357), .Y(n_990) );
BUFx6f_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
BUFx3_ASAP7_75t_L g696 ( .A(n_358), .Y(n_696) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g680 ( .A1(n_360), .A2(n_663), .B1(n_665), .B2(n_681), .C(n_682), .Y(n_680) );
HB1xp67_ASAP7_75t_L g793 ( .A(n_360), .Y(n_793) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_360), .B(n_920), .Y(n_919) );
AND2x4_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .Y(n_360) );
INVx1_ASAP7_75t_L g879 ( .A(n_361), .Y(n_879) );
OR2x2_ASAP7_75t_L g1120 ( .A(n_361), .B(n_711), .Y(n_1120) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g539 ( .A(n_362), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_362), .B(n_580), .Y(n_671) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_366), .B1(n_369), .B2(n_370), .Y(n_364) );
OAI22xp33_ASAP7_75t_L g399 ( .A1(n_365), .A2(n_390), .B1(n_400), .B2(n_406), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g1254 ( .A1(n_366), .A2(n_1255), .B1(n_1256), .B2(n_1257), .C(n_1258), .Y(n_1254) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
BUFx6f_ASAP7_75t_L g660 ( .A(n_368), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g789 ( .A1(n_368), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_789) );
OAI22x1_ASAP7_75t_SL g795 ( .A1(n_368), .A2(n_771), .B1(n_792), .B2(n_796), .Y(n_795) );
BUFx3_ASAP7_75t_L g1095 ( .A(n_368), .Y(n_1095) );
OAI22xp5_ASAP7_75t_L g437 ( .A1(n_369), .A2(n_391), .B1(n_438), .B2(n_440), .Y(n_437) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx4_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g638 ( .A(n_373), .Y(n_638) );
INVx2_ASAP7_75t_L g792 ( .A(n_373), .Y(n_792) );
BUFx6f_ASAP7_75t_L g874 ( .A(n_373), .Y(n_874) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_373), .Y(n_1020) );
INVx1_ASAP7_75t_L g1098 ( .A(n_373), .Y(n_1098) );
INVx8_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OR2x2_ASAP7_75t_L g494 ( .A(n_374), .B(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g679 ( .A(n_374), .Y(n_679) );
BUFx6f_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_388), .Y(n_382) );
AND2x4_ASAP7_75t_L g797 ( .A(n_383), .B(n_388), .Y(n_797) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OR2x2_ASAP7_75t_L g395 ( .A(n_385), .B(n_396), .Y(n_395) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_385), .Y(n_477) );
OR2x2_ASAP7_75t_L g564 ( .A(n_385), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_SL g667 ( .A(n_385), .B(n_388), .Y(n_667) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
BUFx2_ASAP7_75t_L g515 ( .A(n_386), .Y(n_515) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx4_ASAP7_75t_L g608 ( .A(n_388), .Y(n_608) );
INVx1_ASAP7_75t_SL g856 ( .A(n_388), .Y(n_856) );
INVx4_ASAP7_75t_L g1087 ( .A(n_388), .Y(n_1087) );
OAI33xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_399), .A3(n_414), .B1(n_424), .B2(n_429), .B3(n_437), .Y(n_392) );
BUFx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
OAI22xp5_ASAP7_75t_SL g955 ( .A1(n_394), .A2(n_956), .B1(n_964), .B2(n_966), .Y(n_955) );
BUFx4f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx2_ASAP7_75t_L g1043 ( .A(n_395), .Y(n_1043) );
BUFx4f_ASAP7_75t_L g1066 ( .A(n_395), .Y(n_1066) );
BUFx8_ASAP7_75t_L g1335 ( .A(n_395), .Y(n_1335) );
BUFx2_ASAP7_75t_L g718 ( .A(n_396), .Y(n_718) );
NAND2xp33_ASAP7_75t_SL g396 ( .A(n_397), .B(n_398), .Y(n_396) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_397), .Y(n_475) );
INVx1_ASAP7_75t_L g530 ( .A(n_397), .Y(n_530) );
AND3x4_ASAP7_75t_L g538 ( .A(n_397), .B(n_461), .C(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g902 ( .A(n_397), .B(n_461), .Y(n_902) );
INVx3_ASAP7_75t_L g433 ( .A(n_398), .Y(n_433) );
BUFx3_ASAP7_75t_L g461 ( .A(n_398), .Y(n_461) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g439 ( .A(n_401), .Y(n_439) );
OAI22xp5_ASAP7_75t_L g895 ( .A1(n_401), .A2(n_896), .B1(n_897), .B2(n_898), .Y(n_895) );
OAI22xp5_ASAP7_75t_L g1633 ( .A1(n_401), .A2(n_1634), .B1(n_1635), .B2(n_1636), .Y(n_1633) );
BUFx4f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OR2x4_ASAP7_75t_L g445 ( .A(n_402), .B(n_446), .Y(n_445) );
OR2x4_ASAP7_75t_L g470 ( .A(n_402), .B(n_433), .Y(n_470) );
INVx2_ASAP7_75t_L g561 ( .A(n_402), .Y(n_561) );
OR2x2_ASAP7_75t_L g402 ( .A(n_403), .B(n_404), .Y(n_402) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_403), .Y(n_413) );
INVx2_ASAP7_75t_L g419 ( .A(n_403), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_403), .B(n_412), .Y(n_423) );
AND2x4_ASAP7_75t_L g454 ( .A(n_403), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g544 ( .A(n_404), .Y(n_544) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVxp67_ASAP7_75t_L g418 ( .A(n_405), .Y(n_418) );
INVx2_ASAP7_75t_SL g406 ( .A(n_407), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OR2x2_ASAP7_75t_L g588 ( .A(n_409), .B(n_564), .Y(n_588) );
INVx3_ASAP7_75t_L g781 ( .A(n_409), .Y(n_781) );
INVx4_ASAP7_75t_L g1630 ( .A(n_409), .Y(n_1630) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
BUFx3_ASAP7_75t_L g428 ( .A(n_410), .Y(n_428) );
BUFx2_ASAP7_75t_L g739 ( .A(n_410), .Y(n_739) );
NAND2x1p5_ASAP7_75t_L g410 ( .A(n_411), .B(n_413), .Y(n_410) );
BUFx2_ASAP7_75t_L g466 ( .A(n_411), .Y(n_466) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g455 ( .A(n_412), .Y(n_455) );
BUFx2_ASAP7_75t_L g462 ( .A(n_413), .Y(n_462) );
INVx2_ASAP7_75t_L g526 ( .A(n_413), .Y(n_526) );
AND2x4_ASAP7_75t_L g551 ( .A(n_413), .B(n_536), .Y(n_551) );
INVx1_ASAP7_75t_L g1268 ( .A(n_415), .Y(n_1268) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_416), .Y(n_426) );
AND2x4_ASAP7_75t_L g472 ( .A(n_416), .B(n_446), .Y(n_472) );
BUFx6f_ASAP7_75t_L g829 ( .A(n_416), .Y(n_829) );
INVx2_ASAP7_75t_L g967 ( .A(n_416), .Y(n_967) );
INVx2_ASAP7_75t_L g1042 ( .A(n_416), .Y(n_1042) );
BUFx6f_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
BUFx8_ASAP7_75t_L g549 ( .A(n_417), .Y(n_549) );
INVx2_ASAP7_75t_L g708 ( .A(n_417), .Y(n_708) );
BUFx6f_ASAP7_75t_L g717 ( .A(n_417), .Y(n_717) );
AND2x4_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
AND2x4_ASAP7_75t_L g543 ( .A(n_419), .B(n_544), .Y(n_543) );
OAI22xp5_ASAP7_75t_L g903 ( .A1(n_420), .A2(n_904), .B1(n_905), .B2(n_906), .Y(n_903) );
OAI22xp33_ASAP7_75t_L g1336 ( .A1(n_420), .A2(n_1046), .B1(n_1337), .B2(n_1338), .Y(n_1336) );
OAI22xp5_ASAP7_75t_L g1344 ( .A1(n_420), .A2(n_1345), .B1(n_1346), .B2(n_1347), .Y(n_1344) );
INVx3_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx3_ASAP7_75t_L g440 ( .A(n_421), .Y(n_440) );
INVx3_ASAP7_75t_L g897 ( .A(n_421), .Y(n_897) );
CKINVDCx8_ASAP7_75t_R g969 ( .A(n_421), .Y(n_969) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g577 ( .A(n_422), .Y(n_577) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g450 ( .A(n_423), .Y(n_450) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
OAI33xp33_ASAP7_75t_L g1334 ( .A1(n_429), .A2(n_1335), .A3(n_1336), .B1(n_1339), .B2(n_1344), .B3(n_1348), .Y(n_1334) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g1159 ( .A(n_430), .B(n_1160), .C(n_1161), .Y(n_1159) );
AOI33xp33_ASAP7_75t_L g1264 ( .A1(n_430), .A2(n_538), .A3(n_1265), .B1(n_1267), .B2(n_1269), .B3(n_1270), .Y(n_1264) );
BUFx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g553 ( .A(n_431), .Y(n_553) );
BUFx2_ASAP7_75t_L g834 ( .A(n_431), .Y(n_834) );
BUFx2_ASAP7_75t_L g1294 ( .A(n_431), .Y(n_1294) );
INVx3_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx3_ASAP7_75t_L g965 ( .A(n_432), .Y(n_965) );
NAND3x1_ASAP7_75t_L g432 ( .A(n_433), .B(n_434), .C(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g446 ( .A(n_433), .Y(n_446) );
OR2x6_ASAP7_75t_L g449 ( .A(n_433), .B(n_450), .Y(n_449) );
AND2x4_ASAP7_75t_L g453 ( .A(n_433), .B(n_454), .Y(n_453) );
AND2x4_ASAP7_75t_L g529 ( .A(n_433), .B(n_530), .Y(n_529) );
NAND2x1p5_ASAP7_75t_L g711 ( .A(n_433), .B(n_436), .Y(n_711) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g528 ( .A(n_435), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_435), .B(n_598), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g1044 ( .A1(n_438), .A2(n_1028), .B1(n_1045), .B2(n_1046), .Y(n_1044) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
OAI22xp5_ASAP7_75t_L g1040 ( .A1(n_440), .A2(n_1018), .B1(n_1041), .B2(n_1042), .Y(n_1040) );
OAI31xp33_ASAP7_75t_L g441 ( .A1(n_442), .A2(n_451), .A3(n_467), .B(n_473), .Y(n_441) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g960 ( .A(n_450), .Y(n_960) );
BUFx3_ASAP7_75t_L g1051 ( .A(n_450), .Y(n_1051) );
CKINVDCx8_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
BUFx3_ASAP7_75t_L g545 ( .A(n_454), .Y(n_545) );
BUFx2_ASAP7_75t_L g572 ( .A(n_454), .Y(n_572) );
INVx2_ASAP7_75t_L g714 ( .A(n_454), .Y(n_714) );
AND2x2_ASAP7_75t_L g728 ( .A(n_454), .B(n_726), .Y(n_728) );
BUFx2_ASAP7_75t_L g839 ( .A(n_454), .Y(n_839) );
BUFx2_ASAP7_75t_L g963 ( .A(n_454), .Y(n_963) );
BUFx2_ASAP7_75t_L g1266 ( .A(n_454), .Y(n_1266) );
INVx1_ASAP7_75t_L g536 ( .A(n_455), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B1(n_463), .B2(n_464), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_457), .A2(n_503), .B1(n_506), .B2(n_507), .Y(n_502) );
BUFx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_462), .Y(n_459) );
AND2x4_ASAP7_75t_L g465 ( .A(n_460), .B(n_466), .Y(n_465) );
INVx3_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
BUFx6f_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_SL g473 ( .A(n_474), .B(n_476), .Y(n_473) );
INVx1_ASAP7_75t_SL g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OAI31xp33_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_487), .A3(n_496), .B(n_512), .Y(n_478) );
INVx3_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g606 ( .A(n_485), .Y(n_606) );
INVx2_ASAP7_75t_L g645 ( .A(n_485), .Y(n_645) );
BUFx3_ASAP7_75t_L g788 ( .A(n_485), .Y(n_788) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x4_ASAP7_75t_L g504 ( .A(n_495), .B(n_505), .Y(n_504) );
INVx3_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_500), .Y(n_498) );
BUFx6f_ASAP7_75t_L g602 ( .A(n_500), .Y(n_602) );
AND2x6_ASAP7_75t_L g614 ( .A(n_500), .B(n_580), .Y(n_614) );
AND2x4_ASAP7_75t_SL g627 ( .A(n_500), .B(n_598), .Y(n_627) );
BUFx3_ASAP7_75t_L g641 ( .A(n_500), .Y(n_641) );
BUFx3_ASAP7_75t_L g787 ( .A(n_500), .Y(n_787) );
BUFx3_ASAP7_75t_L g1023 ( .A(n_500), .Y(n_1023) );
INVx1_ASAP7_75t_L g1186 ( .A(n_500), .Y(n_1186) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g853 ( .A(n_501), .Y(n_853) );
BUFx3_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g630 ( .A(n_505), .Y(n_630) );
INVx1_ASAP7_75t_L g673 ( .A(n_505), .Y(n_673) );
BUFx2_ASAP7_75t_L g1140 ( .A(n_505), .Y(n_1140) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_510), .B(n_580), .Y(n_587) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx3_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
OR2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_587), .Y(n_586) );
INVxp67_ASAP7_75t_L g591 ( .A(n_515), .Y(n_591) );
OR2x2_ASAP7_75t_L g674 ( .A(n_515), .B(n_587), .Y(n_674) );
INVx1_ASAP7_75t_L g703 ( .A(n_515), .Y(n_703) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_519), .B(n_573), .C(n_592), .Y(n_518) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_558), .C(n_569), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_521), .B(n_537), .Y(n_520) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_522), .A2(n_523), .B1(n_531), .B2(n_532), .Y(n_521) );
AOI22xp5_ASAP7_75t_L g1282 ( .A1(n_523), .A2(n_532), .B1(n_1283), .B2(n_1284), .Y(n_1282) );
AOI221xp5_ASAP7_75t_L g1597 ( .A1(n_523), .A2(n_532), .B1(n_1598), .B2(n_1599), .C(n_1600), .Y(n_1597) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
NAND2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
AND2x6_ASAP7_75t_L g735 ( .A(n_525), .B(n_529), .Y(n_735) );
AND2x2_ASAP7_75t_L g815 ( .A(n_525), .B(n_527), .Y(n_815) );
AND2x2_ASAP7_75t_L g1081 ( .A(n_525), .B(n_527), .Y(n_1081) );
AND2x4_ASAP7_75t_SL g1116 ( .A(n_525), .B(n_527), .Y(n_1116) );
INVx3_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x4_ASAP7_75t_L g532 ( .A(n_527), .B(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g571 ( .A(n_527), .B(n_572), .Y(n_571) );
AND2x4_ASAP7_75t_SL g974 ( .A(n_527), .B(n_533), .Y(n_974) );
AND2x4_ASAP7_75t_L g527 ( .A(n_528), .B(n_529), .Y(n_527) );
OR2x2_ASAP7_75t_L g578 ( .A(n_528), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g685 ( .A(n_528), .Y(n_685) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_529), .B(n_543), .Y(n_590) );
AND2x2_ASAP7_75t_L g737 ( .A(n_529), .B(n_535), .Y(n_737) );
INVx1_ASAP7_75t_L g740 ( .A(n_529), .Y(n_740) );
AO22x1_ASAP7_75t_L g813 ( .A1(n_532), .A2(n_814), .B1(n_815), .B2(n_816), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_532), .A2(n_815), .B1(n_1006), .B2(n_1007), .Y(n_1005) );
AOI22xp33_ASAP7_75t_L g1165 ( .A1(n_532), .A2(n_815), .B1(n_1166), .B2(n_1167), .Y(n_1165) );
AOI22xp33_ASAP7_75t_L g1198 ( .A1(n_532), .A2(n_815), .B1(n_1199), .B2(n_1200), .Y(n_1198) );
AOI22xp33_ASAP7_75t_L g1272 ( .A1(n_532), .A2(n_1081), .B1(n_1273), .B2(n_1274), .Y(n_1272) );
HB1xp67_ASAP7_75t_L g1332 ( .A(n_532), .Y(n_1332) );
INVx2_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AOI33xp33_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_540), .A3(n_546), .B1(n_552), .B2(n_553), .B3(n_554), .Y(n_537) );
BUFx3_ASAP7_75t_L g824 ( .A(n_538), .Y(n_824) );
INVx1_ASAP7_75t_L g1123 ( .A(n_538), .Y(n_1123) );
AOI33xp33_ASAP7_75t_L g1287 ( .A1(n_538), .A2(n_1288), .A3(n_1289), .B1(n_1292), .B2(n_1293), .B3(n_1294), .Y(n_1287) );
INVx2_ASAP7_75t_SL g648 ( .A(n_539), .Y(n_648) );
INVx1_ASAP7_75t_L g748 ( .A(n_539), .Y(n_748) );
OAI31xp33_ASAP7_75t_SL g761 ( .A1(n_539), .A2(n_762), .A3(n_763), .B(n_767), .Y(n_761) );
OAI31xp33_ASAP7_75t_L g892 ( .A1(n_539), .A2(n_893), .A3(n_894), .B(n_910), .Y(n_892) );
INVx8_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
CKINVDCx5p33_ASAP7_75t_R g773 ( .A(n_542), .Y(n_773) );
INVx3_ASAP7_75t_L g836 ( .A(n_542), .Y(n_836) );
INVx2_ASAP7_75t_L g844 ( .A(n_542), .Y(n_844) );
INVx2_ASAP7_75t_L g1053 ( .A(n_542), .Y(n_1053) );
INVx8_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
BUFx3_ASAP7_75t_L g557 ( .A(n_543), .Y(n_557) );
BUFx3_ASAP7_75t_L g721 ( .A(n_543), .Y(n_721) );
AND2x2_ASAP7_75t_L g725 ( .A(n_543), .B(n_726), .Y(n_725) );
HB1xp67_ASAP7_75t_L g1070 ( .A(n_543), .Y(n_1070) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
INVx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g567 ( .A(n_549), .B(n_568), .Y(n_567) );
HB1xp67_ASAP7_75t_L g1154 ( .A(n_549), .Y(n_1154) );
INVx2_ASAP7_75t_SL g1345 ( .A(n_549), .Y(n_1345) );
INVx2_ASAP7_75t_SL g1672 ( .A(n_549), .Y(n_1672) );
BUFx3_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
BUFx2_ASAP7_75t_L g709 ( .A(n_551), .Y(n_709) );
BUFx12f_ASAP7_75t_L g722 ( .A(n_551), .Y(n_722) );
AND2x4_ASAP7_75t_L g746 ( .A(n_551), .B(n_744), .Y(n_746) );
INVx5_ASAP7_75t_L g831 ( .A(n_551), .Y(n_831) );
BUFx3_ASAP7_75t_L g1155 ( .A(n_551), .Y(n_1155) );
AOI33xp33_ASAP7_75t_L g1201 ( .A1(n_553), .A2(n_824), .A3(n_1202), .B1(n_1203), .B2(n_1206), .B3(n_1208), .Y(n_1201) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx2_ASAP7_75t_SL g827 ( .A(n_557), .Y(n_827) );
NAND2xp5_ASAP7_75t_L g1591 ( .A(n_559), .B(n_701), .Y(n_1591) );
OR2x6_ASAP7_75t_L g559 ( .A(n_560), .B(n_562), .Y(n_559) );
OR2x2_ASAP7_75t_L g1303 ( .A(n_560), .B(n_562), .Y(n_1303) );
INVx2_ASAP7_75t_SL g1341 ( .A(n_560), .Y(n_1341) );
INVx2_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
INVx3_ASAP7_75t_L g1628 ( .A(n_561), .Y(n_1628) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
AND2x2_ASAP7_75t_L g1144 ( .A(n_563), .B(n_1075), .Y(n_1144) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g568 ( .A(n_564), .Y(n_568) );
OR2x2_ASAP7_75t_L g576 ( .A(n_564), .B(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g726 ( .A(n_565), .Y(n_726) );
INVx1_ASAP7_75t_L g744 ( .A(n_565), .Y(n_744) );
INVxp67_ASAP7_75t_L g1107 ( .A(n_566), .Y(n_1107) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_567), .A2(n_842), .B1(n_843), .B2(n_845), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g994 ( .A1(n_567), .A2(n_843), .B1(n_984), .B2(n_986), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_567), .A2(n_843), .B1(n_1171), .B2(n_1172), .Y(n_1191) );
INVx2_ASAP7_75t_L g1263 ( .A(n_567), .Y(n_1263) );
AOI22xp33_ASAP7_75t_L g1684 ( .A1(n_567), .A2(n_843), .B1(n_1658), .B2(n_1659), .Y(n_1684) );
AND2x4_ASAP7_75t_L g843 ( .A(n_568), .B(n_844), .Y(n_843) );
AND2x4_ASAP7_75t_L g1143 ( .A(n_568), .B(n_844), .Y(n_1143) );
NOR4xp25_ASAP7_75t_L g1329 ( .A(n_569), .B(n_1330), .C(n_1333), .D(n_1334), .Y(n_1329) );
INVx2_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
NAND5xp2_ASAP7_75t_L g1004 ( .A(n_570), .B(n_1005), .C(n_1008), .D(n_1011), .E(n_1012), .Y(n_1004) );
NAND3xp33_ASAP7_75t_SL g1113 ( .A(n_570), .B(n_1114), .C(n_1118), .Y(n_1113) );
AND4x1_ASAP7_75t_L g1260 ( .A(n_570), .B(n_1261), .C(n_1264), .D(n_1272), .Y(n_1260) );
INVx3_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
INVx3_ASAP7_75t_L g822 ( .A(n_571), .Y(n_822) );
HB1xp67_ASAP7_75t_L g954 ( .A(n_571), .Y(n_954) );
NOR3xp33_ASAP7_75t_SL g1064 ( .A(n_571), .B(n_1065), .C(n_1079), .Y(n_1064) );
AOI221xp5_ASAP7_75t_L g1623 ( .A1(n_571), .A2(n_824), .B1(n_965), .B2(n_1624), .C(n_1631), .Y(n_1623) );
NOR3xp33_ASAP7_75t_L g1669 ( .A(n_571), .B(n_1670), .C(n_1680), .Y(n_1669) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_572), .Y(n_1158) );
AOI21xp33_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_583), .B(n_584), .Y(n_573) );
AOI211x1_ASAP7_75t_L g809 ( .A1(n_574), .A2(n_810), .B(n_811), .C(n_840), .Y(n_809) );
AOI21xp5_ASAP7_75t_L g949 ( .A1(n_574), .A2(n_950), .B(n_951), .Y(n_949) );
AOI221xp5_ASAP7_75t_L g1110 ( .A1(n_574), .A2(n_1010), .B1(n_1111), .B2(n_1112), .C(n_1113), .Y(n_1110) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_574), .B(n_1193), .Y(n_1192) );
AOI21xp5_ASAP7_75t_L g1210 ( .A1(n_574), .A2(n_1211), .B(n_1212), .Y(n_1210) );
AOI21xp33_ASAP7_75t_L g1240 ( .A1(n_574), .A2(n_1241), .B(n_1242), .Y(n_1240) );
NAND2xp33_ASAP7_75t_L g1295 ( .A(n_574), .B(n_1296), .Y(n_1295) );
AOI21xp33_ASAP7_75t_L g1364 ( .A1(n_574), .A2(n_1365), .B(n_1366), .Y(n_1364) );
AOI21xp5_ASAP7_75t_L g1681 ( .A1(n_574), .A2(n_1682), .B(n_1683), .Y(n_1681) );
INVx8_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_578), .Y(n_575) );
BUFx3_ASAP7_75t_L g770 ( .A(n_577), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_578), .B(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g686 ( .A(n_579), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_580), .B(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g631 ( .A(n_580), .Y(n_631) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_580), .B(n_1140), .Y(n_1139) );
HB1xp67_ASAP7_75t_L g1611 ( .A(n_580), .Y(n_1611) );
INVx3_ASAP7_75t_L g611 ( .A(n_581), .Y(n_611) );
AND2x2_ASAP7_75t_L g619 ( .A(n_581), .B(n_598), .Y(n_619) );
BUFx6f_ASAP7_75t_L g982 ( .A(n_581), .Y(n_982) );
INVx2_ASAP7_75t_L g1037 ( .A(n_585), .Y(n_1037) );
HB1xp67_ASAP7_75t_L g1367 ( .A(n_585), .Y(n_1367) );
AND2x4_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
INVx2_ASAP7_75t_SL g801 ( .A(n_586), .Y(n_801) );
AND2x4_ASAP7_75t_L g952 ( .A(n_586), .B(n_588), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g939 ( .A(n_589), .B(n_940), .Y(n_939) );
OR2x2_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx2_ASAP7_75t_L g732 ( .A(n_590), .Y(n_732) );
OR2x6_ASAP7_75t_L g821 ( .A(n_590), .B(n_591), .Y(n_821) );
OAI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_623), .B(n_648), .Y(n_592) );
INVx2_ASAP7_75t_SL g594 ( .A(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_R g861 ( .A(n_595), .B(n_819), .Y(n_861) );
INVx3_ASAP7_75t_L g1034 ( .A(n_595), .Y(n_1034) );
AOI221xp5_ASAP7_75t_SL g1173 ( .A1(n_595), .A2(n_614), .B1(n_1164), .B2(n_1174), .C(n_1177), .Y(n_1173) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_596), .Y(n_1178) );
BUFx6f_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
BUFx3_ASAP7_75t_L g613 ( .A(n_597), .Y(n_613) );
INVx2_ASAP7_75t_L g692 ( .A(n_597), .Y(n_692) );
BUFx3_ASAP7_75t_L g935 ( .A(n_597), .Y(n_935) );
AND2x4_ASAP7_75t_L g622 ( .A(n_598), .B(n_606), .Y(n_622) );
AND2x2_ASAP7_75t_L g752 ( .A(n_598), .B(n_606), .Y(n_752) );
AND2x2_ASAP7_75t_L g1085 ( .A(n_598), .B(n_691), .Y(n_1085) );
AOI21xp5_ASAP7_75t_SL g599 ( .A1(n_600), .A2(n_609), .B(n_614), .Y(n_599) );
BUFx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
HB1xp67_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g1218 ( .A(n_604), .Y(n_1218) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g1182 ( .A(n_605), .Y(n_1182) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
BUFx6f_ASAP7_75t_L g855 ( .A(n_606), .Y(n_855) );
INVx1_ASAP7_75t_L g1655 ( .A(n_606), .Y(n_1655) );
HB1xp67_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_SL g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g858 ( .A(n_611), .Y(n_858) );
INVx2_ASAP7_75t_L g923 ( .A(n_611), .Y(n_923) );
INVx2_ASAP7_75t_L g1133 ( .A(n_611), .Y(n_1133) );
INVx1_ASAP7_75t_L g1137 ( .A(n_611), .Y(n_1137) );
INVx1_ASAP7_75t_L g1359 ( .A(n_611), .Y(n_1359) );
BUFx3_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_SL g860 ( .A(n_613), .Y(n_860) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_614), .A2(n_850), .B(n_857), .Y(n_849) );
AOI21xp5_ASAP7_75t_L g977 ( .A1(n_614), .A2(n_978), .B(n_979), .Y(n_977) );
INVx1_ASAP7_75t_L g1024 ( .A(n_614), .Y(n_1024) );
AOI221xp5_ASAP7_75t_L g1084 ( .A1(n_614), .A2(n_1063), .B1(n_1085), .B2(n_1086), .C(n_1088), .Y(n_1084) );
AOI221xp5_ASAP7_75t_L g1130 ( .A1(n_614), .A2(n_1085), .B1(n_1111), .B2(n_1131), .C(n_1132), .Y(n_1130) );
AOI21xp5_ASAP7_75t_L g1215 ( .A1(n_614), .A2(n_1216), .B(n_1219), .Y(n_1215) );
AOI21xp5_ASAP7_75t_L g1248 ( .A1(n_614), .A2(n_1249), .B(n_1252), .Y(n_1248) );
AOI21xp5_ASAP7_75t_L g1306 ( .A1(n_614), .A2(n_1307), .B(n_1308), .Y(n_1306) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_614), .A2(n_1357), .B(n_1358), .Y(n_1356) );
AOI21xp5_ASAP7_75t_L g1652 ( .A1(n_614), .A2(n_1653), .B(n_1656), .Y(n_1652) );
AOI22xp33_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B1(n_620), .B2(n_621), .Y(n_615) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_617), .A2(n_622), .B1(n_842), .B2(n_845), .Y(n_848) );
AOI22xp33_ASAP7_75t_L g1220 ( .A1(n_617), .A2(n_1221), .B1(n_1222), .B2(n_1223), .Y(n_1220) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_617), .A2(n_1361), .B1(n_1362), .B2(n_1363), .Y(n_1360) );
INVx2_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_619), .Y(n_618) );
AND2x4_ASAP7_75t_L g702 ( .A(n_619), .B(n_703), .Y(n_702) );
BUFx6f_ASAP7_75t_L g985 ( .A(n_619), .Y(n_985) );
AOI22xp33_ASAP7_75t_L g1657 ( .A1(n_619), .A2(n_622), .B1(n_1658), .B2(n_1659), .Y(n_1657) );
INVxp67_ASAP7_75t_SL g1026 ( .A(n_621), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g1245 ( .A1(n_621), .A2(n_985), .B1(n_1246), .B2(n_1247), .Y(n_1245) );
BUFx6f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_622), .A2(n_984), .B1(n_985), .B2(n_986), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g1090 ( .A1(n_622), .A2(n_985), .B1(n_1091), .B2(n_1092), .Y(n_1090) );
AOI22xp5_ASAP7_75t_L g1127 ( .A1(n_622), .A2(n_985), .B1(n_1128), .B2(n_1129), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g1170 ( .A1(n_622), .A2(n_985), .B1(n_1171), .B2(n_1172), .Y(n_1170) );
INVx1_ASAP7_75t_L g1224 ( .A(n_622), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1310 ( .A1(n_622), .A2(n_985), .B1(n_1311), .B2(n_1312), .Y(n_1310) );
HB1xp67_ASAP7_75t_L g1363 ( .A(n_622), .Y(n_1363) );
INVx2_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
INVx1_ASAP7_75t_L g863 ( .A(n_625), .Y(n_863) );
AOI22xp33_ASAP7_75t_L g1231 ( .A1(n_625), .A2(n_629), .B1(n_1199), .B2(n_1200), .Y(n_1231) );
INVx2_ASAP7_75t_L g1314 ( .A(n_625), .Y(n_1314) );
INVx4_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
BUFx3_ASAP7_75t_L g1135 ( .A(n_627), .Y(n_1135) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g876 ( .A(n_629), .Y(n_876) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
OAI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_636), .B1(n_637), .B2(n_639), .C(n_640), .Y(n_632) );
OAI22xp5_ASAP7_75t_L g870 ( .A1(n_633), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_870) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx6f_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g658 ( .A(n_637), .Y(n_658) );
BUFx2_ASAP7_75t_L g1256 ( .A(n_637), .Y(n_1256) );
BUFx6f_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g1175 ( .A(n_643), .Y(n_1175) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
HB1xp67_ASAP7_75t_L g1228 ( .A(n_644), .Y(n_1228) );
INVx1_ASAP7_75t_L g1251 ( .A(n_644), .Y(n_1251) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx2_ASAP7_75t_L g921 ( .A(n_645), .Y(n_921) );
INVx2_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OAI221xp5_ASAP7_75t_L g864 ( .A1(n_647), .A2(n_665), .B1(n_865), .B2(n_866), .C(n_869), .Y(n_864) );
INVx3_ASAP7_75t_L g1031 ( .A(n_647), .Y(n_1031) );
INVx2_ASAP7_75t_L g1104 ( .A(n_647), .Y(n_1104) );
INVx1_ASAP7_75t_L g1666 ( .A(n_647), .Y(n_1666) );
AOI21xp5_ASAP7_75t_SL g1168 ( .A1(n_648), .A2(n_1169), .B(n_1190), .Y(n_1168) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
BUFx2_ASAP7_75t_SL g805 ( .A(n_651), .Y(n_805) );
INVxp67_ASAP7_75t_SL g651 ( .A(n_652), .Y(n_651) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_653), .B(n_754), .Y(n_652) );
XNOR2x1_ASAP7_75t_L g653 ( .A(n_654), .B(n_753), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_704), .Y(n_654) );
NAND3xp33_ASAP7_75t_SL g655 ( .A(n_656), .B(n_683), .C(n_698), .Y(n_655) );
AOI211xp5_ASAP7_75t_SL g656 ( .A1(n_657), .A2(n_661), .B(n_668), .C(n_677), .Y(n_656) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g1017 ( .A1(n_660), .A2(n_1018), .B1(n_1019), .B2(n_1021), .C(n_1022), .Y(n_1017) );
OAI221xp5_ASAP7_75t_L g1027 ( .A1(n_660), .A2(n_679), .B1(n_1028), .B2(n_1029), .C(n_1030), .Y(n_1027) );
OAI221xp5_ASAP7_75t_SL g1353 ( .A1(n_660), .A2(n_1256), .B1(n_1342), .B2(n_1349), .C(n_1354), .Y(n_1353) );
INVx2_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
OAI21xp5_ASAP7_75t_L g930 ( .A1(n_666), .A2(n_675), .B(n_931), .Y(n_930) );
INVx2_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g800 ( .A(n_669), .Y(n_800) );
INVx2_ASAP7_75t_SL g927 ( .A(n_669), .Y(n_927) );
NAND2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_672), .Y(n_669) );
INVx1_ASAP7_75t_L g676 ( .A(n_670), .Y(n_676) );
INVx2_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx2_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_SL g925 ( .A(n_674), .Y(n_925) );
CKINVDCx5p33_ASAP7_75t_R g804 ( .A(n_675), .Y(n_804) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
AOI222xp33_ASAP7_75t_L g683 ( .A1(n_684), .A2(n_687), .B1(n_688), .B2(n_693), .C1(n_694), .C2(n_697), .Y(n_683) );
AOI21xp33_ASAP7_75t_SL g802 ( .A1(n_684), .A2(n_803), .B(n_804), .Y(n_802) );
AND2x4_ASAP7_75t_L g684 ( .A(n_685), .B(n_686), .Y(n_684) );
AOI222xp33_ASAP7_75t_L g798 ( .A1(n_688), .A2(n_765), .B1(n_777), .B2(n_799), .C1(n_800), .C2(n_801), .Y(n_798) );
INVx1_ASAP7_75t_L g940 ( .A(n_688), .Y(n_940) );
AND2x4_ASAP7_75t_L g688 ( .A(n_689), .B(n_691), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g695 ( .A(n_690), .B(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g929 ( .A(n_690), .B(n_696), .Y(n_929) );
INVx3_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g993 ( .A(n_692), .Y(n_993) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_693), .A2(n_730), .B(n_733), .C(n_741), .Y(n_729) );
AOI222xp33_ASAP7_75t_L g785 ( .A1(n_694), .A2(n_766), .B1(n_786), .B2(n_793), .C1(n_794), .C2(n_797), .Y(n_785) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx2_ASAP7_75t_SL g1664 ( .A(n_696), .Y(n_1664) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx3_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_702), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_702), .A2(n_751), .B1(n_890), .B2(n_891), .Y(n_889) );
AND2x4_ASAP7_75t_L g751 ( .A(n_703), .B(n_752), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_729), .B(n_747), .C(n_749), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_706), .A2(n_710), .B1(n_712), .B2(n_719), .C(n_723), .Y(n_705) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
OR2x6_ASAP7_75t_SL g742 ( .A(n_708), .B(n_743), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g956 ( .A1(n_708), .A2(n_957), .B1(n_958), .B2(n_961), .C(n_962), .Y(n_956) );
INVx3_ASAP7_75t_L g1075 ( .A(n_708), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1205 ( .A(n_708), .Y(n_1205) );
INVx3_ASAP7_75t_L g775 ( .A(n_711), .Y(n_775) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g913 ( .A(n_714), .Y(n_913) );
INVx1_ASAP7_75t_L g1054 ( .A(n_714), .Y(n_1054) );
INVx1_ASAP7_75t_L g1271 ( .A(n_714), .Y(n_1271) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI221xp5_ASAP7_75t_L g768 ( .A1(n_716), .A2(n_769), .B1(n_770), .B2(n_771), .C(n_772), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g899 ( .A1(n_716), .A2(n_739), .B1(n_900), .B2(n_901), .C(n_902), .Y(n_899) );
INVx3_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_SL g904 ( .A(n_717), .Y(n_904) );
INVx5_ASAP7_75t_L g1049 ( .A(n_717), .Y(n_1049) );
INVx2_ASAP7_75t_SL g1291 ( .A(n_717), .Y(n_1291) );
BUFx2_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx2_ASAP7_75t_L g833 ( .A(n_722), .Y(n_833) );
INVx2_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AOI22xp5_ASAP7_75t_L g776 ( .A1(n_725), .A2(n_728), .B1(n_757), .B2(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx4_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_735), .A2(n_737), .B1(n_765), .B2(n_766), .Y(n_764) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
OAI221xp5_ASAP7_75t_L g894 ( .A1(n_738), .A2(n_895), .B1(n_899), .B2(n_903), .C(n_907), .Y(n_894) );
OR2x6_ASAP7_75t_L g738 ( .A(n_739), .B(n_740), .Y(n_738) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
HB1xp67_ASAP7_75t_L g915 ( .A(n_744), .Y(n_915) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_746), .B(n_879), .Y(n_944) );
INVx1_ASAP7_75t_L g1233 ( .A(n_747), .Y(n_1233) );
HB1xp67_ASAP7_75t_L g1622 ( .A(n_747), .Y(n_1622) );
BUFx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx2_ASAP7_75t_L g1668 ( .A(n_748), .Y(n_1668) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_751), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_L g1595 ( .A(n_751), .Y(n_1595) );
AOI211x1_ASAP7_75t_L g755 ( .A1(n_756), .A2(n_757), .B(n_758), .C(n_784), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_761), .Y(n_758) );
NAND3xp33_ASAP7_75t_L g767 ( .A(n_768), .B(n_776), .C(n_778), .Y(n_767) );
INVx3_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_782), .C(n_783), .Y(n_778) );
OAI21xp5_ASAP7_75t_SL g907 ( .A1(n_780), .A2(n_908), .B(n_909), .Y(n_907) );
INVx3_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx2_ASAP7_75t_L g1046 ( .A(n_781), .Y(n_1046) );
INVx2_ASAP7_75t_L g1636 ( .A(n_781), .Y(n_1636) );
NAND3xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_798), .C(n_802), .Y(n_784) );
INVx1_ASAP7_75t_L g1320 ( .A(n_788), .Y(n_1320) );
INVx1_ASAP7_75t_L g997 ( .A(n_806), .Y(n_997) );
AOI22xp5_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_881), .B1(n_882), .B2(n_996), .Y(n_806) );
INVx2_ASAP7_75t_L g996 ( .A(n_807), .Y(n_996) );
XOR2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_880), .Y(n_807) );
NAND2xp5_ASAP7_75t_SL g808 ( .A(n_809), .B(n_846), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_823), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g812 ( .A(n_813), .B(n_817), .Y(n_812) );
NAND2xp5_ASAP7_75t_SL g817 ( .A(n_818), .B(n_822), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_819), .B(n_820), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g1285 ( .A(n_820), .B(n_1286), .Y(n_1285) );
INVx5_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx3_ASAP7_75t_L g1010 ( .A(n_821), .Y(n_1010) );
NAND3xp33_ASAP7_75t_L g1162 ( .A(n_822), .B(n_1163), .C(n_1165), .Y(n_1162) );
NAND4xp25_ASAP7_75t_SL g1281 ( .A(n_822), .B(n_1282), .C(n_1285), .D(n_1287), .Y(n_1281) );
AOI33xp33_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_825), .A3(n_828), .B1(n_832), .B2(n_834), .B3(n_835), .Y(n_823) );
NAND2xp5_ASAP7_75t_L g1156 ( .A(n_824), .B(n_1157), .Y(n_1156) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_843), .B(n_1013), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1106 ( .A1(n_843), .A2(n_1091), .B1(n_1092), .B2(n_1107), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_844), .A2(n_890), .B1(n_912), .B2(n_913), .Y(n_911) );
OAI21xp5_ASAP7_75t_L g846 ( .A1(n_847), .A2(n_862), .B(n_877), .Y(n_846) );
NAND3xp33_ASAP7_75t_SL g847 ( .A(n_848), .B(n_849), .C(n_861), .Y(n_847) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
INVx2_ASAP7_75t_L g1176 ( .A(n_852), .Y(n_1176) );
BUFx2_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_L g1103 ( .A(n_853), .Y(n_1103) );
BUFx3_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_SL g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
INVx4_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx5_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
BUFx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
OAI21xp5_ASAP7_75t_L g975 ( .A1(n_877), .A2(n_976), .B(n_987), .Y(n_975) );
AOI21xp5_ASAP7_75t_L g1125 ( .A1(n_877), .A2(n_1126), .B(n_1141), .Y(n_1125) );
OAI21xp5_ASAP7_75t_L g1304 ( .A1(n_877), .A2(n_1305), .B(n_1313), .Y(n_1304) );
INVx2_ASAP7_75t_L g877 ( .A(n_878), .Y(n_877) );
INVx1_ASAP7_75t_L g1105 ( .A(n_878), .Y(n_1105) );
BUFx2_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g1035 ( .A(n_879), .Y(n_1035) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_883), .A2(n_884), .B1(n_945), .B2(n_995), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
HB1xp67_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
XNOR2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
NOR2x1_ASAP7_75t_L g887 ( .A(n_888), .B(n_916), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_892), .Y(n_888) );
OAI211xp5_ASAP7_75t_L g931 ( .A1(n_900), .A2(n_932), .B(n_934), .C(n_936), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g1067 ( .A1(n_904), .A2(n_1068), .B(n_1069), .C(n_1071), .Y(n_1067) );
AOI22xp5_ASAP7_75t_L g924 ( .A1(n_912), .A2(n_925), .B1(n_926), .B2(n_927), .Y(n_924) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
NAND3xp33_ASAP7_75t_L g916 ( .A(n_917), .B(n_937), .C(n_941), .Y(n_916) );
NOR3xp33_ASAP7_75t_SL g917 ( .A(n_918), .B(n_928), .C(n_930), .Y(n_917) );
OAI21xp5_ASAP7_75t_SL g918 ( .A1(n_919), .A2(n_922), .B(n_924), .Y(n_918) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g937 ( .A(n_938), .B(n_939), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g941 ( .A(n_942), .B(n_943), .Y(n_941) );
INVx1_ASAP7_75t_L g995 ( .A(n_945), .Y(n_995) );
INVx1_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
AND4x1_ASAP7_75t_L g948 ( .A(n_949), .B(n_953), .C(n_975), .D(n_994), .Y(n_948) );
INVx1_ASAP7_75t_SL g1062 ( .A(n_952), .Y(n_1062) );
NOR3xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .C(n_972), .Y(n_953) );
NOR3xp33_ASAP7_75t_L g1196 ( .A(n_954), .B(n_1197), .C(n_1209), .Y(n_1196) );
OAI221xp5_ASAP7_75t_L g1671 ( .A1(n_958), .A2(n_1672), .B1(n_1673), .B2(n_1674), .C(n_1675), .Y(n_1671) );
INVx3_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
BUFx2_ASAP7_75t_L g959 ( .A(n_960), .Y(n_959) );
INVx2_ASAP7_75t_L g964 ( .A(n_965), .Y(n_964) );
INVx2_ASAP7_75t_L g1072 ( .A(n_965), .Y(n_1072) );
CKINVDCx5p33_ASAP7_75t_R g1676 ( .A(n_965), .Y(n_1676) );
OAI221xp5_ASAP7_75t_L g966 ( .A1(n_967), .A2(n_968), .B1(n_969), .B2(n_970), .C(n_971), .Y(n_966) );
OAI211xp5_ASAP7_75t_L g988 ( .A1(n_968), .A2(n_989), .B(n_991), .C(n_992), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g1677 ( .A1(n_969), .A2(n_1662), .B1(n_1672), .B2(n_1678), .C(n_1679), .Y(n_1677) );
INVx1_ASAP7_75t_L g973 ( .A(n_974), .Y(n_973) );
AOI22xp5_ASAP7_75t_L g1114 ( .A1(n_974), .A2(n_1115), .B1(n_1116), .B2(n_1117), .Y(n_1114) );
INVx2_ASAP7_75t_SL g980 ( .A(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g1089 ( .A(n_981), .Y(n_1089) );
INVx3_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
BUFx6f_ASAP7_75t_L g1309 ( .A(n_982), .Y(n_1309) );
INVx1_ASAP7_75t_L g1033 ( .A(n_985), .Y(n_1033) );
OAI211xp5_ASAP7_75t_L g1612 ( .A1(n_989), .A2(n_1613), .B(n_1614), .C(n_1615), .Y(n_1612) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx2_ASAP7_75t_L g1317 ( .A(n_990), .Y(n_1317) );
INVx1_ASAP7_75t_L g1606 ( .A(n_990), .Y(n_1606) );
INVxp67_ASAP7_75t_SL g1369 ( .A(n_998), .Y(n_1369) );
XOR2x2_ASAP7_75t_L g998 ( .A(n_999), .B(n_1235), .Y(n_998) );
XOR2xp5_ASAP7_75t_L g999 ( .A(n_1000), .B(n_1146), .Y(n_999) );
AOI22xp5_ASAP7_75t_L g1000 ( .A1(n_1001), .A2(n_1002), .B1(n_1056), .B2(n_1145), .Y(n_1000) );
INVx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
XNOR2x1_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1055), .Y(n_1002) );
NOR2x1_ASAP7_75t_L g1003 ( .A(n_1004), .B(n_1014), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1010), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g1060 ( .A1(n_1010), .A2(n_1061), .B1(n_1062), .B2(n_1063), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1163 ( .A(n_1010), .B(n_1164), .Y(n_1163) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1036), .Y(n_1014) );
OAI31xp33_ASAP7_75t_L g1015 ( .A1(n_1016), .A2(n_1025), .A3(n_1032), .B(n_1035), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
OAI221xp5_ASAP7_75t_L g1047 ( .A1(n_1021), .A2(n_1048), .B1(n_1050), .B2(n_1051), .C(n_1052), .Y(n_1047) );
OAI21xp5_ASAP7_75t_L g1243 ( .A1(n_1035), .A2(n_1244), .B(n_1253), .Y(n_1243) );
AOI21xp5_ASAP7_75t_SL g1036 ( .A1(n_1037), .A2(n_1038), .B(n_1039), .Y(n_1036) );
AOI21xp5_ASAP7_75t_L g1300 ( .A1(n_1037), .A2(n_1301), .B(n_1302), .Y(n_1300) );
OAI22xp33_ASAP7_75t_L g1348 ( .A1(n_1046), .A2(n_1340), .B1(n_1349), .B2(n_1350), .Y(n_1348) );
OAI22xp5_ASAP7_75t_L g1339 ( .A1(n_1048), .A2(n_1340), .B1(n_1342), .B2(n_1343), .Y(n_1339) );
BUFx3_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
INVx8_ASAP7_75t_L g1207 ( .A(n_1049), .Y(n_1207) );
OAI221xp5_ASAP7_75t_L g1073 ( .A1(n_1051), .A2(n_1074), .B1(n_1076), .B2(n_1077), .C(n_1078), .Y(n_1073) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1056), .Y(n_1145) );
XNOR2x1_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1108), .Y(n_1056) );
NAND4xp75_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1064), .C(n_1082), .D(n_1106), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1067), .B1(n_1072), .B2(n_1073), .Y(n_1065) );
INVx2_ASAP7_75t_L g1074 ( .A(n_1075), .Y(n_1074) );
INVx1_ASAP7_75t_L g1080 ( .A(n_1081), .Y(n_1080) );
OAI21xp5_ASAP7_75t_L g1082 ( .A1(n_1083), .A2(n_1093), .B(n_1105), .Y(n_1082) );
NAND2xp5_ASAP7_75t_L g1083 ( .A(n_1084), .B(n_1090), .Y(n_1083) );
INVx2_ASAP7_75t_L g1621 ( .A(n_1085), .Y(n_1621) );
OAI221xp5_ASAP7_75t_L g1094 ( .A1(n_1095), .A2(n_1096), .B1(n_1097), .B2(n_1099), .C(n_1100), .Y(n_1094) );
BUFx3_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx2_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
INVx1_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_1110), .B(n_1125), .Y(n_1109) );
AOI222xp33_ASAP7_75t_L g1134 ( .A1(n_1115), .A2(n_1117), .B1(n_1135), .B2(n_1136), .C1(n_1138), .C2(n_1139), .Y(n_1134) );
AOI22xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1121), .B1(n_1122), .B2(n_1124), .Y(n_1118) );
NAND3xp33_ASAP7_75t_L g1126 ( .A(n_1127), .B(n_1130), .C(n_1134), .Y(n_1126) );
AOI22xp33_ASAP7_75t_L g1142 ( .A1(n_1128), .A2(n_1129), .B1(n_1143), .B2(n_1144), .Y(n_1142) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1135), .Y(n_1188) );
INVx1_ASAP7_75t_L g1189 ( .A(n_1139), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1607 ( .A1(n_1140), .A2(n_1598), .B1(n_1608), .B2(n_1609), .Y(n_1607) );
INVx2_ASAP7_75t_SL g1594 ( .A(n_1144), .Y(n_1594) );
OAI22x1_ASAP7_75t_L g1146 ( .A1(n_1147), .A2(n_1148), .B1(n_1194), .B2(n_1234), .Y(n_1146) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1148), .Y(n_1147) );
XNOR2x1_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1150), .Y(n_1148) );
AND3x2_ASAP7_75t_L g1150 ( .A(n_1151), .B(n_1168), .C(n_1192), .Y(n_1150) );
NOR2xp33_ASAP7_75t_SL g1151 ( .A(n_1152), .B(n_1162), .Y(n_1151) );
OAI21xp5_ASAP7_75t_SL g1152 ( .A1(n_1153), .A2(n_1156), .B(n_1159), .Y(n_1152) );
NAND3xp33_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1173), .C(n_1179), .Y(n_1169) );
AOI31xp33_ASAP7_75t_L g1179 ( .A1(n_1180), .A2(n_1183), .A3(n_1184), .B(n_1187), .Y(n_1179) );
BUFx2_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1186), .Y(n_1259) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1194), .Y(n_1234) );
NAND3xp33_ASAP7_75t_L g1195 ( .A(n_1196), .B(n_1210), .C(n_1213), .Y(n_1195) );
NAND2xp5_ASAP7_75t_L g1197 ( .A(n_1198), .B(n_1201), .Y(n_1197) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g1213 ( .A1(n_1214), .A2(n_1225), .B(n_1232), .Y(n_1213) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_1227), .B(n_1229), .Y(n_1226) );
OAI21xp5_ASAP7_75t_L g1351 ( .A1(n_1232), .A2(n_1352), .B(n_1355), .Y(n_1351) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
XNOR2x1_ASAP7_75t_L g1235 ( .A(n_1236), .B(n_1326), .Y(n_1235) );
OAI22x1_ASAP7_75t_L g1236 ( .A1(n_1237), .A2(n_1276), .B1(n_1277), .B2(n_1325), .Y(n_1236) );
INVx2_ASAP7_75t_L g1325 ( .A(n_1237), .Y(n_1325) );
AO21x2_ASAP7_75t_L g1237 ( .A1(n_1238), .A2(n_1239), .B(n_1275), .Y(n_1237) );
NAND3xp33_ASAP7_75t_SL g1239 ( .A(n_1240), .B(n_1243), .C(n_1260), .Y(n_1239) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1261 ( .A(n_1262), .Y(n_1261) );
INVx2_ASAP7_75t_L g1276 ( .A(n_1277), .Y(n_1276) );
NAND2x1p5_ASAP7_75t_L g1277 ( .A(n_1278), .B(n_1297), .Y(n_1277) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_1280), .B(n_1295), .Y(n_1279) );
INVxp67_ASAP7_75t_L g1280 ( .A(n_1281), .Y(n_1280) );
NOR2xp33_ASAP7_75t_SL g1322 ( .A(n_1281), .B(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1295), .B(n_1324), .Y(n_1323) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
NAND2xp5_ASAP7_75t_L g1299 ( .A(n_1300), .B(n_1304), .Y(n_1299) );
A2O1A1Ixp33_ASAP7_75t_L g1603 ( .A1(n_1309), .A2(n_1604), .B(n_1605), .C(n_1611), .Y(n_1603) );
OAI211xp5_ASAP7_75t_L g1315 ( .A1(n_1316), .A2(n_1317), .B(n_1318), .C(n_1321), .Y(n_1315) );
OAI211xp5_ASAP7_75t_L g1616 ( .A1(n_1317), .A2(n_1617), .B(n_1618), .C(n_1619), .Y(n_1616) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1320), .Y(n_1319) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1328), .Y(n_1327) );
AND3x2_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1351), .C(n_1364), .Y(n_1328) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1332), .Y(n_1331) );
OAI22xp5_ASAP7_75t_SL g1670 ( .A1(n_1335), .A2(n_1671), .B1(n_1676), .B2(n_1677), .Y(n_1670) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1341), .Y(n_1340) );
INVx1_ASAP7_75t_L g1632 ( .A(n_1345), .Y(n_1632) );
OAI221xp5_ASAP7_75t_SL g1370 ( .A1(n_1371), .A2(n_1581), .B1(n_1585), .B2(n_1637), .C(n_1640), .Y(n_1370) );
AND5x1_ASAP7_75t_L g1371 ( .A(n_1372), .B(n_1537), .C(n_1554), .D(n_1563), .E(n_1574), .Y(n_1371) );
OAI33xp33_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1465), .A3(n_1482), .B1(n_1491), .B2(n_1518), .B3(n_1532), .Y(n_1372) );
OAI211xp5_ASAP7_75t_SL g1373 ( .A1(n_1374), .A2(n_1395), .B(n_1412), .C(n_1455), .Y(n_1373) );
CKINVDCx5p33_ASAP7_75t_R g1472 ( .A(n_1374), .Y(n_1472) );
OR2x2_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1390), .Y(n_1374) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_1375), .A2(n_1422), .B1(n_1425), .B2(n_1428), .Y(n_1421) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1375), .B(n_1429), .Y(n_1428) );
OR2x2_ASAP7_75t_L g1464 ( .A(n_1375), .B(n_1391), .Y(n_1464) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1375), .Y(n_1475) );
INVx2_ASAP7_75t_L g1493 ( .A(n_1375), .Y(n_1493) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1375), .B(n_1431), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1553 ( .A(n_1375), .B(n_1430), .Y(n_1553) );
AND2x2_ASAP7_75t_L g1562 ( .A(n_1375), .B(n_1431), .Y(n_1562) );
INVx2_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1414 ( .A(n_1376), .B(n_1390), .Y(n_1414) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1384), .Y(n_1376) );
AND2x6_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1380), .Y(n_1378) );
AND2x2_ASAP7_75t_L g1382 ( .A(n_1379), .B(n_1383), .Y(n_1382) );
AND2x4_ASAP7_75t_L g1385 ( .A(n_1379), .B(n_1386), .Y(n_1385) );
AND2x6_ASAP7_75t_L g1388 ( .A(n_1379), .B(n_1389), .Y(n_1388) );
AND2x2_ASAP7_75t_L g1393 ( .A(n_1379), .B(n_1383), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1434 ( .A(n_1379), .B(n_1383), .Y(n_1434) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1379), .B(n_1386), .Y(n_1443) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1381), .B(n_1387), .Y(n_1386) );
OAI21xp5_ASAP7_75t_L g1687 ( .A1(n_1383), .A2(n_1688), .B(n_1689), .Y(n_1687) );
INVx2_ASAP7_75t_L g1445 ( .A(n_1388), .Y(n_1445) );
INVx1_ASAP7_75t_L g1436 ( .A(n_1390), .Y(n_1436) );
NOR2xp33_ASAP7_75t_L g1550 ( .A(n_1390), .B(n_1477), .Y(n_1550) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1391), .Y(n_1429) );
NAND2xp5_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1394), .Y(n_1391) );
OR2x2_ASAP7_75t_L g1395 ( .A(n_1396), .B(n_1400), .Y(n_1395) );
NOR2xp33_ASAP7_75t_L g1422 ( .A(n_1396), .B(n_1423), .Y(n_1422) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1396), .B(n_1458), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1490 ( .A(n_1396), .B(n_1472), .Y(n_1490) );
CKINVDCx5p33_ASAP7_75t_R g1517 ( .A(n_1396), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1396), .B(n_1426), .Y(n_1524) );
NAND2xp5_ASAP7_75t_L g1533 ( .A(n_1396), .B(n_1439), .Y(n_1533) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1396), .B(n_1436), .Y(n_1566) );
INVx4_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
O2A1O1Ixp33_ASAP7_75t_L g1448 ( .A1(n_1397), .A2(n_1449), .B(n_1451), .C(n_1454), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1452 ( .A(n_1397), .B(n_1453), .Y(n_1452) );
INVx4_ASAP7_75t_L g1468 ( .A(n_1397), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1470 ( .A(n_1397), .B(n_1471), .Y(n_1470) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1397), .B(n_1418), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1476 ( .A(n_1397), .B(n_1466), .Y(n_1476) );
NAND2xp5_ASAP7_75t_SL g1481 ( .A(n_1397), .B(n_1418), .Y(n_1481) );
NOR2xp33_ASAP7_75t_L g1488 ( .A(n_1397), .B(n_1419), .Y(n_1488) );
NOR3xp33_ASAP7_75t_L g1510 ( .A(n_1397), .B(n_1507), .C(n_1511), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1397), .B(n_1460), .Y(n_1561) );
AND2x4_ASAP7_75t_SL g1397 ( .A(n_1398), .B(n_1399), .Y(n_1397) );
NOR2xp33_ASAP7_75t_L g1536 ( .A(n_1400), .B(n_1499), .Y(n_1536) );
OR2x2_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1404), .Y(n_1400) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_1401), .B(n_1406), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1504 ( .A(n_1401), .B(n_1505), .Y(n_1504) );
AND2x2_ASAP7_75t_L g1512 ( .A(n_1401), .B(n_1453), .Y(n_1512) );
NAND2xp5_ASAP7_75t_L g1578 ( .A(n_1401), .B(n_1488), .Y(n_1578) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1403), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1402), .B(n_1403), .Y(n_1418) );
OR2x2_ASAP7_75t_L g1528 ( .A(n_1404), .B(n_1417), .Y(n_1528) );
NAND2xp5_ASAP7_75t_L g1575 ( .A(n_1404), .B(n_1576), .Y(n_1575) );
NAND2xp5_ASAP7_75t_L g1404 ( .A(n_1405), .B(n_1409), .Y(n_1404) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
OR2x2_ASAP7_75t_L g1419 ( .A(n_1406), .B(n_1409), .Y(n_1419) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1406), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1406), .B(n_1409), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1453 ( .A(n_1406), .B(n_1427), .Y(n_1453) );
NAND2xp5_ASAP7_75t_L g1497 ( .A(n_1406), .B(n_1418), .Y(n_1497) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1407), .B(n_1408), .Y(n_1406) );
INVx2_ASAP7_75t_L g1427 ( .A(n_1409), .Y(n_1427) );
NAND2x1p5_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1411), .Y(n_1409) );
AOI211xp5_ASAP7_75t_L g1412 ( .A1(n_1413), .A2(n_1415), .B(n_1420), .C(n_1448), .Y(n_1412) );
NAND2xp5_ASAP7_75t_L g1516 ( .A(n_1413), .B(n_1517), .Y(n_1516) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_1414), .Y(n_1413) );
OR2x2_ASAP7_75t_L g1580 ( .A(n_1414), .B(n_1430), .Y(n_1580) );
INVx1_ASAP7_75t_L g1415 ( .A(n_1416), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1508 ( .A(n_1416), .B(n_1462), .Y(n_1508) );
OR2x2_ASAP7_75t_L g1416 ( .A(n_1417), .B(n_1419), .Y(n_1416) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1417), .B(n_1427), .Y(n_1426) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1417), .B(n_1453), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1417), .B(n_1479), .Y(n_1514) );
A2O1A1Ixp33_ASAP7_75t_L g1574 ( .A1(n_1417), .A2(n_1575), .B(n_1577), .C(n_1579), .Y(n_1574) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_1418), .B(n_1424), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1438 ( .A(n_1418), .B(n_1439), .Y(n_1438) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1418), .B(n_1424), .Y(n_1450) );
OR2x2_ASAP7_75t_L g1471 ( .A(n_1418), .B(n_1427), .Y(n_1471) );
AND2x2_ASAP7_75t_L g1547 ( .A(n_1418), .B(n_1427), .Y(n_1547) );
INVx1_ASAP7_75t_L g1479 ( .A(n_1419), .Y(n_1479) );
OR2x2_ASAP7_75t_L g1540 ( .A(n_1419), .B(n_1474), .Y(n_1540) );
OAI221xp5_ASAP7_75t_SL g1420 ( .A1(n_1421), .A2(n_1430), .B1(n_1435), .B2(n_1437), .C(n_1440), .Y(n_1420) );
HB1xp67_ASAP7_75t_L g1425 ( .A(n_1426), .Y(n_1425) );
INVx1_ASAP7_75t_L g1521 ( .A(n_1428), .Y(n_1521) );
OR2x2_ASAP7_75t_L g1454 ( .A(n_1429), .B(n_1430), .Y(n_1454) );
INVx2_ASAP7_75t_L g1466 ( .A(n_1429), .Y(n_1466) );
OAI221xp5_ASAP7_75t_L g1482 ( .A1(n_1429), .A2(n_1475), .B1(n_1483), .B2(n_1487), .C(n_1489), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1498 ( .A(n_1429), .B(n_1499), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1526 ( .A(n_1429), .B(n_1468), .Y(n_1526) );
A2O1A1Ixp33_ASAP7_75t_L g1554 ( .A1(n_1429), .A2(n_1555), .B(n_1561), .C(n_1562), .Y(n_1554) );
OR2x2_ASAP7_75t_L g1435 ( .A(n_1430), .B(n_1436), .Y(n_1435) );
A2O1A1Ixp33_ASAP7_75t_L g1469 ( .A1(n_1430), .A2(n_1470), .B(n_1472), .C(n_1473), .Y(n_1469) );
CKINVDCx14_ASAP7_75t_R g1531 ( .A(n_1430), .Y(n_1531) );
INVx3_ASAP7_75t_L g1430 ( .A(n_1431), .Y(n_1430) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1431), .Y(n_1463) );
AOI221xp5_ASAP7_75t_L g1537 ( .A1(n_1431), .A2(n_1466), .B1(n_1538), .B2(n_1541), .C(n_1548), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1543 ( .A(n_1431), .B(n_1475), .Y(n_1543) );
OAI21xp33_ASAP7_75t_L g1548 ( .A1(n_1431), .A2(n_1549), .B(n_1551), .Y(n_1548) );
AND2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
HB1xp67_ASAP7_75t_L g1584 ( .A(n_1434), .Y(n_1584) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1436), .Y(n_1485) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
NAND2x1_ASAP7_75t_L g1467 ( .A(n_1438), .B(n_1468), .Y(n_1467) );
OAI21xp33_ASAP7_75t_L g1551 ( .A1(n_1438), .A2(n_1552), .B(n_1553), .Y(n_1551) );
OAI321xp33_ASAP7_75t_L g1473 ( .A1(n_1439), .A2(n_1449), .A3(n_1474), .B1(n_1475), .B2(n_1476), .C(n_1477), .Y(n_1473) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1439), .Y(n_1505) );
OAI21xp5_ASAP7_75t_L g1513 ( .A1(n_1439), .A2(n_1514), .B(n_1515), .Y(n_1513) );
AND2x2_ASAP7_75t_L g1545 ( .A(n_1439), .B(n_1480), .Y(n_1545) );
AOI211xp5_ASAP7_75t_L g1522 ( .A1(n_1440), .A2(n_1523), .B(n_1524), .C(n_1525), .Y(n_1522) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1441), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1530 ( .A(n_1441), .B(n_1531), .Y(n_1530) );
INVx1_ASAP7_75t_L g1441 ( .A(n_1442), .Y(n_1441) );
OAI221xp5_ASAP7_75t_L g1442 ( .A1(n_1443), .A2(n_1444), .B1(n_1445), .B2(n_1446), .C(n_1447), .Y(n_1442) );
NAND2xp5_ASAP7_75t_SL g1503 ( .A(n_1449), .B(n_1504), .Y(n_1503) );
O2A1O1Ixp33_ASAP7_75t_L g1518 ( .A1(n_1449), .A2(n_1519), .B(n_1522), .C(n_1529), .Y(n_1518) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
NAND2xp5_ASAP7_75t_L g1489 ( .A(n_1450), .B(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1576 ( .A(n_1453), .Y(n_1576) );
OAI322xp33_ASAP7_75t_L g1532 ( .A1(n_1454), .A2(n_1459), .A3(n_1463), .B1(n_1472), .B2(n_1533), .C1(n_1534), .C2(n_1535), .Y(n_1532) );
OAI21xp33_ASAP7_75t_L g1455 ( .A1(n_1456), .A2(n_1460), .B(n_1461), .Y(n_1455) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1457), .Y(n_1456) );
INVxp67_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g1486 ( .A(n_1459), .B(n_1468), .Y(n_1486) );
NAND2xp5_ASAP7_75t_L g1501 ( .A(n_1460), .B(n_1472), .Y(n_1501) );
INVx1_ASAP7_75t_L g1571 ( .A(n_1460), .Y(n_1571) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1462), .Y(n_1461) );
OR2x2_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1464), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1565 ( .A(n_1463), .B(n_1566), .Y(n_1565) );
OAI21xp33_ASAP7_75t_L g1465 ( .A1(n_1466), .A2(n_1467), .B(n_1469), .Y(n_1465) );
OR2x2_ASAP7_75t_L g1534 ( .A(n_1466), .B(n_1507), .Y(n_1534) );
CKINVDCx5p33_ASAP7_75t_R g1499 ( .A(n_1468), .Y(n_1499) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_1472), .B(n_1517), .Y(n_1573) );
NOR2xp33_ASAP7_75t_L g1494 ( .A(n_1475), .B(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1475), .Y(n_1523) );
INVx1_ASAP7_75t_L g1477 ( .A(n_1478), .Y(n_1477) );
AOI211xp5_ASAP7_75t_L g1492 ( .A1(n_1478), .A2(n_1493), .B(n_1494), .C(n_1500), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1570 ( .A(n_1478), .B(n_1485), .Y(n_1570) );
AND2x2_ASAP7_75t_L g1478 ( .A(n_1479), .B(n_1480), .Y(n_1478) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVxp67_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
AND2x2_ASAP7_75t_L g1484 ( .A(n_1485), .B(n_1486), .Y(n_1484) );
AND2x2_ASAP7_75t_L g1538 ( .A(n_1485), .B(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
O2A1O1Ixp33_ASAP7_75t_L g1563 ( .A1(n_1490), .A2(n_1564), .B(n_1567), .C(n_1569), .Y(n_1563) );
NAND4xp25_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1502), .C(n_1509), .D(n_1513), .Y(n_1491) );
INVxp33_ASAP7_75t_L g1552 ( .A(n_1495), .Y(n_1552) );
NAND2xp5_ASAP7_75t_L g1495 ( .A(n_1496), .B(n_1498), .Y(n_1495) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
OR2x2_ASAP7_75t_L g1558 ( .A(n_1497), .B(n_1517), .Y(n_1558) );
AOI31xp33_ASAP7_75t_L g1502 ( .A1(n_1499), .A2(n_1503), .A3(n_1506), .B(n_1508), .Y(n_1502) );
NOR2xp33_ASAP7_75t_L g1520 ( .A(n_1499), .B(n_1521), .Y(n_1520) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
CKINVDCx14_ASAP7_75t_R g1506 ( .A(n_1507), .Y(n_1506) );
OAI22xp5_ASAP7_75t_L g1541 ( .A1(n_1507), .A2(n_1542), .B1(n_1544), .B2(n_1546), .Y(n_1541) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1510), .Y(n_1509) );
AND2x2_ASAP7_75t_L g1568 ( .A(n_1511), .B(n_1560), .Y(n_1568) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1560 ( .A(n_1514), .Y(n_1560) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVxp67_ASAP7_75t_SL g1519 ( .A(n_1520), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1569 ( .A1(n_1523), .A2(n_1570), .B1(n_1571), .B2(n_1572), .Y(n_1569) );
INVx1_ASAP7_75t_L g1559 ( .A(n_1524), .Y(n_1559) );
AND2x2_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1527), .Y(n_1525) );
INVx1_ASAP7_75t_L g1527 ( .A(n_1528), .Y(n_1527) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
INVx1_ASAP7_75t_L g1539 ( .A(n_1540), .Y(n_1539) );
INVx1_ASAP7_75t_L g1542 ( .A(n_1543), .Y(n_1542) );
INVx1_ASAP7_75t_L g1544 ( .A(n_1545), .Y(n_1544) );
CKINVDCx14_ASAP7_75t_R g1546 ( .A(n_1547), .Y(n_1546) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
NAND2xp5_ASAP7_75t_L g1555 ( .A(n_1556), .B(n_1560), .Y(n_1555) );
INVxp67_ASAP7_75t_SL g1556 ( .A(n_1557), .Y(n_1556) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_1558), .B(n_1559), .Y(n_1557) );
INVx1_ASAP7_75t_L g1564 ( .A(n_1565), .Y(n_1564) );
INVxp67_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1578), .Y(n_1577) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
CKINVDCx20_ASAP7_75t_R g1581 ( .A(n_1582), .Y(n_1581) );
CKINVDCx20_ASAP7_75t_R g1582 ( .A(n_1583), .Y(n_1582) );
INVx4_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
INVxp67_ASAP7_75t_SL g1585 ( .A(n_1586), .Y(n_1585) );
XNOR2x1_ASAP7_75t_L g1586 ( .A(n_1587), .B(n_1588), .Y(n_1586) );
NOR2x1_ASAP7_75t_L g1588 ( .A(n_1589), .B(n_1596), .Y(n_1588) );
INVxp67_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
NAND2x1_ASAP7_75t_L g1593 ( .A(n_1594), .B(n_1595), .Y(n_1593) );
NAND3xp33_ASAP7_75t_SL g1596 ( .A(n_1597), .B(n_1601), .C(n_1623), .Y(n_1596) );
OAI21xp5_ASAP7_75t_L g1601 ( .A1(n_1602), .A2(n_1620), .B(n_1622), .Y(n_1601) );
NAND3xp33_ASAP7_75t_L g1602 ( .A(n_1603), .B(n_1612), .C(n_1616), .Y(n_1602) );
NAND2xp5_ASAP7_75t_SL g1605 ( .A(n_1606), .B(n_1607), .Y(n_1605) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
OAI22xp5_ASAP7_75t_L g1625 ( .A1(n_1617), .A2(n_1626), .B1(n_1627), .B2(n_1629), .Y(n_1625) );
BUFx4f_ASAP7_75t_SL g1627 ( .A(n_1628), .Y(n_1627) );
INVx2_ASAP7_75t_L g1629 ( .A(n_1630), .Y(n_1629) );
INVx2_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1641 ( .A(n_1642), .Y(n_1641) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_1644), .Y(n_1643) );
BUFx3_ASAP7_75t_L g1644 ( .A(n_1645), .Y(n_1644) );
INVxp33_ASAP7_75t_L g1646 ( .A(n_1647), .Y(n_1646) );
HB1xp67_ASAP7_75t_L g1648 ( .A(n_1649), .Y(n_1648) );
AND4x1_ASAP7_75t_L g1649 ( .A(n_1650), .B(n_1669), .C(n_1681), .D(n_1684), .Y(n_1649) );
OAI21xp5_ASAP7_75t_L g1650 ( .A1(n_1651), .A2(n_1660), .B(n_1668), .Y(n_1650) );
INVx2_ASAP7_75t_SL g1654 ( .A(n_1655), .Y(n_1654) );
OAI211xp5_ASAP7_75t_L g1661 ( .A1(n_1662), .A2(n_1663), .B(n_1665), .C(n_1667), .Y(n_1661) );
INVx5_ASAP7_75t_L g1663 ( .A(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1685 ( .A(n_1686), .Y(n_1685) );
INVx1_ASAP7_75t_L g1686 ( .A(n_1687), .Y(n_1686) );
INVx1_ASAP7_75t_L g1689 ( .A(n_1690), .Y(n_1689) );
endmodule