module fake_jpeg_10993_n_149 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_149);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_149;

wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_93;
wire n_54;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_6),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_14),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_11),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_17),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_10),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_24),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_0),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_12),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_35),
.Y(n_66)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_8),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_49),
.B(n_0),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_72),
.Y(n_89)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_70),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_73),
.A2(n_77),
.B(n_5),
.Y(n_88)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_26),
.B1(n_45),
.B2(n_44),
.Y(n_74)
);

AO21x1_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_68),
.B(n_57),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_1),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_78),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_62),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_77),
.B(n_47),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_83),
.B(n_85),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_60),
.B1(n_54),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_87),
.B1(n_79),
.B2(n_90),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_75),
.B(n_63),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_88),
.A2(n_5),
.B(n_6),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_91),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_69),
.Y(n_91)
);

O2A1O1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_88),
.A2(n_52),
.B(n_61),
.C(n_59),
.Y(n_92)
);

AO21x1_ASAP7_75t_L g122 ( 
.A1(n_92),
.A2(n_105),
.B(n_108),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx13_ASAP7_75t_L g94 ( 
.A(n_79),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

NOR2x1_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_98),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_58),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_97),
.B(n_102),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_87),
.A2(n_58),
.B1(n_56),
.B2(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_99),
.A2(n_106),
.B1(n_19),
.B2(n_22),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_29),
.C(n_41),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_100),
.B(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_51),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_101),
.B(n_107),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_103),
.A2(n_30),
.B(n_31),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_80),
.B(n_66),
.Y(n_104)
);

A2O1A1Ixp33_ASAP7_75t_L g105 ( 
.A1(n_80),
.A2(n_7),
.B(n_9),
.C(n_10),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_81),
.A2(n_56),
.B1(n_55),
.B2(n_7),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_90),
.B(n_9),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_15),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_110),
.B(n_114),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_113),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_25),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_97),
.A2(n_27),
.B(n_28),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_123),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_92),
.B(n_34),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_117),
.B(n_118),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_102),
.A2(n_36),
.B1(n_38),
.B2(n_42),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_105),
.A2(n_43),
.B(n_46),
.Y(n_119)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_119),
.A2(n_100),
.B(n_121),
.C(n_115),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_93),
.B(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_124),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_94),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_125),
.Y(n_133)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_120),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_134),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_136),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_131),
.B(n_122),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_117),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_137),
.B(n_136),
.Y(n_144)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_133),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_141),
.Y(n_142)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_135),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_128),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_143),
.B(n_144),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_145),
.A2(n_126),
.B(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_146),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_147),
.A2(n_142),
.B(n_132),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_148),
.B(n_129),
.C(n_139),
.Y(n_149)
);


endmodule