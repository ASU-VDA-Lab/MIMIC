module fake_netlist_5_156_n_2933 (n_137, n_294, n_431, n_318, n_380, n_419, n_444, n_469, n_82, n_194, n_316, n_389, n_549, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_408, n_61, n_376, n_503, n_127, n_75, n_235, n_226, n_74, n_515, n_57, n_353, n_351, n_367, n_452, n_397, n_493, n_111, n_525, n_483, n_544, n_155, n_552, n_547, n_43, n_116, n_22, n_467, n_564, n_423, n_284, n_46, n_245, n_21, n_501, n_139, n_38, n_105, n_280, n_590, n_4, n_378, n_551, n_17, n_581, n_382, n_554, n_254, n_33, n_23, n_583, n_302, n_265, n_526, n_293, n_372, n_443, n_244, n_47, n_173, n_198, n_447, n_247, n_314, n_368, n_433, n_8, n_321, n_292, n_100, n_455, n_417, n_212, n_385, n_498, n_516, n_507, n_119, n_497, n_559, n_275, n_252, n_26, n_295, n_133, n_330, n_508, n_506, n_2, n_6, n_509, n_568, n_39, n_147, n_373, n_67, n_307, n_439, n_87, n_150, n_530, n_556, n_106, n_209, n_259, n_448, n_375, n_301, n_576, n_68, n_93, n_186, n_537, n_134, n_191, n_587, n_51, n_63, n_492, n_563, n_171, n_153, n_524, n_399, n_341, n_204, n_394, n_250, n_579, n_548, n_543, n_260, n_298, n_320, n_518, n_505, n_286, n_122, n_282, n_331, n_10, n_24, n_406, n_519, n_470, n_325, n_449, n_132, n_90, n_546, n_101, n_281, n_240, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_31, n_456, n_13, n_371, n_481, n_535, n_152, n_540, n_317, n_9, n_323, n_569, n_195, n_42, n_356, n_227, n_592, n_45, n_271, n_94, n_335, n_123, n_370, n_167, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_297, n_156, n_5, n_225, n_377, n_484, n_219, n_442, n_157, n_131, n_192, n_223, n_392, n_158, n_138, n_264, n_109, n_472, n_454, n_387, n_374, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_398, n_396, n_347, n_169, n_59, n_522, n_550, n_255, n_215, n_350, n_196, n_459, n_211, n_218, n_400, n_181, n_436, n_3, n_290, n_580, n_221, n_178, n_386, n_578, n_287, n_344, n_555, n_473, n_422, n_475, n_72, n_104, n_41, n_415, n_56, n_141, n_485, n_496, n_355, n_486, n_15, n_336, n_584, n_591, n_145, n_48, n_521, n_50, n_337, n_430, n_313, n_88, n_479, n_528, n_510, n_216, n_168, n_395, n_164, n_432, n_553, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_369, n_296, n_241, n_357, n_184, n_446, n_445, n_65, n_78, n_144, n_114, n_96, n_165, n_468, n_499, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_363, n_402, n_413, n_197, n_107, n_573, n_69, n_236, n_388, n_1, n_249, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_309, n_30, n_512, n_14, n_84, n_462, n_130, n_322, n_567, n_258, n_29, n_79, n_151, n_25, n_306, n_458, n_288, n_188, n_190, n_201, n_263, n_471, n_44, n_224, n_40, n_34, n_228, n_283, n_383, n_474, n_112, n_542, n_85, n_463, n_488, n_502, n_239, n_466, n_420, n_489, n_55, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_586, n_465, n_76, n_358, n_362, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_440, n_478, n_545, n_441, n_450, n_312, n_476, n_429, n_534, n_345, n_210, n_494, n_365, n_91, n_176, n_557, n_182, n_143, n_83, n_354, n_575, n_480, n_237, n_425, n_513, n_407, n_527, n_180, n_560, n_340, n_207, n_561, n_37, n_346, n_393, n_229, n_108, n_487, n_495, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_16, n_0, n_58, n_405, n_18, n_359, n_490, n_117, n_326, n_233, n_404, n_205, n_366, n_572, n_113, n_246, n_179, n_125, n_410, n_558, n_269, n_529, n_128, n_285, n_412, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_491, n_427, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_409, n_589, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_435, n_159, n_334, n_541, n_391, n_434, n_539, n_175, n_538, n_262, n_238, n_99, n_411, n_414, n_319, n_364, n_20, n_536, n_531, n_121, n_242, n_360, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_438, n_115, n_324, n_416, n_199, n_187, n_32, n_401, n_103, n_348, n_97, n_166, n_11, n_424, n_7, n_256, n_305, n_533, n_52, n_278, n_110, n_2933);

input n_137;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_444;
input n_469;
input n_82;
input n_194;
input n_316;
input n_389;
input n_549;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_408;
input n_61;
input n_376;
input n_503;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_515;
input n_57;
input n_353;
input n_351;
input n_367;
input n_452;
input n_397;
input n_493;
input n_111;
input n_525;
input n_483;
input n_544;
input n_155;
input n_552;
input n_547;
input n_43;
input n_116;
input n_22;
input n_467;
input n_564;
input n_423;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_139;
input n_38;
input n_105;
input n_280;
input n_590;
input n_4;
input n_378;
input n_551;
input n_17;
input n_581;
input n_382;
input n_554;
input n_254;
input n_33;
input n_23;
input n_583;
input n_302;
input n_265;
input n_526;
input n_293;
input n_372;
input n_443;
input n_244;
input n_47;
input n_173;
input n_198;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_8;
input n_321;
input n_292;
input n_100;
input n_455;
input n_417;
input n_212;
input n_385;
input n_498;
input n_516;
input n_507;
input n_119;
input n_497;
input n_559;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_508;
input n_506;
input n_2;
input n_6;
input n_509;
input n_568;
input n_39;
input n_147;
input n_373;
input n_67;
input n_307;
input n_439;
input n_87;
input n_150;
input n_530;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_375;
input n_301;
input n_576;
input n_68;
input n_93;
input n_186;
input n_537;
input n_134;
input n_191;
input n_587;
input n_51;
input n_63;
input n_492;
input n_563;
input n_171;
input n_153;
input n_524;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_548;
input n_543;
input n_260;
input n_298;
input n_320;
input n_518;
input n_505;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_406;
input n_519;
input n_470;
input n_325;
input n_449;
input n_132;
input n_90;
input n_546;
input n_101;
input n_281;
input n_240;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_31;
input n_456;
input n_13;
input n_371;
input n_481;
input n_535;
input n_152;
input n_540;
input n_317;
input n_9;
input n_323;
input n_569;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_370;
input n_167;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_297;
input n_156;
input n_5;
input n_225;
input n_377;
input n_484;
input n_219;
input n_442;
input n_157;
input n_131;
input n_192;
input n_223;
input n_392;
input n_158;
input n_138;
input n_264;
input n_109;
input n_472;
input n_454;
input n_387;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_347;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_215;
input n_350;
input n_196;
input n_459;
input n_211;
input n_218;
input n_400;
input n_181;
input n_436;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_386;
input n_578;
input n_287;
input n_344;
input n_555;
input n_473;
input n_422;
input n_475;
input n_72;
input n_104;
input n_41;
input n_415;
input n_56;
input n_141;
input n_485;
input n_496;
input n_355;
input n_486;
input n_15;
input n_336;
input n_584;
input n_591;
input n_145;
input n_48;
input n_521;
input n_50;
input n_337;
input n_430;
input n_313;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_168;
input n_395;
input n_164;
input n_432;
input n_553;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_369;
input n_296;
input n_241;
input n_357;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_468;
input n_499;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_363;
input n_402;
input n_413;
input n_197;
input n_107;
input n_573;
input n_69;
input n_236;
input n_388;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_309;
input n_30;
input n_512;
input n_14;
input n_84;
input n_462;
input n_130;
input n_322;
input n_567;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_458;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_471;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_383;
input n_474;
input n_112;
input n_542;
input n_85;
input n_463;
input n_488;
input n_502;
input n_239;
input n_466;
input n_420;
input n_489;
input n_55;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_586;
input n_465;
input n_76;
input n_358;
input n_362;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_440;
input n_478;
input n_545;
input n_441;
input n_450;
input n_312;
input n_476;
input n_429;
input n_534;
input n_345;
input n_210;
input n_494;
input n_365;
input n_91;
input n_176;
input n_557;
input n_182;
input n_143;
input n_83;
input n_354;
input n_575;
input n_480;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_180;
input n_560;
input n_340;
input n_207;
input n_561;
input n_37;
input n_346;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_16;
input n_0;
input n_58;
input n_405;
input n_18;
input n_359;
input n_490;
input n_117;
input n_326;
input n_233;
input n_404;
input n_205;
input n_366;
input n_572;
input n_113;
input n_246;
input n_179;
input n_125;
input n_410;
input n_558;
input n_269;
input n_529;
input n_128;
input n_285;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_409;
input n_589;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_435;
input n_159;
input n_334;
input n_541;
input n_391;
input n_434;
input n_539;
input n_175;
input n_538;
input n_262;
input n_238;
input n_99;
input n_411;
input n_414;
input n_319;
input n_364;
input n_20;
input n_536;
input n_531;
input n_121;
input n_242;
input n_360;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_438;
input n_115;
input n_324;
input n_416;
input n_199;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_424;
input n_7;
input n_256;
input n_305;
input n_533;
input n_52;
input n_278;
input n_110;

output n_2933;

wire n_924;
wire n_1263;
wire n_1378;
wire n_977;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_785;
wire n_2617;
wire n_2200;
wire n_1161;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_1780;
wire n_1488;
wire n_667;
wire n_2899;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_2395;
wire n_880;
wire n_1007;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1198;
wire n_1360;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_2391;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_1695;
wire n_688;
wire n_2487;
wire n_1353;
wire n_800;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_2001;
wire n_1494;
wire n_625;
wire n_1462;
wire n_854;
wire n_2069;
wire n_1799;
wire n_2396;
wire n_1580;
wire n_674;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_2244;
wire n_933;
wire n_2257;
wire n_1152;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_1118;
wire n_755;
wire n_1686;
wire n_947;
wire n_1285;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2076;
wire n_2031;
wire n_2482;
wire n_2677;
wire n_1230;
wire n_668;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_2770;
wire n_1124;
wire n_2127;
wire n_1818;
wire n_1576;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2142;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_1016;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_2761;
wire n_731;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_2306;
wire n_920;
wire n_2515;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_2715;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_976;
wire n_1449;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_1146;
wire n_882;
wire n_2384;
wire n_1036;
wire n_1749;
wire n_1097;
wire n_696;
wire n_897;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_926;
wire n_2180;
wire n_2249;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_1070;
wire n_1547;
wire n_777;
wire n_2089;
wire n_1030;
wire n_2470;
wire n_1755;
wire n_1561;
wire n_1165;
wire n_1267;
wire n_1071;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_1600;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_1880;
wire n_888;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_2118;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_2932;
wire n_2753;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_889;
wire n_2358;
wire n_973;
wire n_1700;
wire n_2833;
wire n_1585;
wire n_2684;
wire n_2712;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_2855;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_2370;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_736;
wire n_892;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_2258;
wire n_748;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_793;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_1527;
wire n_2042;
wire n_1882;
wire n_884;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_647;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_832;
wire n_857;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_2154;
wire n_1951;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_2798;
wire n_2331;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_2808;
wire n_1276;
wire n_702;
wire n_2548;
wire n_1412;
wire n_822;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_728;
wire n_1162;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_2698;
wire n_809;
wire n_1711;
wire n_870;
wire n_599;
wire n_1891;
wire n_1662;
wire n_931;
wire n_1481;
wire n_2626;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_1876;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_1477;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_1189;
wire n_2690;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_2621;
wire n_851;
wire n_615;
wire n_1759;
wire n_843;
wire n_2177;
wire n_1788;
wire n_2491;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_649;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_1734;
wire n_744;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_1767;
wire n_2913;
wire n_2336;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_677;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_604;
wire n_2007;
wire n_949;
wire n_2539;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_1380;
wire n_624;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_1500;
wire n_1090;
wire n_2796;
wire n_757;
wire n_2342;
wire n_633;
wire n_2856;
wire n_1832;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_906;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_2846;
wire n_724;
wire n_2084;
wire n_1781;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_959;
wire n_2459;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_1017;
wire n_2481;
wire n_2171;
wire n_978;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2339;
wire n_1045;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2473;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_1033;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_742;
wire n_2029;
wire n_750;
wire n_995;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_1989;
wire n_2359;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_662;
wire n_2312;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_2812;
wire n_2048;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_2729;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_2909;
wire n_2111;
wire n_1724;
wire n_2521;
wire n_1237;
wire n_700;
wire n_1420;
wire n_1132;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_2681;
wire n_1562;
wire n_834;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_874;
wire n_2464;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_1846;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_860;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_729;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_2645;
wire n_2467;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1044;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_1552;
wire n_2508;
wire n_602;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_2088;
wire n_824;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_1684;
wire n_921;
wire n_2658;
wire n_1717;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_1821;
wire n_2929;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_1229;
wire n_1437;
wire n_701;
wire n_1023;
wire n_2075;
wire n_645;
wire n_803;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_2216;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_2647;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_1519;
wire n_950;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_1346;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_2465;
wire n_2824;
wire n_2650;
wire n_912;
wire n_968;
wire n_619;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_2333;
wire n_885;
wire n_2916;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_1305;
wire n_873;
wire n_1826;
wire n_1112;
wire n_2304;
wire n_1283;
wire n_1644;
wire n_762;
wire n_2334;
wire n_2637;
wire n_690;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_2289;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_1966;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_1312;
wire n_1439;
wire n_804;
wire n_2827;
wire n_1688;
wire n_945;
wire n_1504;
wire n_943;
wire n_992;
wire n_1932;
wire n_2755;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_883;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_2364;
wire n_2533;
wire n_618;
wire n_896;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_2291;
wire n_2596;
wire n_1636;
wire n_894;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_2318;
wire n_833;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2707;
wire n_2751;
wire n_2793;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_2758;
wire n_1458;
wire n_669;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_2600;
wire n_849;
wire n_2795;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2002;
wire n_2282;
wire n_2800;
wire n_2371;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_2444;
wire n_2068;
wire n_875;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_749;
wire n_1895;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_1401;
wire n_969;
wire n_2492;
wire n_1998;
wire n_1105;
wire n_1019;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_778;
wire n_1122;
wire n_2608;
wire n_2657;
wire n_770;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_2097;
wire n_1834;
wire n_2313;
wire n_2542;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_876;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_726;
wire n_982;
wire n_2575;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_1584;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_1125;
wire n_2547;
wire n_708;
wire n_1812;
wire n_735;
wire n_2501;
wire n_1915;
wire n_1109;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_2665;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_1067;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_2003;
wire n_1457;
wire n_766;
wire n_2692;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_2245;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_1011;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_827;
wire n_1703;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_676;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_855;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_620;
wire n_643;
wire n_2363;
wire n_2430;
wire n_916;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_2332;
wire n_1235;
wire n_703;
wire n_1115;
wire n_698;
wire n_980;
wire n_2433;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2601;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_823;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_2773;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_1120;
wire n_719;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_909;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_2884;
wire n_1268;
wire n_825;
wire n_2819;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_737;
wire n_986;
wire n_2315;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_792;
wire n_1429;
wire n_756;
wire n_1238;
wire n_2448;
wire n_812;
wire n_2104;
wire n_2748;
wire n_2057;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_2889;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_1675;
wire n_1924;
wire n_2573;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_1221;
wire n_2345;
wire n_654;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_1641;
wire n_1361;
wire n_2382;
wire n_1707;
wire n_853;
wire n_2317;
wire n_751;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_786;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_930;
wire n_1873;
wire n_1411;
wire n_1962;
wire n_622;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_1567;
wire n_682;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_922;
wire n_816;
wire n_1648;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_631;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_2360;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_1842;
wire n_871;
wire n_2442;
wire n_685;
wire n_598;
wire n_1367;
wire n_608;
wire n_928;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_2834;
wire n_2531;
wire n_1589;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_2208;
wire n_1404;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_2321;
wire n_1226;
wire n_1277;
wire n_722;
wire n_2591;
wire n_2146;
wire n_844;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1601;
wire n_1028;
wire n_781;
wire n_1546;
wire n_595;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_1627;
wire n_2918;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_1739;
wire n_616;
wire n_2278;
wire n_2594;
wire n_2394;
wire n_1914;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_1654;
wire n_2569;
wire n_2349;
wire n_1103;
wire n_648;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_712;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_2013;
wire n_927;
wire n_1089;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_1693;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g594 ( 
.A(n_334),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_132),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_505),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_384),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_535),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_99),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_367),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_565),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_266),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_322),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_152),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_13),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_208),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_393),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_99),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_382),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_153),
.Y(n_610)
);

BUFx2_ASAP7_75t_L g611 ( 
.A(n_591),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_341),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_224),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_552),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_313),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_82),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_43),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_214),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_165),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_456),
.Y(n_620)
);

CKINVDCx14_ASAP7_75t_R g621 ( 
.A(n_589),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_555),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_432),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_68),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_113),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_119),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_345),
.Y(n_628)
);

BUFx5_ASAP7_75t_L g629 ( 
.A(n_199),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_98),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_175),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_269),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_527),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_199),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_198),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_279),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_539),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_456),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_386),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_326),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_521),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_217),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_359),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_188),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_507),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_592),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_396),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_60),
.Y(n_648)
);

BUFx3_ASAP7_75t_L g649 ( 
.A(n_390),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_564),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_281),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_161),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_577),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_416),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_230),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_141),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_556),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_582),
.Y(n_658)
);

CKINVDCx5p33_ASAP7_75t_R g659 ( 
.A(n_347),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_204),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_141),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_440),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_201),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_451),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_479),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_106),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_230),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_527),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_435),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_157),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_253),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_450),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_101),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_536),
.Y(n_674)
);

BUFx10_ASAP7_75t_L g675 ( 
.A(n_512),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_41),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_441),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_370),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_122),
.Y(n_679)
);

CKINVDCx16_ASAP7_75t_R g680 ( 
.A(n_544),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_280),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_119),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_313),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_452),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_253),
.Y(n_685)
);

BUFx8_ASAP7_75t_SL g686 ( 
.A(n_528),
.Y(n_686)
);

BUFx5_ASAP7_75t_L g687 ( 
.A(n_29),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_492),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_391),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_70),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_264),
.Y(n_691)
);

INVx1_ASAP7_75t_SL g692 ( 
.A(n_254),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_495),
.Y(n_693)
);

BUFx2_ASAP7_75t_L g694 ( 
.A(n_41),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_272),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_306),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_90),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_533),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_39),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_110),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_383),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_461),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_194),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_59),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_568),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_553),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_91),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_404),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_392),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_261),
.Y(n_710)
);

BUFx3_ASAP7_75t_L g711 ( 
.A(n_399),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_492),
.Y(n_712)
);

BUFx10_ASAP7_75t_L g713 ( 
.A(n_537),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_12),
.Y(n_714)
);

CKINVDCx20_ASAP7_75t_R g715 ( 
.A(n_448),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_593),
.Y(n_716)
);

CKINVDCx20_ASAP7_75t_R g717 ( 
.A(n_385),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_411),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_586),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_523),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_60),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_556),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_368),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_443),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_346),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_376),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_188),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_374),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_265),
.Y(n_729)
);

CKINVDCx20_ASAP7_75t_R g730 ( 
.A(n_551),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_559),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_101),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_581),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_475),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_350),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_167),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_512),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_465),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_86),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_268),
.Y(n_740)
);

INVx1_ASAP7_75t_SL g741 ( 
.A(n_558),
.Y(n_741)
);

BUFx3_ASAP7_75t_L g742 ( 
.A(n_182),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_337),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_378),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_415),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_583),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_160),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_439),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_516),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_391),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_31),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_70),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_501),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_228),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_424),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_126),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_359),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_422),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_376),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_525),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_177),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_315),
.Y(n_762)
);

INVxp67_ASAP7_75t_L g763 ( 
.A(n_56),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_249),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_439),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_242),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_147),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_531),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_429),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_229),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_314),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_559),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_22),
.Y(n_773)
);

CKINVDCx20_ASAP7_75t_R g774 ( 
.A(n_346),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_580),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_111),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_451),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_270),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_357),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_11),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_277),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_409),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_546),
.Y(n_783)
);

INVx1_ASAP7_75t_SL g784 ( 
.A(n_548),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_57),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_1),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_195),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_524),
.Y(n_788)
);

BUFx3_ASAP7_75t_L g789 ( 
.A(n_550),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_315),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_311),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_62),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_53),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_38),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_197),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_348),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_365),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_126),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_326),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_560),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_163),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_312),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_96),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_361),
.Y(n_804)
);

INVx3_ASAP7_75t_L g805 ( 
.A(n_153),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_557),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_337),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_382),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_368),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_18),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_534),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_214),
.Y(n_812)
);

INVx1_ASAP7_75t_SL g813 ( 
.A(n_203),
.Y(n_813)
);

BUFx2_ASAP7_75t_L g814 ( 
.A(n_561),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_256),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_262),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_163),
.Y(n_817)
);

CKINVDCx5p33_ASAP7_75t_R g818 ( 
.A(n_268),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_579),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_425),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_454),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_281),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_587),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_535),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_478),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_302),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_520),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_526),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_338),
.Y(n_829)
);

BUFx2_ASAP7_75t_L g830 ( 
.A(n_562),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_169),
.Y(n_831)
);

CKINVDCx5p33_ASAP7_75t_R g832 ( 
.A(n_555),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_329),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_365),
.Y(n_834)
);

CKINVDCx5p33_ASAP7_75t_R g835 ( 
.A(n_145),
.Y(n_835)
);

INVx1_ASAP7_75t_SL g836 ( 
.A(n_4),
.Y(n_836)
);

INVxp67_ASAP7_75t_SL g837 ( 
.A(n_563),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_90),
.Y(n_838)
);

BUFx10_ASAP7_75t_L g839 ( 
.A(n_98),
.Y(n_839)
);

CKINVDCx14_ASAP7_75t_R g840 ( 
.A(n_423),
.Y(n_840)
);

INVx2_ASAP7_75t_SL g841 ( 
.A(n_26),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_218),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_134),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_121),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_345),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_165),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_481),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_167),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_11),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_538),
.Y(n_850)
);

BUFx10_ASAP7_75t_L g851 ( 
.A(n_574),
.Y(n_851)
);

INVx1_ASAP7_75t_SL g852 ( 
.A(n_18),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_159),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_263),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_0),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_108),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_543),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_329),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_300),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_404),
.Y(n_860)
);

BUFx8_ASAP7_75t_SL g861 ( 
.A(n_157),
.Y(n_861)
);

CKINVDCx16_ASAP7_75t_R g862 ( 
.A(n_526),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_220),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_274),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_107),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_283),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_571),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_181),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_300),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_409),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_388),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_578),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_78),
.Y(n_873)
);

CKINVDCx5p33_ASAP7_75t_R g874 ( 
.A(n_530),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_560),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_78),
.Y(n_876)
);

BUFx8_ASAP7_75t_SL g877 ( 
.A(n_107),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_532),
.Y(n_878)
);

INVx1_ASAP7_75t_SL g879 ( 
.A(n_48),
.Y(n_879)
);

CKINVDCx14_ASAP7_75t_R g880 ( 
.A(n_455),
.Y(n_880)
);

BUFx2_ASAP7_75t_SL g881 ( 
.A(n_241),
.Y(n_881)
);

BUFx10_ASAP7_75t_L g882 ( 
.A(n_554),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_255),
.Y(n_883)
);

BUFx5_ASAP7_75t_L g884 ( 
.A(n_144),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_575),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_418),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_73),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_212),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_171),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_453),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_390),
.Y(n_891)
);

CKINVDCx20_ASAP7_75t_R g892 ( 
.A(n_518),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_549),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_191),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_135),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_534),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_542),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_244),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_10),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_433),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_108),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_352),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_244),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_457),
.Y(n_904)
);

CKINVDCx20_ASAP7_75t_R g905 ( 
.A(n_304),
.Y(n_905)
);

CKINVDCx20_ASAP7_75t_R g906 ( 
.A(n_474),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_187),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_541),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_32),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_490),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_111),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_106),
.Y(n_912)
);

CKINVDCx16_ASAP7_75t_R g913 ( 
.A(n_302),
.Y(n_913)
);

CKINVDCx5p33_ASAP7_75t_R g914 ( 
.A(n_434),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_570),
.Y(n_915)
);

CKINVDCx16_ASAP7_75t_R g916 ( 
.A(n_289),
.Y(n_916)
);

CKINVDCx5p33_ASAP7_75t_R g917 ( 
.A(n_335),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_474),
.Y(n_918)
);

CKINVDCx20_ASAP7_75t_R g919 ( 
.A(n_425),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_547),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_431),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_482),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_371),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_271),
.Y(n_924)
);

BUFx2_ASAP7_75t_L g925 ( 
.A(n_354),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_291),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_58),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_257),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_269),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_117),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_242),
.Y(n_931)
);

CKINVDCx5p33_ASAP7_75t_R g932 ( 
.A(n_532),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_259),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_573),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_533),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_159),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_355),
.Y(n_937)
);

CKINVDCx5p33_ASAP7_75t_R g938 ( 
.A(n_55),
.Y(n_938)
);

INVx2_ASAP7_75t_SL g939 ( 
.A(n_572),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_566),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_58),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_364),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_104),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_47),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_71),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_459),
.B(n_286),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_481),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_388),
.Y(n_948)
);

CKINVDCx20_ASAP7_75t_R g949 ( 
.A(n_272),
.Y(n_949)
);

CKINVDCx20_ASAP7_75t_R g950 ( 
.A(n_348),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_432),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_493),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_364),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_590),
.Y(n_954)
);

CKINVDCx5p33_ASAP7_75t_R g955 ( 
.A(n_344),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_545),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_453),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_468),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_112),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_30),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_50),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_386),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_158),
.Y(n_963)
);

CKINVDCx16_ASAP7_75t_R g964 ( 
.A(n_110),
.Y(n_964)
);

BUFx6f_ASAP7_75t_L g965 ( 
.A(n_515),
.Y(n_965)
);

CKINVDCx5p33_ASAP7_75t_R g966 ( 
.A(n_246),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_445),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_506),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_428),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_562),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_333),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_31),
.Y(n_972)
);

CKINVDCx20_ASAP7_75t_R g973 ( 
.A(n_92),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_234),
.Y(n_974)
);

CKINVDCx16_ASAP7_75t_R g975 ( 
.A(n_440),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_252),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_437),
.Y(n_977)
);

CKINVDCx20_ASAP7_75t_R g978 ( 
.A(n_529),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_540),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_207),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_172),
.Y(n_981)
);

BUFx3_ASAP7_75t_L g982 ( 
.A(n_360),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_236),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_211),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_238),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_198),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_331),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_485),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_470),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_361),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_554),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_406),
.Y(n_992)
);

CKINVDCx5p33_ASAP7_75t_R g993 ( 
.A(n_518),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_263),
.Y(n_994)
);

BUFx5_ASAP7_75t_L g995 ( 
.A(n_501),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_170),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_381),
.Y(n_997)
);

INVx1_ASAP7_75t_SL g998 ( 
.A(n_220),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_517),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_422),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_548),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_584),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_341),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_279),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_113),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_338),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_122),
.Y(n_1007)
);

CKINVDCx20_ASAP7_75t_R g1008 ( 
.A(n_189),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_389),
.Y(n_1009)
);

BUFx10_ASAP7_75t_L g1010 ( 
.A(n_349),
.Y(n_1010)
);

INVx1_ASAP7_75t_SL g1011 ( 
.A(n_354),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_411),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_27),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_576),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_83),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_109),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_340),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_470),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_135),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_56),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_486),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_234),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_541),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_266),
.Y(n_1024)
);

BUFx10_ASAP7_75t_L g1025 ( 
.A(n_208),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_40),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_429),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_384),
.Y(n_1028)
);

BUFx3_ASAP7_75t_L g1029 ( 
.A(n_585),
.Y(n_1029)
);

BUFx10_ASAP7_75t_L g1030 ( 
.A(n_133),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_298),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_174),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_686),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_629),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_629),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_629),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_629),
.Y(n_1037)
);

BUFx2_ASAP7_75t_L g1038 ( 
.A(n_694),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_621),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_629),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_629),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_872),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_861),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_629),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_629),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_629),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_687),
.Y(n_1047)
);

CKINVDCx16_ASAP7_75t_R g1048 ( 
.A(n_680),
.Y(n_1048)
);

HB1xp67_ASAP7_75t_L g1049 ( 
.A(n_694),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_687),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_687),
.Y(n_1051)
);

BUFx8_ASAP7_75t_SL g1052 ( 
.A(n_877),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_687),
.Y(n_1053)
);

INVxp67_ASAP7_75t_SL g1054 ( 
.A(n_611),
.Y(n_1054)
);

NOR2xp67_ASAP7_75t_L g1055 ( 
.A(n_805),
.B(n_0),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_653),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_687),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_687),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_687),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_687),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_814),
.Y(n_1061)
);

INVxp67_ASAP7_75t_SL g1062 ( 
.A(n_611),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_687),
.Y(n_1063)
);

INVx1_ASAP7_75t_SL g1064 ( 
.A(n_814),
.Y(n_1064)
);

CKINVDCx16_ASAP7_75t_R g1065 ( 
.A(n_680),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_884),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_840),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_884),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_884),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_884),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_884),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_884),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_884),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_830),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_658),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_705),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_884),
.Y(n_1077)
);

INVx3_ASAP7_75t_L g1078 ( 
.A(n_628),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_884),
.Y(n_1079)
);

INVxp67_ASAP7_75t_L g1080 ( 
.A(n_830),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_934),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_872),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_995),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_995),
.Y(n_1084)
);

INVxp33_ASAP7_75t_SL g1085 ( 
.A(n_793),
.Y(n_1085)
);

CKINVDCx20_ASAP7_75t_R g1086 ( 
.A(n_880),
.Y(n_1086)
);

INVxp33_ASAP7_75t_SL g1087 ( 
.A(n_803),
.Y(n_1087)
);

NOR2xp67_ASAP7_75t_L g1088 ( 
.A(n_805),
.B(n_1),
.Y(n_1088)
);

INVx1_ASAP7_75t_L g1089 ( 
.A(n_995),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_940),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_849),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_995),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_954),
.Y(n_1093)
);

CKINVDCx20_ASAP7_75t_R g1094 ( 
.A(n_1002),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_995),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_995),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_995),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_1014),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_995),
.Y(n_1099)
);

HB1xp67_ASAP7_75t_L g1100 ( 
.A(n_849),
.Y(n_1100)
);

CKINVDCx14_ASAP7_75t_R g1101 ( 
.A(n_925),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1029),
.Y(n_1102)
);

INVxp67_ASAP7_75t_SL g1103 ( 
.A(n_805),
.Y(n_1103)
);

INVxp67_ASAP7_75t_SL g1104 ( 
.A(n_805),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_596),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_995),
.Y(n_1106)
);

INVxp33_ASAP7_75t_L g1107 ( 
.A(n_925),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_SL g1108 ( 
.A1(n_1101),
.A2(n_602),
.B1(n_622),
.B2(n_600),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1034),
.Y(n_1109)
);

CKINVDCx6p67_ASAP7_75t_R g1110 ( 
.A(n_1039),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1078),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1103),
.B(n_1104),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1078),
.Y(n_1113)
);

AND2x6_ASAP7_75t_L g1114 ( 
.A(n_1035),
.B(n_946),
.Y(n_1114)
);

BUFx6f_ASAP7_75t_L g1115 ( 
.A(n_1078),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1082),
.B(n_946),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1034),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_1105),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_1056),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1035),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1036),
.A2(n_819),
.B(n_719),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_1075),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_1066),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1082),
.B(n_628),
.Y(n_1124)
);

INVx2_ASAP7_75t_L g1125 ( 
.A(n_1068),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1082),
.B(n_628),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1082),
.B(n_628),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_1048),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1082),
.B(n_628),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1102),
.B(n_628),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1042),
.B(n_1054),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1036),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1037),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1062),
.B(n_939),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_1069),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_1096),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1037),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_1040),
.Y(n_1138)
);

AOI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_1085),
.A2(n_895),
.B1(n_913),
.B2(n_862),
.Y(n_1139)
);

AOI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1087),
.A2(n_895),
.B1(n_913),
.B2(n_862),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1065),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1102),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1040),
.Y(n_1143)
);

BUFx8_ASAP7_75t_L g1144 ( 
.A(n_1038),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1041),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1041),
.Y(n_1146)
);

AND2x6_ASAP7_75t_L g1147 ( 
.A(n_1044),
.B(n_719),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1044),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1045),
.Y(n_1149)
);

XNOR2xp5_ASAP7_75t_L g1150 ( 
.A(n_1064),
.B(n_650),
.Y(n_1150)
);

INVx3_ASAP7_75t_L g1151 ( 
.A(n_1045),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1055),
.B(n_1088),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_1046),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1102),
.B(n_631),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1047),
.A2(n_646),
.B(n_627),
.Y(n_1155)
);

INVx2_ASAP7_75t_L g1156 ( 
.A(n_1047),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_1050),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1102),
.B(n_631),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_1102),
.B(n_631),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1050),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1051),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1051),
.Y(n_1162)
);

BUFx6f_ASAP7_75t_L g1163 ( 
.A(n_1053),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1053),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1057),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_1057),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1076),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1058),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1132),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1132),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_1110),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1133),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1133),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_1110),
.Y(n_1174)
);

CKINVDCx20_ASAP7_75t_R g1175 ( 
.A(n_1110),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_1119),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1115),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_1122),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1137),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1137),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_1167),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1118),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_1150),
.Y(n_1183)
);

CKINVDCx20_ASAP7_75t_R g1184 ( 
.A(n_1128),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_1150),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1161),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_1144),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_1144),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1161),
.Y(n_1189)
);

HB1xp67_ASAP7_75t_L g1190 ( 
.A(n_1141),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_1144),
.Y(n_1191)
);

CKINVDCx16_ASAP7_75t_R g1192 ( 
.A(n_1108),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_1144),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1131),
.B(n_1042),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1165),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1108),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1165),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_1142),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1131),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_1139),
.Y(n_1200)
);

CKINVDCx20_ASAP7_75t_R g1201 ( 
.A(n_1139),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_1140),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1140),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1152),
.B(n_1112),
.Y(n_1204)
);

CKINVDCx16_ASAP7_75t_R g1205 ( 
.A(n_1152),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1134),
.Y(n_1206)
);

CKINVDCx20_ASAP7_75t_R g1207 ( 
.A(n_1112),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1109),
.Y(n_1208)
);

CKINVDCx20_ASAP7_75t_R g1209 ( 
.A(n_1116),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_R g1210 ( 
.A(n_1116),
.B(n_1081),
.Y(n_1210)
);

AND2x4_ASAP7_75t_L g1211 ( 
.A(n_1152),
.B(n_1029),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1109),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_1152),
.Y(n_1213)
);

CKINVDCx16_ASAP7_75t_R g1214 ( 
.A(n_1142),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_1142),
.Y(n_1215)
);

NOR2xp67_ASAP7_75t_L g1216 ( 
.A(n_1111),
.B(n_1098),
.Y(n_1216)
);

INVxp33_ASAP7_75t_SL g1217 ( 
.A(n_1124),
.Y(n_1217)
);

INVxp67_ASAP7_75t_L g1218 ( 
.A(n_1124),
.Y(n_1218)
);

CKINVDCx20_ASAP7_75t_R g1219 ( 
.A(n_1126),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1114),
.B(n_1093),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1147),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1147),
.Y(n_1222)
);

NOR2xp33_ASAP7_75t_R g1223 ( 
.A(n_1151),
.B(n_1090),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1147),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1147),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1147),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_1181),
.Y(n_1227)
);

NAND2x1p5_ASAP7_75t_L g1228 ( 
.A(n_1198),
.B(n_1155),
.Y(n_1228)
);

INVx4_ASAP7_75t_L g1229 ( 
.A(n_1177),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1209),
.Y(n_1230)
);

INVx4_ASAP7_75t_L g1231 ( 
.A(n_1177),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_SL g1232 ( 
.A(n_1213),
.B(n_1094),
.Y(n_1232)
);

AND2x2_ASAP7_75t_SL g1233 ( 
.A(n_1192),
.B(n_968),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_SL g1234 ( 
.A(n_1206),
.B(n_939),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1169),
.Y(n_1235)
);

INVxp33_ASAP7_75t_L g1236 ( 
.A(n_1194),
.Y(n_1236)
);

NOR2xp33_ASAP7_75t_L g1237 ( 
.A(n_1206),
.B(n_1067),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1204),
.B(n_1218),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_1207),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_L g1240 ( 
.A(n_1199),
.B(n_1086),
.Y(n_1240)
);

INVx1_ASAP7_75t_SL g1241 ( 
.A(n_1184),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1170),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1213),
.B(n_733),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_1176),
.Y(n_1244)
);

BUFx8_ASAP7_75t_SL g1245 ( 
.A(n_1175),
.Y(n_1245)
);

AND2x4_ASAP7_75t_L g1246 ( 
.A(n_1204),
.B(n_627),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1198),
.Y(n_1247)
);

INVxp67_ASAP7_75t_L g1248 ( 
.A(n_1190),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1217),
.B(n_1114),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_SL g1250 ( 
.A(n_1205),
.B(n_851),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1194),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1172),
.Y(n_1252)
);

BUFx3_ASAP7_75t_L g1253 ( 
.A(n_1219),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_SL g1254 ( 
.A(n_1223),
.B(n_851),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1173),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1182),
.Y(n_1256)
);

BUFx6f_ASAP7_75t_L g1257 ( 
.A(n_1177),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1179),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1180),
.B(n_1114),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1186),
.A2(n_1114),
.B1(n_1153),
.B2(n_1151),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1214),
.B(n_1107),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_1189),
.B(n_1033),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_L g1263 ( 
.A(n_1195),
.B(n_1043),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1208),
.Y(n_1264)
);

OR2x2_ASAP7_75t_L g1265 ( 
.A(n_1183),
.B(n_1038),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_L g1266 ( 
.A(n_1197),
.B(n_1074),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1208),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1210),
.B(n_851),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1211),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1211),
.B(n_1114),
.Y(n_1270)
);

NAND2x1p5_ASAP7_75t_L g1271 ( 
.A(n_1177),
.B(n_1155),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1212),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1211),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1177),
.Y(n_1274)
);

OR2x2_ASAP7_75t_L g1275 ( 
.A(n_1185),
.B(n_1049),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1212),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_SL g1277 ( 
.A(n_1216),
.B(n_851),
.Y(n_1277)
);

AND2x6_ASAP7_75t_L g1278 ( 
.A(n_1220),
.B(n_646),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1215),
.B(n_1080),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_R g1280 ( 
.A(n_1176),
.B(n_916),
.Y(n_1280)
);

HB1xp67_ASAP7_75t_L g1281 ( 
.A(n_1202),
.Y(n_1281)
);

INVx3_ASAP7_75t_L g1282 ( 
.A(n_1221),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1215),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1226),
.B(n_1114),
.Y(n_1284)
);

INVx2_ASAP7_75t_SL g1285 ( 
.A(n_1221),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1222),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1222),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1178),
.Y(n_1288)
);

INVx4_ASAP7_75t_L g1289 ( 
.A(n_1224),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_L g1290 ( 
.A(n_1224),
.B(n_1114),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1171),
.Y(n_1291)
);

INVx2_ASAP7_75t_L g1292 ( 
.A(n_1225),
.Y(n_1292)
);

INVx3_ASAP7_75t_L g1293 ( 
.A(n_1225),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1202),
.B(n_1061),
.Y(n_1294)
);

BUFx3_ASAP7_75t_L g1295 ( 
.A(n_1226),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1200),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1201),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1196),
.B(n_1114),
.Y(n_1298)
);

INVx4_ASAP7_75t_L g1299 ( 
.A(n_1187),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1188),
.B(n_1114),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1191),
.B(n_916),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1203),
.Y(n_1302)
);

AND2x4_ASAP7_75t_L g1303 ( 
.A(n_1193),
.B(n_716),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1171),
.B(n_1091),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1238),
.B(n_1151),
.Y(n_1305)
);

INVx2_ASAP7_75t_SL g1306 ( 
.A(n_1253),
.Y(n_1306)
);

INVxp33_ASAP7_75t_L g1307 ( 
.A(n_1261),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1235),
.Y(n_1308)
);

BUFx6f_ASAP7_75t_L g1309 ( 
.A(n_1247),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_SL g1310 ( 
.A(n_1298),
.B(n_1283),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1270),
.A2(n_1162),
.B(n_1143),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_SL g1312 ( 
.A(n_1283),
.B(n_1151),
.Y(n_1312)
);

BUFx6f_ASAP7_75t_SL g1313 ( 
.A(n_1299),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1246),
.B(n_1153),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1242),
.Y(n_1315)
);

AOI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1246),
.A2(n_1273),
.B1(n_1269),
.B2(n_1251),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1253),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1252),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_1255),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1246),
.B(n_1153),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1264),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1258),
.Y(n_1322)
);

INVx5_ASAP7_75t_L g1323 ( 
.A(n_1257),
.Y(n_1323)
);

NAND2x1p5_ASAP7_75t_L g1324 ( 
.A(n_1295),
.B(n_1155),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1264),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1251),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_1288),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1236),
.B(n_964),
.Y(n_1328)
);

BUFx6f_ASAP7_75t_L g1329 ( 
.A(n_1247),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1285),
.B(n_1153),
.Y(n_1330)
);

INVx2_ASAP7_75t_L g1331 ( 
.A(n_1267),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1282),
.A2(n_746),
.B1(n_775),
.B2(n_716),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1267),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1294),
.B(n_1100),
.C(n_1174),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1236),
.B(n_964),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_SL g1336 ( 
.A(n_1249),
.B(n_1160),
.Y(n_1336)
);

NAND2xp5_ASAP7_75t_SL g1337 ( 
.A(n_1287),
.B(n_1160),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1279),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1285),
.B(n_1160),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1279),
.B(n_1174),
.Y(n_1340)
);

NOR2xp33_ASAP7_75t_L g1341 ( 
.A(n_1266),
.B(n_975),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1256),
.B(n_975),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1282),
.B(n_1160),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1272),
.Y(n_1344)
);

INVx2_ASAP7_75t_L g1345 ( 
.A(n_1272),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_SL g1346 ( 
.A(n_1287),
.B(n_1168),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1282),
.B(n_1168),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1293),
.B(n_1168),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1276),
.Y(n_1349)
);

HB1xp67_ASAP7_75t_L g1350 ( 
.A(n_1230),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1248),
.B(n_702),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1293),
.B(n_1168),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1230),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_SL g1354 ( 
.A(n_1280),
.B(n_746),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1247),
.Y(n_1355)
);

OR2x2_ASAP7_75t_L g1356 ( 
.A(n_1265),
.B(n_692),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1247),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1232),
.B(n_715),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1247),
.B(n_837),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1237),
.B(n_968),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1257),
.Y(n_1361)
);

AND2x2_ASAP7_75t_SL g1362 ( 
.A(n_1233),
.B(n_775),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1233),
.A2(n_1027),
.B1(n_996),
.B2(n_742),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_SL g1364 ( 
.A(n_1292),
.B(n_1163),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1257),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1257),
.Y(n_1366)
);

NAND3xp33_ASAP7_75t_L g1367 ( 
.A(n_1240),
.B(n_1027),
.C(n_996),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1257),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1293),
.B(n_1295),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1286),
.Y(n_1370)
);

NAND2xp33_ASAP7_75t_SL g1371 ( 
.A(n_1227),
.B(n_717),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1271),
.Y(n_1372)
);

AOI221xp5_ASAP7_75t_L g1373 ( 
.A1(n_1234),
.A2(n_741),
.B1(n_759),
.B2(n_728),
.C(n_709),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1292),
.B(n_1138),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1229),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1227),
.Y(n_1376)
);

OR2x2_ASAP7_75t_L g1377 ( 
.A(n_1265),
.B(n_784),
.Y(n_1377)
);

NOR3xp33_ASAP7_75t_L g1378 ( 
.A(n_1301),
.B(n_763),
.C(n_806),
.Y(n_1378)
);

INVx2_ASAP7_75t_SL g1379 ( 
.A(n_1239),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_L g1380 ( 
.A(n_1289),
.B(n_1138),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1289),
.B(n_1138),
.Y(n_1381)
);

NOR2xp33_ASAP7_75t_L g1382 ( 
.A(n_1243),
.B(n_1250),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_1288),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1289),
.B(n_1143),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1239),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1259),
.B(n_1163),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1271),
.Y(n_1387)
);

INVx2_ASAP7_75t_L g1388 ( 
.A(n_1228),
.Y(n_1388)
);

O2A1O1Ixp33_ASAP7_75t_L g1389 ( 
.A1(n_1300),
.A2(n_1127),
.B(n_1129),
.C(n_1126),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1271),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1228),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1228),
.Y(n_1392)
);

AOI22xp5_ASAP7_75t_L g1393 ( 
.A1(n_1278),
.A2(n_1125),
.B1(n_1136),
.B2(n_1135),
.Y(n_1393)
);

A2O1A1Ixp33_ASAP7_75t_L g1394 ( 
.A1(n_1234),
.A2(n_867),
.B(n_885),
.C(n_823),
.Y(n_1394)
);

INVx2_ASAP7_75t_SL g1395 ( 
.A(n_1275),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1229),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1229),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1260),
.B(n_1163),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1231),
.B(n_1143),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1231),
.B(n_1146),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_SL g1401 ( 
.A(n_1284),
.B(n_1163),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1231),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1274),
.Y(n_1403)
);

INVx3_ASAP7_75t_L g1404 ( 
.A(n_1274),
.Y(n_1404)
);

NOR2xp33_ASAP7_75t_L g1405 ( 
.A(n_1304),
.B(n_725),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1274),
.B(n_1146),
.Y(n_1406)
);

AND2x4_ASAP7_75t_L g1407 ( 
.A(n_1303),
.B(n_823),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1338),
.A2(n_1281),
.B1(n_1291),
.B2(n_1244),
.Y(n_1408)
);

HB1xp67_ASAP7_75t_L g1409 ( 
.A(n_1350),
.Y(n_1409)
);

O2A1O1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1341),
.A2(n_1268),
.B(n_1277),
.C(n_1254),
.Y(n_1410)
);

CKINVDCx10_ASAP7_75t_R g1411 ( 
.A(n_1313),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1376),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1323),
.A2(n_1404),
.B(n_1375),
.Y(n_1413)
);

AOI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1401),
.A2(n_1290),
.B(n_1129),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1323),
.A2(n_1149),
.B(n_1146),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1323),
.A2(n_1156),
.B(n_1149),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_SL g1417 ( 
.A(n_1338),
.B(n_1382),
.Y(n_1417)
);

AOI21xp5_ASAP7_75t_L g1418 ( 
.A1(n_1323),
.A2(n_1156),
.B(n_1149),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_L g1419 ( 
.A1(n_1375),
.A2(n_1157),
.B(n_1156),
.Y(n_1419)
);

OAI21xp5_ASAP7_75t_L g1420 ( 
.A1(n_1336),
.A2(n_1311),
.B(n_1401),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1343),
.A2(n_1121),
.B(n_1127),
.Y(n_1421)
);

AOI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1404),
.A2(n_1162),
.B(n_1157),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1382),
.A2(n_1263),
.B1(n_1262),
.B2(n_1302),
.Y(n_1423)
);

AOI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1380),
.A2(n_1162),
.B(n_1157),
.Y(n_1424)
);

AOI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1381),
.A2(n_1164),
.B(n_1117),
.Y(n_1425)
);

O2A1O1Ixp33_ASAP7_75t_L g1426 ( 
.A1(n_1341),
.A2(n_1303),
.B(n_1304),
.C(n_696),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1308),
.Y(n_1427)
);

INVx4_ASAP7_75t_L g1428 ( 
.A(n_1402),
.Y(n_1428)
);

NAND2xp5_ASAP7_75t_SL g1429 ( 
.A(n_1395),
.B(n_1244),
.Y(n_1429)
);

AOI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1310),
.A2(n_1154),
.B(n_1130),
.Y(n_1430)
);

OAI21xp33_ASAP7_75t_L g1431 ( 
.A1(n_1363),
.A2(n_1275),
.B(n_1302),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1321),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_SL g1433 ( 
.A(n_1359),
.B(n_1291),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1370),
.B(n_1303),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1384),
.A2(n_1164),
.B(n_1117),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1307),
.B(n_1296),
.Y(n_1436)
);

BUFx8_ASAP7_75t_L g1437 ( 
.A(n_1313),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1358),
.A2(n_1297),
.B1(n_1278),
.B2(n_1241),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1315),
.B(n_1278),
.Y(n_1439)
);

AOI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1347),
.A2(n_1164),
.B(n_1117),
.Y(n_1440)
);

NOR2xp33_ASAP7_75t_L g1441 ( 
.A(n_1405),
.B(n_1299),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1348),
.A2(n_1121),
.B(n_1130),
.Y(n_1442)
);

AND2x2_ASAP7_75t_L g1443 ( 
.A(n_1360),
.B(n_1299),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1325),
.Y(n_1444)
);

INVxp67_ASAP7_75t_L g1445 ( 
.A(n_1350),
.Y(n_1445)
);

OAI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1336),
.A2(n_1278),
.B(n_1121),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1318),
.B(n_1278),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1319),
.Y(n_1448)
);

OAI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1386),
.A2(n_1278),
.B(n_1158),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_L g1450 ( 
.A1(n_1352),
.A2(n_1109),
.B(n_1120),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1322),
.Y(n_1451)
);

AOI21xp5_ASAP7_75t_L g1452 ( 
.A1(n_1402),
.A2(n_1145),
.B(n_1120),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1359),
.B(n_1111),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1328),
.B(n_1113),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_SL g1455 ( 
.A(n_1402),
.B(n_729),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1333),
.Y(n_1456)
);

NOR2xp33_ASAP7_75t_L g1457 ( 
.A(n_1405),
.B(n_1245),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1402),
.A2(n_1145),
.B(n_1120),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1344),
.Y(n_1459)
);

NAND2xp5_ASAP7_75t_L g1460 ( 
.A(n_1328),
.B(n_1113),
.Y(n_1460)
);

BUFx3_ASAP7_75t_L g1461 ( 
.A(n_1327),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1399),
.A2(n_1145),
.B(n_1120),
.Y(n_1462)
);

AOI21xp5_ASAP7_75t_L g1463 ( 
.A1(n_1400),
.A2(n_1145),
.B(n_1120),
.Y(n_1463)
);

AOI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1358),
.A2(n_749),
.B1(n_768),
.B2(n_730),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1353),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1331),
.Y(n_1466)
);

INVx2_ASAP7_75t_SL g1467 ( 
.A(n_1379),
.Y(n_1467)
);

O2A1O1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1394),
.A2(n_696),
.B(n_783),
.C(n_644),
.Y(n_1468)
);

OAI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1386),
.A2(n_1305),
.B(n_1389),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1383),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1335),
.B(n_867),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_L g1472 ( 
.A(n_1306),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1335),
.B(n_885),
.Y(n_1473)
);

AND2x6_ASAP7_75t_L g1474 ( 
.A(n_1391),
.B(n_915),
.Y(n_1474)
);

AOI21xp5_ASAP7_75t_L g1475 ( 
.A1(n_1406),
.A2(n_1145),
.B(n_1120),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1342),
.B(n_626),
.Y(n_1476)
);

BUFx6f_ASAP7_75t_L g1477 ( 
.A(n_1309),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1326),
.B(n_915),
.Y(n_1478)
);

NOR2x1_ASAP7_75t_L g1479 ( 
.A(n_1310),
.B(n_772),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1345),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_L g1481 ( 
.A(n_1351),
.B(n_1245),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1362),
.B(n_626),
.Y(n_1482)
);

OR2x6_ASAP7_75t_L g1483 ( 
.A(n_1317),
.B(n_1385),
.Y(n_1483)
);

AO21x1_ASAP7_75t_L g1484 ( 
.A1(n_1332),
.A2(n_1158),
.B(n_1154),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1362),
.A2(n_774),
.B1(n_792),
.B2(n_787),
.Y(n_1485)
);

A2O1A1Ixp33_ASAP7_75t_L g1486 ( 
.A1(n_1316),
.A2(n_644),
.B(n_841),
.C(n_783),
.Y(n_1486)
);

AOI21xp5_ASAP7_75t_L g1487 ( 
.A1(n_1369),
.A2(n_1145),
.B(n_1120),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1349),
.Y(n_1488)
);

A2O1A1Ixp33_ASAP7_75t_L g1489 ( 
.A1(n_1367),
.A2(n_907),
.B(n_991),
.C(n_841),
.Y(n_1489)
);

INVx5_ASAP7_75t_L g1490 ( 
.A(n_1309),
.Y(n_1490)
);

A2O1A1Ixp33_ASAP7_75t_L g1491 ( 
.A1(n_1314),
.A2(n_991),
.B(n_907),
.C(n_789),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1334),
.B(n_809),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1320),
.A2(n_1148),
.B(n_1145),
.Y(n_1493)
);

AOI21xp5_ASAP7_75t_L g1494 ( 
.A1(n_1330),
.A2(n_1163),
.B(n_1148),
.Y(n_1494)
);

NOR2xp33_ASAP7_75t_L g1495 ( 
.A(n_1351),
.B(n_1052),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1312),
.B(n_1125),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1407),
.B(n_1135),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1361),
.Y(n_1498)
);

AOI21xp5_ASAP7_75t_L g1499 ( 
.A1(n_1339),
.A2(n_1163),
.B(n_1148),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1309),
.B(n_829),
.Y(n_1500)
);

NAND2x1_ASAP7_75t_L g1501 ( 
.A(n_1309),
.B(n_1135),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1329),
.B(n_892),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1385),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1365),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

OAI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1423),
.A2(n_1397),
.B1(n_1396),
.B2(n_1329),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1427),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1441),
.B(n_1417),
.Y(n_1508)
);

NAND3xp33_ASAP7_75t_SL g1509 ( 
.A(n_1464),
.B(n_1373),
.C(n_1378),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1471),
.A2(n_1363),
.B1(n_1378),
.B2(n_1407),
.Y(n_1510)
);

AOI21xp5_ASAP7_75t_L g1511 ( 
.A1(n_1469),
.A2(n_1374),
.B(n_1388),
.Y(n_1511)
);

O2A1O1Ixp33_ASAP7_75t_L g1512 ( 
.A1(n_1426),
.A2(n_1354),
.B(n_1340),
.C(n_1356),
.Y(n_1512)
);

AOI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1469),
.A2(n_1392),
.B(n_1364),
.Y(n_1513)
);

AOI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1413),
.A2(n_1364),
.B(n_1324),
.Y(n_1514)
);

CKINVDCx11_ASAP7_75t_R g1515 ( 
.A(n_1461),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1443),
.B(n_1377),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1448),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_SL g1518 ( 
.A(n_1410),
.B(n_1329),
.Y(n_1518)
);

INVx5_ASAP7_75t_L g1519 ( 
.A(n_1477),
.Y(n_1519)
);

INVx3_ASAP7_75t_L g1520 ( 
.A(n_1428),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1473),
.B(n_1355),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_SL g1522 ( 
.A(n_1479),
.B(n_1329),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1482),
.A2(n_742),
.B1(n_789),
.B2(n_711),
.Y(n_1523)
);

AOI22xp5_ASAP7_75t_L g1524 ( 
.A1(n_1436),
.A2(n_1371),
.B1(n_1357),
.B2(n_906),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1459),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1420),
.A2(n_1324),
.B(n_1398),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1431),
.B(n_1337),
.Y(n_1527)
);

BUFx3_ASAP7_75t_L g1528 ( 
.A(n_1412),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1451),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1466),
.Y(n_1530)
);

AND2x2_ASAP7_75t_L g1531 ( 
.A(n_1476),
.B(n_626),
.Y(n_1531)
);

AOI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1430),
.A2(n_1346),
.B(n_1337),
.Y(n_1532)
);

INVxp67_ASAP7_75t_SL g1533 ( 
.A(n_1477),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_1411),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1434),
.B(n_1372),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_L g1536 ( 
.A1(n_1484),
.A2(n_1346),
.B(n_1390),
.C(n_1387),
.Y(n_1536)
);

AOI21xp5_ASAP7_75t_L g1537 ( 
.A1(n_1420),
.A2(n_1398),
.B(n_1403),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_L g1538 ( 
.A(n_1428),
.B(n_1366),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_SL g1539 ( 
.A(n_1470),
.B(n_905),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1488),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_SL g1541 ( 
.A1(n_1439),
.A2(n_1368),
.B(n_595),
.C(n_598),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1454),
.B(n_1393),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_SL g1543 ( 
.A(n_1438),
.B(n_1159),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1446),
.A2(n_1163),
.B(n_1148),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1432),
.Y(n_1545)
);

BUFx2_ASAP7_75t_L g1546 ( 
.A(n_1409),
.Y(n_1546)
);

INVx3_ASAP7_75t_L g1547 ( 
.A(n_1477),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_SL g1548 ( 
.A1(n_1485),
.A2(n_949),
.B1(n_952),
.B2(n_919),
.Y(n_1548)
);

AOI21xp5_ASAP7_75t_L g1549 ( 
.A1(n_1446),
.A2(n_1166),
.B(n_1148),
.Y(n_1549)
);

AOI22x1_ASAP7_75t_L g1550 ( 
.A1(n_1444),
.A2(n_881),
.B1(n_595),
.B2(n_598),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1424),
.A2(n_1166),
.B(n_1148),
.Y(n_1551)
);

HB1xp67_ASAP7_75t_L g1552 ( 
.A(n_1503),
.Y(n_1552)
);

O2A1O1Ixp33_ASAP7_75t_L g1553 ( 
.A1(n_1489),
.A2(n_826),
.B(n_836),
.C(n_813),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1437),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1408),
.A2(n_973),
.B1(n_978),
.B2(n_950),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1460),
.B(n_843),
.Y(n_1556)
);

BUFx2_ASAP7_75t_L g1557 ( 
.A(n_1445),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_1437),
.Y(n_1558)
);

INVx1_ASAP7_75t_SL g1559 ( 
.A(n_1465),
.Y(n_1559)
);

O2A1O1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1485),
.A2(n_879),
.B(n_941),
.C(n_852),
.Y(n_1560)
);

OAI21x1_ASAP7_75t_L g1561 ( 
.A1(n_1421),
.A2(n_1159),
.B(n_1136),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1480),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1453),
.B(n_998),
.Y(n_1563)
);

INVxp67_ASAP7_75t_SL g1564 ( 
.A(n_1498),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1455),
.B(n_1011),
.Y(n_1565)
);

INVxp67_ASAP7_75t_SL g1566 ( 
.A(n_1504),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1433),
.B(n_881),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1500),
.B(n_626),
.Y(n_1568)
);

BUFx8_ASAP7_75t_SL g1569 ( 
.A(n_1472),
.Y(n_1569)
);

O2A1O1Ixp33_ASAP7_75t_L g1570 ( 
.A1(n_1492),
.A2(n_608),
.B(n_614),
.C(n_594),
.Y(n_1570)
);

O2A1O1Ixp33_ASAP7_75t_L g1571 ( 
.A1(n_1408),
.A2(n_608),
.B(n_614),
.C(n_594),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1502),
.B(n_675),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1478),
.B(n_597),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1447),
.B(n_1123),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1497),
.Y(n_1575)
);

NOR2xp33_ASAP7_75t_L g1576 ( 
.A(n_1457),
.B(n_983),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1467),
.B(n_617),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_L g1578 ( 
.A(n_1486),
.B(n_599),
.Y(n_1578)
);

BUFx6f_ASAP7_75t_SL g1579 ( 
.A(n_1483),
.Y(n_1579)
);

INVx5_ASAP7_75t_L g1580 ( 
.A(n_1490),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_SL g1581 ( 
.A(n_1490),
.B(n_1123),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1483),
.B(n_675),
.Y(n_1582)
);

AO22x1_ASAP7_75t_L g1583 ( 
.A1(n_1495),
.A2(n_1481),
.B1(n_1474),
.B2(n_1490),
.Y(n_1583)
);

O2A1O1Ixp5_ASAP7_75t_SL g1584 ( 
.A1(n_1449),
.A2(n_617),
.B(n_620),
.C(n_618),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1496),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1491),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1501),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1449),
.A2(n_1166),
.B(n_1148),
.Y(n_1588)
);

AND3x1_ASAP7_75t_SL g1589 ( 
.A(n_1429),
.B(n_620),
.C(n_618),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1483),
.B(n_601),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1442),
.Y(n_1591)
);

NAND3xp33_ASAP7_75t_L g1592 ( 
.A(n_1468),
.B(n_604),
.C(n_603),
.Y(n_1592)
);

CKINVDCx5p33_ASAP7_75t_R g1593 ( 
.A(n_1472),
.Y(n_1593)
);

BUFx4f_ASAP7_75t_L g1594 ( 
.A(n_1474),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1490),
.Y(n_1595)
);

O2A1O1Ixp33_ASAP7_75t_L g1596 ( 
.A1(n_1487),
.A2(n_625),
.B(n_640),
.C(n_633),
.Y(n_1596)
);

OAI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1414),
.A2(n_1008),
.B1(n_607),
.B2(n_609),
.Y(n_1597)
);

INVxp67_ASAP7_75t_SL g1598 ( 
.A(n_1452),
.Y(n_1598)
);

AOI21xp5_ASAP7_75t_L g1599 ( 
.A1(n_1462),
.A2(n_1166),
.B(n_1136),
.Y(n_1599)
);

NAND3xp33_ASAP7_75t_SL g1600 ( 
.A(n_1425),
.B(n_612),
.C(n_605),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1474),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1474),
.Y(n_1602)
);

NOR3xp33_ASAP7_75t_L g1603 ( 
.A(n_1493),
.B(n_633),
.C(n_625),
.Y(n_1603)
);

OAI22xp33_ASAP7_75t_L g1604 ( 
.A1(n_1435),
.A2(n_649),
.B1(n_606),
.B2(n_711),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1419),
.B(n_613),
.Y(n_1605)
);

AO31x2_ASAP7_75t_L g1606 ( 
.A1(n_1591),
.A2(n_1526),
.A3(n_1511),
.B(n_1513),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_SL g1607 ( 
.A(n_1534),
.B(n_1569),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_L g1608 ( 
.A1(n_1509),
.A2(n_1499),
.B(n_1494),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1510),
.A2(n_615),
.B1(n_619),
.B2(n_616),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1516),
.B(n_623),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1556),
.B(n_1508),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1528),
.B(n_1458),
.Y(n_1612)
);

NOR2xp67_ASAP7_75t_L g1613 ( 
.A(n_1580),
.B(n_1440),
.Y(n_1613)
);

AOI21xp5_ASAP7_75t_L g1614 ( 
.A1(n_1518),
.A2(n_1475),
.B(n_1463),
.Y(n_1614)
);

CKINVDCx5p33_ASAP7_75t_R g1615 ( 
.A(n_1515),
.Y(n_1615)
);

BUFx6f_ASAP7_75t_L g1616 ( 
.A(n_1528),
.Y(n_1616)
);

INVx4_ASAP7_75t_L g1617 ( 
.A(n_1580),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1510),
.B(n_624),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1561),
.A2(n_1514),
.B(n_1532),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1518),
.A2(n_1450),
.B(n_1422),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1599),
.A2(n_1416),
.B(n_1415),
.Y(n_1621)
);

AOI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1583),
.A2(n_1543),
.B(n_1588),
.Y(n_1622)
);

OAI22x1_ASAP7_75t_L g1623 ( 
.A1(n_1524),
.A2(n_641),
.B1(n_651),
.B2(n_640),
.Y(n_1623)
);

A2O1A1Ixp33_ASAP7_75t_L g1624 ( 
.A1(n_1512),
.A2(n_742),
.B(n_789),
.C(n_711),
.Y(n_1624)
);

INVxp67_ASAP7_75t_L g1625 ( 
.A(n_1552),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_SL g1626 ( 
.A(n_1539),
.B(n_675),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1537),
.A2(n_1418),
.B(n_1166),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1507),
.Y(n_1628)
);

INVx5_ASAP7_75t_L g1629 ( 
.A(n_1580),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1598),
.A2(n_1166),
.B(n_1123),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1573),
.A2(n_666),
.B(n_663),
.Y(n_1631)
);

NAND3x1_ASAP7_75t_L g1632 ( 
.A(n_1576),
.B(n_669),
.C(n_666),
.Y(n_1632)
);

OAI21xp5_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_670),
.B(n_669),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1575),
.B(n_630),
.Y(n_1634)
);

A2O1A1Ixp33_ASAP7_75t_L g1635 ( 
.A1(n_1560),
.A2(n_982),
.B(n_649),
.C(n_606),
.Y(n_1635)
);

INVx3_ASAP7_75t_L g1636 ( 
.A(n_1580),
.Y(n_1636)
);

AOI21xp5_ASAP7_75t_L g1637 ( 
.A1(n_1598),
.A2(n_1166),
.B(n_1123),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1563),
.B(n_634),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1517),
.Y(n_1639)
);

OAI21xp5_ASAP7_75t_L g1640 ( 
.A1(n_1605),
.A2(n_671),
.B(n_670),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_SL g1641 ( 
.A(n_1576),
.B(n_637),
.C(n_636),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1529),
.Y(n_1642)
);

NOR2xp67_ASAP7_75t_L g1643 ( 
.A(n_1600),
.B(n_567),
.Y(n_1643)
);

OAI21xp5_ASAP7_75t_L g1644 ( 
.A1(n_1527),
.A2(n_672),
.B(n_671),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1505),
.Y(n_1645)
);

OAI21x1_ASAP7_75t_L g1646 ( 
.A1(n_1551),
.A2(n_1059),
.B(n_1058),
.Y(n_1646)
);

A2O1A1Ixp33_ASAP7_75t_L g1647 ( 
.A1(n_1553),
.A2(n_982),
.B(n_674),
.C(n_676),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1552),
.B(n_672),
.Y(n_1648)
);

OR2x2_ASAP7_75t_L g1649 ( 
.A(n_1546),
.B(n_1565),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1548),
.A2(n_638),
.B1(n_639),
.B2(n_635),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1543),
.A2(n_1549),
.B(n_1544),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1542),
.A2(n_1123),
.B(n_1060),
.Y(n_1652)
);

NOR2xp33_ASAP7_75t_L g1653 ( 
.A(n_1555),
.B(n_642),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1559),
.B(n_1557),
.Y(n_1654)
);

AOI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1521),
.A2(n_1535),
.B(n_1574),
.Y(n_1655)
);

AO31x2_ASAP7_75t_L g1656 ( 
.A1(n_1527),
.A2(n_632),
.A3(n_678),
.B(n_610),
.Y(n_1656)
);

O2A1O1Ixp5_ASAP7_75t_L g1657 ( 
.A1(n_1522),
.A2(n_676),
.B(n_682),
.C(n_674),
.Y(n_1657)
);

XNOR2xp5_ASAP7_75t_L g1658 ( 
.A(n_1558),
.B(n_643),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1531),
.B(n_645),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1505),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1536),
.A2(n_1060),
.B(n_1059),
.Y(n_1661)
);

NOR2xp67_ASAP7_75t_L g1662 ( 
.A(n_1592),
.B(n_569),
.Y(n_1662)
);

AOI21xp5_ASAP7_75t_SL g1663 ( 
.A1(n_1506),
.A2(n_890),
.B(n_631),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1525),
.Y(n_1664)
);

AO21x2_ASAP7_75t_L g1665 ( 
.A1(n_1574),
.A2(n_683),
.B(n_682),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1581),
.A2(n_1070),
.B(n_1063),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_SL g1667 ( 
.A(n_1567),
.B(n_675),
.Y(n_1667)
);

NOR2xp33_ASAP7_75t_L g1668 ( 
.A(n_1590),
.B(n_647),
.Y(n_1668)
);

AOI21xp5_ASAP7_75t_L g1669 ( 
.A1(n_1564),
.A2(n_1123),
.B(n_1070),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1584),
.A2(n_1071),
.B(n_1063),
.Y(n_1670)
);

OAI21x1_ASAP7_75t_SL g1671 ( 
.A1(n_1596),
.A2(n_632),
.B(n_610),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1520),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1597),
.A2(n_685),
.B(n_683),
.Y(n_1673)
);

CKINVDCx11_ASAP7_75t_R g1674 ( 
.A(n_1554),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1578),
.A2(n_689),
.B(n_685),
.Y(n_1675)
);

OAI21x1_ASAP7_75t_L g1676 ( 
.A1(n_1586),
.A2(n_1587),
.B(n_1581),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1525),
.Y(n_1677)
);

INVx3_ASAP7_75t_L g1678 ( 
.A(n_1520),
.Y(n_1678)
);

BUFx6f_ASAP7_75t_L g1679 ( 
.A(n_1519),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1564),
.A2(n_1072),
.B(n_1071),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1540),
.Y(n_1681)
);

OAI21xp5_ASAP7_75t_L g1682 ( 
.A1(n_1571),
.A2(n_691),
.B(n_689),
.Y(n_1682)
);

AND2x6_ASAP7_75t_L g1683 ( 
.A(n_1601),
.B(n_691),
.Y(n_1683)
);

INVx2_ASAP7_75t_L g1684 ( 
.A(n_1545),
.Y(n_1684)
);

NAND2xp5_ASAP7_75t_L g1685 ( 
.A(n_1568),
.B(n_648),
.Y(n_1685)
);

NAND3xp33_ASAP7_75t_L g1686 ( 
.A(n_1523),
.B(n_654),
.C(n_652),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1639),
.Y(n_1687)
);

CKINVDCx6p67_ASAP7_75t_R g1688 ( 
.A(n_1674),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1619),
.A2(n_1602),
.B(n_1550),
.Y(n_1689)
);

AOI22x1_ASAP7_75t_L g1690 ( 
.A1(n_1633),
.A2(n_1572),
.B1(n_1566),
.B2(n_1593),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1614),
.A2(n_1541),
.B(n_1603),
.Y(n_1691)
);

AOI21x1_ASAP7_75t_L g1692 ( 
.A1(n_1622),
.A2(n_1585),
.B(n_1538),
.Y(n_1692)
);

CKINVDCx16_ASAP7_75t_R g1693 ( 
.A(n_1607),
.Y(n_1693)
);

AND2x4_ASAP7_75t_SL g1694 ( 
.A(n_1616),
.B(n_1547),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1608),
.A2(n_1566),
.B(n_1530),
.Y(n_1695)
);

AOI22xp33_ASAP7_75t_L g1696 ( 
.A1(n_1640),
.A2(n_1523),
.B1(n_839),
.B2(n_882),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.B(n_1562),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1645),
.Y(n_1698)
);

O2A1O1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1631),
.A2(n_1570),
.B(n_1541),
.C(n_1604),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1642),
.Y(n_1700)
);

AOI21xp5_ASAP7_75t_L g1701 ( 
.A1(n_1655),
.A2(n_1594),
.B(n_1533),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1625),
.B(n_1577),
.Y(n_1702)
);

OR2x2_ASAP7_75t_L g1703 ( 
.A(n_1611),
.B(n_1577),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

INVx2_ASAP7_75t_SL g1705 ( 
.A(n_1616),
.Y(n_1705)
);

OAI21x1_ASAP7_75t_L g1706 ( 
.A1(n_1620),
.A2(n_1595),
.B(n_1547),
.Y(n_1706)
);

OAI21x1_ASAP7_75t_L g1707 ( 
.A1(n_1621),
.A2(n_1533),
.B(n_1582),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1630),
.A2(n_695),
.B(n_693),
.Y(n_1708)
);

OR2x2_ASAP7_75t_L g1709 ( 
.A(n_1664),
.B(n_1677),
.Y(n_1709)
);

OA21x2_ASAP7_75t_L g1710 ( 
.A1(n_1637),
.A2(n_695),
.B(n_693),
.Y(n_1710)
);

AND2x4_ASAP7_75t_L g1711 ( 
.A(n_1681),
.B(n_1628),
.Y(n_1711)
);

OAI21x1_ASAP7_75t_SL g1712 ( 
.A1(n_1644),
.A2(n_1589),
.B(n_684),
.Y(n_1712)
);

OAI21x1_ASAP7_75t_L g1713 ( 
.A1(n_1627),
.A2(n_1077),
.B(n_1073),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1618),
.B(n_1604),
.Y(n_1714)
);

BUFx4f_ASAP7_75t_L g1715 ( 
.A(n_1616),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1641),
.A2(n_1579),
.B1(n_1589),
.B2(n_1594),
.Y(n_1716)
);

OAI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1675),
.A2(n_710),
.B1(n_718),
.B2(n_708),
.C(n_703),
.Y(n_1717)
);

AO32x2_ASAP7_75t_L g1718 ( 
.A1(n_1609),
.A2(n_1579),
.A3(n_882),
.B1(n_1010),
.B2(n_839),
.Y(n_1718)
);

AOI21x1_ASAP7_75t_L g1719 ( 
.A1(n_1613),
.A2(n_708),
.B(n_703),
.Y(n_1719)
);

BUFx5_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1684),
.B(n_1519),
.Y(n_1721)
);

NOR2x1_ASAP7_75t_L g1722 ( 
.A(n_1612),
.B(n_982),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1663),
.B(n_1519),
.Y(n_1723)
);

INVx3_ASAP7_75t_L g1724 ( 
.A(n_1679),
.Y(n_1724)
);

OAI21xp5_ASAP7_75t_L g1725 ( 
.A1(n_1653),
.A2(n_1624),
.B(n_1635),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1679),
.Y(n_1726)
);

AOI22x1_ASAP7_75t_L g1727 ( 
.A1(n_1623),
.A2(n_655),
.B1(n_657),
.B2(n_656),
.Y(n_1727)
);

OA21x2_ASAP7_75t_L g1728 ( 
.A1(n_1651),
.A2(n_718),
.B(n_710),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1615),
.Y(n_1729)
);

OAI21x1_ASAP7_75t_L g1730 ( 
.A1(n_1676),
.A2(n_1646),
.B(n_1661),
.Y(n_1730)
);

OA21x2_ASAP7_75t_L g1731 ( 
.A1(n_1652),
.A2(n_727),
.B(n_723),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1656),
.Y(n_1732)
);

OA21x2_ASAP7_75t_L g1733 ( 
.A1(n_1670),
.A2(n_727),
.B(n_723),
.Y(n_1733)
);

NOR2x1_ASAP7_75t_L g1734 ( 
.A(n_1612),
.B(n_732),
.Y(n_1734)
);

OAI21x1_ASAP7_75t_L g1735 ( 
.A1(n_1666),
.A2(n_1079),
.B(n_1077),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1656),
.Y(n_1736)
);

AOI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1650),
.A2(n_660),
.B1(n_662),
.B2(n_661),
.C(n_659),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1654),
.B(n_1519),
.Y(n_1738)
);

O2A1O1Ixp33_ASAP7_75t_SL g1739 ( 
.A1(n_1647),
.A2(n_735),
.B(n_736),
.C(n_732),
.Y(n_1739)
);

BUFx2_ASAP7_75t_L g1740 ( 
.A(n_1672),
.Y(n_1740)
);

AOI221xp5_ASAP7_75t_L g1741 ( 
.A1(n_1673),
.A2(n_665),
.B1(n_668),
.B2(n_667),
.C(n_664),
.Y(n_1741)
);

AOI22xp33_ASAP7_75t_L g1742 ( 
.A1(n_1626),
.A2(n_1682),
.B1(n_1686),
.B2(n_839),
.Y(n_1742)
);

OAI21x1_ASAP7_75t_L g1743 ( 
.A1(n_1669),
.A2(n_1084),
.B(n_1083),
.Y(n_1743)
);

NAND3xp33_ASAP7_75t_L g1744 ( 
.A(n_1668),
.B(n_677),
.C(n_673),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1687),
.Y(n_1745)
);

OAI21x1_ASAP7_75t_L g1746 ( 
.A1(n_1730),
.A2(n_1613),
.B(n_1657),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1698),
.Y(n_1747)
);

O2A1O1Ixp33_ASAP7_75t_L g1748 ( 
.A1(n_1725),
.A2(n_1667),
.B(n_1685),
.C(n_1671),
.Y(n_1748)
);

OAI21xp5_ASAP7_75t_L g1749 ( 
.A1(n_1699),
.A2(n_1632),
.B(n_1643),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1700),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1698),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1711),
.B(n_1606),
.Y(n_1752)
);

OAI21x1_ASAP7_75t_SL g1753 ( 
.A1(n_1712),
.A2(n_1617),
.B(n_1680),
.Y(n_1753)
);

OAI21xp5_ASAP7_75t_L g1754 ( 
.A1(n_1690),
.A2(n_1643),
.B(n_1662),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1711),
.Y(n_1755)
);

AOI21xp5_ASAP7_75t_L g1756 ( 
.A1(n_1695),
.A2(n_1629),
.B(n_1662),
.Y(n_1756)
);

OAI21x1_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1689),
.B(n_1706),
.Y(n_1757)
);

OA21x2_ASAP7_75t_L g1758 ( 
.A1(n_1732),
.A2(n_736),
.B(n_735),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1704),
.Y(n_1760)
);

INVx8_ASAP7_75t_L g1761 ( 
.A(n_1723),
.Y(n_1761)
);

OAI21x1_ASAP7_75t_L g1762 ( 
.A1(n_1689),
.A2(n_1636),
.B(n_1672),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1736),
.B(n_1606),
.Y(n_1763)
);

INVx1_ASAP7_75t_SL g1764 ( 
.A(n_1740),
.Y(n_1764)
);

OAI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1742),
.A2(n_1659),
.B(n_1638),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1707),
.A2(n_748),
.B(n_745),
.Y(n_1766)
);

AO31x2_ASAP7_75t_L g1767 ( 
.A1(n_1701),
.A2(n_1714),
.A3(n_1728),
.B(n_1695),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1695),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1709),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1711),
.Y(n_1770)
);

NAND2x1p5_ASAP7_75t_L g1771 ( 
.A(n_1707),
.B(n_1629),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1716),
.B(n_1703),
.Y(n_1772)
);

OAI21x1_ASAP7_75t_L g1773 ( 
.A1(n_1706),
.A2(n_1636),
.B(n_1678),
.Y(n_1773)
);

OAI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1742),
.A2(n_1634),
.B(n_1610),
.Y(n_1774)
);

AO21x2_ASAP7_75t_L g1775 ( 
.A1(n_1692),
.A2(n_1665),
.B(n_748),
.Y(n_1775)
);

NAND2x1p5_ASAP7_75t_L g1776 ( 
.A(n_1734),
.B(n_1629),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1697),
.B(n_1665),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1728),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1722),
.B(n_1678),
.Y(n_1779)
);

AO21x2_ASAP7_75t_L g1780 ( 
.A1(n_1691),
.A2(n_754),
.B(n_745),
.Y(n_1780)
);

AOI21x1_ASAP7_75t_L g1781 ( 
.A1(n_1719),
.A2(n_1648),
.B(n_758),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1728),
.Y(n_1782)
);

AOI22xp33_ASAP7_75t_L g1783 ( 
.A1(n_1696),
.A2(n_1683),
.B1(n_678),
.B2(n_747),
.Y(n_1783)
);

OAI21x1_ASAP7_75t_L g1784 ( 
.A1(n_1713),
.A2(n_758),
.B(n_754),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1708),
.Y(n_1785)
);

HB1xp67_ASAP7_75t_L g1786 ( 
.A(n_1702),
.Y(n_1786)
);

INVx2_ASAP7_75t_L g1787 ( 
.A(n_1733),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1708),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1708),
.Y(n_1789)
);

CKINVDCx5p33_ASAP7_75t_R g1790 ( 
.A(n_1729),
.Y(n_1790)
);

OA21x2_ASAP7_75t_L g1791 ( 
.A1(n_1713),
.A2(n_776),
.B(n_765),
.Y(n_1791)
);

NOR2x1_ASAP7_75t_SL g1792 ( 
.A(n_1723),
.B(n_1679),
.Y(n_1792)
);

HB1xp67_ASAP7_75t_L g1793 ( 
.A(n_1768),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1747),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1752),
.B(n_1710),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1747),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1747),
.Y(n_1797)
);

AO21x2_ASAP7_75t_L g1798 ( 
.A1(n_1768),
.A2(n_1691),
.B(n_1717),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1752),
.B(n_1710),
.Y(n_1799)
);

BUFx3_ASAP7_75t_L g1800 ( 
.A(n_1761),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1768),
.B(n_1710),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1751),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1751),
.B(n_1726),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1770),
.B(n_1733),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1751),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1759),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1770),
.B(n_1733),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1759),
.Y(n_1808)
);

BUFx2_ASAP7_75t_L g1809 ( 
.A(n_1771),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1759),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1760),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1760),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1760),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1745),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1787),
.Y(n_1815)
);

BUFx3_ASAP7_75t_L g1816 ( 
.A(n_1761),
.Y(n_1816)
);

BUFx3_ASAP7_75t_L g1817 ( 
.A(n_1761),
.Y(n_1817)
);

INVx2_ASAP7_75t_L g1818 ( 
.A(n_1787),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1745),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1761),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1769),
.B(n_1731),
.Y(n_1822)
);

OR2x2_ASAP7_75t_L g1823 ( 
.A(n_1767),
.B(n_1731),
.Y(n_1823)
);

AO21x2_ASAP7_75t_L g1824 ( 
.A1(n_1756),
.A2(n_1739),
.B(n_1735),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1750),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1787),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1750),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1758),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1786),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1758),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1785),
.Y(n_1831)
);

BUFx2_ASAP7_75t_L g1832 ( 
.A(n_1771),
.Y(n_1832)
);

BUFx2_ASAP7_75t_L g1833 ( 
.A(n_1771),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1758),
.Y(n_1834)
);

BUFx6f_ASAP7_75t_L g1835 ( 
.A(n_1766),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1766),
.B(n_1720),
.Y(n_1836)
);

AND2x2_ASAP7_75t_L g1837 ( 
.A(n_1766),
.B(n_1720),
.Y(n_1837)
);

OR2x2_ASAP7_75t_L g1838 ( 
.A(n_1767),
.B(n_1738),
.Y(n_1838)
);

BUFx2_ASAP7_75t_L g1839 ( 
.A(n_1762),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1785),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1758),
.Y(n_1841)
);

AND2x4_ASAP7_75t_L g1842 ( 
.A(n_1762),
.B(n_1726),
.Y(n_1842)
);

OR2x6_ASAP7_75t_L g1843 ( 
.A(n_1761),
.B(n_1723),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1758),
.Y(n_1844)
);

HB1xp67_ASAP7_75t_L g1845 ( 
.A(n_1763),
.Y(n_1845)
);

INVx3_ASAP7_75t_L g1846 ( 
.A(n_1762),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1829),
.A2(n_1765),
.B1(n_1774),
.B2(n_1696),
.C(n_778),
.Y(n_1847)
);

OAI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1843),
.A2(n_1749),
.B1(n_1754),
.B2(n_1776),
.Y(n_1848)
);

AOI22xp33_ASAP7_75t_L g1849 ( 
.A1(n_1800),
.A2(n_1772),
.B1(n_1749),
.B2(n_1744),
.Y(n_1849)
);

INVx4_ASAP7_75t_L g1850 ( 
.A(n_1843),
.Y(n_1850)
);

OR2x2_ASAP7_75t_L g1851 ( 
.A(n_1838),
.B(n_1829),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_L g1852 ( 
.A1(n_1800),
.A2(n_1765),
.B1(n_1774),
.B2(n_1754),
.Y(n_1852)
);

AND2x2_ASAP7_75t_SL g1853 ( 
.A(n_1835),
.B(n_1836),
.Y(n_1853)
);

OA21x2_ASAP7_75t_L g1854 ( 
.A1(n_1839),
.A2(n_1757),
.B(n_1756),
.Y(n_1854)
);

OAI221xp5_ASAP7_75t_L g1855 ( 
.A1(n_1838),
.A2(n_1748),
.B1(n_1741),
.B2(n_1783),
.C(n_1737),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1819),
.Y(n_1856)
);

HB1xp67_ASAP7_75t_L g1857 ( 
.A(n_1845),
.Y(n_1857)
);

OAI21xp33_ASAP7_75t_L g1858 ( 
.A1(n_1838),
.A2(n_1777),
.B(n_776),
.Y(n_1858)
);

OAI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1843),
.A2(n_1776),
.B1(n_1755),
.B2(n_1748),
.Y(n_1859)
);

AOI222xp33_ASAP7_75t_L g1860 ( 
.A1(n_1836),
.A2(n_796),
.B1(n_778),
.B2(n_798),
.C1(n_790),
.C2(n_765),
.Y(n_1860)
);

AOI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1800),
.A2(n_1727),
.B1(n_1753),
.B2(n_1720),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1845),
.Y(n_1862)
);

AOI222xp33_ASAP7_75t_L g1863 ( 
.A1(n_1836),
.A2(n_802),
.B1(n_796),
.B2(n_812),
.C1(n_798),
.C2(n_790),
.Y(n_1863)
);

OAI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1838),
.A2(n_1776),
.B1(n_1658),
.B2(n_816),
.C(n_817),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1795),
.B(n_1755),
.Y(n_1865)
);

OAI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1843),
.A2(n_1761),
.B1(n_1693),
.B2(n_1764),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1819),
.Y(n_1867)
);

INVx3_ASAP7_75t_SL g1868 ( 
.A(n_1843),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1794),
.B(n_1767),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1794),
.Y(n_1870)
);

AOI22xp33_ASAP7_75t_L g1871 ( 
.A1(n_1800),
.A2(n_1753),
.B1(n_1720),
.B2(n_1779),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1803),
.B(n_1764),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1795),
.B(n_1767),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1816),
.A2(n_1720),
.B1(n_1779),
.B2(n_1777),
.Y(n_1874)
);

AOI222xp33_ASAP7_75t_L g1875 ( 
.A1(n_1836),
.A2(n_817),
.B1(n_812),
.B2(n_824),
.C1(n_816),
.C2(n_802),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1803),
.B(n_1767),
.Y(n_1876)
);

AO21x2_ASAP7_75t_L g1877 ( 
.A1(n_1828),
.A2(n_1757),
.B(n_1778),
.Y(n_1877)
);

AOI221xp5_ASAP7_75t_L g1878 ( 
.A1(n_1822),
.A2(n_831),
.B1(n_838),
.B2(n_828),
.C(n_824),
.Y(n_1878)
);

BUFx6f_ASAP7_75t_L g1879 ( 
.A(n_1868),
.Y(n_1879)
);

INVx2_ASAP7_75t_L g1880 ( 
.A(n_1870),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1870),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1857),
.Y(n_1882)
);

AND2x2_ASAP7_75t_L g1883 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1883)
);

HB1xp67_ASAP7_75t_L g1884 ( 
.A(n_1862),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1869),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1886)
);

OR2x2_ASAP7_75t_L g1887 ( 
.A(n_1851),
.B(n_1876),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1856),
.Y(n_1888)
);

AOI22xp33_ASAP7_75t_L g1889 ( 
.A1(n_1847),
.A2(n_1855),
.B1(n_1852),
.B2(n_1864),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1856),
.Y(n_1890)
);

AOI22xp33_ASAP7_75t_L g1891 ( 
.A1(n_1848),
.A2(n_1817),
.B1(n_1821),
.B2(n_1816),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1853),
.B(n_1832),
.Y(n_1892)
);

INVxp67_ASAP7_75t_SL g1893 ( 
.A(n_1869),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1851),
.B(n_1873),
.Y(n_1894)
);

OAI22xp5_ASAP7_75t_L g1895 ( 
.A1(n_1849),
.A2(n_1835),
.B1(n_1823),
.B2(n_1843),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1867),
.B(n_1814),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1867),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1877),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1865),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1865),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1872),
.B(n_1790),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1858),
.A2(n_1835),
.B1(n_1823),
.B2(n_1843),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1850),
.B(n_1688),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1877),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1873),
.B(n_1814),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1868),
.B(n_1820),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1877),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1868),
.B(n_1833),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1850),
.B(n_1820),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1890),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1890),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1888),
.Y(n_1912)
);

NAND2xp5_ASAP7_75t_L g1913 ( 
.A(n_1888),
.B(n_1897),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1897),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1883),
.B(n_1850),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1898),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1879),
.B(n_1809),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1896),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1905),
.B(n_1793),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1883),
.B(n_1809),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1898),
.Y(n_1921)
);

INVx2_ASAP7_75t_L g1922 ( 
.A(n_1898),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1909),
.B(n_1820),
.Y(n_1923)
);

INVx1_ASAP7_75t_SL g1924 ( 
.A(n_1882),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1886),
.B(n_1809),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1886),
.B(n_1833),
.Y(n_1926)
);

NAND2x1p5_ASAP7_75t_SL g1927 ( 
.A(n_1889),
.B(n_1718),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1896),
.Y(n_1928)
);

INVx2_ASAP7_75t_L g1929 ( 
.A(n_1907),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1907),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1892),
.B(n_1833),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1907),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1879),
.B(n_1892),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1880),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1880),
.Y(n_1935)
);

INVx1_ASAP7_75t_L g1936 ( 
.A(n_1880),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1884),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1905),
.B(n_1793),
.Y(n_1938)
);

INVxp67_ASAP7_75t_L g1939 ( 
.A(n_1903),
.Y(n_1939)
);

AND2x2_ASAP7_75t_L g1940 ( 
.A(n_1908),
.B(n_1842),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1881),
.Y(n_1941)
);

AND2x2_ASAP7_75t_SL g1942 ( 
.A(n_1891),
.B(n_1835),
.Y(n_1942)
);

BUFx6f_ASAP7_75t_L g1943 ( 
.A(n_1933),
.Y(n_1943)
);

OAI211xp5_ASAP7_75t_L g1944 ( 
.A1(n_1924),
.A2(n_1863),
.B(n_1875),
.C(n_1860),
.Y(n_1944)
);

INVx1_ASAP7_75t_L g1945 ( 
.A(n_1912),
.Y(n_1945)
);

HB1xp67_ASAP7_75t_L g1946 ( 
.A(n_1937),
.Y(n_1946)
);

AND4x1_ASAP7_75t_L g1947 ( 
.A(n_1927),
.B(n_1878),
.C(n_1861),
.D(n_1901),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1912),
.Y(n_1948)
);

AND2x2_ASAP7_75t_L g1949 ( 
.A(n_1933),
.B(n_1908),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1916),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1916),
.Y(n_1951)
);

AND2x4_ASAP7_75t_L g1952 ( 
.A(n_1933),
.B(n_1879),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1933),
.B(n_1879),
.Y(n_1953)
);

NAND2x1_ASAP7_75t_L g1954 ( 
.A(n_1917),
.B(n_1879),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1916),
.Y(n_1955)
);

NOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1924),
.B(n_1879),
.Y(n_1956)
);

HB1xp67_ASAP7_75t_L g1957 ( 
.A(n_1937),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1921),
.Y(n_1958)
);

INVx1_ASAP7_75t_L g1959 ( 
.A(n_1914),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1914),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1915),
.B(n_1906),
.Y(n_1961)
);

AOI33xp33_ASAP7_75t_L g1962 ( 
.A1(n_1927),
.A2(n_1911),
.A3(n_1910),
.B1(n_1928),
.B2(n_1918),
.B3(n_842),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1915),
.B(n_1906),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1910),
.Y(n_1964)
);

INVx2_ASAP7_75t_L g1965 ( 
.A(n_1921),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1931),
.B(n_1909),
.Y(n_1966)
);

INVx1_ASAP7_75t_SL g1967 ( 
.A(n_1917),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1927),
.B(n_1893),
.Y(n_1968)
);

AND2x2_ASAP7_75t_L g1969 ( 
.A(n_1931),
.B(n_1899),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1923),
.B(n_1887),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1911),
.Y(n_1971)
);

NOR2xp33_ASAP7_75t_L g1972 ( 
.A(n_1939),
.B(n_1729),
.Y(n_1972)
);

OAI31xp33_ASAP7_75t_L g1973 ( 
.A1(n_1939),
.A2(n_1895),
.A3(n_1902),
.B(n_1859),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1949),
.B(n_1931),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1946),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1943),
.Y(n_1976)
);

INVx2_ASAP7_75t_SL g1977 ( 
.A(n_1943),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1949),
.B(n_1917),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_L g1979 ( 
.A(n_1962),
.B(n_1942),
.Y(n_1979)
);

HB1xp67_ASAP7_75t_L g1980 ( 
.A(n_1946),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1957),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_L g1982 ( 
.A(n_1967),
.B(n_1942),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1956),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1973),
.B(n_1942),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_L g1985 ( 
.A(n_1967),
.B(n_1920),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1947),
.B(n_1920),
.Y(n_1986)
);

AND2x4_ASAP7_75t_L g1987 ( 
.A(n_1956),
.B(n_1917),
.Y(n_1987)
);

OR2x2_ASAP7_75t_L g1988 ( 
.A(n_1968),
.B(n_1913),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1968),
.B(n_1913),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1947),
.B(n_1925),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1953),
.B(n_1943),
.Y(n_1991)
);

INVx2_ASAP7_75t_L g1992 ( 
.A(n_1943),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1953),
.B(n_1952),
.Y(n_1993)
);

CKINVDCx5p33_ASAP7_75t_R g1994 ( 
.A(n_1972),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1943),
.B(n_1952),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1952),
.B(n_1925),
.Y(n_1996)
);

OAI21xp5_ASAP7_75t_SL g1997 ( 
.A1(n_1944),
.A2(n_1895),
.B(n_1902),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1945),
.Y(n_1998)
);

NAND2xp5_ASAP7_75t_L g1999 ( 
.A(n_1943),
.B(n_1952),
.Y(n_1999)
);

INVx4_ASAP7_75t_SL g2000 ( 
.A(n_1964),
.Y(n_2000)
);

AND2x2_ASAP7_75t_L g2001 ( 
.A(n_1961),
.B(n_1926),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1950),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1950),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1961),
.B(n_1926),
.Y(n_2004)
);

INVx2_ASAP7_75t_L g2005 ( 
.A(n_1950),
.Y(n_2005)
);

AND2x2_ASAP7_75t_L g2006 ( 
.A(n_1963),
.B(n_1940),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1945),
.Y(n_2007)
);

AOI22xp33_ASAP7_75t_L g2008 ( 
.A1(n_1973),
.A2(n_1866),
.B1(n_1940),
.B2(n_1816),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1948),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1963),
.B(n_1918),
.Y(n_2010)
);

OR2x2_ASAP7_75t_L g2011 ( 
.A(n_1970),
.B(n_1964),
.Y(n_2011)
);

INVx2_ASAP7_75t_L g2012 ( 
.A(n_1951),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1966),
.B(n_1928),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1951),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1948),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1959),
.Y(n_2016)
);

INVx2_ASAP7_75t_L g2017 ( 
.A(n_1951),
.Y(n_2017)
);

INVxp67_ASAP7_75t_SL g2018 ( 
.A(n_1983),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1980),
.B(n_1971),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1975),
.Y(n_2020)
);

INVx1_ASAP7_75t_SL g2021 ( 
.A(n_1993),
.Y(n_2021)
);

AOI22xp33_ASAP7_75t_L g2022 ( 
.A1(n_1984),
.A2(n_1954),
.B1(n_1971),
.B2(n_1960),
.Y(n_2022)
);

INVx2_ASAP7_75t_L g2023 ( 
.A(n_1987),
.Y(n_2023)
);

AND2x2_ASAP7_75t_L g2024 ( 
.A(n_1993),
.B(n_1978),
.Y(n_2024)
);

AND2x2_ASAP7_75t_L g2025 ( 
.A(n_1978),
.B(n_1966),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1996),
.B(n_1969),
.Y(n_2026)
);

INVx2_ASAP7_75t_L g2027 ( 
.A(n_1987),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1987),
.Y(n_2028)
);

NOR2x1_ASAP7_75t_L g2029 ( 
.A(n_1975),
.B(n_1954),
.Y(n_2029)
);

NOR2xp33_ASAP7_75t_L g2030 ( 
.A(n_1994),
.B(n_1944),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_2011),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1996),
.B(n_1969),
.Y(n_2032)
);

OAI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1997),
.A2(n_1960),
.B(n_1959),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_2011),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1987),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1998),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1974),
.B(n_1970),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1998),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1981),
.B(n_1986),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1974),
.B(n_1899),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_2007),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2001),
.B(n_1900),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_2007),
.Y(n_2043)
);

OR2x2_ASAP7_75t_L g2044 ( 
.A(n_1985),
.B(n_1923),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1981),
.B(n_1955),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2009),
.Y(n_2046)
);

CKINVDCx5p33_ASAP7_75t_R g2047 ( 
.A(n_1995),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1990),
.B(n_1955),
.Y(n_2048)
);

AND2x4_ASAP7_75t_L g2049 ( 
.A(n_1977),
.B(n_1976),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_2001),
.B(n_1900),
.Y(n_2050)
);

NOR2xp33_ASAP7_75t_L g2051 ( 
.A(n_1979),
.B(n_1991),
.Y(n_2051)
);

INVx2_ASAP7_75t_L g2052 ( 
.A(n_1977),
.Y(n_2052)
);

INVx4_ASAP7_75t_L g2053 ( 
.A(n_1976),
.Y(n_2053)
);

OR2x2_ASAP7_75t_L g2054 ( 
.A(n_2004),
.B(n_1894),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1999),
.B(n_1894),
.Y(n_2055)
);

CKINVDCx16_ASAP7_75t_R g2056 ( 
.A(n_1976),
.Y(n_2056)
);

NAND2x1p5_ASAP7_75t_L g2057 ( 
.A(n_1992),
.B(n_1715),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_2006),
.B(n_1887),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_L g2059 ( 
.A(n_1992),
.B(n_1955),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_2009),
.Y(n_2060)
);

INVxp33_ASAP7_75t_L g2061 ( 
.A(n_1982),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2015),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1992),
.B(n_1958),
.Y(n_2063)
);

NAND2x1p5_ASAP7_75t_L g2064 ( 
.A(n_2002),
.B(n_1715),
.Y(n_2064)
);

INVxp67_ASAP7_75t_L g2065 ( 
.A(n_2015),
.Y(n_2065)
);

INVx1_ASAP7_75t_L g2066 ( 
.A(n_2016),
.Y(n_2066)
);

INVx1_ASAP7_75t_L g2067 ( 
.A(n_2016),
.Y(n_2067)
);

INVx1_ASAP7_75t_SL g2068 ( 
.A(n_2010),
.Y(n_2068)
);

AND2x2_ASAP7_75t_L g2069 ( 
.A(n_2006),
.B(n_2010),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2000),
.Y(n_2070)
);

OR2x2_ASAP7_75t_L g2071 ( 
.A(n_2013),
.B(n_1919),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2000),
.Y(n_2072)
);

AND2x2_ASAP7_75t_L g2073 ( 
.A(n_2008),
.B(n_1958),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2000),
.B(n_1958),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_L g2075 ( 
.A(n_2000),
.B(n_1965),
.Y(n_2075)
);

OR2x2_ASAP7_75t_L g2076 ( 
.A(n_1988),
.B(n_1919),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_2000),
.B(n_1965),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1988),
.B(n_1965),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1997),
.B(n_1934),
.Y(n_2079)
);

AOI22xp5_ASAP7_75t_L g2080 ( 
.A1(n_1989),
.A2(n_1874),
.B1(n_1871),
.B2(n_1843),
.Y(n_2080)
);

OR2x2_ASAP7_75t_L g2081 ( 
.A(n_1989),
.B(n_1938),
.Y(n_2081)
);

OAI21xp33_ASAP7_75t_L g2082 ( 
.A1(n_2030),
.A2(n_2003),
.B(n_2002),
.Y(n_2082)
);

AND2x2_ASAP7_75t_L g2083 ( 
.A(n_2024),
.B(n_2002),
.Y(n_2083)
);

OAI21xp33_ASAP7_75t_L g2084 ( 
.A1(n_2030),
.A2(n_2005),
.B(n_2003),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2021),
.B(n_2003),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2068),
.Y(n_2086)
);

NAND2x1p5_ASAP7_75t_L g2087 ( 
.A(n_2029),
.B(n_2005),
.Y(n_2087)
);

NAND2xp5_ASAP7_75t_L g2088 ( 
.A(n_2056),
.B(n_2005),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_2035),
.Y(n_2089)
);

AO221x1_ASAP7_75t_L g2090 ( 
.A1(n_2023),
.A2(n_2017),
.B1(n_2014),
.B2(n_2012),
.C(n_1936),
.Y(n_2090)
);

AND2x4_ASAP7_75t_L g2091 ( 
.A(n_2027),
.B(n_2012),
.Y(n_2091)
);

OR2x2_ASAP7_75t_L g2092 ( 
.A(n_2039),
.B(n_2079),
.Y(n_2092)
);

OAI21xp5_ASAP7_75t_SL g2093 ( 
.A1(n_2022),
.A2(n_831),
.B(n_828),
.Y(n_2093)
);

AOI211xp5_ASAP7_75t_L g2094 ( 
.A1(n_2033),
.A2(n_893),
.B(n_902),
.C(n_869),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2018),
.Y(n_2095)
);

AOI21xp33_ASAP7_75t_L g2096 ( 
.A1(n_2061),
.A2(n_2014),
.B(n_2012),
.Y(n_2096)
);

OR2x2_ASAP7_75t_L g2097 ( 
.A(n_2039),
.B(n_2014),
.Y(n_2097)
);

AND2x4_ASAP7_75t_L g2098 ( 
.A(n_2028),
.B(n_2017),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_2018),
.Y(n_2099)
);

AOI22xp33_ASAP7_75t_L g2100 ( 
.A1(n_2073),
.A2(n_2017),
.B1(n_1816),
.B2(n_1821),
.Y(n_2100)
);

O2A1O1Ixp33_ASAP7_75t_L g2101 ( 
.A1(n_2022),
.A2(n_842),
.B(n_848),
.C(n_838),
.Y(n_2101)
);

AND2x4_ASAP7_75t_SL g2102 ( 
.A(n_2037),
.B(n_1705),
.Y(n_2102)
);

OR2x2_ASAP7_75t_L g2103 ( 
.A(n_2079),
.B(n_1938),
.Y(n_2103)
);

INVx1_ASAP7_75t_SL g2104 ( 
.A(n_2069),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2048),
.B(n_1934),
.Y(n_2105)
);

OAI21xp33_ASAP7_75t_L g2106 ( 
.A1(n_2061),
.A2(n_1941),
.B(n_1936),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2026),
.B(n_1941),
.Y(n_2107)
);

AOI22xp5_ASAP7_75t_L g2108 ( 
.A1(n_2051),
.A2(n_850),
.B1(n_854),
.B2(n_848),
.Y(n_2108)
);

AOI22xp5_ASAP7_75t_L g2109 ( 
.A1(n_2051),
.A2(n_854),
.B1(n_855),
.B2(n_850),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2031),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_2034),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2052),
.B(n_1935),
.Y(n_2112)
);

INVx1_ASAP7_75t_L g2113 ( 
.A(n_2049),
.Y(n_2113)
);

AND2x2_ASAP7_75t_L g2114 ( 
.A(n_2032),
.B(n_1935),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2049),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_2048),
.B(n_1935),
.Y(n_2116)
);

AOI32xp33_ASAP7_75t_L g2117 ( 
.A1(n_2025),
.A2(n_1893),
.A3(n_1904),
.B1(n_1885),
.B2(n_1921),
.Y(n_2117)
);

INVx1_ASAP7_75t_SL g2118 ( 
.A(n_2047),
.Y(n_2118)
);

AOI21xp5_ASAP7_75t_L g2119 ( 
.A1(n_2019),
.A2(n_856),
.B(n_855),
.Y(n_2119)
);

AND2x4_ASAP7_75t_SL g2120 ( 
.A(n_2053),
.B(n_2070),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_2053),
.Y(n_2121)
);

NAND2xp5_ASAP7_75t_SL g2122 ( 
.A(n_2044),
.B(n_1881),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2059),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_2058),
.B(n_1885),
.Y(n_2124)
);

INVx1_ASAP7_75t_SL g2125 ( 
.A(n_2078),
.Y(n_2125)
);

INVxp33_ASAP7_75t_L g2126 ( 
.A(n_2055),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2059),
.Y(n_2127)
);

AOI21xp5_ASAP7_75t_L g2128 ( 
.A1(n_2019),
.A2(n_2045),
.B(n_2065),
.Y(n_2128)
);

INVx1_ASAP7_75t_L g2129 ( 
.A(n_2063),
.Y(n_2129)
);

AOI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_2054),
.A2(n_1817),
.B1(n_1821),
.B2(n_1835),
.Y(n_2130)
);

INVxp67_ASAP7_75t_L g2131 ( 
.A(n_2074),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2080),
.A2(n_1885),
.B1(n_1821),
.B2(n_1817),
.Y(n_2132)
);

NAND2xp5_ASAP7_75t_L g2133 ( 
.A(n_2020),
.B(n_1881),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2072),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2042),
.A2(n_1929),
.B(n_1922),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2050),
.B(n_856),
.Y(n_2136)
);

OAI21xp33_ASAP7_75t_L g2137 ( 
.A1(n_2040),
.A2(n_1929),
.B(n_1922),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_2063),
.Y(n_2138)
);

OAI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_2064),
.A2(n_1835),
.B1(n_1854),
.B2(n_1823),
.Y(n_2139)
);

INVx1_ASAP7_75t_SL g2140 ( 
.A(n_2057),
.Y(n_2140)
);

OAI221xp5_ASAP7_75t_SL g2141 ( 
.A1(n_2071),
.A2(n_2076),
.B1(n_2081),
.B2(n_2065),
.C(n_2045),
.Y(n_2141)
);

NAND3xp33_ASAP7_75t_SL g2142 ( 
.A(n_2064),
.B(n_681),
.C(n_679),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_2036),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2038),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2041),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2057),
.B(n_2043),
.Y(n_2146)
);

AND2x2_ASAP7_75t_L g2147 ( 
.A(n_2046),
.B(n_1922),
.Y(n_2147)
);

OAI322xp33_ASAP7_75t_L g2148 ( 
.A1(n_2060),
.A2(n_1932),
.A3(n_1929),
.B1(n_1930),
.B2(n_1904),
.C1(n_868),
.C2(n_866),
.Y(n_2148)
);

AOI322xp5_ASAP7_75t_L g2149 ( 
.A1(n_2062),
.A2(n_866),
.A3(n_863),
.B1(n_868),
.B2(n_869),
.C1(n_865),
.C2(n_859),
.Y(n_2149)
);

NOR2xp33_ASAP7_75t_L g2150 ( 
.A(n_2066),
.B(n_859),
.Y(n_2150)
);

INVx2_ASAP7_75t_L g2151 ( 
.A(n_2077),
.Y(n_2151)
);

AND2x2_ASAP7_75t_L g2152 ( 
.A(n_2067),
.B(n_1930),
.Y(n_2152)
);

INVx1_ASAP7_75t_L g2153 ( 
.A(n_2075),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2075),
.Y(n_2154)
);

AOI21xp33_ASAP7_75t_SL g2155 ( 
.A1(n_2077),
.A2(n_865),
.B(n_863),
.Y(n_2155)
);

OR2x2_ASAP7_75t_L g2156 ( 
.A(n_2039),
.B(n_1930),
.Y(n_2156)
);

INVx1_ASAP7_75t_SL g2157 ( 
.A(n_2024),
.Y(n_2157)
);

O2A1O1Ixp33_ASAP7_75t_L g2158 ( 
.A1(n_2039),
.A2(n_875),
.B(n_878),
.C(n_873),
.Y(n_2158)
);

AOI31xp33_ASAP7_75t_L g2159 ( 
.A1(n_2022),
.A2(n_875),
.A3(n_878),
.B(n_873),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2018),
.Y(n_2160)
);

OAI21xp33_ASAP7_75t_L g2161 ( 
.A1(n_2030),
.A2(n_1932),
.B(n_1842),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2021),
.B(n_886),
.Y(n_2162)
);

AOI21xp33_ASAP7_75t_SL g2163 ( 
.A1(n_2030),
.A2(n_887),
.B(n_886),
.Y(n_2163)
);

NOR2xp33_ASAP7_75t_L g2164 ( 
.A(n_2030),
.B(n_887),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2021),
.B(n_889),
.Y(n_2165)
);

AOI22xp5_ASAP7_75t_L g2166 ( 
.A1(n_2030),
.A2(n_1842),
.B1(n_1854),
.B2(n_1779),
.Y(n_2166)
);

AOI22xp5_ASAP7_75t_SL g2167 ( 
.A1(n_2018),
.A2(n_891),
.B1(n_893),
.B2(n_889),
.Y(n_2167)
);

OR2x2_ASAP7_75t_L g2168 ( 
.A(n_2039),
.B(n_1932),
.Y(n_2168)
);

OAI21xp5_ASAP7_75t_SL g2169 ( 
.A1(n_2126),
.A2(n_902),
.B(n_891),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_2157),
.B(n_2104),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2113),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2118),
.B(n_1817),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_2087),
.Y(n_2173)
);

NAND4xp25_ASAP7_75t_SL g2174 ( 
.A(n_2086),
.B(n_904),
.C(n_911),
.D(n_903),
.Y(n_2174)
);

CKINVDCx14_ASAP7_75t_R g2175 ( 
.A(n_2095),
.Y(n_2175)
);

AOI22xp5_ASAP7_75t_L g2176 ( 
.A1(n_2125),
.A2(n_1842),
.B1(n_1854),
.B2(n_1779),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_L g2177 ( 
.A(n_2115),
.Y(n_2177)
);

AND2x2_ASAP7_75t_L g2178 ( 
.A(n_2089),
.B(n_1842),
.Y(n_2178)
);

INVx1_ASAP7_75t_SL g2179 ( 
.A(n_2083),
.Y(n_2179)
);

OAI22xp33_ASAP7_75t_L g2180 ( 
.A1(n_2159),
.A2(n_1854),
.B1(n_1835),
.B2(n_1823),
.Y(n_2180)
);

AOI21xp33_ASAP7_75t_L g2181 ( 
.A1(n_2092),
.A2(n_904),
.B(n_903),
.Y(n_2181)
);

AOI21xp5_ASAP7_75t_L g2182 ( 
.A1(n_2128),
.A2(n_921),
.B(n_911),
.Y(n_2182)
);

OAI22xp5_ASAP7_75t_L g2183 ( 
.A1(n_2100),
.A2(n_1839),
.B1(n_1842),
.B2(n_1835),
.Y(n_2183)
);

OAI22xp5_ASAP7_75t_L g2184 ( 
.A1(n_2141),
.A2(n_1839),
.B1(n_1835),
.B2(n_1846),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_2099),
.A2(n_1846),
.B1(n_1825),
.B2(n_1827),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_L g2186 ( 
.A(n_2131),
.B(n_2120),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_2091),
.Y(n_2187)
);

AND2x2_ASAP7_75t_L g2188 ( 
.A(n_2102),
.B(n_921),
.Y(n_2188)
);

INVxp67_ASAP7_75t_L g2189 ( 
.A(n_2088),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_2091),
.Y(n_2190)
);

INVx1_ASAP7_75t_L g2191 ( 
.A(n_2098),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2160),
.B(n_923),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_2140),
.B(n_1803),
.Y(n_2193)
);

INVx2_ASAP7_75t_SL g2194 ( 
.A(n_2121),
.Y(n_2194)
);

NOR2x1_ASAP7_75t_L g2195 ( 
.A(n_2093),
.B(n_923),
.Y(n_2195)
);

INVx3_ASAP7_75t_SL g2196 ( 
.A(n_2167),
.Y(n_2196)
);

AOI22xp33_ASAP7_75t_L g2197 ( 
.A1(n_2164),
.A2(n_1720),
.B1(n_1837),
.B2(n_1798),
.Y(n_2197)
);

NAND2xp5_ASAP7_75t_L g2198 ( 
.A(n_2134),
.B(n_926),
.Y(n_2198)
);

OAI22xp5_ASAP7_75t_L g2199 ( 
.A1(n_2130),
.A2(n_2103),
.B1(n_2094),
.B2(n_2108),
.Y(n_2199)
);

AOI31xp33_ASAP7_75t_L g2200 ( 
.A1(n_2085),
.A2(n_927),
.A3(n_928),
.B(n_926),
.Y(n_2200)
);

AOI221xp5_ASAP7_75t_L g2201 ( 
.A1(n_2082),
.A2(n_929),
.B1(n_942),
.B2(n_928),
.C(n_927),
.Y(n_2201)
);

XOR2x2_ASAP7_75t_L g2202 ( 
.A(n_2142),
.B(n_2),
.Y(n_2202)
);

OR2x2_ASAP7_75t_L g2203 ( 
.A(n_2110),
.B(n_929),
.Y(n_2203)
);

AOI22xp5_ASAP7_75t_L g2204 ( 
.A1(n_2132),
.A2(n_943),
.B1(n_945),
.B2(n_942),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2098),
.Y(n_2205)
);

NAND2xp5_ASAP7_75t_SL g2206 ( 
.A(n_2146),
.B(n_1803),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_2151),
.Y(n_2207)
);

OAI221xp5_ASAP7_75t_SL g2208 ( 
.A1(n_2084),
.A2(n_948),
.B1(n_951),
.B2(n_945),
.C(n_943),
.Y(n_2208)
);

OAI221xp5_ASAP7_75t_L g2209 ( 
.A1(n_2101),
.A2(n_958),
.B1(n_959),
.B2(n_951),
.C(n_948),
.Y(n_2209)
);

AOI222xp33_ASAP7_75t_L g2210 ( 
.A1(n_2090),
.A2(n_958),
.B1(n_977),
.B2(n_985),
.C1(n_984),
.C2(n_959),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2153),
.Y(n_2211)
);

AOI22x1_ASAP7_75t_L g2212 ( 
.A1(n_2111),
.A2(n_684),
.B1(n_764),
.B2(n_747),
.Y(n_2212)
);

AOI22xp5_ASAP7_75t_L g2213 ( 
.A1(n_2161),
.A2(n_984),
.B1(n_985),
.B2(n_977),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2154),
.Y(n_2214)
);

OAI221xp5_ASAP7_75t_L g2215 ( 
.A1(n_2096),
.A2(n_1001),
.B1(n_1004),
.B2(n_999),
.C(n_997),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2097),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_2136),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_2143),
.B(n_1803),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_2124),
.B(n_997),
.Y(n_2219)
);

AOI22xp5_ASAP7_75t_L g2220 ( 
.A1(n_2114),
.A2(n_2107),
.B1(n_2106),
.B2(n_2108),
.Y(n_2220)
);

AOI22xp5_ASAP7_75t_L g2221 ( 
.A1(n_2109),
.A2(n_1001),
.B1(n_1004),
.B2(n_999),
.Y(n_2221)
);

NAND3xp33_ASAP7_75t_L g2222 ( 
.A(n_2149),
.B(n_2109),
.C(n_2117),
.Y(n_2222)
);

AOI22xp5_ASAP7_75t_L g2223 ( 
.A1(n_2166),
.A2(n_1019),
.B1(n_1023),
.B2(n_1015),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_2112),
.Y(n_2224)
);

O2A1O1Ixp33_ASAP7_75t_L g2225 ( 
.A1(n_2158),
.A2(n_1019),
.B(n_1031),
.C(n_1024),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2147),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_2122),
.A2(n_1023),
.B1(n_1024),
.B2(n_1015),
.Y(n_2227)
);

AOI22xp5_ASAP7_75t_L g2228 ( 
.A1(n_2123),
.A2(n_1032),
.B1(n_1031),
.B2(n_1846),
.Y(n_2228)
);

OAI22xp33_ASAP7_75t_L g2229 ( 
.A1(n_2156),
.A2(n_1846),
.B1(n_1828),
.B2(n_1834),
.Y(n_2229)
);

AOI221xp5_ASAP7_75t_L g2230 ( 
.A1(n_2148),
.A2(n_1032),
.B1(n_785),
.B2(n_808),
.C(n_773),
.Y(n_2230)
);

AOI22xp5_ASAP7_75t_L g2231 ( 
.A1(n_2127),
.A2(n_2129),
.B1(n_2138),
.B2(n_2144),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_2162),
.B(n_688),
.Y(n_2232)
);

OAI32xp33_ASAP7_75t_L g2233 ( 
.A1(n_2168),
.A2(n_785),
.A3(n_808),
.B1(n_773),
.B2(n_764),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2152),
.Y(n_2234)
);

OAI22xp5_ASAP7_75t_L g2235 ( 
.A1(n_2116),
.A2(n_1846),
.B1(n_1814),
.B2(n_1827),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_2145),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_2165),
.B(n_690),
.Y(n_2237)
);

AOI22xp5_ASAP7_75t_L g2238 ( 
.A1(n_2150),
.A2(n_1846),
.B1(n_876),
.B2(n_953),
.Y(n_2238)
);

O2A1O1Ixp33_ASAP7_75t_L g2239 ( 
.A1(n_2163),
.A2(n_918),
.B(n_953),
.C(n_876),
.Y(n_2239)
);

NOR2xp67_ASAP7_75t_L g2240 ( 
.A(n_2105),
.B(n_3),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2133),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_2155),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2155),
.Y(n_2243)
);

OR2x2_ASAP7_75t_L g2244 ( 
.A(n_2119),
.B(n_2),
.Y(n_2244)
);

OAI32xp33_ASAP7_75t_L g2245 ( 
.A1(n_2135),
.A2(n_986),
.A3(n_976),
.B1(n_918),
.B2(n_1718),
.Y(n_2245)
);

OAI21xp5_ASAP7_75t_L g2246 ( 
.A1(n_2163),
.A2(n_986),
.B(n_976),
.Y(n_2246)
);

INVxp67_ASAP7_75t_L g2247 ( 
.A(n_2137),
.Y(n_2247)
);

O2A1O1Ixp33_ASAP7_75t_L g2248 ( 
.A1(n_2139),
.A2(n_1739),
.B(n_1718),
.C(n_839),
.Y(n_2248)
);

OAI33xp33_ASAP7_75t_L g2249 ( 
.A1(n_2092),
.A2(n_700),
.A3(n_698),
.B1(n_701),
.B2(n_699),
.B3(n_697),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2157),
.B(n_1803),
.Y(n_2250)
);

NOR2xp33_ASAP7_75t_L g2251 ( 
.A(n_2118),
.B(n_704),
.Y(n_2251)
);

AND2x2_ASAP7_75t_L g2252 ( 
.A(n_2157),
.B(n_1795),
.Y(n_2252)
);

OA21x2_ASAP7_75t_L g2253 ( 
.A1(n_2128),
.A2(n_707),
.B(n_706),
.Y(n_2253)
);

INVx1_ASAP7_75t_L g2254 ( 
.A(n_2113),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_2157),
.B(n_712),
.Y(n_2255)
);

O2A1O1Ixp33_ASAP7_75t_SL g2256 ( 
.A1(n_2092),
.A2(n_1718),
.B(n_882),
.C(n_1010),
.Y(n_2256)
);

INVx1_ASAP7_75t_L g2257 ( 
.A(n_2113),
.Y(n_2257)
);

INVx1_ASAP7_75t_L g2258 ( 
.A(n_2113),
.Y(n_2258)
);

INVx1_ASAP7_75t_L g2259 ( 
.A(n_2113),
.Y(n_2259)
);

NOR2xp33_ASAP7_75t_L g2260 ( 
.A(n_2118),
.B(n_714),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_2118),
.B(n_720),
.Y(n_2261)
);

INVxp67_ASAP7_75t_L g2262 ( 
.A(n_2088),
.Y(n_2262)
);

AND2x2_ASAP7_75t_L g2263 ( 
.A(n_2157),
.B(n_1795),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_2113),
.Y(n_2264)
);

OAI22xp33_ASAP7_75t_L g2265 ( 
.A1(n_2087),
.A2(n_1828),
.B1(n_1834),
.B2(n_1830),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2113),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2157),
.B(n_1799),
.Y(n_2267)
);

OR2x2_ASAP7_75t_L g2268 ( 
.A(n_2104),
.B(n_3),
.Y(n_2268)
);

AOI21xp33_ASAP7_75t_SL g2269 ( 
.A1(n_2159),
.A2(n_722),
.B(n_721),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2118),
.B(n_724),
.Y(n_2270)
);

AOI22xp5_ASAP7_75t_SL g2271 ( 
.A1(n_2087),
.A2(n_726),
.B1(n_734),
.B2(n_731),
.Y(n_2271)
);

AOI22xp5_ASAP7_75t_L g2272 ( 
.A1(n_2157),
.A2(n_713),
.B1(n_1010),
.B2(n_882),
.Y(n_2272)
);

OAI31xp33_ASAP7_75t_L g2273 ( 
.A1(n_2087),
.A2(n_1837),
.A3(n_1694),
.B(n_1724),
.Y(n_2273)
);

INVxp67_ASAP7_75t_L g2274 ( 
.A(n_2088),
.Y(n_2274)
);

NAND2x1_ASAP7_75t_SL g2275 ( 
.A(n_2113),
.B(n_1724),
.Y(n_2275)
);

AOI222xp33_ASAP7_75t_L g2276 ( 
.A1(n_2090),
.A2(n_1030),
.B1(n_713),
.B2(n_1025),
.C1(n_1010),
.C2(n_738),
.Y(n_2276)
);

INVx1_ASAP7_75t_L g2277 ( 
.A(n_2113),
.Y(n_2277)
);

OAI22xp33_ASAP7_75t_SL g2278 ( 
.A1(n_2087),
.A2(n_737),
.B1(n_740),
.B2(n_739),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_2087),
.Y(n_2279)
);

OAI32xp33_ASAP7_75t_L g2280 ( 
.A1(n_2087),
.A2(n_1830),
.A3(n_1841),
.B1(n_1834),
.B2(n_1828),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2157),
.B(n_1799),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2113),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_2087),
.A2(n_1825),
.B1(n_1827),
.B2(n_1837),
.Y(n_2283)
);

AOI332xp33_ASAP7_75t_L g2284 ( 
.A1(n_2095),
.A2(n_1025),
.A3(n_1030),
.B1(n_713),
.B2(n_10),
.B3(n_6),
.C1(n_9),
.C2(n_8),
.Y(n_2284)
);

INVxp67_ASAP7_75t_L g2285 ( 
.A(n_2088),
.Y(n_2285)
);

INVx1_ASAP7_75t_L g2286 ( 
.A(n_2113),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2113),
.Y(n_2287)
);

NOR2xp33_ASAP7_75t_L g2288 ( 
.A(n_2118),
.B(n_743),
.Y(n_2288)
);

INVx1_ASAP7_75t_L g2289 ( 
.A(n_2113),
.Y(n_2289)
);

HB1xp67_ASAP7_75t_L g2290 ( 
.A(n_2087),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2157),
.B(n_1799),
.Y(n_2291)
);

OR2x2_ASAP7_75t_L g2292 ( 
.A(n_2104),
.B(n_4),
.Y(n_2292)
);

INVx1_ASAP7_75t_L g2293 ( 
.A(n_2113),
.Y(n_2293)
);

OR2x2_ASAP7_75t_L g2294 ( 
.A(n_2104),
.B(n_5),
.Y(n_2294)
);

NAND3xp33_ASAP7_75t_L g2295 ( 
.A(n_2094),
.B(n_890),
.C(n_631),
.Y(n_2295)
);

INVx1_ASAP7_75t_SL g2296 ( 
.A(n_2157),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2113),
.Y(n_2297)
);

INVx1_ASAP7_75t_L g2298 ( 
.A(n_2113),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2157),
.B(n_744),
.Y(n_2299)
);

AOI21xp33_ASAP7_75t_SL g2300 ( 
.A1(n_2087),
.A2(n_5),
.B(n_6),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2113),
.Y(n_2301)
);

NAND2xp5_ASAP7_75t_L g2302 ( 
.A(n_2157),
.B(n_750),
.Y(n_2302)
);

OAI21xp5_ASAP7_75t_L g2303 ( 
.A1(n_2128),
.A2(n_752),
.B(n_751),
.Y(n_2303)
);

AOI22xp5_ASAP7_75t_L g2304 ( 
.A1(n_2157),
.A2(n_713),
.B1(n_1030),
.B2(n_1025),
.Y(n_2304)
);

OAI21xp5_ASAP7_75t_L g2305 ( 
.A1(n_2128),
.A2(n_755),
.B(n_753),
.Y(n_2305)
);

INVx1_ASAP7_75t_L g2306 ( 
.A(n_2113),
.Y(n_2306)
);

AOI22xp5_ASAP7_75t_L g2307 ( 
.A1(n_2157),
.A2(n_1025),
.B1(n_1030),
.B2(n_756),
.Y(n_2307)
);

INVxp67_ASAP7_75t_L g2308 ( 
.A(n_2088),
.Y(n_2308)
);

A2O1A1Ixp33_ASAP7_75t_L g2309 ( 
.A1(n_2128),
.A2(n_757),
.B(n_761),
.C(n_760),
.Y(n_2309)
);

NAND2xp5_ASAP7_75t_L g2310 ( 
.A(n_2157),
.B(n_762),
.Y(n_2310)
);

AOI21xp33_ASAP7_75t_SL g2311 ( 
.A1(n_2159),
.A2(n_767),
.B(n_766),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_2113),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_2113),
.Y(n_2313)
);

OR2x2_ASAP7_75t_L g2314 ( 
.A(n_2104),
.B(n_7),
.Y(n_2314)
);

O2A1O1Ixp33_ASAP7_75t_L g2315 ( 
.A1(n_2159),
.A2(n_1780),
.B(n_1837),
.C(n_1721),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2159),
.A2(n_770),
.B(n_769),
.Y(n_2316)
);

INVxp67_ASAP7_75t_SL g2317 ( 
.A(n_2087),
.Y(n_2317)
);

INVx1_ASAP7_75t_L g2318 ( 
.A(n_2113),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2179),
.B(n_771),
.Y(n_2319)
);

AOI322xp5_ASAP7_75t_L g2320 ( 
.A1(n_2175),
.A2(n_780),
.A3(n_777),
.B1(n_781),
.B2(n_786),
.C1(n_782),
.C2(n_779),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_2177),
.Y(n_2321)
);

OR2x2_ASAP7_75t_L g2322 ( 
.A(n_2296),
.B(n_7),
.Y(n_2322)
);

INVxp67_ASAP7_75t_L g2323 ( 
.A(n_2290),
.Y(n_2323)
);

OAI21xp33_ASAP7_75t_L g2324 ( 
.A1(n_2186),
.A2(n_811),
.B(n_795),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2187),
.Y(n_2325)
);

OAI31xp33_ASAP7_75t_L g2326 ( 
.A1(n_2222),
.A2(n_1694),
.A3(n_1834),
.B(n_1830),
.Y(n_2326)
);

NAND2xp5_ASAP7_75t_L g2327 ( 
.A(n_2170),
.B(n_788),
.Y(n_2327)
);

AOI221xp5_ASAP7_75t_L g2328 ( 
.A1(n_2247),
.A2(n_794),
.B1(n_799),
.B2(n_797),
.C(n_791),
.Y(n_2328)
);

AOI22xp5_ASAP7_75t_L g2329 ( 
.A1(n_2196),
.A2(n_2317),
.B1(n_2210),
.B2(n_2279),
.Y(n_2329)
);

NOR2x1p5_ASAP7_75t_L g2330 ( 
.A(n_2279),
.B(n_2171),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2276),
.A2(n_800),
.B1(n_804),
.B2(n_801),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_2190),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2191),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_L g2334 ( 
.A(n_2205),
.B(n_807),
.Y(n_2334)
);

INVx1_ASAP7_75t_SL g2335 ( 
.A(n_2275),
.Y(n_2335)
);

OAI31xp33_ASAP7_75t_L g2336 ( 
.A1(n_2256),
.A2(n_1841),
.A3(n_1844),
.B(n_1830),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2194),
.Y(n_2337)
);

OAI21xp5_ASAP7_75t_L g2338 ( 
.A1(n_2240),
.A2(n_835),
.B(n_820),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_2268),
.Y(n_2339)
);

BUFx3_ASAP7_75t_L g2340 ( 
.A(n_2172),
.Y(n_2340)
);

OAI22xp33_ASAP7_75t_L g2341 ( 
.A1(n_2300),
.A2(n_1841),
.B1(n_1844),
.B2(n_1822),
.Y(n_2341)
);

NAND2xp5_ASAP7_75t_L g2342 ( 
.A(n_2254),
.B(n_810),
.Y(n_2342)
);

AOI21xp33_ASAP7_75t_L g2343 ( 
.A1(n_2278),
.A2(n_818),
.B(n_815),
.Y(n_2343)
);

NAND2xp5_ASAP7_75t_L g2344 ( 
.A(n_2257),
.B(n_821),
.Y(n_2344)
);

AOI22xp5_ASAP7_75t_L g2345 ( 
.A1(n_2202),
.A2(n_822),
.B1(n_827),
.B2(n_825),
.Y(n_2345)
);

NAND2xp5_ASAP7_75t_L g2346 ( 
.A(n_2258),
.B(n_832),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2292),
.Y(n_2347)
);

OAI32xp33_ASAP7_75t_SL g2348 ( 
.A1(n_2295),
.A2(n_12),
.A3(n_8),
.B1(n_9),
.B2(n_13),
.Y(n_2348)
);

AOI22xp5_ASAP7_75t_L g2349 ( 
.A1(n_2189),
.A2(n_2262),
.B1(n_2285),
.B2(n_2274),
.Y(n_2349)
);

INVx1_ASAP7_75t_SL g2350 ( 
.A(n_2294),
.Y(n_2350)
);

XOR2x2_ASAP7_75t_L g2351 ( 
.A(n_2271),
.B(n_14),
.Y(n_2351)
);

OAI22xp33_ASAP7_75t_L g2352 ( 
.A1(n_2173),
.A2(n_1844),
.B1(n_1841),
.B2(n_1831),
.Y(n_2352)
);

INVx1_ASAP7_75t_SL g2353 ( 
.A(n_2314),
.Y(n_2353)
);

NAND2xp5_ASAP7_75t_L g2354 ( 
.A(n_2318),
.B(n_833),
.Y(n_2354)
);

OAI211xp5_ASAP7_75t_L g2355 ( 
.A1(n_2284),
.A2(n_834),
.B(n_845),
.C(n_844),
.Y(n_2355)
);

INVx1_ASAP7_75t_L g2356 ( 
.A(n_2259),
.Y(n_2356)
);

INVx1_ASAP7_75t_L g2357 ( 
.A(n_2264),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2308),
.A2(n_1825),
.B1(n_1840),
.B2(n_1831),
.Y(n_2358)
);

AND2x2_ASAP7_75t_L g2359 ( 
.A(n_2266),
.B(n_1799),
.Y(n_2359)
);

NOR2x1_ASAP7_75t_SL g2360 ( 
.A(n_2216),
.B(n_1780),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2277),
.B(n_846),
.Y(n_2361)
);

INVx1_ASAP7_75t_SL g2362 ( 
.A(n_2282),
.Y(n_2362)
);

INVx1_ASAP7_75t_L g2363 ( 
.A(n_2286),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_L g2364 ( 
.A(n_2287),
.B(n_847),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2289),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_2293),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2297),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2298),
.Y(n_2368)
);

INVxp67_ASAP7_75t_SL g2369 ( 
.A(n_2253),
.Y(n_2369)
);

AOI22xp5_ASAP7_75t_SL g2370 ( 
.A1(n_2253),
.A2(n_853),
.B1(n_858),
.B2(n_857),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_2301),
.Y(n_2371)
);

INVx2_ASAP7_75t_L g2372 ( 
.A(n_2306),
.Y(n_2372)
);

NAND2xp5_ASAP7_75t_SL g2373 ( 
.A(n_2269),
.B(n_631),
.Y(n_2373)
);

INVxp33_ASAP7_75t_L g2374 ( 
.A(n_2251),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_2312),
.B(n_860),
.Y(n_2375)
);

OAI21xp5_ASAP7_75t_L g2376 ( 
.A1(n_2220),
.A2(n_896),
.B(n_864),
.Y(n_2376)
);

NOR2x1_ASAP7_75t_L g2377 ( 
.A(n_2174),
.B(n_890),
.Y(n_2377)
);

AND2x2_ASAP7_75t_L g2378 ( 
.A(n_2313),
.B(n_870),
.Y(n_2378)
);

AOI211x1_ASAP7_75t_L g2379 ( 
.A1(n_2193),
.A2(n_1840),
.B(n_1831),
.C(n_1802),
.Y(n_2379)
);

AND2x2_ASAP7_75t_L g2380 ( 
.A(n_2207),
.B(n_871),
.Y(n_2380)
);

OAI21xp33_ASAP7_75t_L g2381 ( 
.A1(n_2250),
.A2(n_2206),
.B(n_2204),
.Y(n_2381)
);

AOI21xp5_ASAP7_75t_L g2382 ( 
.A1(n_2303),
.A2(n_900),
.B(n_874),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2226),
.B(n_883),
.Y(n_2383)
);

OAI21xp33_ASAP7_75t_L g2384 ( 
.A1(n_2252),
.A2(n_894),
.B(n_888),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2234),
.Y(n_2385)
);

AOI21xp33_ASAP7_75t_SL g2386 ( 
.A1(n_2200),
.A2(n_14),
.B(n_15),
.Y(n_2386)
);

INVx2_ASAP7_75t_L g2387 ( 
.A(n_2219),
.Y(n_2387)
);

OAI21xp33_ASAP7_75t_L g2388 ( 
.A1(n_2263),
.A2(n_898),
.B(n_897),
.Y(n_2388)
);

OAI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2223),
.A2(n_1844),
.B1(n_1840),
.B2(n_899),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2242),
.B(n_901),
.Y(n_2390)
);

NOR2xp33_ASAP7_75t_L g2391 ( 
.A(n_2243),
.B(n_908),
.Y(n_2391)
);

INVx1_ASAP7_75t_L g2392 ( 
.A(n_2211),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2214),
.Y(n_2393)
);

AOI211xp5_ASAP7_75t_L g2394 ( 
.A1(n_2199),
.A2(n_909),
.B(n_944),
.C(n_930),
.Y(n_2394)
);

OAI221xp5_ASAP7_75t_SL g2395 ( 
.A1(n_2273),
.A2(n_1801),
.B1(n_1804),
.B2(n_1807),
.C(n_1805),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_2198),
.Y(n_2396)
);

NOR2xp67_ASAP7_75t_L g2397 ( 
.A(n_2231),
.B(n_15),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2217),
.B(n_910),
.Y(n_2398)
);

INVx2_ASAP7_75t_L g2399 ( 
.A(n_2188),
.Y(n_2399)
);

OAI31xp33_ASAP7_75t_SL g2400 ( 
.A1(n_2180),
.A2(n_19),
.A3(n_16),
.B(n_17),
.Y(n_2400)
);

NAND2xp5_ASAP7_75t_L g2401 ( 
.A(n_2269),
.B(n_912),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2305),
.A2(n_936),
.B(n_917),
.Y(n_2402)
);

NAND2x1_ASAP7_75t_L g2403 ( 
.A(n_2218),
.B(n_1683),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2203),
.Y(n_2404)
);

OAI31xp33_ASAP7_75t_L g2405 ( 
.A1(n_2309),
.A2(n_1801),
.A3(n_19),
.B(n_16),
.Y(n_2405)
);

NAND2x1_ASAP7_75t_L g2406 ( 
.A(n_2218),
.B(n_1683),
.Y(n_2406)
);

AOI221xp5_ASAP7_75t_L g2407 ( 
.A1(n_2208),
.A2(n_2315),
.B1(n_2236),
.B2(n_2230),
.C(n_2245),
.Y(n_2407)
);

OAI21xp5_ASAP7_75t_L g2408 ( 
.A1(n_2182),
.A2(n_955),
.B(n_924),
.Y(n_2408)
);

OR2x2_ASAP7_75t_L g2409 ( 
.A(n_2224),
.B(n_17),
.Y(n_2409)
);

OAI22xp33_ASAP7_75t_L g2410 ( 
.A1(n_2244),
.A2(n_914),
.B1(n_922),
.B2(n_920),
.Y(n_2410)
);

NAND3xp33_ASAP7_75t_SL g2411 ( 
.A(n_2311),
.B(n_932),
.C(n_931),
.Y(n_2411)
);

NOR2xp67_ASAP7_75t_SL g2412 ( 
.A(n_2169),
.B(n_947),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2192),
.Y(n_2413)
);

AND2x2_ASAP7_75t_L g2414 ( 
.A(n_2260),
.B(n_933),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2261),
.B(n_935),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2221),
.A2(n_937),
.B1(n_956),
.B2(n_938),
.Y(n_2416)
);

OR2x2_ASAP7_75t_L g2417 ( 
.A(n_2255),
.B(n_2299),
.Y(n_2417)
);

OAI321xp33_ASAP7_75t_L g2418 ( 
.A1(n_2183),
.A2(n_965),
.A3(n_979),
.B1(n_890),
.B2(n_1781),
.C(n_1804),
.Y(n_2418)
);

AND2x2_ASAP7_75t_L g2419 ( 
.A(n_2270),
.B(n_957),
.Y(n_2419)
);

AOI32xp33_ASAP7_75t_L g2420 ( 
.A1(n_2178),
.A2(n_1026),
.A3(n_1012),
.B1(n_993),
.B2(n_962),
.Y(n_2420)
);

INVx2_ASAP7_75t_L g2421 ( 
.A(n_2212),
.Y(n_2421)
);

INVx1_ASAP7_75t_SL g2422 ( 
.A(n_2302),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_SL g2423 ( 
.A(n_2311),
.B(n_890),
.Y(n_2423)
);

AOI21xp5_ASAP7_75t_L g2424 ( 
.A1(n_2310),
.A2(n_980),
.B(n_966),
.Y(n_2424)
);

OAI21xp5_ASAP7_75t_L g2425 ( 
.A1(n_2225),
.A2(n_987),
.B(n_967),
.Y(n_2425)
);

AOI21xp5_ASAP7_75t_L g2426 ( 
.A1(n_2288),
.A2(n_989),
.B(n_969),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2267),
.B(n_960),
.Y(n_2427)
);

INVx1_ASAP7_75t_SL g2428 ( 
.A(n_2195),
.Y(n_2428)
);

INVx1_ASAP7_75t_L g2429 ( 
.A(n_2241),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2239),
.Y(n_2430)
);

O2A1O1Ixp5_ASAP7_75t_L g2431 ( 
.A1(n_2184),
.A2(n_1781),
.B(n_1796),
.C(n_1794),
.Y(n_2431)
);

OAI22xp5_ASAP7_75t_L g2432 ( 
.A1(n_2307),
.A2(n_1805),
.B1(n_1806),
.B2(n_1802),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2227),
.Y(n_2433)
);

OR2x2_ASAP7_75t_L g2434 ( 
.A(n_2272),
.B(n_20),
.Y(n_2434)
);

NAND3xp33_ASAP7_75t_L g2435 ( 
.A(n_2201),
.B(n_963),
.C(n_961),
.Y(n_2435)
);

INVx1_ASAP7_75t_L g2436 ( 
.A(n_2246),
.Y(n_2436)
);

OR2x2_ASAP7_75t_L g2437 ( 
.A(n_2304),
.B(n_20),
.Y(n_2437)
);

OAI211xp5_ASAP7_75t_L g2438 ( 
.A1(n_2329),
.A2(n_2213),
.B(n_2228),
.C(n_2238),
.Y(n_2438)
);

INVxp67_ASAP7_75t_L g2439 ( 
.A(n_2321),
.Y(n_2439)
);

AOI22xp5_ASAP7_75t_L g2440 ( 
.A1(n_2323),
.A2(n_2281),
.B1(n_2291),
.B2(n_2249),
.Y(n_2440)
);

OAI21xp33_ASAP7_75t_L g2441 ( 
.A1(n_2329),
.A2(n_2176),
.B(n_2197),
.Y(n_2441)
);

OAI221xp5_ASAP7_75t_L g2442 ( 
.A1(n_2326),
.A2(n_2248),
.B1(n_2209),
.B2(n_2181),
.C(n_2215),
.Y(n_2442)
);

AOI211xp5_ASAP7_75t_L g2443 ( 
.A1(n_2397),
.A2(n_2233),
.B(n_2237),
.C(n_2232),
.Y(n_2443)
);

AOI22xp33_ASAP7_75t_L g2444 ( 
.A1(n_2340),
.A2(n_2283),
.B1(n_2265),
.B2(n_2185),
.Y(n_2444)
);

AOI21xp33_ASAP7_75t_L g2445 ( 
.A1(n_2374),
.A2(n_2280),
.B(n_2235),
.Y(n_2445)
);

AOI211xp5_ASAP7_75t_L g2446 ( 
.A1(n_2400),
.A2(n_2316),
.B(n_2229),
.C(n_971),
.Y(n_2446)
);

OR2x2_ASAP7_75t_L g2447 ( 
.A(n_2322),
.B(n_21),
.Y(n_2447)
);

AOI22xp33_ASAP7_75t_L g2448 ( 
.A1(n_2337),
.A2(n_1798),
.B1(n_965),
.B2(n_979),
.Y(n_2448)
);

NAND2xp5_ASAP7_75t_L g2449 ( 
.A(n_2330),
.B(n_970),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2325),
.Y(n_2450)
);

AOI21xp33_ASAP7_75t_L g2451 ( 
.A1(n_2350),
.A2(n_974),
.B(n_972),
.Y(n_2451)
);

OAI21xp5_ASAP7_75t_SL g2452 ( 
.A1(n_2349),
.A2(n_965),
.B(n_890),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2332),
.Y(n_2453)
);

AOI21xp5_ASAP7_75t_L g2454 ( 
.A1(n_2369),
.A2(n_988),
.B(n_981),
.Y(n_2454)
);

OAI211xp5_ASAP7_75t_L g2455 ( 
.A1(n_2349),
.A2(n_992),
.B(n_994),
.C(n_990),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2353),
.B(n_1000),
.Y(n_2456)
);

OAI21xp33_ASAP7_75t_L g2457 ( 
.A1(n_2381),
.A2(n_1005),
.B(n_1003),
.Y(n_2457)
);

AOI21xp33_ASAP7_75t_SL g2458 ( 
.A1(n_2339),
.A2(n_1007),
.B(n_1006),
.Y(n_2458)
);

AOI322xp5_ASAP7_75t_L g2459 ( 
.A1(n_2362),
.A2(n_1013),
.A3(n_1017),
.B1(n_1016),
.B2(n_1020),
.C1(n_1018),
.C2(n_1009),
.Y(n_2459)
);

OAI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2345),
.A2(n_1022),
.B1(n_1028),
.B2(n_1021),
.Y(n_2460)
);

AOI21xp5_ASAP7_75t_L g2461 ( 
.A1(n_2338),
.A2(n_2355),
.B(n_2373),
.Y(n_2461)
);

NAND2xp5_ASAP7_75t_SL g2462 ( 
.A(n_2386),
.B(n_965),
.Y(n_2462)
);

AOI22xp33_ASAP7_75t_L g2463 ( 
.A1(n_2433),
.A2(n_1798),
.B1(n_979),
.B2(n_965),
.Y(n_2463)
);

AOI211xp5_ASAP7_75t_L g2464 ( 
.A1(n_2335),
.A2(n_979),
.B(n_965),
.C(n_23),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_L g2465 ( 
.A(n_2347),
.B(n_21),
.Y(n_2465)
);

OAI211xp5_ASAP7_75t_SL g2466 ( 
.A1(n_2394),
.A2(n_24),
.B(n_22),
.C(n_23),
.Y(n_2466)
);

NOR3xp33_ASAP7_75t_L g2467 ( 
.A(n_2376),
.B(n_1089),
.C(n_1084),
.Y(n_2467)
);

AOI21xp5_ASAP7_75t_L g2468 ( 
.A1(n_2423),
.A2(n_979),
.B(n_1792),
.Y(n_2468)
);

INVx1_ASAP7_75t_L g2469 ( 
.A(n_2333),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2399),
.B(n_24),
.Y(n_2470)
);

AOI211xp5_ASAP7_75t_L g2471 ( 
.A1(n_2428),
.A2(n_979),
.B(n_27),
.C(n_25),
.Y(n_2471)
);

NAND3xp33_ASAP7_75t_SL g2472 ( 
.A(n_2405),
.B(n_28),
.C(n_26),
.Y(n_2472)
);

NAND3xp33_ASAP7_75t_L g2473 ( 
.A(n_2328),
.B(n_25),
.C(n_28),
.Y(n_2473)
);

AOI322xp5_ASAP7_75t_L g2474 ( 
.A1(n_2407),
.A2(n_1801),
.A3(n_1804),
.B1(n_1807),
.B2(n_1789),
.C1(n_1788),
.C2(n_1805),
.Y(n_2474)
);

AOI22xp5_ASAP7_75t_L g2475 ( 
.A1(n_2345),
.A2(n_1780),
.B1(n_1798),
.B2(n_1802),
.Y(n_2475)
);

AND2x2_ASAP7_75t_L g2476 ( 
.A(n_2387),
.B(n_1792),
.Y(n_2476)
);

AOI21xp5_ASAP7_75t_L g2477 ( 
.A1(n_2351),
.A2(n_1780),
.B(n_1766),
.Y(n_2477)
);

AOI221xp5_ASAP7_75t_L g2478 ( 
.A1(n_2348),
.A2(n_1798),
.B1(n_32),
.B2(n_29),
.C(n_30),
.Y(n_2478)
);

AOI22xp5_ASAP7_75t_L g2479 ( 
.A1(n_2385),
.A2(n_1798),
.B1(n_1810),
.B2(n_1806),
.Y(n_2479)
);

OAI22xp5_ASAP7_75t_L g2480 ( 
.A1(n_2422),
.A2(n_1810),
.B1(n_1811),
.B2(n_1806),
.Y(n_2480)
);

OAI21xp5_ASAP7_75t_SL g2481 ( 
.A1(n_2331),
.A2(n_33),
.B(n_34),
.Y(n_2481)
);

AOI22xp5_ASAP7_75t_L g2482 ( 
.A1(n_2359),
.A2(n_1811),
.B1(n_1812),
.B2(n_1810),
.Y(n_2482)
);

A2O1A1Ixp33_ASAP7_75t_L g2483 ( 
.A1(n_2370),
.A2(n_2391),
.B(n_2331),
.C(n_2336),
.Y(n_2483)
);

AOI221xp5_ASAP7_75t_L g2484 ( 
.A1(n_2341),
.A2(n_35),
.B1(n_33),
.B2(n_34),
.C(n_36),
.Y(n_2484)
);

NAND4xp25_ASAP7_75t_SL g2485 ( 
.A(n_2420),
.B(n_37),
.C(n_35),
.D(n_36),
.Y(n_2485)
);

AOI211xp5_ASAP7_75t_L g2486 ( 
.A1(n_2389),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2486)
);

OAI21xp33_ASAP7_75t_L g2487 ( 
.A1(n_2384),
.A2(n_1801),
.B(n_1804),
.Y(n_2487)
);

AOI221xp5_ASAP7_75t_L g2488 ( 
.A1(n_2356),
.A2(n_43),
.B1(n_40),
.B2(n_42),
.C(n_44),
.Y(n_2488)
);

OAI21xp5_ASAP7_75t_L g2489 ( 
.A1(n_2367),
.A2(n_1784),
.B(n_1773),
.Y(n_2489)
);

AOI221x1_ASAP7_75t_L g2490 ( 
.A1(n_2324),
.A2(n_45),
.B1(n_42),
.B2(n_44),
.C(n_46),
.Y(n_2490)
);

AOI221xp5_ASAP7_75t_L g2491 ( 
.A1(n_2357),
.A2(n_47),
.B1(n_45),
.B2(n_46),
.C(n_48),
.Y(n_2491)
);

OR2x2_ASAP7_75t_L g2492 ( 
.A(n_2372),
.B(n_49),
.Y(n_2492)
);

AND2x2_ASAP7_75t_L g2493 ( 
.A(n_2404),
.B(n_49),
.Y(n_2493)
);

AOI22xp5_ASAP7_75t_L g2494 ( 
.A1(n_2363),
.A2(n_1811),
.B1(n_1813),
.B2(n_1812),
.Y(n_2494)
);

OAI221xp5_ASAP7_75t_L g2495 ( 
.A1(n_2324),
.A2(n_1766),
.B1(n_1813),
.B2(n_1812),
.C(n_1796),
.Y(n_2495)
);

AOI22xp33_ASAP7_75t_L g2496 ( 
.A1(n_2436),
.A2(n_1824),
.B1(n_1807),
.B2(n_1789),
.Y(n_2496)
);

OAI21xp5_ASAP7_75t_SL g2497 ( 
.A1(n_2365),
.A2(n_50),
.B(n_51),
.Y(n_2497)
);

AOI22xp33_ASAP7_75t_L g2498 ( 
.A1(n_2430),
.A2(n_1824),
.B1(n_1807),
.B2(n_1788),
.Y(n_2498)
);

OAI22xp5_ASAP7_75t_L g2499 ( 
.A1(n_2366),
.A2(n_1813),
.B1(n_1794),
.B2(n_1797),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_2327),
.A2(n_1092),
.B(n_1089),
.Y(n_2500)
);

AOI221xp5_ASAP7_75t_L g2501 ( 
.A1(n_2368),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_2501)
);

OR2x2_ASAP7_75t_L g2502 ( 
.A(n_2371),
.B(n_52),
.Y(n_2502)
);

AOI22xp5_ASAP7_75t_L g2503 ( 
.A1(n_2396),
.A2(n_1818),
.B1(n_1826),
.B2(n_1815),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_2409),
.Y(n_2504)
);

OA22x2_ASAP7_75t_L g2505 ( 
.A1(n_2429),
.A2(n_1796),
.B1(n_1808),
.B2(n_1797),
.Y(n_2505)
);

OAI21xp33_ASAP7_75t_SL g2506 ( 
.A1(n_2392),
.A2(n_2393),
.B(n_2320),
.Y(n_2506)
);

AOI211xp5_ASAP7_75t_L g2507 ( 
.A1(n_2410),
.A2(n_57),
.B(n_54),
.C(n_55),
.Y(n_2507)
);

OR2x2_ASAP7_75t_L g2508 ( 
.A(n_2417),
.B(n_59),
.Y(n_2508)
);

AOI221xp5_ASAP7_75t_L g2509 ( 
.A1(n_2388),
.A2(n_2413),
.B1(n_2432),
.B2(n_2421),
.C(n_2418),
.Y(n_2509)
);

AOI211xp5_ASAP7_75t_L g2510 ( 
.A1(n_2411),
.A2(n_63),
.B(n_61),
.C(n_62),
.Y(n_2510)
);

OAI21xp33_ASAP7_75t_L g2511 ( 
.A1(n_2390),
.A2(n_1818),
.B(n_1815),
.Y(n_2511)
);

AOI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2319),
.A2(n_1095),
.B(n_1092),
.Y(n_2512)
);

OAI221xp5_ASAP7_75t_L g2513 ( 
.A1(n_2403),
.A2(n_1808),
.B1(n_1797),
.B2(n_1796),
.C(n_64),
.Y(n_2513)
);

OAI321xp33_ASAP7_75t_L g2514 ( 
.A1(n_2395),
.A2(n_64),
.A3(n_66),
.B1(n_61),
.B2(n_63),
.C(n_65),
.Y(n_2514)
);

AOI321xp33_ASAP7_75t_L g2515 ( 
.A1(n_2427),
.A2(n_67),
.A3(n_69),
.B1(n_65),
.B2(n_66),
.C(n_68),
.Y(n_2515)
);

AOI22xp33_ASAP7_75t_L g2516 ( 
.A1(n_2406),
.A2(n_1824),
.B1(n_1775),
.B2(n_1818),
.Y(n_2516)
);

AOI211xp5_ASAP7_75t_L g2517 ( 
.A1(n_2334),
.A2(n_71),
.B(n_67),
.C(n_69),
.Y(n_2517)
);

INVxp67_ASAP7_75t_L g2518 ( 
.A(n_2412),
.Y(n_2518)
);

INVx2_ASAP7_75t_SL g2519 ( 
.A(n_2434),
.Y(n_2519)
);

NAND2xp5_ASAP7_75t_SL g2520 ( 
.A(n_2437),
.B(n_1797),
.Y(n_2520)
);

AOI22xp5_ASAP7_75t_L g2521 ( 
.A1(n_2398),
.A2(n_1815),
.B1(n_1826),
.B2(n_1818),
.Y(n_2521)
);

AND3x1_ASAP7_75t_L g2522 ( 
.A(n_2377),
.B(n_72),
.C(n_73),
.Y(n_2522)
);

AOI221xp5_ASAP7_75t_L g2523 ( 
.A1(n_2342),
.A2(n_75),
.B1(n_72),
.B2(n_74),
.C(n_76),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_SL g2524 ( 
.A(n_2414),
.B(n_1815),
.Y(n_2524)
);

AOI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_2415),
.A2(n_1826),
.B1(n_1808),
.B2(n_1824),
.Y(n_2525)
);

AOI21xp5_ASAP7_75t_L g2526 ( 
.A1(n_2401),
.A2(n_1097),
.B(n_1095),
.Y(n_2526)
);

NOR3xp33_ASAP7_75t_L g2527 ( 
.A(n_2344),
.B(n_1099),
.C(n_1097),
.Y(n_2527)
);

AOI222xp33_ASAP7_75t_L g2528 ( 
.A1(n_2360),
.A2(n_76),
.B1(n_79),
.B2(n_74),
.C1(n_75),
.C2(n_77),
.Y(n_2528)
);

INVx1_ASAP7_75t_L g2529 ( 
.A(n_2383),
.Y(n_2529)
);

AOI221xp5_ASAP7_75t_L g2530 ( 
.A1(n_2346),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.C(n_81),
.Y(n_2530)
);

NOR2xp33_ASAP7_75t_SL g2531 ( 
.A(n_2419),
.B(n_1826),
.Y(n_2531)
);

NOR3xp33_ASAP7_75t_SL g2532 ( 
.A(n_2354),
.B(n_2364),
.C(n_2361),
.Y(n_2532)
);

NOR2xp33_ASAP7_75t_L g2533 ( 
.A(n_2375),
.B(n_80),
.Y(n_2533)
);

AOI21xp5_ASAP7_75t_L g2534 ( 
.A1(n_2424),
.A2(n_1106),
.B(n_1099),
.Y(n_2534)
);

AOI211xp5_ASAP7_75t_L g2535 ( 
.A1(n_2380),
.A2(n_83),
.B(n_81),
.C(n_82),
.Y(n_2535)
);

OAI21xp5_ASAP7_75t_L g2536 ( 
.A1(n_2416),
.A2(n_1784),
.B(n_1773),
.Y(n_2536)
);

NOR2xp33_ASAP7_75t_L g2537 ( 
.A(n_2378),
.B(n_84),
.Y(n_2537)
);

OAI22xp5_ASAP7_75t_L g2538 ( 
.A1(n_2416),
.A2(n_1808),
.B1(n_1763),
.B2(n_1782),
.Y(n_2538)
);

AOI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2352),
.A2(n_2358),
.B1(n_2435),
.B2(n_2408),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2431),
.A2(n_1784),
.B(n_1773),
.Y(n_2540)
);

OAI21xp33_ASAP7_75t_L g2541 ( 
.A1(n_2425),
.A2(n_1782),
.B(n_1778),
.Y(n_2541)
);

NOR3x1_ASAP7_75t_L g2542 ( 
.A(n_2343),
.B(n_84),
.C(n_85),
.Y(n_2542)
);

OAI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2382),
.A2(n_87),
.B1(n_85),
.B2(n_86),
.C(n_88),
.Y(n_2543)
);

NOR2xp33_ASAP7_75t_SL g2544 ( 
.A(n_2426),
.B(n_1106),
.Y(n_2544)
);

AOI322xp5_ASAP7_75t_L g2545 ( 
.A1(n_2379),
.A2(n_93),
.A3(n_92),
.B1(n_89),
.B2(n_87),
.C1(n_88),
.C2(n_91),
.Y(n_2545)
);

AOI321xp33_ASAP7_75t_L g2546 ( 
.A1(n_2402),
.A2(n_94),
.A3(n_96),
.B1(n_89),
.B2(n_93),
.C(n_95),
.Y(n_2546)
);

OAI22xp33_ASAP7_75t_L g2547 ( 
.A1(n_2329),
.A2(n_1791),
.B1(n_97),
.B2(n_94),
.Y(n_2547)
);

AND2x2_ASAP7_75t_SL g2548 ( 
.A(n_2322),
.B(n_1791),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2321),
.Y(n_2549)
);

INVx1_ASAP7_75t_L g2550 ( 
.A(n_2321),
.Y(n_2550)
);

NAND3xp33_ASAP7_75t_L g2551 ( 
.A(n_2329),
.B(n_95),
.C(n_97),
.Y(n_2551)
);

XNOR2x1_ASAP7_75t_L g2552 ( 
.A(n_2351),
.B(n_100),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_L g2553 ( 
.A(n_2321),
.B(n_100),
.Y(n_2553)
);

AOI22xp33_ASAP7_75t_SL g2554 ( 
.A1(n_2340),
.A2(n_1824),
.B1(n_1791),
.B2(n_1775),
.Y(n_2554)
);

NAND2xp5_ASAP7_75t_L g2555 ( 
.A(n_2321),
.B(n_102),
.Y(n_2555)
);

AOI222xp33_ASAP7_75t_L g2556 ( 
.A1(n_2369),
.A2(n_104),
.B1(n_109),
.B2(n_102),
.C1(n_103),
.C2(n_105),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2321),
.B(n_103),
.Y(n_2557)
);

OAI32xp33_ASAP7_75t_L g2558 ( 
.A1(n_2335),
.A2(n_114),
.A3(n_105),
.B1(n_112),
.B2(n_115),
.Y(n_2558)
);

INVx2_ASAP7_75t_L g2559 ( 
.A(n_2330),
.Y(n_2559)
);

NOR3xp33_ASAP7_75t_L g2560 ( 
.A(n_2355),
.B(n_114),
.C(n_115),
.Y(n_2560)
);

NAND2xp33_ASAP7_75t_SL g2561 ( 
.A(n_2330),
.B(n_1775),
.Y(n_2561)
);

OAI32xp33_ASAP7_75t_L g2562 ( 
.A1(n_2335),
.A2(n_118),
.A3(n_116),
.B1(n_117),
.B2(n_120),
.Y(n_2562)
);

NAND3xp33_ASAP7_75t_SL g2563 ( 
.A(n_2329),
.B(n_116),
.C(n_118),
.Y(n_2563)
);

OAI21xp33_ASAP7_75t_L g2564 ( 
.A1(n_2329),
.A2(n_1757),
.B(n_1746),
.Y(n_2564)
);

AOI322xp5_ASAP7_75t_L g2565 ( 
.A1(n_2362),
.A2(n_127),
.A3(n_125),
.B1(n_123),
.B2(n_120),
.C1(n_121),
.C2(n_124),
.Y(n_2565)
);

AOI22xp33_ASAP7_75t_L g2566 ( 
.A1(n_2340),
.A2(n_1824),
.B1(n_1775),
.B2(n_1791),
.Y(n_2566)
);

NAND4xp25_ASAP7_75t_L g2567 ( 
.A(n_2329),
.B(n_125),
.C(n_123),
.D(n_124),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2321),
.B(n_127),
.Y(n_2568)
);

NOR3xp33_ASAP7_75t_L g2569 ( 
.A(n_2355),
.B(n_128),
.C(n_129),
.Y(n_2569)
);

AOI221xp5_ASAP7_75t_L g2570 ( 
.A1(n_2323),
.A2(n_130),
.B1(n_128),
.B2(n_129),
.C(n_131),
.Y(n_2570)
);

NAND2xp5_ASAP7_75t_L g2571 ( 
.A(n_2321),
.B(n_130),
.Y(n_2571)
);

AOI21xp5_ASAP7_75t_L g2572 ( 
.A1(n_2369),
.A2(n_1791),
.B(n_131),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2321),
.Y(n_2573)
);

AOI21xp5_ASAP7_75t_L g2574 ( 
.A1(n_2369),
.A2(n_132),
.B(n_133),
.Y(n_2574)
);

NAND4xp75_ASAP7_75t_L g2575 ( 
.A(n_2397),
.B(n_137),
.C(n_134),
.D(n_136),
.Y(n_2575)
);

OAI221xp5_ASAP7_75t_L g2576 ( 
.A1(n_2329),
.A2(n_138),
.B1(n_136),
.B2(n_137),
.C(n_139),
.Y(n_2576)
);

OA22x2_ASAP7_75t_L g2577 ( 
.A1(n_2329),
.A2(n_140),
.B1(n_138),
.B2(n_139),
.Y(n_2577)
);

HB1xp67_ASAP7_75t_L g2578 ( 
.A(n_2330),
.Y(n_2578)
);

OAI211xp5_ASAP7_75t_L g2579 ( 
.A1(n_2329),
.A2(n_143),
.B(n_140),
.C(n_142),
.Y(n_2579)
);

BUFx2_ASAP7_75t_L g2580 ( 
.A(n_2321),
.Y(n_2580)
);

AOI21xp5_ASAP7_75t_L g2581 ( 
.A1(n_2369),
.A2(n_142),
.B(n_143),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2321),
.B(n_144),
.Y(n_2582)
);

AOI21xp5_ASAP7_75t_L g2583 ( 
.A1(n_2369),
.A2(n_145),
.B(n_146),
.Y(n_2583)
);

OAI211xp5_ASAP7_75t_L g2584 ( 
.A1(n_2329),
.A2(n_148),
.B(n_146),
.C(n_147),
.Y(n_2584)
);

NAND4xp25_ASAP7_75t_L g2585 ( 
.A(n_2329),
.B(n_150),
.C(n_148),
.D(n_149),
.Y(n_2585)
);

OAI22xp5_ASAP7_75t_L g2586 ( 
.A1(n_2329),
.A2(n_151),
.B1(n_149),
.B2(n_150),
.Y(n_2586)
);

AOI21xp33_ASAP7_75t_L g2587 ( 
.A1(n_2578),
.A2(n_151),
.B(n_152),
.Y(n_2587)
);

AOI222xp33_ASAP7_75t_L g2588 ( 
.A1(n_2563),
.A2(n_156),
.B1(n_160),
.B2(n_154),
.C1(n_155),
.C2(n_158),
.Y(n_2588)
);

OAI32xp33_ASAP7_75t_L g2589 ( 
.A1(n_2506),
.A2(n_156),
.A3(n_154),
.B1(n_155),
.B2(n_161),
.Y(n_2589)
);

OAI211xp5_ASAP7_75t_SL g2590 ( 
.A1(n_2440),
.A2(n_2441),
.B(n_2439),
.C(n_2559),
.Y(n_2590)
);

OAI22xp5_ASAP7_75t_L g2591 ( 
.A1(n_2551),
.A2(n_166),
.B1(n_162),
.B2(n_164),
.Y(n_2591)
);

OAI22xp33_ASAP7_75t_L g2592 ( 
.A1(n_2567),
.A2(n_166),
.B1(n_162),
.B2(n_164),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2580),
.Y(n_2593)
);

AOI22xp5_ASAP7_75t_L g2594 ( 
.A1(n_2560),
.A2(n_1746),
.B1(n_170),
.B2(n_168),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_SL g2595 ( 
.A(n_2522),
.B(n_1746),
.Y(n_2595)
);

AOI211xp5_ASAP7_75t_L g2596 ( 
.A1(n_2586),
.A2(n_2576),
.B(n_2584),
.C(n_2579),
.Y(n_2596)
);

INVx1_ASAP7_75t_SL g2597 ( 
.A(n_2575),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2447),
.Y(n_2598)
);

AOI22xp5_ASAP7_75t_L g2599 ( 
.A1(n_2569),
.A2(n_171),
.B1(n_168),
.B2(n_169),
.Y(n_2599)
);

OAI21xp5_ASAP7_75t_L g2600 ( 
.A1(n_2552),
.A2(n_172),
.B(n_173),
.Y(n_2600)
);

AND3x1_ASAP7_75t_L g2601 ( 
.A(n_2446),
.B(n_173),
.C(n_174),
.Y(n_2601)
);

AOI32xp33_ASAP7_75t_L g2602 ( 
.A1(n_2478),
.A2(n_2547),
.A3(n_2476),
.B1(n_2550),
.B2(n_2549),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2493),
.B(n_175),
.Y(n_2603)
);

AND2x2_ASAP7_75t_L g2604 ( 
.A(n_2519),
.B(n_176),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_SL g2605 ( 
.A(n_2514),
.B(n_176),
.Y(n_2605)
);

INVx1_ASAP7_75t_L g2606 ( 
.A(n_2577),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2472),
.A2(n_179),
.B1(n_177),
.B2(n_178),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_L g2608 ( 
.A(n_2556),
.B(n_178),
.Y(n_2608)
);

AO21x1_ASAP7_75t_L g2609 ( 
.A1(n_2574),
.A2(n_179),
.B(n_180),
.Y(n_2609)
);

O2A1O1Ixp33_ASAP7_75t_SL g2610 ( 
.A1(n_2483),
.A2(n_182),
.B(n_180),
.C(n_181),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2581),
.B(n_183),
.Y(n_2611)
);

O2A1O1Ixp33_ASAP7_75t_L g2612 ( 
.A1(n_2567),
.A2(n_185),
.B(n_183),
.C(n_184),
.Y(n_2612)
);

OAI22xp5_ASAP7_75t_L g2613 ( 
.A1(n_2444),
.A2(n_186),
.B1(n_184),
.B2(n_185),
.Y(n_2613)
);

OAI21xp33_ASAP7_75t_SL g2614 ( 
.A1(n_2585),
.A2(n_186),
.B(n_187),
.Y(n_2614)
);

OAI21xp33_ASAP7_75t_SL g2615 ( 
.A1(n_2585),
.A2(n_189),
.B(n_190),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2502),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2515),
.B(n_190),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2508),
.Y(n_2618)
);

AOI21xp33_ASAP7_75t_L g2619 ( 
.A1(n_2528),
.A2(n_191),
.B(n_192),
.Y(n_2619)
);

AOI21xp5_ASAP7_75t_L g2620 ( 
.A1(n_2583),
.A2(n_2454),
.B(n_2449),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2492),
.Y(n_2621)
);

AOI221x1_ASAP7_75t_L g2622 ( 
.A1(n_2457),
.A2(n_194),
.B1(n_192),
.B2(n_193),
.C(n_195),
.Y(n_2622)
);

OAI221xp5_ASAP7_75t_L g2623 ( 
.A1(n_2573),
.A2(n_197),
.B1(n_193),
.B2(n_196),
.C(n_200),
.Y(n_2623)
);

XNOR2xp5_ASAP7_75t_L g2624 ( 
.A(n_2535),
.B(n_196),
.Y(n_2624)
);

AOI32xp33_ASAP7_75t_L g2625 ( 
.A1(n_2466),
.A2(n_2453),
.A3(n_2469),
.B1(n_2450),
.B2(n_2529),
.Y(n_2625)
);

O2A1O1Ixp33_ASAP7_75t_L g2626 ( 
.A1(n_2481),
.A2(n_202),
.B(n_200),
.C(n_201),
.Y(n_2626)
);

O2A1O1Ixp5_ASAP7_75t_SL g2627 ( 
.A1(n_2455),
.A2(n_204),
.B(n_202),
.C(n_203),
.Y(n_2627)
);

AOI21xp5_ASAP7_75t_L g2628 ( 
.A1(n_2461),
.A2(n_205),
.B(n_206),
.Y(n_2628)
);

INVx1_ASAP7_75t_L g2629 ( 
.A(n_2553),
.Y(n_2629)
);

OAI211xp5_ASAP7_75t_SL g2630 ( 
.A1(n_2509),
.A2(n_207),
.B(n_205),
.C(n_206),
.Y(n_2630)
);

OAI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2490),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2631)
);

AOI21xp5_ASAP7_75t_L g2632 ( 
.A1(n_2462),
.A2(n_209),
.B(n_210),
.Y(n_2632)
);

AOI321xp33_ASAP7_75t_L g2633 ( 
.A1(n_2504),
.A2(n_215),
.A3(n_217),
.B1(n_212),
.B2(n_213),
.C(n_216),
.Y(n_2633)
);

AOI211xp5_ASAP7_75t_L g2634 ( 
.A1(n_2481),
.A2(n_216),
.B(n_213),
.C(n_215),
.Y(n_2634)
);

OAI22xp5_ASAP7_75t_L g2635 ( 
.A1(n_2518),
.A2(n_221),
.B1(n_218),
.B2(n_219),
.Y(n_2635)
);

OAI21xp33_ASAP7_75t_SL g2636 ( 
.A1(n_2474),
.A2(n_219),
.B(n_221),
.Y(n_2636)
);

OAI221xp5_ASAP7_75t_L g2637 ( 
.A1(n_2445),
.A2(n_224),
.B1(n_222),
.B2(n_223),
.C(n_225),
.Y(n_2637)
);

AOI22xp5_ASAP7_75t_L g2638 ( 
.A1(n_2485),
.A2(n_225),
.B1(n_222),
.B2(n_223),
.Y(n_2638)
);

OA22x2_ASAP7_75t_L g2639 ( 
.A1(n_2497),
.A2(n_2564),
.B1(n_2555),
.B2(n_2557),
.Y(n_2639)
);

AOI221xp5_ASAP7_75t_L g2640 ( 
.A1(n_2442),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2640)
);

AOI211x1_ASAP7_75t_L g2641 ( 
.A1(n_2438),
.A2(n_231),
.B(n_226),
.C(n_227),
.Y(n_2641)
);

INVx2_ASAP7_75t_SL g2642 ( 
.A(n_2568),
.Y(n_2642)
);

AOI211xp5_ASAP7_75t_L g2643 ( 
.A1(n_2558),
.A2(n_233),
.B(n_231),
.C(n_232),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2571),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2465),
.B(n_232),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2582),
.Y(n_2646)
);

NOR2xp67_ASAP7_75t_L g2647 ( 
.A(n_2468),
.B(n_233),
.Y(n_2647)
);

NOR2xp67_ASAP7_75t_L g2648 ( 
.A(n_2458),
.B(n_235),
.Y(n_2648)
);

AOI21xp33_ASAP7_75t_L g2649 ( 
.A1(n_2456),
.A2(n_235),
.B(n_236),
.Y(n_2649)
);

OAI21xp33_ASAP7_75t_L g2650 ( 
.A1(n_2532),
.A2(n_237),
.B(n_238),
.Y(n_2650)
);

AOI22xp5_ASAP7_75t_L g2651 ( 
.A1(n_2484),
.A2(n_240),
.B1(n_237),
.B2(n_239),
.Y(n_2651)
);

NAND3xp33_ASAP7_75t_SL g2652 ( 
.A(n_2471),
.B(n_239),
.C(n_240),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_SL g2653 ( 
.A1(n_2548),
.A2(n_245),
.B1(n_241),
.B2(n_243),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2470),
.Y(n_2654)
);

OAI22xp33_ASAP7_75t_L g2655 ( 
.A1(n_2524),
.A2(n_246),
.B1(n_243),
.B2(n_245),
.Y(n_2655)
);

OAI21xp33_ASAP7_75t_L g2656 ( 
.A1(n_2487),
.A2(n_247),
.B(n_248),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_SL g2657 ( 
.A(n_2562),
.B(n_247),
.Y(n_2657)
);

OAI211xp5_ASAP7_75t_SL g2658 ( 
.A1(n_2443),
.A2(n_250),
.B(n_248),
.C(n_249),
.Y(n_2658)
);

AOI221xp5_ASAP7_75t_L g2659 ( 
.A1(n_2513),
.A2(n_252),
.B1(n_250),
.B2(n_251),
.C(n_254),
.Y(n_2659)
);

OAI21xp33_ASAP7_75t_L g2660 ( 
.A1(n_2539),
.A2(n_251),
.B(n_255),
.Y(n_2660)
);

OAI222xp33_ASAP7_75t_L g2661 ( 
.A1(n_2495),
.A2(n_256),
.B1(n_257),
.B2(n_258),
.C1(n_259),
.C2(n_260),
.Y(n_2661)
);

AOI21xp5_ASAP7_75t_L g2662 ( 
.A1(n_2451),
.A2(n_258),
.B(n_260),
.Y(n_2662)
);

INVx1_ASAP7_75t_L g2663 ( 
.A(n_2537),
.Y(n_2663)
);

AOI221xp5_ASAP7_75t_L g2664 ( 
.A1(n_2570),
.A2(n_264),
.B1(n_261),
.B2(n_262),
.C(n_265),
.Y(n_2664)
);

OAI21xp33_ASAP7_75t_L g2665 ( 
.A1(n_2531),
.A2(n_267),
.B(n_270),
.Y(n_2665)
);

AND2x2_ASAP7_75t_L g2666 ( 
.A(n_2542),
.B(n_267),
.Y(n_2666)
);

AOI21xp5_ASAP7_75t_L g2667 ( 
.A1(n_2460),
.A2(n_271),
.B(n_273),
.Y(n_2667)
);

OAI22xp5_ASAP7_75t_L g2668 ( 
.A1(n_2473),
.A2(n_2510),
.B1(n_2517),
.B2(n_2507),
.Y(n_2668)
);

O2A1O1Ixp5_ASAP7_75t_L g2669 ( 
.A1(n_2561),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_2669)
);

AOI21xp5_ASAP7_75t_L g2670 ( 
.A1(n_2520),
.A2(n_275),
.B(n_276),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2533),
.Y(n_2671)
);

AOI222xp33_ASAP7_75t_L g2672 ( 
.A1(n_2541),
.A2(n_276),
.B1(n_277),
.B2(n_278),
.C1(n_280),
.C2(n_282),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2464),
.B(n_278),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_SL g2674 ( 
.A(n_2546),
.B(n_2545),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_2606),
.B(n_2486),
.Y(n_2675)
);

OAI22xp5_ASAP7_75t_L g2676 ( 
.A1(n_2638),
.A2(n_2543),
.B1(n_2477),
.B2(n_2498),
.Y(n_2676)
);

OAI211xp5_ASAP7_75t_L g2677 ( 
.A1(n_2614),
.A2(n_2452),
.B(n_2565),
.C(n_2491),
.Y(n_2677)
);

OAI22xp5_ASAP7_75t_L g2678 ( 
.A1(n_2593),
.A2(n_2516),
.B1(n_2463),
.B2(n_2523),
.Y(n_2678)
);

NAND5xp2_ASAP7_75t_L g2679 ( 
.A(n_2602),
.B(n_2488),
.C(n_2501),
.D(n_2530),
.E(n_2459),
.Y(n_2679)
);

AOI211xp5_ASAP7_75t_L g2680 ( 
.A1(n_2589),
.A2(n_2572),
.B(n_2467),
.C(n_2527),
.Y(n_2680)
);

OAI221xp5_ASAP7_75t_L g2681 ( 
.A1(n_2615),
.A2(n_2448),
.B1(n_2536),
.B2(n_2511),
.C(n_2475),
.Y(n_2681)
);

O2A1O1Ixp33_ASAP7_75t_L g2682 ( 
.A1(n_2610),
.A2(n_2613),
.B(n_2617),
.C(n_2605),
.Y(n_2682)
);

AOI211xp5_ASAP7_75t_L g2683 ( 
.A1(n_2619),
.A2(n_2500),
.B(n_2512),
.C(n_2526),
.Y(n_2683)
);

AND2x2_ASAP7_75t_L g2684 ( 
.A(n_2666),
.B(n_2544),
.Y(n_2684)
);

OAI21xp33_ASAP7_75t_SL g2685 ( 
.A1(n_2674),
.A2(n_2505),
.B(n_2494),
.Y(n_2685)
);

A2O1A1Ixp33_ASAP7_75t_L g2686 ( 
.A1(n_2612),
.A2(n_2534),
.B(n_2489),
.C(n_2538),
.Y(n_2686)
);

OAI21xp5_ASAP7_75t_L g2687 ( 
.A1(n_2636),
.A2(n_2540),
.B(n_2525),
.Y(n_2687)
);

NOR2xp33_ASAP7_75t_L g2688 ( 
.A(n_2658),
.B(n_2480),
.Y(n_2688)
);

NOR2xp67_ASAP7_75t_SL g2689 ( 
.A(n_2618),
.B(n_282),
.Y(n_2689)
);

NOR2xp67_ASAP7_75t_L g2690 ( 
.A(n_2652),
.B(n_2499),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2609),
.Y(n_2691)
);

NAND3x1_ASAP7_75t_L g2692 ( 
.A(n_2608),
.B(n_2611),
.C(n_2600),
.Y(n_2692)
);

NAND2xp33_ASAP7_75t_SL g2693 ( 
.A(n_2604),
.B(n_2496),
.Y(n_2693)
);

AOI22xp5_ASAP7_75t_L g2694 ( 
.A1(n_2657),
.A2(n_2479),
.B1(n_2554),
.B2(n_2521),
.Y(n_2694)
);

OAI221xp5_ASAP7_75t_L g2695 ( 
.A1(n_2625),
.A2(n_2660),
.B1(n_2653),
.B2(n_2656),
.C(n_2637),
.Y(n_2695)
);

AOI322xp5_ASAP7_75t_L g2696 ( 
.A1(n_2597),
.A2(n_2566),
.A3(n_2482),
.B1(n_2503),
.B2(n_286),
.C1(n_287),
.C2(n_288),
.Y(n_2696)
);

OAI221xp5_ASAP7_75t_L g2697 ( 
.A1(n_2596),
.A2(n_285),
.B1(n_283),
.B2(n_284),
.C(n_287),
.Y(n_2697)
);

AOI22xp5_ASAP7_75t_L g2698 ( 
.A1(n_2590),
.A2(n_288),
.B1(n_284),
.B2(n_285),
.Y(n_2698)
);

INVx1_ASAP7_75t_SL g2699 ( 
.A(n_2603),
.Y(n_2699)
);

AOI22xp5_ASAP7_75t_L g2700 ( 
.A1(n_2630),
.A2(n_291),
.B1(n_289),
.B2(n_290),
.Y(n_2700)
);

AOI22xp5_ASAP7_75t_L g2701 ( 
.A1(n_2668),
.A2(n_293),
.B1(n_290),
.B2(n_292),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2624),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2645),
.Y(n_2703)
);

NAND2xp33_ASAP7_75t_SL g2704 ( 
.A(n_2598),
.B(n_292),
.Y(n_2704)
);

OAI22xp33_ASAP7_75t_SL g2705 ( 
.A1(n_2616),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_2705)
);

OAI22xp5_ASAP7_75t_SL g2706 ( 
.A1(n_2641),
.A2(n_296),
.B1(n_294),
.B2(n_295),
.Y(n_2706)
);

AOI21xp33_ASAP7_75t_SL g2707 ( 
.A1(n_2631),
.A2(n_296),
.B(n_297),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2639),
.Y(n_2708)
);

NOR3xp33_ASAP7_75t_L g2709 ( 
.A(n_2640),
.B(n_297),
.C(n_298),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_SL g2710 ( 
.A(n_2643),
.B(n_299),
.Y(n_2710)
);

INVxp67_ASAP7_75t_SL g2711 ( 
.A(n_2643),
.Y(n_2711)
);

AOI221xp5_ASAP7_75t_L g2712 ( 
.A1(n_2601),
.A2(n_303),
.B1(n_299),
.B2(n_301),
.C(n_304),
.Y(n_2712)
);

AOI221xp5_ASAP7_75t_L g2713 ( 
.A1(n_2592),
.A2(n_305),
.B1(n_301),
.B2(n_303),
.C(n_306),
.Y(n_2713)
);

OAI221xp5_ASAP7_75t_L g2714 ( 
.A1(n_2607),
.A2(n_308),
.B1(n_305),
.B2(n_307),
.C(n_309),
.Y(n_2714)
);

AOI21xp5_ASAP7_75t_L g2715 ( 
.A1(n_2626),
.A2(n_307),
.B(n_308),
.Y(n_2715)
);

AOI322xp5_ASAP7_75t_L g2716 ( 
.A1(n_2673),
.A2(n_309),
.A3(n_310),
.B1(n_311),
.B2(n_312),
.C1(n_314),
.C2(n_316),
.Y(n_2716)
);

AOI22xp5_ASAP7_75t_L g2717 ( 
.A1(n_2650),
.A2(n_317),
.B1(n_310),
.B2(n_316),
.Y(n_2717)
);

CKINVDCx5p33_ASAP7_75t_R g2718 ( 
.A(n_2621),
.Y(n_2718)
);

XNOR2xp5_ASAP7_75t_L g2719 ( 
.A(n_2599),
.B(n_317),
.Y(n_2719)
);

HB1xp67_ASAP7_75t_L g2720 ( 
.A(n_2648),
.Y(n_2720)
);

AND2x2_ASAP7_75t_L g2721 ( 
.A(n_2642),
.B(n_2588),
.Y(n_2721)
);

AND4x1_ASAP7_75t_L g2722 ( 
.A(n_2634),
.B(n_320),
.C(n_318),
.D(n_319),
.Y(n_2722)
);

OAI22xp5_ASAP7_75t_L g2723 ( 
.A1(n_2651),
.A2(n_320),
.B1(n_318),
.B2(n_319),
.Y(n_2723)
);

O2A1O1Ixp33_ASAP7_75t_L g2724 ( 
.A1(n_2634),
.A2(n_323),
.B(n_321),
.C(n_322),
.Y(n_2724)
);

OAI311xp33_ASAP7_75t_L g2725 ( 
.A1(n_2672),
.A2(n_321),
.A3(n_323),
.B1(n_324),
.C1(n_325),
.Y(n_2725)
);

A2O1A1Ixp33_ASAP7_75t_L g2726 ( 
.A1(n_2628),
.A2(n_327),
.B(n_324),
.C(n_325),
.Y(n_2726)
);

OAI22xp5_ASAP7_75t_L g2727 ( 
.A1(n_2594),
.A2(n_330),
.B1(n_327),
.B2(n_328),
.Y(n_2727)
);

AOI211xp5_ASAP7_75t_SL g2728 ( 
.A1(n_2647),
.A2(n_331),
.B(n_328),
.C(n_330),
.Y(n_2728)
);

AOI22xp5_ASAP7_75t_L g2729 ( 
.A1(n_2591),
.A2(n_334),
.B1(n_332),
.B2(n_333),
.Y(n_2729)
);

OAI21xp5_ASAP7_75t_L g2730 ( 
.A1(n_2670),
.A2(n_332),
.B(n_335),
.Y(n_2730)
);

CKINVDCx20_ASAP7_75t_R g2731 ( 
.A(n_2671),
.Y(n_2731)
);

INVx1_ASAP7_75t_L g2732 ( 
.A(n_2635),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_SL g2733 ( 
.A1(n_2711),
.A2(n_2629),
.B1(n_2646),
.B2(n_2644),
.Y(n_2733)
);

NAND4xp75_ASAP7_75t_L g2734 ( 
.A(n_2698),
.B(n_2663),
.C(n_2620),
.D(n_2654),
.Y(n_2734)
);

AOI22xp5_ASAP7_75t_L g2735 ( 
.A1(n_2731),
.A2(n_2665),
.B1(n_2664),
.B2(n_2659),
.Y(n_2735)
);

A2O1A1Ixp33_ASAP7_75t_L g2736 ( 
.A1(n_2724),
.A2(n_2669),
.B(n_2633),
.C(n_2662),
.Y(n_2736)
);

AOI222xp33_ASAP7_75t_L g2737 ( 
.A1(n_2708),
.A2(n_2691),
.B1(n_2685),
.B2(n_2693),
.C1(n_2690),
.C2(n_2675),
.Y(n_2737)
);

OAI221xp5_ASAP7_75t_L g2738 ( 
.A1(n_2695),
.A2(n_2632),
.B1(n_2587),
.B2(n_2667),
.C(n_2649),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2699),
.B(n_2655),
.Y(n_2739)
);

NAND2xp5_ASAP7_75t_L g2740 ( 
.A(n_2699),
.B(n_2622),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2720),
.Y(n_2741)
);

AOI211xp5_ASAP7_75t_L g2742 ( 
.A1(n_2707),
.A2(n_2706),
.B(n_2725),
.C(n_2677),
.Y(n_2742)
);

OAI21xp5_ASAP7_75t_L g2743 ( 
.A1(n_2715),
.A2(n_2692),
.B(n_2682),
.Y(n_2743)
);

OAI21xp5_ASAP7_75t_L g2744 ( 
.A1(n_2710),
.A2(n_2627),
.B(n_2661),
.Y(n_2744)
);

OAI221xp5_ASAP7_75t_L g2745 ( 
.A1(n_2687),
.A2(n_2595),
.B1(n_2623),
.B2(n_340),
.C(n_342),
.Y(n_2745)
);

AOI22xp33_ASAP7_75t_SL g2746 ( 
.A1(n_2718),
.A2(n_342),
.B1(n_336),
.B2(n_339),
.Y(n_2746)
);

AO22x2_ASAP7_75t_L g2747 ( 
.A1(n_2732),
.A2(n_343),
.B1(n_336),
.B2(n_339),
.Y(n_2747)
);

AOI22xp5_ASAP7_75t_L g2748 ( 
.A1(n_2721),
.A2(n_347),
.B1(n_343),
.B2(n_344),
.Y(n_2748)
);

AOI222xp33_ASAP7_75t_L g2749 ( 
.A1(n_2688),
.A2(n_349),
.B1(n_350),
.B2(n_351),
.C1(n_352),
.C2(n_353),
.Y(n_2749)
);

AOI22xp5_ASAP7_75t_L g2750 ( 
.A1(n_2709),
.A2(n_2676),
.B1(n_2702),
.B2(n_2700),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2689),
.Y(n_2751)
);

AOI21xp33_ASAP7_75t_L g2752 ( 
.A1(n_2680),
.A2(n_351),
.B(n_353),
.Y(n_2752)
);

AOI22xp5_ASAP7_75t_SL g2753 ( 
.A1(n_2705),
.A2(n_357),
.B1(n_355),
.B2(n_356),
.Y(n_2753)
);

NOR2x1_ASAP7_75t_L g2754 ( 
.A(n_2697),
.B(n_356),
.Y(n_2754)
);

NAND4xp25_ASAP7_75t_SL g2755 ( 
.A(n_2694),
.B(n_362),
.C(n_358),
.D(n_360),
.Y(n_2755)
);

NOR2x1_ASAP7_75t_L g2756 ( 
.A(n_2726),
.B(n_358),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2728),
.B(n_362),
.Y(n_2757)
);

INVx1_ASAP7_75t_L g2758 ( 
.A(n_2722),
.Y(n_2758)
);

A2O1A1Ixp33_ASAP7_75t_L g2759 ( 
.A1(n_2704),
.A2(n_367),
.B(n_363),
.C(n_366),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2719),
.Y(n_2760)
);

INVx1_ASAP7_75t_SL g2761 ( 
.A(n_2684),
.Y(n_2761)
);

OA22x2_ASAP7_75t_L g2762 ( 
.A1(n_2717),
.A2(n_369),
.B1(n_363),
.B2(n_366),
.Y(n_2762)
);

AOI21xp33_ASAP7_75t_L g2763 ( 
.A1(n_2678),
.A2(n_369),
.B(n_370),
.Y(n_2763)
);

AO22x1_ASAP7_75t_L g2764 ( 
.A1(n_2730),
.A2(n_373),
.B1(n_371),
.B2(n_372),
.Y(n_2764)
);

O2A1O1Ixp33_ASAP7_75t_L g2765 ( 
.A1(n_2723),
.A2(n_374),
.B(n_372),
.C(n_373),
.Y(n_2765)
);

HB1xp67_ASAP7_75t_L g2766 ( 
.A(n_2712),
.Y(n_2766)
);

NOR2x1_ASAP7_75t_SL g2767 ( 
.A(n_2727),
.B(n_375),
.Y(n_2767)
);

NAND2xp5_ASAP7_75t_L g2768 ( 
.A(n_2716),
.B(n_375),
.Y(n_2768)
);

NOR2x1_ASAP7_75t_L g2769 ( 
.A(n_2751),
.B(n_2703),
.Y(n_2769)
);

AND2x2_ASAP7_75t_SL g2770 ( 
.A(n_2740),
.B(n_2713),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2747),
.Y(n_2771)
);

AOI22xp5_ASAP7_75t_L g2772 ( 
.A1(n_2755),
.A2(n_2737),
.B1(n_2758),
.B2(n_2761),
.Y(n_2772)
);

AOI22xp5_ASAP7_75t_L g2773 ( 
.A1(n_2741),
.A2(n_2729),
.B1(n_2714),
.B2(n_2681),
.Y(n_2773)
);

NOR2x1_ASAP7_75t_L g2774 ( 
.A(n_2734),
.B(n_2679),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2747),
.Y(n_2775)
);

AOI22xp5_ASAP7_75t_L g2776 ( 
.A1(n_2735),
.A2(n_2701),
.B1(n_2683),
.B2(n_2686),
.Y(n_2776)
);

INVxp67_ASAP7_75t_SL g2777 ( 
.A(n_2753),
.Y(n_2777)
);

OAI22xp5_ASAP7_75t_L g2778 ( 
.A1(n_2748),
.A2(n_2750),
.B1(n_2742),
.B2(n_2736),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2757),
.Y(n_2779)
);

AOI22xp5_ASAP7_75t_L g2780 ( 
.A1(n_2739),
.A2(n_2696),
.B1(n_379),
.B2(n_377),
.Y(n_2780)
);

AND2x2_ASAP7_75t_SL g2781 ( 
.A(n_2768),
.B(n_377),
.Y(n_2781)
);

AO22x2_ASAP7_75t_L g2782 ( 
.A1(n_2760),
.A2(n_380),
.B1(n_378),
.B2(n_379),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2762),
.Y(n_2783)
);

NOR2x1_ASAP7_75t_L g2784 ( 
.A(n_2759),
.B(n_2743),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2744),
.B(n_380),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2767),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2754),
.B(n_381),
.Y(n_2787)
);

OA22x2_ASAP7_75t_L g2788 ( 
.A1(n_2766),
.A2(n_387),
.B1(n_383),
.B2(n_385),
.Y(n_2788)
);

CKINVDCx20_ASAP7_75t_R g2789 ( 
.A(n_2776),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2788),
.Y(n_2790)
);

INVx2_ASAP7_75t_SL g2791 ( 
.A(n_2786),
.Y(n_2791)
);

INVx1_ASAP7_75t_L g2792 ( 
.A(n_2771),
.Y(n_2792)
);

AND2x2_ASAP7_75t_SL g2793 ( 
.A(n_2770),
.B(n_2764),
.Y(n_2793)
);

NOR2x1_ASAP7_75t_L g2794 ( 
.A(n_2775),
.B(n_2756),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2782),
.Y(n_2795)
);

NOR2xp33_ASAP7_75t_L g2796 ( 
.A(n_2777),
.B(n_2738),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2782),
.Y(n_2797)
);

NAND2xp5_ASAP7_75t_L g2798 ( 
.A(n_2785),
.B(n_2746),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2787),
.Y(n_2799)
);

AO22x2_ASAP7_75t_L g2800 ( 
.A1(n_2778),
.A2(n_2763),
.B1(n_2733),
.B2(n_2752),
.Y(n_2800)
);

BUFx2_ASAP7_75t_L g2801 ( 
.A(n_2769),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2772),
.A2(n_2745),
.B1(n_2765),
.B2(n_2749),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2783),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2780),
.B(n_2779),
.Y(n_2804)
);

NOR2x1_ASAP7_75t_L g2805 ( 
.A(n_2784),
.B(n_387),
.Y(n_2805)
);

OAI211xp5_ASAP7_75t_SL g2806 ( 
.A1(n_2794),
.A2(n_2773),
.B(n_2774),
.C(n_2781),
.Y(n_2806)
);

O2A1O1Ixp33_ASAP7_75t_L g2807 ( 
.A1(n_2801),
.A2(n_2797),
.B(n_2795),
.C(n_2791),
.Y(n_2807)
);

A2O1A1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_2796),
.A2(n_393),
.B(n_389),
.C(n_392),
.Y(n_2808)
);

AOI221xp5_ASAP7_75t_L g2809 ( 
.A1(n_2802),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.C(n_397),
.Y(n_2809)
);

NAND2x1p5_ASAP7_75t_L g2810 ( 
.A(n_2793),
.B(n_1743),
.Y(n_2810)
);

AO22x2_ASAP7_75t_L g2811 ( 
.A1(n_2792),
.A2(n_397),
.B1(n_394),
.B2(n_395),
.Y(n_2811)
);

AOI221xp5_ASAP7_75t_L g2812 ( 
.A1(n_2800),
.A2(n_398),
.B1(n_399),
.B2(n_400),
.C(n_401),
.Y(n_2812)
);

AOI221xp5_ASAP7_75t_L g2813 ( 
.A1(n_2800),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.C(n_402),
.Y(n_2813)
);

OAI21xp33_ASAP7_75t_L g2814 ( 
.A1(n_2803),
.A2(n_402),
.B(n_403),
.Y(n_2814)
);

XNOR2x1_ASAP7_75t_L g2815 ( 
.A(n_2804),
.B(n_403),
.Y(n_2815)
);

NAND3xp33_ASAP7_75t_SL g2816 ( 
.A(n_2789),
.B(n_405),
.C(n_406),
.Y(n_2816)
);

AOI22xp5_ASAP7_75t_L g2817 ( 
.A1(n_2790),
.A2(n_408),
.B1(n_405),
.B2(n_407),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2805),
.Y(n_2818)
);

AOI221xp5_ASAP7_75t_L g2819 ( 
.A1(n_2798),
.A2(n_407),
.B1(n_408),
.B2(n_410),
.C(n_412),
.Y(n_2819)
);

NAND2xp5_ASAP7_75t_SL g2820 ( 
.A(n_2799),
.B(n_410),
.Y(n_2820)
);

AOI221xp5_ASAP7_75t_L g2821 ( 
.A1(n_2802),
.A2(n_412),
.B1(n_413),
.B2(n_414),
.C(n_415),
.Y(n_2821)
);

NAND3xp33_ASAP7_75t_L g2822 ( 
.A(n_2801),
.B(n_413),
.C(n_414),
.Y(n_2822)
);

AOI221xp5_ASAP7_75t_L g2823 ( 
.A1(n_2802),
.A2(n_416),
.B1(n_417),
.B2(n_418),
.C(n_419),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2797),
.B(n_417),
.Y(n_2824)
);

BUFx2_ASAP7_75t_L g2825 ( 
.A(n_2811),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2812),
.B(n_419),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2824),
.Y(n_2827)
);

AND2x2_ASAP7_75t_L g2828 ( 
.A(n_2815),
.B(n_420),
.Y(n_2828)
);

BUFx2_ASAP7_75t_L g2829 ( 
.A(n_2811),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2818),
.B(n_420),
.Y(n_2830)
);

OAI22xp33_ASAP7_75t_L g2831 ( 
.A1(n_2822),
.A2(n_2817),
.B1(n_2816),
.B2(n_2813),
.Y(n_2831)
);

INVx2_ASAP7_75t_SL g2832 ( 
.A(n_2820),
.Y(n_2832)
);

XOR2x2_ASAP7_75t_L g2833 ( 
.A(n_2809),
.B(n_421),
.Y(n_2833)
);

NAND3x1_ASAP7_75t_L g2834 ( 
.A(n_2821),
.B(n_421),
.C(n_423),
.Y(n_2834)
);

XNOR2xp5_ASAP7_75t_L g2835 ( 
.A(n_2823),
.B(n_424),
.Y(n_2835)
);

NAND2xp5_ASAP7_75t_L g2836 ( 
.A(n_2814),
.B(n_426),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2807),
.Y(n_2837)
);

AND2x4_ASAP7_75t_L g2838 ( 
.A(n_2808),
.B(n_2806),
.Y(n_2838)
);

NAND4xp25_ASAP7_75t_L g2839 ( 
.A(n_2819),
.B(n_426),
.C(n_427),
.D(n_428),
.Y(n_2839)
);

NOR2x1_ASAP7_75t_L g2840 ( 
.A(n_2810),
.B(n_427),
.Y(n_2840)
);

XOR2xp5_ASAP7_75t_L g2841 ( 
.A(n_2815),
.B(n_430),
.Y(n_2841)
);

BUFx2_ASAP7_75t_L g2842 ( 
.A(n_2811),
.Y(n_2842)
);

AOI21x1_ASAP7_75t_L g2843 ( 
.A1(n_2818),
.A2(n_430),
.B(n_431),
.Y(n_2843)
);

XOR2x2_ASAP7_75t_L g2844 ( 
.A(n_2815),
.B(n_433),
.Y(n_2844)
);

AND2x4_ASAP7_75t_L g2845 ( 
.A(n_2818),
.B(n_434),
.Y(n_2845)
);

AND2x2_ASAP7_75t_L g2846 ( 
.A(n_2828),
.B(n_435),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2825),
.Y(n_2847)
);

XNOR2xp5_ASAP7_75t_L g2848 ( 
.A(n_2841),
.B(n_436),
.Y(n_2848)
);

AOI22x1_ASAP7_75t_L g2849 ( 
.A1(n_2829),
.A2(n_436),
.B1(n_437),
.B2(n_438),
.Y(n_2849)
);

INVx4_ASAP7_75t_L g2850 ( 
.A(n_2842),
.Y(n_2850)
);

OAI22x1_ASAP7_75t_L g2851 ( 
.A1(n_2837),
.A2(n_2835),
.B1(n_2838),
.B2(n_2832),
.Y(n_2851)
);

HB1xp67_ASAP7_75t_L g2852 ( 
.A(n_2843),
.Y(n_2852)
);

INVx1_ASAP7_75t_L g2853 ( 
.A(n_2830),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2845),
.Y(n_2854)
);

XOR2x1_ASAP7_75t_L g2855 ( 
.A(n_2844),
.B(n_438),
.Y(n_2855)
);

NOR2xp67_ASAP7_75t_L g2856 ( 
.A(n_2839),
.B(n_441),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2840),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2833),
.Y(n_2858)
);

AOI22xp5_ASAP7_75t_L g2859 ( 
.A1(n_2831),
.A2(n_442),
.B1(n_443),
.B2(n_444),
.Y(n_2859)
);

XNOR2xp5_ASAP7_75t_L g2860 ( 
.A(n_2834),
.B(n_442),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2848),
.Y(n_2861)
);

AOI22xp5_ASAP7_75t_L g2862 ( 
.A1(n_2847),
.A2(n_2836),
.B1(n_2827),
.B2(n_2835),
.Y(n_2862)
);

INVx1_ASAP7_75t_SL g2863 ( 
.A(n_2846),
.Y(n_2863)
);

NOR2xp67_ASAP7_75t_SL g2864 ( 
.A(n_2852),
.B(n_2826),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2860),
.Y(n_2865)
);

AOI22xp5_ASAP7_75t_L g2866 ( 
.A1(n_2856),
.A2(n_444),
.B1(n_445),
.B2(n_446),
.Y(n_2866)
);

AOI221xp5_ASAP7_75t_L g2867 ( 
.A1(n_2850),
.A2(n_446),
.B1(n_447),
.B2(n_448),
.C(n_449),
.Y(n_2867)
);

OAI211xp5_ASAP7_75t_L g2868 ( 
.A1(n_2849),
.A2(n_447),
.B(n_449),
.C(n_450),
.Y(n_2868)
);

OAI21x1_ASAP7_75t_L g2869 ( 
.A1(n_2855),
.A2(n_1743),
.B(n_452),
.Y(n_2869)
);

BUFx2_ASAP7_75t_L g2870 ( 
.A(n_2857),
.Y(n_2870)
);

AOI22x1_ASAP7_75t_L g2871 ( 
.A1(n_2851),
.A2(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_2871)
);

HB1xp67_ASAP7_75t_L g2872 ( 
.A(n_2853),
.Y(n_2872)
);

CKINVDCx20_ASAP7_75t_R g2873 ( 
.A(n_2858),
.Y(n_2873)
);

NAND3xp33_ASAP7_75t_L g2874 ( 
.A(n_2854),
.B(n_458),
.C(n_459),
.Y(n_2874)
);

INVx2_ASAP7_75t_L g2875 ( 
.A(n_2871),
.Y(n_2875)
);

INVx1_ASAP7_75t_L g2876 ( 
.A(n_2872),
.Y(n_2876)
);

INVx1_ASAP7_75t_L g2877 ( 
.A(n_2866),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2870),
.A2(n_2859),
.B(n_458),
.Y(n_2878)
);

HB1xp67_ASAP7_75t_L g2879 ( 
.A(n_2874),
.Y(n_2879)
);

OAI22xp5_ASAP7_75t_L g2880 ( 
.A1(n_2873),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.Y(n_2880)
);

NOR3xp33_ASAP7_75t_L g2881 ( 
.A(n_2865),
.B(n_460),
.C(n_462),
.Y(n_2881)
);

AO22x1_ASAP7_75t_L g2882 ( 
.A1(n_2863),
.A2(n_463),
.B1(n_464),
.B2(n_465),
.Y(n_2882)
);

OAI22xp33_ASAP7_75t_L g2883 ( 
.A1(n_2862),
.A2(n_463),
.B1(n_464),
.B2(n_466),
.Y(n_2883)
);

AOI22xp33_ASAP7_75t_L g2884 ( 
.A1(n_2864),
.A2(n_466),
.B1(n_467),
.B2(n_468),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2868),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2861),
.Y(n_2886)
);

HB1xp67_ASAP7_75t_L g2887 ( 
.A(n_2869),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2867),
.Y(n_2888)
);

AO22x2_ASAP7_75t_L g2889 ( 
.A1(n_2863),
.A2(n_467),
.B1(n_469),
.B2(n_471),
.Y(n_2889)
);

BUFx12f_ASAP7_75t_L g2890 ( 
.A(n_2870),
.Y(n_2890)
);

AOI22x1_ASAP7_75t_L g2891 ( 
.A1(n_2890),
.A2(n_469),
.B1(n_471),
.B2(n_472),
.Y(n_2891)
);

AOI22xp5_ASAP7_75t_L g2892 ( 
.A1(n_2876),
.A2(n_472),
.B1(n_473),
.B2(n_475),
.Y(n_2892)
);

OAI22xp5_ASAP7_75t_SL g2893 ( 
.A1(n_2875),
.A2(n_473),
.B1(n_476),
.B2(n_477),
.Y(n_2893)
);

AOI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2886),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_2894)
);

AOI22xp5_ASAP7_75t_L g2895 ( 
.A1(n_2885),
.A2(n_479),
.B1(n_480),
.B2(n_482),
.Y(n_2895)
);

OAI22xp5_ASAP7_75t_SL g2896 ( 
.A1(n_2887),
.A2(n_480),
.B1(n_483),
.B2(n_484),
.Y(n_2896)
);

BUFx2_ASAP7_75t_L g2897 ( 
.A(n_2889),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2881),
.B(n_483),
.Y(n_2898)
);

INVx1_ASAP7_75t_L g2899 ( 
.A(n_2889),
.Y(n_2899)
);

NAND2xp5_ASAP7_75t_L g2900 ( 
.A(n_2884),
.B(n_484),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2882),
.Y(n_2901)
);

OAI22xp5_ASAP7_75t_SL g2902 ( 
.A1(n_2877),
.A2(n_485),
.B1(n_486),
.B2(n_487),
.Y(n_2902)
);

OAI22xp5_ASAP7_75t_L g2903 ( 
.A1(n_2900),
.A2(n_2888),
.B1(n_2879),
.B2(n_2878),
.Y(n_2903)
);

OAI22xp5_ASAP7_75t_L g2904 ( 
.A1(n_2901),
.A2(n_2883),
.B1(n_2880),
.B2(n_489),
.Y(n_2904)
);

OR2x2_ASAP7_75t_L g2905 ( 
.A(n_2898),
.B(n_487),
.Y(n_2905)
);

AOI22xp5_ASAP7_75t_L g2906 ( 
.A1(n_2899),
.A2(n_488),
.B1(n_489),
.B2(n_490),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2897),
.A2(n_488),
.B1(n_491),
.B2(n_493),
.Y(n_2907)
);

INVxp33_ASAP7_75t_SL g2908 ( 
.A(n_2895),
.Y(n_2908)
);

OAI22xp5_ASAP7_75t_L g2909 ( 
.A1(n_2891),
.A2(n_491),
.B1(n_494),
.B2(n_495),
.Y(n_2909)
);

AOI221xp5_ASAP7_75t_L g2910 ( 
.A1(n_2896),
.A2(n_494),
.B1(n_496),
.B2(n_497),
.C(n_498),
.Y(n_2910)
);

AOI22xp5_ASAP7_75t_L g2911 ( 
.A1(n_2893),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.Y(n_2911)
);

AOI22xp5_ASAP7_75t_SL g2912 ( 
.A1(n_2902),
.A2(n_499),
.B1(n_500),
.B2(n_502),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2892),
.Y(n_2913)
);

AOI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2908),
.A2(n_2894),
.B1(n_500),
.B2(n_502),
.Y(n_2914)
);

AOI221xp5_ASAP7_75t_L g2915 ( 
.A1(n_2904),
.A2(n_2909),
.B1(n_2903),
.B2(n_2913),
.C(n_2910),
.Y(n_2915)
);

OAI21xp33_ASAP7_75t_L g2916 ( 
.A1(n_2911),
.A2(n_499),
.B(n_503),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2905),
.A2(n_2912),
.B1(n_2906),
.B2(n_2907),
.Y(n_2917)
);

INVx1_ASAP7_75t_L g2918 ( 
.A(n_2905),
.Y(n_2918)
);

OAI21xp5_ASAP7_75t_L g2919 ( 
.A1(n_2904),
.A2(n_503),
.B(n_504),
.Y(n_2919)
);

OAI21xp33_ASAP7_75t_L g2920 ( 
.A1(n_2908),
.A2(n_504),
.B(n_505),
.Y(n_2920)
);

OAI21xp5_ASAP7_75t_L g2921 ( 
.A1(n_2904),
.A2(n_506),
.B(n_507),
.Y(n_2921)
);

AO221x1_ASAP7_75t_L g2922 ( 
.A1(n_2909),
.A2(n_508),
.B1(n_509),
.B2(n_510),
.C(n_511),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2903),
.A2(n_508),
.B(n_509),
.Y(n_2923)
);

AOI22x1_ASAP7_75t_L g2924 ( 
.A1(n_2919),
.A2(n_510),
.B1(n_511),
.B2(n_513),
.Y(n_2924)
);

AOI22xp33_ASAP7_75t_SL g2925 ( 
.A1(n_2922),
.A2(n_513),
.B1(n_514),
.B2(n_515),
.Y(n_2925)
);

BUFx3_ASAP7_75t_L g2926 ( 
.A(n_2918),
.Y(n_2926)
);

OAI21xp5_ASAP7_75t_L g2927 ( 
.A1(n_2914),
.A2(n_514),
.B(n_516),
.Y(n_2927)
);

AOI222xp33_ASAP7_75t_L g2928 ( 
.A1(n_2915),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.C1(n_521),
.C2(n_522),
.Y(n_2928)
);

AOI22xp33_ASAP7_75t_L g2929 ( 
.A1(n_2926),
.A2(n_2916),
.B1(n_2917),
.B2(n_2921),
.Y(n_2929)
);

AOI22xp33_ASAP7_75t_L g2930 ( 
.A1(n_2925),
.A2(n_2923),
.B1(n_2920),
.B2(n_523),
.Y(n_2930)
);

OR2x6_ASAP7_75t_L g2931 ( 
.A(n_2929),
.B(n_2927),
.Y(n_2931)
);

O2A1O1Ixp33_ASAP7_75t_R g2932 ( 
.A1(n_2931),
.A2(n_2930),
.B(n_2924),
.C(n_2928),
.Y(n_2932)
);

AOI211xp5_ASAP7_75t_L g2933 ( 
.A1(n_2932),
.A2(n_519),
.B(n_522),
.C(n_524),
.Y(n_2933)
);


endmodule