module fake_netlist_1_9647_n_694 (n_117, n_44, n_133, n_149, n_81, n_69, n_185, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_125, n_9, n_161, n_10, n_177, n_130, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_154, n_7, n_29, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_139, n_16, n_13, n_169, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_38, n_64, n_142, n_184, n_46, n_31, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_96, n_39, n_694);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_185;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_125;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_154;
input n_7;
input n_29;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_139;
input n_16;
input n_13;
input n_169;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_38;
input n_64;
input n_142;
input n_184;
input n_46;
input n_31;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_96;
input n_39;
output n_694;
wire n_663;
wire n_361;
wire n_513;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_607;
wire n_431;
wire n_484;
wire n_496;
wire n_667;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_202;
wire n_386;
wire n_432;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_227;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_568;
wire n_357;
wire n_245;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_673;
wire n_669;
wire n_616;
wire n_365;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_295;
wire n_654;
wire n_263;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_300;
wire n_524;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_602;
wire n_198;
wire n_424;
wire n_629;
wire n_569;
wire n_297;
wire n_410;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_375;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_421;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g189 ( .A(n_20), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_151), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_113), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g192 ( .A(n_30), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g193 ( .A(n_140), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_81), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_111), .Y(n_195) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_15), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_69), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_115), .Y(n_198) );
BUFx3_ASAP7_75t_L g199 ( .A(n_165), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_183), .Y(n_200) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_38), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_86), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_49), .Y(n_205) );
BUFx5_ASAP7_75t_L g206 ( .A(n_137), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_146), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_142), .Y(n_208) );
CKINVDCx5p33_ASAP7_75t_R g209 ( .A(n_166), .Y(n_209) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_175), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_157), .Y(n_211) );
CKINVDCx5p33_ASAP7_75t_R g212 ( .A(n_32), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_133), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_22), .Y(n_214) );
CKINVDCx20_ASAP7_75t_R g215 ( .A(n_29), .Y(n_215) );
BUFx5_ASAP7_75t_L g216 ( .A(n_20), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_138), .B(n_59), .Y(n_217) );
BUFx5_ASAP7_75t_L g218 ( .A(n_126), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_181), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_176), .Y(n_220) );
INVxp67_ASAP7_75t_L g221 ( .A(n_128), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_44), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_5), .Y(n_223) );
INVxp67_ASAP7_75t_L g224 ( .A(n_159), .Y(n_224) );
INVx2_ASAP7_75t_L g225 ( .A(n_89), .Y(n_225) );
CKINVDCx5p33_ASAP7_75t_R g226 ( .A(n_188), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_43), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_108), .Y(n_228) );
CKINVDCx5p33_ASAP7_75t_R g229 ( .A(n_129), .Y(n_229) );
INVx1_ASAP7_75t_SL g230 ( .A(n_45), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_118), .Y(n_231) );
INVx2_ASAP7_75t_SL g232 ( .A(n_155), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_182), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_54), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_41), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_99), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_70), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_73), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_109), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_27), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_172), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g243 ( .A(n_3), .Y(n_243) );
INVx1_ASAP7_75t_L g244 ( .A(n_173), .Y(n_244) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_52), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_167), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_82), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_17), .B(n_147), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_114), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_150), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_130), .Y(n_251) );
BUFx10_ASAP7_75t_L g252 ( .A(n_60), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_83), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_67), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_3), .Y(n_255) );
CKINVDCx16_ASAP7_75t_R g256 ( .A(n_121), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g257 ( .A(n_13), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_18), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_9), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_40), .Y(n_260) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_76), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_174), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_15), .Y(n_263) );
BUFx2_ASAP7_75t_L g264 ( .A(n_106), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_34), .Y(n_265) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_95), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_94), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_28), .Y(n_268) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_1), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_162), .B(n_149), .Y(n_270) );
CKINVDCx5p33_ASAP7_75t_R g271 ( .A(n_48), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_180), .Y(n_272) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_37), .Y(n_273) );
HB1xp67_ASAP7_75t_L g274 ( .A(n_47), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_148), .Y(n_275) );
CKINVDCx5p33_ASAP7_75t_R g276 ( .A(n_13), .Y(n_276) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_4), .Y(n_277) );
CKINVDCx5p33_ASAP7_75t_R g278 ( .A(n_156), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_186), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_80), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_39), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_187), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_33), .Y(n_283) );
HB1xp67_ASAP7_75t_L g284 ( .A(n_65), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_184), .Y(n_285) );
BUFx3_ASAP7_75t_L g286 ( .A(n_170), .Y(n_286) );
CKINVDCx5p33_ASAP7_75t_R g287 ( .A(n_68), .Y(n_287) );
CKINVDCx5p33_ASAP7_75t_R g288 ( .A(n_66), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_17), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g290 ( .A(n_134), .Y(n_290) );
INVx1_ASAP7_75t_L g291 ( .A(n_4), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_139), .Y(n_292) );
INVxp67_ASAP7_75t_L g293 ( .A(n_5), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_71), .Y(n_294) );
CKINVDCx16_ASAP7_75t_R g295 ( .A(n_185), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_122), .Y(n_296) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_210), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_272), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_274), .Y(n_299) );
OA21x2_ASAP7_75t_L g300 ( .A1(n_190), .A2(n_194), .B(n_191), .Y(n_300) );
BUFx8_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
AND2x4_ASAP7_75t_SL g302 ( .A(n_252), .B(n_23), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_216), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_216), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_272), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_256), .B(n_0), .Y(n_306) );
INVx3_ASAP7_75t_L g307 ( .A(n_252), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_206), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_284), .B(n_0), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_293), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_216), .Y(n_311) );
INVx2_ASAP7_75t_L g312 ( .A(n_206), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_232), .B(n_1), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_295), .A2(n_2), .B1(n_6), .B2(n_7), .Y(n_314) );
CKINVDCx5p33_ASAP7_75t_R g315 ( .A(n_215), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_283), .B(n_2), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_216), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_189), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_195), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_225), .B(n_7), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_223), .B(n_8), .Y(n_321) );
OA21x2_ASAP7_75t_L g322 ( .A1(n_197), .A2(n_25), .B(n_24), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_206), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_255), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_258), .Y(n_325) );
INVx4_ASAP7_75t_SL g326 ( .A(n_316), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g327 ( .A1(n_319), .A2(n_263), .B1(n_289), .B2(n_259), .Y(n_327) );
CKINVDCx20_ASAP7_75t_R g328 ( .A(n_301), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_316), .Y(n_329) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_297), .Y(n_330) );
OR2x6_ASAP7_75t_L g331 ( .A(n_314), .B(n_291), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_307), .B(n_221), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_311), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_311), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_310), .A2(n_196), .B1(n_277), .B2(n_243), .Y(n_335) );
INVx8_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
NAND2xp5_ASAP7_75t_SL g337 ( .A(n_307), .B(n_224), .Y(n_337) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_319), .B(n_238), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_306), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_317), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_297), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_299), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_303), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_303), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_200), .B1(n_202), .B2(n_198), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_317), .Y(n_347) );
AND2x6_ASAP7_75t_L g348 ( .A(n_321), .B(n_204), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
INVx3_ASAP7_75t_L g350 ( .A(n_298), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_304), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_308), .Y(n_352) );
INVx3_ASAP7_75t_L g353 ( .A(n_298), .Y(n_353) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_343), .A2(n_306), .B1(n_301), .B2(n_309), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_350), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_348), .A2(n_301), .B1(n_321), .B2(n_302), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_340), .B(n_318), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_348), .B(n_324), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_340), .B(n_315), .Y(n_359) );
OAI22x1_ASAP7_75t_SL g360 ( .A1(n_328), .A2(n_315), .B1(n_247), .B2(n_257), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_337), .B(n_325), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_348), .B(n_313), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_350), .Y(n_363) );
INVx2_ASAP7_75t_L g364 ( .A(n_353), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_348), .B(n_320), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g366 ( .A1(n_329), .A2(n_269), .B1(n_276), .B2(n_214), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_332), .B(n_292), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_335), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_353), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_336), .B(n_305), .Y(n_370) );
INVx8_ASAP7_75t_L g371 ( .A(n_336), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_336), .B(n_192), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_326), .B(n_193), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_339), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g375 ( .A1(n_327), .A2(n_323), .B1(n_312), .B2(n_253), .C(n_250), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_344), .B(n_323), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_326), .B(n_201), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_326), .B(n_203), .Y(n_378) );
INVxp67_ASAP7_75t_SL g379 ( .A(n_345), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_352), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_351), .Y(n_381) );
OR2x6_ASAP7_75t_L g382 ( .A(n_331), .B(n_322), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_346), .B(n_205), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_327), .B(n_208), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_335), .B(n_209), .Y(n_385) );
AOI21xp5_ASAP7_75t_L g386 ( .A1(n_362), .A2(n_341), .B(n_334), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_374), .A2(n_346), .B1(n_349), .B2(n_347), .Y(n_387) );
O2A1O1Ixp33_ASAP7_75t_SL g388 ( .A1(n_383), .A2(n_207), .B(n_219), .C(n_213), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_357), .B(n_333), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_357), .B(n_333), .Y(n_390) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_379), .A2(n_333), .B1(n_220), .B2(n_222), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_371), .Y(n_392) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_385), .B(n_248), .Y(n_393) );
O2A1O1Ixp5_ASAP7_75t_L g394 ( .A1(n_383), .A2(n_367), .B(n_373), .C(n_365), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_382), .A2(n_333), .B(n_228), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_382), .A2(n_233), .B(n_227), .Y(n_396) );
BUFx3_ASAP7_75t_L g397 ( .A(n_371), .Y(n_397) );
OAI21xp5_ASAP7_75t_L g398 ( .A1(n_376), .A2(n_235), .B(n_234), .Y(n_398) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_371), .B(n_211), .Y(n_399) );
INVx3_ASAP7_75t_L g400 ( .A(n_381), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_361), .B(n_212), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_355), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_368), .A2(n_237), .B1(n_239), .B2(n_236), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_363), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_359), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_354), .B(n_230), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
NAND2xp5_ASAP7_75t_SL g408 ( .A(n_356), .B(n_226), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_366), .B(n_229), .Y(n_409) );
OAI21x1_ASAP7_75t_L g410 ( .A1(n_358), .A2(n_242), .B(n_241), .Y(n_410) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_380), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_384), .B(n_231), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_364), .Y(n_413) );
AO21x1_ASAP7_75t_L g414 ( .A1(n_385), .A2(n_246), .B(n_244), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_372), .B(n_240), .Y(n_415) );
OAI22xp5_ASAP7_75t_L g416 ( .A1(n_375), .A2(n_279), .B1(n_275), .B2(n_251), .Y(n_416) );
OAI22xp33_ASAP7_75t_L g417 ( .A1(n_369), .A2(n_281), .B1(n_280), .B2(n_282), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_378), .B(n_260), .Y(n_419) );
AND2x4_ASAP7_75t_L g420 ( .A(n_397), .B(n_262), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g421 ( .A1(n_386), .A2(n_285), .B(n_268), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g422 ( .A(n_392), .B(n_245), .Y(n_422) );
NAND2x1p5_ASAP7_75t_L g423 ( .A(n_400), .B(n_360), .Y(n_423) );
INVx3_ASAP7_75t_L g424 ( .A(n_419), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_405), .Y(n_425) );
AOI21xp5_ASAP7_75t_L g426 ( .A1(n_396), .A2(n_296), .B(n_270), .Y(n_426) );
OAI21x1_ASAP7_75t_L g427 ( .A1(n_395), .A2(n_217), .B(n_206), .Y(n_427) );
AOI22xp5_ASAP7_75t_L g428 ( .A1(n_406), .A2(n_271), .B1(n_265), .B2(n_273), .Y(n_428) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_394), .A2(n_287), .B(n_278), .Y(n_429) );
AOI21xp5_ASAP7_75t_L g430 ( .A1(n_389), .A2(n_290), .B(n_288), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_411), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_418), .B(n_199), .Y(n_432) );
A2O1A1Ixp33_ASAP7_75t_L g433 ( .A1(n_398), .A2(n_254), .B(n_267), .C(n_249), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_390), .A2(n_294), .B(n_286), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_407), .B(n_8), .Y(n_435) );
OAI22xp5_ASAP7_75t_L g436 ( .A1(n_387), .A2(n_210), .B1(n_261), .B2(n_266), .Y(n_436) );
OAI21x1_ASAP7_75t_SL g437 ( .A1(n_414), .A2(n_402), .B(n_403), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_411), .Y(n_438) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_388), .A2(n_9), .B(n_10), .C(n_11), .Y(n_439) );
NOR2x1_ASAP7_75t_SL g440 ( .A(n_399), .B(n_261), .Y(n_440) );
AO31x2_ASAP7_75t_L g441 ( .A1(n_416), .A2(n_218), .A3(n_206), .B(n_297), .Y(n_441) );
OAI21x1_ASAP7_75t_L g442 ( .A1(n_410), .A2(n_218), .B(n_266), .Y(n_442) );
AOI221xp5_ASAP7_75t_SL g443 ( .A1(n_417), .A2(n_297), .B1(n_338), .B2(n_330), .C(n_342), .Y(n_443) );
AO31x2_ASAP7_75t_L g444 ( .A1(n_391), .A2(n_218), .A3(n_338), .B(n_330), .Y(n_444) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_413), .Y(n_445) );
INVxp67_ASAP7_75t_SL g446 ( .A(n_417), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_403), .B(n_10), .Y(n_447) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_415), .A2(n_342), .B(n_218), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_404), .Y(n_449) );
INVx8_ASAP7_75t_L g450 ( .A(n_419), .Y(n_450) );
AO31x2_ASAP7_75t_L g451 ( .A1(n_412), .A2(n_342), .A3(n_12), .B(n_14), .Y(n_451) );
OAI21x1_ASAP7_75t_L g452 ( .A1(n_408), .A2(n_31), .B(n_26), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_424), .B(n_409), .Y(n_453) );
OA21x2_ASAP7_75t_L g454 ( .A1(n_443), .A2(n_401), .B(n_393), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_449), .Y(n_455) );
OAI21x1_ASAP7_75t_L g456 ( .A1(n_442), .A2(n_393), .B(n_35), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_431), .Y(n_457) );
INVx2_ASAP7_75t_L g458 ( .A(n_438), .Y(n_458) );
OAI21x1_ASAP7_75t_L g459 ( .A1(n_427), .A2(n_107), .B(n_178), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_450), .B(n_11), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_435), .B(n_12), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_425), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_448), .A2(n_110), .B(n_177), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_446), .B(n_16), .Y(n_464) );
OAI21x1_ASAP7_75t_SL g465 ( .A1(n_437), .A2(n_19), .B(n_21), .Y(n_465) );
OAI21x1_ASAP7_75t_SL g466 ( .A1(n_437), .A2(n_22), .B(n_36), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_439), .A2(n_42), .B(n_46), .C(n_50), .Y(n_467) );
NAND2xp5_ASAP7_75t_SL g468 ( .A(n_445), .B(n_51), .Y(n_468) );
AND2x4_ASAP7_75t_L g469 ( .A(n_420), .B(n_53), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_451), .Y(n_470) );
AO31x2_ASAP7_75t_L g471 ( .A1(n_436), .A2(n_55), .A3(n_56), .B(n_57), .Y(n_471) );
A2O1A1Ixp33_ASAP7_75t_L g472 ( .A1(n_426), .A2(n_58), .B(n_61), .C(n_62), .Y(n_472) );
OAI21x1_ASAP7_75t_SL g473 ( .A1(n_440), .A2(n_63), .B(n_64), .Y(n_473) );
BUFx6f_ASAP7_75t_L g474 ( .A(n_452), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_451), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_441), .Y(n_476) );
AOI21xp5_ASAP7_75t_L g477 ( .A1(n_421), .A2(n_72), .B(n_74), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_447), .Y(n_478) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_429), .A2(n_75), .B(n_77), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g480 ( .A1(n_434), .A2(n_78), .B(n_79), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_432), .Y(n_481) );
AND2x6_ASAP7_75t_L g482 ( .A(n_428), .B(n_84), .Y(n_482) );
AND2x4_ASAP7_75t_L g483 ( .A(n_422), .B(n_85), .Y(n_483) );
BUFx2_ASAP7_75t_SL g484 ( .A(n_430), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g485 ( .A1(n_444), .A2(n_87), .B(n_88), .Y(n_485) );
OAI21xp5_ASAP7_75t_L g486 ( .A1(n_433), .A2(n_90), .B(n_91), .Y(n_486) );
OAI21x1_ASAP7_75t_L g487 ( .A1(n_442), .A2(n_92), .B(n_93), .Y(n_487) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_423), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_446), .B(n_171), .Y(n_489) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_450), .Y(n_490) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_450), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_476), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_462), .Y(n_493) );
OR2x6_ASAP7_75t_L g494 ( .A(n_469), .B(n_96), .Y(n_494) );
AO21x2_ASAP7_75t_L g495 ( .A1(n_470), .A2(n_97), .B(n_98), .Y(n_495) );
HB1xp67_ASAP7_75t_L g496 ( .A(n_464), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_455), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_490), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_487), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_457), .Y(n_500) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_464), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_491), .B(n_100), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_460), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_481), .Y(n_504) );
BUFx3_ASAP7_75t_L g505 ( .A(n_488), .Y(n_505) );
HB1xp67_ASAP7_75t_L g506 ( .A(n_475), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_482), .A2(n_101), .B1(n_102), .B2(n_103), .Y(n_508) );
OA21x2_ASAP7_75t_L g509 ( .A1(n_456), .A2(n_104), .B(n_105), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_461), .Y(n_510) );
AND2x4_ASAP7_75t_L g511 ( .A(n_478), .B(n_112), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_453), .B(n_116), .Y(n_512) );
OA21x2_ASAP7_75t_L g513 ( .A1(n_485), .A2(n_117), .B(n_119), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_453), .B(n_120), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_489), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_465), .Y(n_516) );
OR2x6_ASAP7_75t_L g517 ( .A(n_483), .B(n_123), .Y(n_517) );
INVx2_ASAP7_75t_L g518 ( .A(n_459), .Y(n_518) );
INVx3_ASAP7_75t_L g519 ( .A(n_482), .Y(n_519) );
HB1xp67_ASAP7_75t_SL g520 ( .A(n_482), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_466), .Y(n_521) );
AND2x4_ASAP7_75t_L g522 ( .A(n_486), .B(n_124), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_484), .B(n_125), .Y(n_523) );
BUFx6f_ASAP7_75t_L g524 ( .A(n_474), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_474), .Y(n_525) );
INVx3_ASAP7_75t_L g526 ( .A(n_454), .Y(n_526) );
AOI21x1_ASAP7_75t_L g527 ( .A1(n_454), .A2(n_169), .B(n_131), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_473), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_467), .A2(n_127), .B1(n_132), .B2(n_135), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_471), .Y(n_530) );
AND2x4_ASAP7_75t_L g531 ( .A(n_471), .B(n_136), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_471), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_479), .Y(n_533) );
AO21x2_ASAP7_75t_L g534 ( .A1(n_463), .A2(n_141), .B(n_143), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_468), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_472), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_480), .B(n_144), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_474), .Y(n_539) );
BUFx3_ASAP7_75t_L g540 ( .A(n_490), .Y(n_540) );
HB1xp67_ASAP7_75t_L g541 ( .A(n_464), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_462), .Y(n_542) );
OR2x2_ASAP7_75t_L g543 ( .A(n_458), .B(n_152), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_464), .Y(n_544) );
INVx3_ASAP7_75t_L g545 ( .A(n_494), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_493), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_496), .B(n_153), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_542), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_500), .Y(n_550) );
INVx2_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
NAND2x1_ASAP7_75t_L g552 ( .A(n_519), .B(n_494), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_503), .B(n_154), .Y(n_553) );
INVxp67_ASAP7_75t_L g554 ( .A(n_520), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_504), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_496), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_501), .Y(n_557) );
OR2x2_ASAP7_75t_L g558 ( .A(n_501), .B(n_164), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_515), .B(n_158), .Y(n_559) );
HB1xp67_ASAP7_75t_L g560 ( .A(n_506), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_507), .B(n_163), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_541), .Y(n_562) );
INVx1_ASAP7_75t_L g563 ( .A(n_541), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_492), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_544), .B(n_160), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g566 ( .A1(n_519), .A2(n_161), .B(n_508), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_544), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_515), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_543), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
BUFx3_ASAP7_75t_L g571 ( .A(n_505), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_506), .Y(n_572) );
INVx5_ASAP7_75t_L g573 ( .A(n_517), .Y(n_573) );
AND2x4_ASAP7_75t_L g574 ( .A(n_519), .B(n_517), .Y(n_574) );
OR2x2_ASAP7_75t_L g575 ( .A(n_498), .B(n_540), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_516), .B(n_521), .Y(n_576) );
INVx3_ASAP7_75t_L g577 ( .A(n_511), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_511), .B(n_530), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_502), .B(n_514), .Y(n_579) );
INVxp67_ASAP7_75t_SL g580 ( .A(n_531), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_498), .B(n_512), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_528), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_523), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_536), .B(n_532), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g585 ( .A(n_538), .B(n_535), .C(n_526), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_522), .B(n_526), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_495), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_495), .Y(n_588) );
HB1xp67_ASAP7_75t_L g589 ( .A(n_525), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_522), .B(n_534), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_525), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_529), .A2(n_537), .B1(n_513), .B2(n_509), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_499), .B(n_518), .Y(n_593) );
INVx3_ASAP7_75t_L g594 ( .A(n_524), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_564), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_549), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_550), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_546), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_551), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
INVx1_ASAP7_75t_SL g601 ( .A(n_571), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_568), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_570), .Y(n_603) );
BUFx2_ASAP7_75t_SL g604 ( .A(n_571), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_584), .B(n_539), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_560), .B(n_539), .Y(n_606) );
INVxp67_ASAP7_75t_SL g607 ( .A(n_572), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_556), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g609 ( .A(n_573), .B(n_527), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_572), .B(n_533), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_557), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_583), .B(n_562), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_563), .B(n_567), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_581), .B(n_579), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_569), .B(n_545), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_576), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_554), .B(n_547), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_575), .B(n_574), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_582), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_586), .B(n_580), .Y(n_620) );
HB1xp67_ASAP7_75t_L g621 ( .A(n_589), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_591), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_591), .B(n_578), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_578), .B(n_590), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_552), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_593), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_559), .Y(n_627) );
OR2x2_ASAP7_75t_L g628 ( .A(n_577), .B(n_548), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_604), .Y(n_629) );
INVx2_ASAP7_75t_L g630 ( .A(n_626), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_596), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_597), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_603), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_598), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_599), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_618), .B(n_594), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_614), .B(n_594), .Y(n_637) );
HB1xp67_ASAP7_75t_L g638 ( .A(n_621), .Y(n_638) );
INVx2_ASAP7_75t_L g639 ( .A(n_622), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_600), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_619), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_602), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_616), .B(n_585), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_624), .B(n_565), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_622), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_612), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_608), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_611), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_613), .Y(n_649) );
INVx1_ASAP7_75t_SL g650 ( .A(n_601), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_615), .B(n_566), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_607), .B(n_559), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_595), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_639), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_631), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_646), .B(n_620), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_632), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_649), .B(n_623), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_637), .B(n_617), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_636), .B(n_620), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_633), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_634), .B(n_627), .Y(n_663) );
INVx2_ASAP7_75t_SL g664 ( .A(n_629), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_635), .B(n_621), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_642), .Y(n_666) );
INVxp67_ASAP7_75t_L g667 ( .A(n_638), .Y(n_667) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_638), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_654), .Y(n_669) );
AOI21xp5_ASAP7_75t_SL g670 ( .A1(n_664), .A2(n_651), .B(n_625), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_668), .Y(n_671) );
NOR4xp25_ASAP7_75t_L g672 ( .A(n_664), .B(n_650), .C(n_647), .D(n_648), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_656), .B(n_640), .Y(n_673) );
BUFx2_ASAP7_75t_L g674 ( .A(n_668), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_659), .B(n_644), .Y(n_675) );
OAI21xp5_ASAP7_75t_L g676 ( .A1(n_672), .A2(n_667), .B(n_665), .Y(n_676) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_671), .A2(n_667), .B(n_663), .C(n_661), .Y(n_677) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_670), .A2(n_656), .B(n_655), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g679 ( .A1(n_674), .A2(n_662), .B1(n_657), .B2(n_666), .C(n_658), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_673), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_669), .A2(n_652), .B(n_643), .Y(n_681) );
NOR2xp33_ASAP7_75t_L g682 ( .A(n_675), .B(n_660), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_677), .A2(n_679), .B1(n_676), .B2(n_678), .C(n_681), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_680), .B(n_682), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_684), .B(n_561), .C(n_553), .Y(n_685) );
NAND4xp75_ASAP7_75t_L g686 ( .A(n_683), .B(n_561), .C(n_592), .D(n_605), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_686), .B(n_685), .C(n_558), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_687), .Y(n_688) );
OAI22xp33_ASAP7_75t_L g689 ( .A1(n_688), .A2(n_609), .B1(n_628), .B2(n_630), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_689), .Y(n_690) );
XOR2xp5_ASAP7_75t_L g691 ( .A(n_690), .B(n_609), .Y(n_691) );
XNOR2xp5_ASAP7_75t_L g692 ( .A(n_691), .B(n_606), .Y(n_692) );
OA21x2_ASAP7_75t_L g693 ( .A1(n_692), .A2(n_587), .B(n_588), .Y(n_693) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_693), .A2(n_610), .B1(n_653), .B2(n_645), .Y(n_694) );
endmodule