module fake_netlist_5_1732_n_1091 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_46, n_233, n_21, n_94, n_203, n_245, n_205, n_113, n_38, n_123, n_139, n_105, n_246, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_234, n_17, n_92, n_19, n_149, n_120, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_247, n_188, n_190, n_8, n_201, n_158, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_243, n_239, n_175, n_252, n_169, n_59, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_230, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_253, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_250, n_52, n_88, n_110, n_216, n_1091);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_234;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_175;
input n_252;
input n_169;
input n_59;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_88;
input n_110;
input n_216;

output n_1091;

wire n_924;
wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_977;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_1060;
wire n_316;
wire n_785;
wire n_389;
wire n_855;
wire n_843;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_968;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_913;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_967;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_620;
wire n_643;
wire n_367;
wire n_1055;
wire n_916;
wire n_452;
wire n_885;
wire n_1081;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_980;
wire n_483;
wire n_544;
wire n_683;
wire n_1007;
wire n_780;
wire n_649;
wire n_552;
wire n_1057;
wire n_1051;
wire n_547;
wire n_1066;
wire n_1085;
wire n_721;
wire n_998;
wire n_841;
wire n_1050;
wire n_956;
wire n_564;
wire n_467;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_823;
wire n_725;
wire n_983;
wire n_280;
wire n_744;
wire n_1021;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_690;
wire n_1013;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_1022;
wire n_526;
wire n_915;
wire n_719;
wire n_443;
wire n_372;
wire n_293;
wire n_677;
wire n_864;
wire n_859;
wire n_951;
wire n_821;
wire n_714;
wire n_447;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_321;
wire n_292;
wire n_909;
wire n_625;
wire n_854;
wire n_949;
wire n_621;
wire n_753;
wire n_997;
wire n_455;
wire n_674;
wire n_1008;
wire n_946;
wire n_417;
wire n_932;
wire n_1048;
wire n_612;
wire n_1001;
wire n_498;
wire n_516;
wire n_385;
wire n_933;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_912;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_624;
wire n_825;
wire n_295;
wire n_1010;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_972;
wire n_692;
wire n_986;
wire n_755;
wire n_568;
wire n_509;
wire n_936;
wire n_373;
wire n_820;
wire n_757;
wire n_947;
wire n_1090;
wire n_307;
wire n_633;
wire n_530;
wire n_439;
wire n_1063;
wire n_556;
wire n_1024;
wire n_259;
wire n_448;
wire n_758;
wire n_999;
wire n_668;
wire n_733;
wire n_991;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_941;
wire n_929;
wire n_981;
wire n_1032;
wire n_804;
wire n_867;
wire n_537;
wire n_902;
wire n_587;
wire n_945;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_943;
wire n_399;
wire n_579;
wire n_394;
wire n_341;
wire n_1049;
wire n_992;
wire n_938;
wire n_741;
wire n_548;
wire n_543;
wire n_1068;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_984;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_906;
wire n_905;
wire n_406;
wire n_519;
wire n_470;
wire n_908;
wire n_782;
wire n_919;
wire n_325;
wire n_449;
wire n_1073;
wire n_862;
wire n_900;
wire n_724;
wire n_856;
wire n_546;
wire n_1016;
wire n_760;
wire n_658;
wire n_281;
wire n_918;
wire n_942;
wire n_381;
wire n_291;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_959;
wire n_1077;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_940;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_592;
wire n_920;
wire n_894;
wire n_1046;
wire n_271;
wire n_934;
wire n_1017;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_978;
wire n_964;
wire n_1054;
wire n_654;
wire n_370;
wire n_976;
wire n_343;
wire n_428;
wire n_379;
wire n_308;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_1045;
wire n_1079;
wire n_853;
wire n_603;
wire n_377;
wire n_1078;
wire n_751;
wire n_484;
wire n_775;
wire n_1033;
wire n_988;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_1083;
wire n_600;
wire n_660;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_1009;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_961;
wire n_995;
wire n_955;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_398;
wire n_396;
wire n_1036;
wire n_635;
wire n_347;
wire n_763;
wire n_522;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_1062;
wire n_662;
wire n_459;
wire n_1020;
wire n_646;
wire n_400;
wire n_930;
wire n_436;
wire n_962;
wire n_290;
wire n_580;
wire n_622;
wire n_1040;
wire n_1087;
wire n_723;
wire n_1065;
wire n_1035;
wire n_386;
wire n_578;
wire n_994;
wire n_926;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_1043;
wire n_1071;
wire n_496;
wire n_355;
wire n_958;
wire n_849;
wire n_1034;
wire n_670;
wire n_486;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_922;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_337;
wire n_430;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_528;
wire n_479;
wire n_510;
wire n_680;
wire n_974;
wire n_395;
wire n_553;
wire n_432;
wire n_727;
wire n_839;
wire n_901;
wire n_311;
wire n_813;
wire n_957;
wire n_830;
wire n_773;
wire n_743;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_829;
wire n_749;
wire n_928;
wire n_858;
wire n_1064;
wire n_923;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_939;
wire n_482;
wire n_342;
wire n_517;
wire n_1088;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_1086;
wire n_700;
wire n_796;
wire n_573;
wire n_866;
wire n_969;
wire n_1069;
wire n_1075;
wire n_388;
wire n_761;
wire n_1012;
wire n_1019;
wire n_903;
wire n_1006;
wire n_740;
wire n_304;
wire n_329;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_973;
wire n_277;
wire n_1061;
wire n_338;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_477;
wire n_309;
wire n_512;
wire n_836;
wire n_990;
wire n_462;
wire n_975;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_907;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_1031;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_989;
wire n_1041;
wire n_1039;
wire n_1028;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_893;
wire n_892;
wire n_1015;
wire n_1000;
wire n_891;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_979;
wire n_1002;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_1058;
wire n_362;
wire n_876;
wire n_332;
wire n_1053;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_953;
wire n_601;
wire n_279;
wire n_917;
wire n_1014;
wire n_966;
wire n_987;
wire n_261;
wire n_289;
wire n_745;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_767;
wire n_993;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_982;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_948;
wire n_1076;
wire n_884;
wire n_899;
wire n_345;
wire n_944;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_729;
wire n_730;
wire n_1059;
wire n_1084;
wire n_970;
wire n_911;
wire n_557;
wire n_1005;
wire n_354;
wire n_647;
wire n_575;
wire n_607;
wire n_679;
wire n_513;
wire n_710;
wire n_425;
wire n_527;
wire n_707;
wire n_407;
wire n_480;
wire n_795;
wire n_695;
wire n_832;
wire n_857;
wire n_1072;
wire n_560;
wire n_656;
wire n_340;
wire n_561;
wire n_1044;
wire n_346;
wire n_937;
wire n_393;
wire n_487;
wire n_495;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_910;
wire n_971;
wire n_490;
wire n_805;
wire n_1027;
wire n_326;
wire n_794;
wire n_768;
wire n_921;
wire n_996;
wire n_404;
wire n_686;
wire n_572;
wire n_366;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_596;
wire n_410;
wire n_1042;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_1037;
wire n_1080;
wire n_266;
wire n_272;
wire n_491;
wire n_1074;
wire n_427;
wire n_791;
wire n_732;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_1038;
wire n_1025;
wire n_1082;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_1067;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_931;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_952;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_1023;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_639;
wire n_799;
wire n_914;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_1026;
wire n_319;
wire n_364;
wire n_965;
wire n_927;
wire n_1089;
wire n_536;
wire n_531;
wire n_935;
wire n_1004;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_890;
wire n_1056;
wire n_960;
wire n_759;
wire n_1018;
wire n_438;
wire n_806;
wire n_713;
wire n_1011;
wire n_904;
wire n_985;
wire n_1047;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_827;
wire n_401;
wire n_348;
wire n_1029;
wire n_626;
wire n_925;
wire n_424;
wire n_1003;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_950;
wire n_747;
wire n_278;
wire n_784;

INVx2_ASAP7_75t_SL g256 ( 
.A(n_235),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_21),
.Y(n_257)
);

BUFx2_ASAP7_75t_SL g258 ( 
.A(n_25),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_56),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_229),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_90),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_109),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_45),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_141),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_162),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_151),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_217),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_69),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_254),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_107),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_113),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_191),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_148),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_121),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_13),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_241),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_165),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_203),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_224),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_253),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_227),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_150),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_23),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_185),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_216),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_108),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_99),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_50),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_159),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_129),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_147),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_210),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_87),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_111),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_206),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_237),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_182),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_91),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_167),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_139),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_175),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_146),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_238),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_218),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_200),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_116),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g309 ( 
.A(n_67),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_193),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_144),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g312 ( 
.A(n_222),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_64),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_242),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_9),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_177),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_11),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_112),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_176),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_243),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_184),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_157),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_42),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_160),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_122),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_212),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_201),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_246),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_51),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_173),
.Y(n_330)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_155),
.B(n_138),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_154),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_52),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_40),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_41),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_202),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_239),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_45),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_4),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_60),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_85),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_70),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_230),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_171),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_62),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_10),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_204),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_134),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_194),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_16),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_245),
.Y(n_351)
);

INVx1_ASAP7_75t_SL g352 ( 
.A(n_248),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_247),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_88),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_187),
.Y(n_355)
);

CKINVDCx14_ASAP7_75t_R g356 ( 
.A(n_169),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_226),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_199),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_156),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_0),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_128),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_49),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_36),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_255),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_37),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_101),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_149),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_142),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_68),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_161),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_166),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g372 ( 
.A(n_95),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_140),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_133),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_34),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_49),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_126),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_97),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_164),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_127),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_30),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_211),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_183),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_152),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_195),
.Y(n_385)
);

BUFx6f_ASAP7_75t_L g386 ( 
.A(n_223),
.Y(n_386)
);

INVxp33_ASAP7_75t_SL g387 ( 
.A(n_13),
.Y(n_387)
);

NOR2xp67_ASAP7_75t_L g388 ( 
.A(n_115),
.B(n_17),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_205),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_192),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_43),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_104),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_31),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_50),
.Y(n_394)
);

INVx1_ASAP7_75t_SL g395 ( 
.A(n_215),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_209),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_84),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_136),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_153),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_231),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_189),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_66),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_145),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_119),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_15),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_219),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_197),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_3),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_114),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_36),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_190),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_123),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_221),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_170),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_110),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_3),
.Y(n_416)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_125),
.Y(n_417)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_27),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_96),
.Y(n_419)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_14),
.Y(n_420)
);

BUFx10_ASAP7_75t_L g421 ( 
.A(n_172),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_234),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_236),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_106),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_179),
.Y(n_425)
);

INVx1_ASAP7_75t_SL g426 ( 
.A(n_117),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_174),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_33),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_220),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_198),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_259),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_278),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g433 ( 
.A(n_421),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_418),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_259),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_421),
.Y(n_436)
);

INVx5_ASAP7_75t_L g437 ( 
.A(n_278),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_259),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_259),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_356),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_410),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_292),
.B(n_5),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_410),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_410),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_410),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_278),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_307),
.B(n_5),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_260),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_282),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_276),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_284),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_317),
.Y(n_452)
);

BUFx8_ASAP7_75t_L g453 ( 
.A(n_364),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g454 ( 
.A(n_307),
.B(n_6),
.Y(n_454)
);

INVx5_ASAP7_75t_L g455 ( 
.A(n_282),
.Y(n_455)
);

BUFx12f_ASAP7_75t_L g456 ( 
.A(n_267),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_282),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_330),
.B(n_6),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_262),
.Y(n_459)
);

INVx5_ASAP7_75t_L g460 ( 
.A(n_289),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_360),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_365),
.Y(n_462)
);

OA21x2_ASAP7_75t_L g463 ( 
.A1(n_265),
.A2(n_7),
.B(n_8),
.Y(n_463)
);

HB1xp67_ASAP7_75t_L g464 ( 
.A(n_290),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_289),
.Y(n_465)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_289),
.B(n_57),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_375),
.Y(n_467)
);

AND2x6_ASAP7_75t_L g468 ( 
.A(n_289),
.B(n_386),
.Y(n_468)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_315),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_312),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_275),
.Y(n_472)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_329),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_256),
.B(n_11),
.Y(n_474)
);

BUFx12f_ASAP7_75t_L g475 ( 
.A(n_334),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_386),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_405),
.Y(n_477)
);

OAI22x1_ASAP7_75t_L g478 ( 
.A1(n_335),
.A2(n_12),
.B1(n_14),
.B2(n_16),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_401),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_401),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_401),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_338),
.Y(n_482)
);

BUFx12f_ASAP7_75t_L g483 ( 
.A(n_339),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_320),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_264),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_401),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_266),
.Y(n_487)
);

BUFx8_ASAP7_75t_SL g488 ( 
.A(n_257),
.Y(n_488)
);

INVx5_ASAP7_75t_L g489 ( 
.A(n_354),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_273),
.B(n_18),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_377),
.Y(n_491)
);

INVx5_ASAP7_75t_L g492 ( 
.A(n_377),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_387),
.A2(n_19),
.B1(n_20),
.B2(n_22),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_416),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_427),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_263),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_427),
.Y(n_497)
);

BUFx3_ASAP7_75t_L g498 ( 
.A(n_268),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_393),
.B(n_396),
.Y(n_499)
);

BUFx12f_ASAP7_75t_L g500 ( 
.A(n_346),
.Y(n_500)
);

BUFx12f_ASAP7_75t_L g501 ( 
.A(n_350),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_391),
.B(n_19),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g503 ( 
.A(n_265),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_263),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_294),
.Y(n_505)
);

BUFx2_ASAP7_75t_L g506 ( 
.A(n_363),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_294),
.B(n_20),
.Y(n_507)
);

BUFx8_ASAP7_75t_SL g508 ( 
.A(n_362),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_301),
.B(n_22),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_423),
.B(n_23),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_323),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_323),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_301),
.B(n_313),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_269),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_381),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_313),
.B(n_24),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_333),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_333),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_258),
.Y(n_519)
);

BUFx2_ASAP7_75t_L g520 ( 
.A(n_394),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_408),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_325),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_325),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_270),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_420),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_428),
.Y(n_526)
);

BUFx12f_ASAP7_75t_L g527 ( 
.A(n_271),
.Y(n_527)
);

OAI22x1_ASAP7_75t_SL g528 ( 
.A1(n_314),
.A2(n_327),
.B1(n_328),
.B2(n_321),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_272),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_274),
.Y(n_530)
);

OA21x2_ASAP7_75t_L g531 ( 
.A1(n_379),
.A2(n_26),
.B(n_27),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_279),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_388),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_SL g534 ( 
.A(n_379),
.B(n_28),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_283),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_261),
.B(n_29),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_406),
.Y(n_537)
);

INVx2_ASAP7_75t_SL g538 ( 
.A(n_280),
.Y(n_538)
);

CKINVDCx6p67_ASAP7_75t_R g539 ( 
.A(n_378),
.Y(n_539)
);

INVx5_ASAP7_75t_L g540 ( 
.A(n_406),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_285),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_419),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_419),
.B(n_32),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_287),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_288),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_343),
.Y(n_546)
);

INVx5_ASAP7_75t_L g547 ( 
.A(n_281),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_286),
.Y(n_548)
);

AOI22x1_ASAP7_75t_SL g549 ( 
.A1(n_380),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_291),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_308),
.B(n_58),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_299),
.A2(n_37),
.B(n_38),
.Y(n_552)
);

BUFx8_ASAP7_75t_SL g553 ( 
.A(n_424),
.Y(n_553)
);

AND2x6_ASAP7_75t_L g554 ( 
.A(n_309),
.B(n_59),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_303),
.Y(n_555)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_351),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_304),
.B(n_39),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_311),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_277),
.B(n_42),
.Y(n_559)
);

INVx3_ASAP7_75t_L g560 ( 
.A(n_316),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_326),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_332),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_352),
.B(n_44),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_336),
.Y(n_564)
);

NOR2xp67_ASAP7_75t_L g565 ( 
.A(n_337),
.B(n_46),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_340),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g567 ( 
.A(n_331),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_464),
.B(n_395),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_553),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_472),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_448),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_459),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_443),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_485),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_487),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_530),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_443),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_548),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_527),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_567),
.A2(n_372),
.B1(n_374),
.B2(n_318),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_488),
.Y(n_581)
);

CKINVDCx5p33_ASAP7_75t_R g582 ( 
.A(n_508),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_526),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_438),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_469),
.B(n_397),
.Y(n_585)
);

NAND2xp33_ASAP7_75t_R g586 ( 
.A(n_506),
.B(n_46),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_528),
.B(n_47),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_539),
.Y(n_588)
);

INVx2_ASAP7_75t_SL g589 ( 
.A(n_433),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_442),
.B(n_417),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_498),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_514),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_529),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_439),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_444),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_453),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_432),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_456),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_475),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_436),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_432),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_538),
.B(n_345),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_483),
.Y(n_603)
);

CKINVDCx20_ASAP7_75t_R g604 ( 
.A(n_453),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_473),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_500),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_501),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_432),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_532),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_532),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_445),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_431),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_435),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_R g614 ( 
.A(n_547),
.B(n_293),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_547),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_482),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_534),
.B(n_426),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_441),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_506),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_520),
.Y(n_620)
);

HB1xp67_ASAP7_75t_L g621 ( 
.A(n_515),
.Y(n_621)
);

CKINVDCx5p33_ASAP7_75t_R g622 ( 
.A(n_520),
.Y(n_622)
);

HB1xp67_ASAP7_75t_L g623 ( 
.A(n_495),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_521),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_521),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_491),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_503),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_R g628 ( 
.A(n_555),
.B(n_295),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_497),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_446),
.Y(n_630)
);

BUFx6f_ASAP7_75t_L g631 ( 
.A(n_446),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_505),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_449),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_505),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_449),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_505),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_519),
.Y(n_637)
);

INVxp33_ASAP7_75t_SL g638 ( 
.A(n_563),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_489),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_489),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_R g641 ( 
.A(n_563),
.B(n_296),
.Y(n_641)
);

NOR2xp33_ASAP7_75t_R g642 ( 
.A(n_560),
.B(n_297),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_492),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_492),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_522),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_522),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_466),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_492),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_457),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_555),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_474),
.B(n_348),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_522),
.Y(n_652)
);

NOR3xp33_ASAP7_75t_L g653 ( 
.A(n_580),
.B(n_440),
.C(n_490),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_590),
.B(n_502),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_651),
.B(n_537),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_635),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_617),
.B(n_499),
.Y(n_657)
);

BUFx6f_ASAP7_75t_SL g658 ( 
.A(n_589),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_568),
.B(n_447),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_597),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_585),
.B(n_458),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_627),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_632),
.B(n_634),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_636),
.B(n_437),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_597),
.Y(n_665)
);

INVx5_ASAP7_75t_L g666 ( 
.A(n_597),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_637),
.B(n_559),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_609),
.B(n_510),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_610),
.B(n_536),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_602),
.B(n_550),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_628),
.B(n_507),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_630),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_621),
.B(n_454),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_645),
.B(n_437),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_646),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_647),
.A2(n_557),
.B(n_543),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_652),
.B(n_455),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_633),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_649),
.B(n_455),
.Y(n_679)
);

AND2x6_ASAP7_75t_L g680 ( 
.A(n_584),
.B(n_507),
.Y(n_680)
);

INVxp33_ASAP7_75t_L g681 ( 
.A(n_621),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_650),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_595),
.B(n_455),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_623),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_612),
.B(n_460),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_647),
.B(n_513),
.C(n_509),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_613),
.B(n_460),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_618),
.B(n_460),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_626),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_601),
.B(n_537),
.Y(n_690)
);

INVx3_ASAP7_75t_L g691 ( 
.A(n_601),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_641),
.B(n_516),
.Y(n_692)
);

INVxp67_ASAP7_75t_L g693 ( 
.A(n_600),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_601),
.B(n_540),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_601),
.B(n_540),
.Y(n_695)
);

NOR3xp33_ASAP7_75t_L g696 ( 
.A(n_619),
.B(n_484),
.C(n_471),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_608),
.B(n_540),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_L g698 ( 
.A(n_571),
.B(n_535),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_608),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_572),
.B(n_574),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_608),
.B(n_631),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_608),
.B(n_542),
.Y(n_702)
);

OA21x2_ASAP7_75t_L g703 ( 
.A1(n_594),
.A2(n_544),
.B(n_541),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_575),
.B(n_545),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_631),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_576),
.B(n_578),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_611),
.B(n_551),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_620),
.B(n_561),
.Y(n_708)
);

AO221x1_ASAP7_75t_L g709 ( 
.A1(n_577),
.A2(n_478),
.B1(n_359),
.B2(n_366),
.C(n_353),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_629),
.B(n_546),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_573),
.Y(n_711)
);

INVxp67_ASAP7_75t_L g712 ( 
.A(n_622),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_642),
.B(n_551),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_591),
.B(n_298),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_592),
.B(n_593),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_639),
.B(n_546),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_640),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_624),
.B(n_300),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_625),
.B(n_562),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_643),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_644),
.B(n_564),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_648),
.B(n_546),
.Y(n_722)
);

OAI21xp5_ASAP7_75t_L g723 ( 
.A1(n_686),
.A2(n_552),
.B(n_531),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_700),
.Y(n_724)
);

BUFx6f_ASAP7_75t_L g725 ( 
.A(n_710),
.Y(n_725)
);

AOI22xp5_ASAP7_75t_SL g726 ( 
.A1(n_667),
.A2(n_638),
.B1(n_587),
.B2(n_616),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_668),
.B(n_554),
.Y(n_727)
);

NAND3xp33_ASAP7_75t_SL g728 ( 
.A(n_653),
.B(n_605),
.C(n_434),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_676),
.A2(n_463),
.B1(n_466),
.B2(n_565),
.Y(n_729)
);

AOI22xp5_ASAP7_75t_L g730 ( 
.A1(n_654),
.A2(n_586),
.B1(n_302),
.B2(n_305),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_SL g731 ( 
.A(n_692),
.B(n_615),
.Y(n_731)
);

HB1xp67_ASAP7_75t_L g732 ( 
.A(n_684),
.Y(n_732)
);

OAI22xp5_ASAP7_75t_L g733 ( 
.A1(n_676),
.A2(n_533),
.B1(n_493),
.B2(n_556),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_710),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_669),
.B(n_588),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_655),
.B(n_614),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_655),
.B(n_466),
.Y(n_737)
);

CKINVDCx6p67_ASAP7_75t_R g738 ( 
.A(n_658),
.Y(n_738)
);

OR2x2_ASAP7_75t_L g739 ( 
.A(n_673),
.B(n_581),
.Y(n_739)
);

INVx5_ASAP7_75t_L g740 ( 
.A(n_682),
.Y(n_740)
);

INVx6_ASAP7_75t_L g741 ( 
.A(n_708),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_719),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_663),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_659),
.A2(n_586),
.B1(n_306),
.B2(n_310),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_711),
.Y(n_745)
);

AND2x4_ASAP7_75t_L g746 ( 
.A(n_689),
.B(n_570),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_L g747 ( 
.A1(n_709),
.A2(n_463),
.B1(n_402),
.B2(n_403),
.Y(n_747)
);

INVx5_ASAP7_75t_L g748 ( 
.A(n_680),
.Y(n_748)
);

AOI221xp5_ASAP7_75t_SL g749 ( 
.A1(n_661),
.A2(n_467),
.B1(n_450),
.B2(n_451),
.C(n_452),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_703),
.Y(n_750)
);

NAND2x2_ASAP7_75t_L g751 ( 
.A(n_716),
.B(n_549),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_670),
.B(n_390),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_671),
.B(n_579),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_657),
.B(n_404),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_SL g755 ( 
.A(n_696),
.B(n_525),
.C(n_582),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_681),
.B(n_583),
.Y(n_756)
);

AND2x6_ASAP7_75t_L g757 ( 
.A(n_707),
.B(n_411),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_672),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_698),
.B(n_414),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_656),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_678),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_706),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_704),
.B(n_415),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_722),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_680),
.B(n_422),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_662),
.B(n_461),
.Y(n_766)
);

INVx5_ASAP7_75t_L g767 ( 
.A(n_660),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_680),
.B(n_429),
.Y(n_768)
);

AOI22xp5_ASAP7_75t_L g769 ( 
.A1(n_713),
.A2(n_322),
.B1(n_324),
.B2(n_319),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_675),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_705),
.B(n_524),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_715),
.B(n_607),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_718),
.B(n_569),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_660),
.Y(n_774)
);

AND2x6_ASAP7_75t_SL g775 ( 
.A(n_721),
.B(n_596),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_691),
.B(n_523),
.Y(n_776)
);

INVx5_ASAP7_75t_L g777 ( 
.A(n_660),
.Y(n_777)
);

NAND2x1p5_ASAP7_75t_L g778 ( 
.A(n_714),
.B(n_462),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_717),
.B(n_598),
.Y(n_779)
);

INVx5_ASAP7_75t_L g780 ( 
.A(n_665),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_701),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_679),
.Y(n_782)
);

OR2x6_ASAP7_75t_L g783 ( 
.A(n_712),
.B(n_470),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_690),
.Y(n_784)
);

AO22x1_ASAP7_75t_L g785 ( 
.A1(n_720),
.A2(n_342),
.B1(n_344),
.B2(n_341),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_694),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_693),
.B(n_599),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_695),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_697),
.Y(n_789)
);

OAI21x1_ASAP7_75t_L g790 ( 
.A1(n_664),
.A2(n_504),
.B(n_496),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_658),
.B(n_603),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_685),
.Y(n_792)
);

OR2x6_ASAP7_75t_L g793 ( 
.A(n_687),
.B(n_477),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_665),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_745),
.B(n_494),
.Y(n_795)
);

NAND2xp33_ASAP7_75t_L g796 ( 
.A(n_748),
.B(n_699),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_770),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_743),
.B(n_699),
.Y(n_798)
);

A2O1A1Ixp33_ASAP7_75t_SL g799 ( 
.A1(n_723),
.A2(n_688),
.B(n_677),
.C(n_674),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_742),
.B(n_604),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_774),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_R g802 ( 
.A(n_724),
.B(n_606),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_740),
.B(n_699),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_R g804 ( 
.A(n_762),
.B(n_347),
.Y(n_804)
);

AOI221xp5_ASAP7_75t_L g805 ( 
.A1(n_733),
.A2(n_566),
.B1(n_512),
.B2(n_517),
.C(n_518),
.Y(n_805)
);

AND2x4_ASAP7_75t_SL g806 ( 
.A(n_732),
.B(n_511),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_735),
.B(n_349),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_729),
.A2(n_683),
.B(n_702),
.Y(n_808)
);

NAND2x1p5_ASAP7_75t_L g809 ( 
.A(n_740),
.B(n_666),
.Y(n_809)
);

BUFx3_ASAP7_75t_L g810 ( 
.A(n_741),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_738),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_783),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_728),
.A2(n_400),
.B1(n_357),
.B2(n_358),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_764),
.B(n_355),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

BUFx2_ASAP7_75t_R g816 ( 
.A(n_751),
.Y(n_816)
);

CKINVDCx14_ASAP7_75t_R g817 ( 
.A(n_756),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_771),
.Y(n_818)
);

BUFx8_ASAP7_75t_L g819 ( 
.A(n_746),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_754),
.B(n_361),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_748),
.A2(n_666),
.B(n_465),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_759),
.B(n_367),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_748),
.A2(n_666),
.B(n_465),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_763),
.B(n_725),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_760),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_752),
.A2(n_399),
.B(n_369),
.C(n_430),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_725),
.B(n_368),
.Y(n_827)
);

AND2x2_ASAP7_75t_SL g828 ( 
.A(n_773),
.B(n_566),
.Y(n_828)
);

AOI22xp33_ASAP7_75t_SL g829 ( 
.A1(n_726),
.A2(n_412),
.B1(n_371),
.B2(n_373),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_734),
.B(n_370),
.Y(n_830)
);

OAI21xp5_ASAP7_75t_L g831 ( 
.A1(n_727),
.A2(n_468),
.B(n_383),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_781),
.B(n_382),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_774),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_761),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_741),
.B(n_384),
.Y(n_835)
);

BUFx6f_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

NAND2x1_ASAP7_75t_L g837 ( 
.A(n_750),
.B(n_468),
.Y(n_837)
);

INVx4_ASAP7_75t_L g838 ( 
.A(n_767),
.Y(n_838)
);

AND3x1_ASAP7_75t_SL g839 ( 
.A(n_755),
.B(n_47),
.C(n_48),
.Y(n_839)
);

XNOR2xp5_ASAP7_75t_L g840 ( 
.A(n_772),
.B(n_385),
.Y(n_840)
);

AO21x1_ASAP7_75t_L g841 ( 
.A1(n_737),
.A2(n_48),
.B(n_51),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_730),
.B(n_558),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_784),
.B(n_389),
.Y(n_843)
);

O2A1O1Ixp33_ASAP7_75t_L g844 ( 
.A1(n_736),
.A2(n_425),
.B(n_398),
.C(n_407),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_758),
.Y(n_845)
);

AOI22xp33_ASAP7_75t_L g846 ( 
.A1(n_757),
.A2(n_747),
.B1(n_789),
.B2(n_788),
.Y(n_846)
);

AND2x2_ASAP7_75t_L g847 ( 
.A(n_744),
.B(n_392),
.Y(n_847)
);

BUFx6f_ASAP7_75t_L g848 ( 
.A(n_777),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_786),
.B(n_409),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_757),
.A2(n_413),
.B1(n_468),
.B2(n_480),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_790),
.Y(n_851)
);

OR2x2_ASAP7_75t_L g852 ( 
.A(n_739),
.B(n_52),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_757),
.Y(n_853)
);

AOI21xp33_ASAP7_75t_L g854 ( 
.A1(n_807),
.A2(n_768),
.B(n_765),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_819),
.Y(n_855)
);

OAI21x1_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_794),
.B(n_776),
.Y(n_856)
);

INVx6_ASAP7_75t_L g857 ( 
.A(n_836),
.Y(n_857)
);

OAI21xp5_ASAP7_75t_L g858 ( 
.A1(n_808),
.A2(n_749),
.B(n_782),
.Y(n_858)
);

BUFx3_ASAP7_75t_L g859 ( 
.A(n_810),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_797),
.Y(n_860)
);

AO21x2_ASAP7_75t_L g861 ( 
.A1(n_799),
.A2(n_731),
.B(n_769),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_836),
.Y(n_862)
);

CKINVDCx16_ASAP7_75t_R g863 ( 
.A(n_802),
.Y(n_863)
);

CKINVDCx20_ASAP7_75t_R g864 ( 
.A(n_811),
.Y(n_864)
);

INVx1_ASAP7_75t_SL g865 ( 
.A(n_806),
.Y(n_865)
);

AOI22x1_ASAP7_75t_L g866 ( 
.A1(n_831),
.A2(n_792),
.B1(n_778),
.B2(n_793),
.Y(n_866)
);

INVx1_ASAP7_75t_SL g867 ( 
.A(n_824),
.Y(n_867)
);

OAI21x1_ASAP7_75t_L g868 ( 
.A1(n_837),
.A2(n_753),
.B(n_779),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_848),
.Y(n_869)
);

OR2x6_ASAP7_75t_L g870 ( 
.A(n_836),
.B(n_787),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_828),
.B(n_791),
.Y(n_871)
);

AOI22x1_ASAP7_75t_L g872 ( 
.A1(n_818),
.A2(n_785),
.B1(n_486),
.B2(n_481),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_804),
.Y(n_873)
);

OA21x2_ASAP7_75t_L g874 ( 
.A1(n_846),
.A2(n_780),
.B(n_777),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_798),
.B(n_780),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_848),
.Y(n_876)
);

INVx3_ASAP7_75t_L g877 ( 
.A(n_848),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_795),
.B(n_780),
.Y(n_878)
);

AOI21x1_ASAP7_75t_L g879 ( 
.A1(n_827),
.A2(n_479),
.B(n_476),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_834),
.B(n_61),
.Y(n_880)
);

NAND3xp33_ASAP7_75t_L g881 ( 
.A(n_813),
.B(n_775),
.C(n_486),
.Y(n_881)
);

INVx4_ASAP7_75t_L g882 ( 
.A(n_801),
.Y(n_882)
);

HB1xp67_ASAP7_75t_L g883 ( 
.A(n_801),
.Y(n_883)
);

AND2x4_ASAP7_75t_L g884 ( 
.A(n_795),
.B(n_63),
.Y(n_884)
);

INVx5_ASAP7_75t_SL g885 ( 
.A(n_801),
.Y(n_885)
);

BUFx12f_ASAP7_75t_L g886 ( 
.A(n_852),
.Y(n_886)
);

INVx1_ASAP7_75t_SL g887 ( 
.A(n_833),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_845),
.Y(n_888)
);

OAI21x1_ASAP7_75t_L g889 ( 
.A1(n_821),
.A2(n_168),
.B(n_252),
.Y(n_889)
);

BUFx3_ASAP7_75t_L g890 ( 
.A(n_833),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_825),
.Y(n_891)
);

OR2x2_ASAP7_75t_L g892 ( 
.A(n_800),
.B(n_814),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_838),
.Y(n_893)
);

HB1xp67_ASAP7_75t_L g894 ( 
.A(n_812),
.Y(n_894)
);

NAND2x1p5_ASAP7_75t_L g895 ( 
.A(n_838),
.B(n_476),
.Y(n_895)
);

OAI21x1_ASAP7_75t_SL g896 ( 
.A1(n_841),
.A2(n_163),
.B(n_251),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_842),
.B(n_65),
.Y(n_897)
);

BUFx2_ASAP7_75t_R g898 ( 
.A(n_840),
.Y(n_898)
);

INVx1_ASAP7_75t_SL g899 ( 
.A(n_830),
.Y(n_899)
);

OAI21x1_ASAP7_75t_L g900 ( 
.A1(n_823),
.A2(n_178),
.B(n_250),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_796),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_832),
.B(n_53),
.Y(n_902)
);

CKINVDCx16_ASAP7_75t_R g903 ( 
.A(n_817),
.Y(n_903)
);

BUFx3_ASAP7_75t_L g904 ( 
.A(n_815),
.Y(n_904)
);

AO21x2_ASAP7_75t_L g905 ( 
.A1(n_820),
.A2(n_158),
.B(n_249),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_867),
.B(n_847),
.Y(n_906)
);

CKINVDCx6p67_ASAP7_75t_R g907 ( 
.A(n_855),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_860),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_869),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_857),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_888),
.Y(n_911)
);

NAND2x1p5_ASAP7_75t_L g912 ( 
.A(n_876),
.B(n_893),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_891),
.Y(n_913)
);

INVx6_ASAP7_75t_L g914 ( 
.A(n_876),
.Y(n_914)
);

BUFx2_ASAP7_75t_R g915 ( 
.A(n_873),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_899),
.B(n_843),
.Y(n_916)
);

AND2x2_ASAP7_75t_L g917 ( 
.A(n_871),
.B(n_829),
.Y(n_917)
);

INVx3_ASAP7_75t_SL g918 ( 
.A(n_863),
.Y(n_918)
);

AOI22xp33_ASAP7_75t_SL g919 ( 
.A1(n_898),
.A2(n_835),
.B1(n_839),
.B2(n_853),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_876),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_876),
.B(n_803),
.Y(n_921)
);

BUFx2_ASAP7_75t_R g922 ( 
.A(n_859),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_880),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_862),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_894),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_902),
.A2(n_805),
.B1(n_822),
.B2(n_849),
.Y(n_926)
);

INVx8_ASAP7_75t_L g927 ( 
.A(n_869),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_883),
.Y(n_928)
);

OR2x6_ASAP7_75t_L g929 ( 
.A(n_870),
.B(n_809),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_884),
.Y(n_930)
);

CKINVDCx14_ASAP7_75t_R g931 ( 
.A(n_864),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_877),
.Y(n_932)
);

OAI22xp33_ASAP7_75t_L g933 ( 
.A1(n_892),
.A2(n_850),
.B1(n_816),
.B2(n_486),
.Y(n_933)
);

OAI21x1_ASAP7_75t_L g934 ( 
.A1(n_856),
.A2(n_844),
.B(n_826),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_877),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_862),
.Y(n_936)
);

CKINVDCx6p67_ASAP7_75t_R g937 ( 
.A(n_903),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_887),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_894),
.Y(n_939)
);

CKINVDCx6p67_ASAP7_75t_R g940 ( 
.A(n_864),
.Y(n_940)
);

CKINVDCx11_ASAP7_75t_R g941 ( 
.A(n_886),
.Y(n_941)
);

HB1xp67_ASAP7_75t_L g942 ( 
.A(n_890),
.Y(n_942)
);

INVx2_ASAP7_75t_L g943 ( 
.A(n_874),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_869),
.Y(n_944)
);

INVx6_ASAP7_75t_L g945 ( 
.A(n_857),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_904),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_874),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_930),
.B(n_878),
.Y(n_948)
);

XNOR2x1_ASAP7_75t_L g949 ( 
.A(n_917),
.B(n_881),
.Y(n_949)
);

AND2x4_ASAP7_75t_SL g950 ( 
.A(n_920),
.B(n_882),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_916),
.B(n_865),
.Y(n_951)
);

NOR3xp33_ASAP7_75t_SL g952 ( 
.A(n_933),
.B(n_897),
.C(n_898),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_916),
.B(n_865),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_906),
.B(n_870),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_908),
.Y(n_955)
);

CKINVDCx16_ASAP7_75t_R g956 ( 
.A(n_931),
.Y(n_956)
);

AOI22xp33_ASAP7_75t_SL g957 ( 
.A1(n_931),
.A2(n_866),
.B1(n_896),
.B2(n_897),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_919),
.B(n_885),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_919),
.B(n_868),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_913),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_918),
.B(n_879),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_927),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_928),
.B(n_895),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_911),
.Y(n_964)
);

AND2x4_ASAP7_75t_L g965 ( 
.A(n_924),
.B(n_901),
.Y(n_965)
);

NAND2x1_ASAP7_75t_L g966 ( 
.A(n_920),
.B(n_875),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_909),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_918),
.B(n_875),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_927),
.B(n_889),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_926),
.A2(n_854),
.B(n_858),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_R g971 ( 
.A(n_940),
.B(n_71),
.Y(n_971)
);

AO31x2_ASAP7_75t_L g972 ( 
.A1(n_943),
.A2(n_861),
.A3(n_872),
.B(n_905),
.Y(n_972)
);

OR2x6_ASAP7_75t_L g973 ( 
.A(n_927),
.B(n_900),
.Y(n_973)
);

INVx2_ASAP7_75t_SL g974 ( 
.A(n_945),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_R g975 ( 
.A(n_936),
.B(n_72),
.Y(n_975)
);

AOI22xp5_ASAP7_75t_L g976 ( 
.A1(n_937),
.A2(n_479),
.B1(n_55),
.B2(n_56),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_929),
.B(n_73),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_909),
.Y(n_978)
);

OAI22xp33_ASAP7_75t_L g979 ( 
.A1(n_946),
.A2(n_54),
.B1(n_55),
.B2(n_74),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_L g980 ( 
.A1(n_923),
.A2(n_75),
.B1(n_76),
.B2(n_77),
.Y(n_980)
);

BUFx4f_ASAP7_75t_SL g981 ( 
.A(n_907),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_929),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_938),
.B(n_925),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_938),
.B(n_81),
.Y(n_984)
);

NOR3xp33_ASAP7_75t_SL g985 ( 
.A(n_939),
.B(n_82),
.C(n_83),
.Y(n_985)
);

AND2x4_ASAP7_75t_SL g986 ( 
.A(n_929),
.B(n_86),
.Y(n_986)
);

INVxp67_ASAP7_75t_L g987 ( 
.A(n_922),
.Y(n_987)
);

NAND2xp33_ASAP7_75t_R g988 ( 
.A(n_932),
.B(n_89),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_L g989 ( 
.A1(n_949),
.A2(n_959),
.B1(n_970),
.B2(n_979),
.Y(n_989)
);

AND2x4_ASAP7_75t_L g990 ( 
.A(n_969),
.B(n_947),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_983),
.B(n_942),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_960),
.B(n_935),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_955),
.Y(n_993)
);

INVx2_ASAP7_75t_L g994 ( 
.A(n_972),
.Y(n_994)
);

INVx2_ASAP7_75t_L g995 ( 
.A(n_964),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_951),
.B(n_944),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_953),
.B(n_954),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_969),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_965),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_973),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_973),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_958),
.B(n_934),
.Y(n_1002)
);

BUFx2_ASAP7_75t_L g1003 ( 
.A(n_968),
.Y(n_1003)
);

NOR2xp33_ASAP7_75t_R g1004 ( 
.A(n_988),
.B(n_941),
.Y(n_1004)
);

AOI221xp5_ASAP7_75t_L g1005 ( 
.A1(n_976),
.A2(n_910),
.B1(n_921),
.B2(n_912),
.C(n_922),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_963),
.B(n_912),
.Y(n_1006)
);

OAI21xp5_ASAP7_75t_SL g1007 ( 
.A1(n_957),
.A2(n_921),
.B(n_915),
.Y(n_1007)
);

BUFx2_ASAP7_75t_SL g1008 ( 
.A(n_977),
.Y(n_1008)
);

BUFx3_ASAP7_75t_L g1009 ( 
.A(n_966),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_948),
.B(n_92),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_948),
.B(n_93),
.Y(n_1011)
);

AND2x2_ASAP7_75t_L g1012 ( 
.A(n_985),
.B(n_94),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_952),
.B(n_98),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_977),
.B(n_100),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_984),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_961),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_967),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_978),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_978),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

AND2x2_ASAP7_75t_L g1021 ( 
.A(n_987),
.B(n_102),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_982),
.Y(n_1022)
);

AND2x2_ASAP7_75t_L g1023 ( 
.A(n_956),
.B(n_103),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_986),
.B(n_105),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_974),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_980),
.Y(n_1026)
);

AND2x4_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_950),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_997),
.B(n_971),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_991),
.B(n_941),
.Y(n_1029)
);

NAND2x1p5_ASAP7_75t_L g1030 ( 
.A(n_1009),
.B(n_975),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_993),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_1015),
.B(n_981),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_1022),
.A2(n_914),
.B1(n_118),
.B2(n_120),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_1016),
.B(n_914),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_1001),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_995),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_998),
.B(n_124),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_SL g1038 ( 
.A(n_1008),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_1002),
.B(n_130),
.Y(n_1039)
);

NAND3xp33_ASAP7_75t_L g1040 ( 
.A(n_989),
.B(n_131),
.C(n_132),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_994),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_1006),
.B(n_244),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_996),
.B(n_135),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_999),
.B(n_137),
.Y(n_1044)
);

AND2x4_ASAP7_75t_L g1045 ( 
.A(n_1000),
.B(n_143),
.Y(n_1045)
);

INVx4_ASAP7_75t_L g1046 ( 
.A(n_1037),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_SL g1047 ( 
.A(n_1030),
.B(n_1004),
.Y(n_1047)
);

NOR2x1_ASAP7_75t_L g1048 ( 
.A(n_1028),
.B(n_1009),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_1031),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1030),
.B(n_1003),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_1031),
.Y(n_1051)
);

HB1xp67_ASAP7_75t_L g1052 ( 
.A(n_1041),
.Y(n_1052)
);

NOR2xp67_ASAP7_75t_L g1053 ( 
.A(n_1032),
.B(n_1035),
.Y(n_1053)
);

AND2x2_ASAP7_75t_SL g1054 ( 
.A(n_1044),
.B(n_1014),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_1027),
.Y(n_1055)
);

BUFx2_ASAP7_75t_L g1056 ( 
.A(n_1027),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_1036),
.B(n_999),
.Y(n_1057)
);

AOI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1047),
.A2(n_1040),
.B1(n_1022),
.B2(n_1026),
.Y(n_1058)
);

AOI211xp5_ASAP7_75t_L g1059 ( 
.A1(n_1050),
.A2(n_1005),
.B(n_1007),
.C(n_1013),
.Y(n_1059)
);

AOI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_1050),
.A2(n_1026),
.B1(n_1008),
.B2(n_1033),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_1049),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_1054),
.A2(n_1038),
.B1(n_1034),
.B2(n_1029),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_1053),
.B(n_990),
.Y(n_1063)
);

OAI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1060),
.A2(n_1046),
.B1(n_1039),
.B2(n_1048),
.Y(n_1064)
);

A2O1A1Ixp33_ASAP7_75t_L g1065 ( 
.A1(n_1059),
.A2(n_1023),
.B(n_1013),
.C(n_1012),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_1061),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1058),
.A2(n_1012),
.B(n_1045),
.Y(n_1067)
);

INVx2_ASAP7_75t_L g1068 ( 
.A(n_1063),
.Y(n_1068)
);

AOI22xp33_ASAP7_75t_L g1069 ( 
.A1(n_1062),
.A2(n_1046),
.B1(n_1023),
.B2(n_1056),
.Y(n_1069)
);

OAI22xp5_ASAP7_75t_L g1070 ( 
.A1(n_1065),
.A2(n_1060),
.B1(n_1038),
.B2(n_1046),
.Y(n_1070)
);

AOI21xp33_ASAP7_75t_L g1071 ( 
.A1(n_1064),
.A2(n_1057),
.B(n_1043),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_1069),
.B(n_1055),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_SL g1073 ( 
.A1(n_1067),
.A2(n_1014),
.B(n_1021),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_1070),
.A2(n_1025),
.B(n_1066),
.C(n_1068),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1073),
.B(n_1042),
.Y(n_1075)
);

AOI21xp33_ASAP7_75t_L g1076 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1071),
.Y(n_1076)
);

AND4x1_ASAP7_75t_L g1077 ( 
.A(n_1075),
.B(n_1024),
.C(n_1010),
.D(n_1011),
.Y(n_1077)
);

OAI221xp5_ASAP7_75t_L g1078 ( 
.A1(n_1077),
.A2(n_1051),
.B1(n_1049),
.B2(n_1020),
.C(n_1019),
.Y(n_1078)
);

AOI211xp5_ASAP7_75t_L g1079 ( 
.A1(n_1076),
.A2(n_1017),
.B(n_992),
.C(n_1018),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_1078),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_1079),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_1080),
.B(n_1052),
.Y(n_1082)
);

AND2x4_ASAP7_75t_L g1083 ( 
.A(n_1082),
.B(n_1081),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1083),
.Y(n_1084)
);

OAI31xp33_ASAP7_75t_L g1085 ( 
.A1(n_1084),
.A2(n_240),
.A3(n_180),
.B(n_181),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1085),
.B(n_186),
.Y(n_1086)
);

OR2x2_ASAP7_75t_L g1087 ( 
.A(n_1086),
.B(n_188),
.Y(n_1087)
);

XNOR2x1_ASAP7_75t_L g1088 ( 
.A(n_1087),
.B(n_196),
.Y(n_1088)
);

AOI22xp5_ASAP7_75t_SL g1089 ( 
.A1(n_1088),
.A2(n_207),
.B1(n_208),
.B2(n_213),
.Y(n_1089)
);

OR2x6_ASAP7_75t_L g1090 ( 
.A(n_1089),
.B(n_225),
.Y(n_1090)
);

AOI22xp33_ASAP7_75t_L g1091 ( 
.A1(n_1090),
.A2(n_228),
.B1(n_232),
.B2(n_233),
.Y(n_1091)
);


endmodule