module fake_jpeg_3616_n_166 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_166);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_166;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

INVx4_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_6),
.B(n_10),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_20),
.Y(n_31)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_19),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_32),
.B(n_11),
.Y(n_65)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_33),
.B(n_37),
.Y(n_64)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g59 ( 
.A(n_34),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_1),
.CON(n_35),
.SN(n_35)
);

NOR2x1_ASAP7_75t_L g66 ( 
.A(n_35),
.B(n_23),
.Y(n_66)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_49),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_47),
.Y(n_58)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_20),
.Y(n_44)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_44),
.Y(n_82)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_5),
.Y(n_84)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_22),
.Y(n_48)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_22),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g50 ( 
.A(n_13),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_51),
.Y(n_61)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_52),
.B(n_53),
.Y(n_74)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_15),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_54),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_55),
.B(n_11),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_32),
.B(n_26),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_56),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_23),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_83),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_52),
.A2(n_18),
.B1(n_27),
.B2(n_14),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_72),
.A2(n_38),
.B1(n_49),
.B2(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_40),
.B(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_79),
.B(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_29),
.B(n_27),
.Y(n_83)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

NOR3xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_91),
.C(n_95),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_94),
.B1(n_97),
.B2(n_82),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_61),
.B(n_34),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_87),
.A2(n_58),
.B(n_57),
.Y(n_107)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_89),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_61),
.B(n_39),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_103),
.C(n_82),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_74),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_68),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_94)
);

INVx13_ASAP7_75t_L g95 ( 
.A(n_59),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_72),
.A2(n_8),
.B1(n_63),
.B2(n_77),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_64),
.B(n_67),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_98),
.B(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_74),
.Y(n_99)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_104),
.Y(n_112)
);

OR2x2_ASAP7_75t_SL g103 ( 
.A(n_66),
.B(n_57),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_58),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_110),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

NAND2xp33_ASAP7_75t_R g122 ( 
.A(n_108),
.B(n_119),
.Y(n_122)
);

MAJx2_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_81),
.C(n_62),
.Y(n_110)
);

AOI32xp33_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_88),
.A3(n_91),
.B1(n_103),
.B2(n_99),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_86),
.B1(n_97),
.B2(n_90),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_100),
.B(n_62),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_96),
.B(n_100),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_121),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_85),
.Y(n_118)
);

INVxp67_ASAP7_75t_SL g124 ( 
.A(n_118),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_69),
.Y(n_121)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_120),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_125),
.B(n_126),
.Y(n_140)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NOR3xp33_ASAP7_75t_SL g129 ( 
.A(n_117),
.B(n_95),
.C(n_87),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_129),
.B(n_113),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_131),
.A2(n_123),
.B1(n_128),
.B2(n_127),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_89),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_109),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_132),
.B(n_108),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_134),
.A2(n_105),
.B(n_116),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_123),
.B(n_130),
.C(n_133),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_141),
.C(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_109),
.A3(n_121),
.B1(n_106),
.B2(n_107),
.C(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_130),
.B(n_90),
.C(n_112),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_124),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_142),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_143),
.B(n_149),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_135),
.B(n_122),
.C(n_129),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_144),
.B(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_131),
.C(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_140),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_102),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_147),
.B(n_138),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_151),
.B(n_152),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_148),
.A2(n_134),
.B1(n_70),
.B2(n_92),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g157 ( 
.A1(n_154),
.A2(n_104),
.B(n_8),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_150),
.A2(n_151),
.B(n_153),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_156),
.B(n_150),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_143),
.B(n_76),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_157),
.B(n_78),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_159),
.B(n_75),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_160),
.B(n_161),
.Y(n_163)
);

OAI21x1_ASAP7_75t_L g161 ( 
.A1(n_158),
.A2(n_69),
.B(n_78),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_75),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_164),
.B(n_70),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g166 ( 
.A(n_165),
.B(n_163),
.Y(n_166)
);


endmodule