module real_aes_5419_n_7 (n_4, n_0, n_3, n_5, n_2, n_6, n_1, n_7);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_6;
input n_1;
output n_7;
wire n_17;
wire n_22;
wire n_13;
wire n_24;
wire n_12;
wire n_19;
wire n_25;
wire n_14;
wire n_11;
wire n_16;
wire n_15;
wire n_23;
wire n_9;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_8;
wire n_10;
NAND3xp33_ASAP7_75t_SL g20 ( .A(n_0), .B(n_21), .C(n_23), .Y(n_20) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_1), .Y(n_22) );
INVx1_ASAP7_75t_L g17 ( .A(n_2), .Y(n_17) );
BUFx6f_ASAP7_75t_L g25 ( .A(n_3), .Y(n_25) );
INVx2_ASAP7_75t_SL g11 ( .A(n_4), .Y(n_11) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
AOI32xp33_ASAP7_75t_L g7 ( .A1(n_8), .A2(n_14), .A3(n_15), .B1(n_16), .B2(n_18), .Y(n_7) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_9), .B(n_12), .Y(n_8) );
OAI21xp33_ASAP7_75t_SL g18 ( .A1(n_9), .A2(n_16), .B(n_19), .Y(n_18) );
AOI21xp5_ASAP7_75t_L g19 ( .A1(n_9), .A2(n_20), .B(n_26), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g26 ( .A(n_9), .B(n_13), .Y(n_26) );
HB1xp67_ASAP7_75t_L g9 ( .A(n_10), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_11), .Y(n_10) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_13), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_15), .Y(n_14) );
INVxp67_ASAP7_75t_L g16 ( .A(n_17), .Y(n_16) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
BUFx2_ASAP7_75t_L g23 ( .A(n_24), .Y(n_23) );
HB1xp67_ASAP7_75t_L g24 ( .A(n_25), .Y(n_24) );
endmodule