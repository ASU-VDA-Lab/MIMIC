module fake_jpeg_11539_n_370 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_370);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_370;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_4),
.B(n_7),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx10_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_0),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_14),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_45),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_46),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_49),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_51),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_26),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_52),
.B(n_84),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_53),
.B(n_40),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_54),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_13),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_55),
.B(n_56),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_34),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_57),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_28),
.Y(n_58)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_58),
.Y(n_104)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_26),
.Y(n_60)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_29),
.Y(n_62)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_62),
.Y(n_89)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_22),
.B(n_12),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_64),
.B(n_74),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_12),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_66),
.B(n_75),
.Y(n_98)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx4f_ASAP7_75t_SL g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx16f_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_72),
.Y(n_103)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_73),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_23),
.B(n_11),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_23),
.B(n_0),
.Y(n_75)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_76),
.Y(n_125)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx11_ASAP7_75t_L g100 ( 
.A(n_77),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_78),
.B(n_83),
.Y(n_121)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_79),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_34),
.B(n_1),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_1),
.Y(n_118)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_32),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_92),
.B(n_93),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_36),
.B1(n_20),
.B2(n_30),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_99),
.A2(n_54),
.B1(n_47),
.B2(n_46),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_69),
.B(n_18),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_128),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_69),
.B(n_18),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_117),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_36),
.B1(n_40),
.B2(n_20),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_112),
.A2(n_113),
.B1(n_124),
.B2(n_126),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_83),
.A2(n_40),
.B1(n_36),
.B2(n_30),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_35),
.Y(n_117)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_123),
.Y(n_162)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_77),
.A2(n_30),
.B1(n_41),
.B2(n_37),
.Y(n_119)
);

AO22x1_ASAP7_75t_SL g168 ( 
.A1(n_119),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_48),
.B(n_35),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_43),
.A2(n_31),
.B1(n_27),
.B2(n_37),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_49),
.A2(n_32),
.B1(n_31),
.B2(n_41),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_78),
.B(n_21),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_137),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_51),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_62),
.B(n_21),
.Y(n_131)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_65),
.B(n_17),
.Y(n_132)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_17),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_139),
.B(n_140),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_134),
.Y(n_140)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_94),
.Y(n_142)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_142),
.Y(n_193)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_111),
.Y(n_143)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_99),
.A2(n_72),
.B1(n_44),
.B2(n_58),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_144),
.A2(n_147),
.B1(n_175),
.B2(n_180),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_100),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_173),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_1),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_148),
.B(n_153),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_70),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_157),
.C(n_171),
.Y(n_215)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_151),
.Y(n_187)
);

INVx4_ASAP7_75t_SL g152 ( 
.A(n_100),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_106),
.B(n_2),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_45),
.B1(n_31),
.B2(n_32),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_155),
.A2(n_181),
.B1(n_157),
.B2(n_164),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_116),
.A2(n_42),
.B1(n_15),
.B2(n_6),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_121),
.A2(n_15),
.B(n_42),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_98),
.B(n_2),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_158),
.B(n_165),
.Y(n_205)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_94),
.Y(n_159)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_133),
.A2(n_15),
.B1(n_5),
.B2(n_6),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_161),
.B(n_166),
.Y(n_192)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_163),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_119),
.B(n_5),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g167 ( 
.A(n_88),
.Y(n_167)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_167),
.Y(n_189)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_168),
.A2(n_183),
.B1(n_122),
.B2(n_111),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_89),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_169),
.A2(n_135),
.B1(n_122),
.B2(n_129),
.Y(n_185)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_89),
.Y(n_170)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_133),
.B(n_9),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_90),
.B(n_9),
.Y(n_172)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_172),
.A2(n_177),
.B(n_182),
.C(n_108),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_112),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_104),
.A2(n_10),
.B1(n_120),
.B2(n_110),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_176),
.Y(n_190)
);

FAx1_ASAP7_75t_SL g177 ( 
.A(n_121),
.B(n_10),
.CI(n_107),
.CON(n_177),
.SN(n_177)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_111),
.Y(n_179)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_179),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_104),
.A2(n_135),
.B1(n_110),
.B2(n_130),
.Y(n_180)
);

OAI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_126),
.A2(n_10),
.B1(n_113),
.B2(n_130),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_102),
.B(n_10),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_95),
.A2(n_97),
.B1(n_115),
.B2(n_91),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_185),
.Y(n_246)
);

OA22x2_ASAP7_75t_L g244 ( 
.A1(n_194),
.A2(n_198),
.B1(n_208),
.B2(n_142),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_174),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_195),
.B(n_209),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_165),
.A2(n_95),
.B1(n_97),
.B2(n_88),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_125),
.B1(n_87),
.B2(n_91),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_201),
.A2(n_219),
.B1(n_167),
.B2(n_159),
.Y(n_241)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_206),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_150),
.B(n_154),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_207),
.B(n_210),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_160),
.B(n_129),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_138),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_211),
.B(n_213),
.Y(n_224)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_183),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_183),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_87),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_216),
.B(n_218),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_153),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_217),
.B(n_172),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_149),
.B(n_108),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_147),
.A2(n_145),
.B1(n_162),
.B2(n_168),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_168),
.B(n_177),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_222),
.A2(n_235),
.B(n_212),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_220),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_225),
.B(n_226),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_220),
.B(n_145),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_227),
.B(n_232),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_215),
.A2(n_177),
.B(n_162),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_228),
.A2(n_239),
.B(n_240),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_229),
.B(n_230),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_204),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_215),
.B(n_171),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_231),
.B(n_234),
.Y(n_268)
);

OAI22x1_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_183),
.B1(n_167),
.B2(n_170),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_188),
.B(n_182),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_236),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_213),
.B(n_171),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_203),
.A2(n_208),
.B(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_158),
.Y(n_236)
);

AOI21xp33_ASAP7_75t_L g237 ( 
.A1(n_205),
.A2(n_148),
.B(n_161),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_237),
.B(n_199),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_192),
.B(n_155),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_245),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_192),
.A2(n_152),
.B(n_108),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_241),
.A2(n_249),
.B1(n_189),
.B2(n_190),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_143),
.Y(n_242)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_242),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_193),
.Y(n_243)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_243),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_244),
.A2(n_202),
.B1(n_199),
.B2(n_193),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_190),
.B(n_209),
.C(n_187),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_200),
.A2(n_208),
.B1(n_198),
.B2(n_189),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_197),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_187),
.B(n_179),
.Y(n_251)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_251),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_252),
.A2(n_260),
.B1(n_253),
.B2(n_259),
.Y(n_296)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_247),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_255),
.Y(n_281)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_259),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_238),
.A2(n_202),
.B1(n_186),
.B2(n_206),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_261),
.A2(n_267),
.B1(n_249),
.B2(n_250),
.Y(n_283)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_251),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_265),
.B(n_248),
.Y(n_288)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_224),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_272),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_242),
.A2(n_186),
.B1(n_184),
.B2(n_211),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_240),
.B(n_235),
.Y(n_279)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_224),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_273),
.B(n_230),
.Y(n_280)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_275),
.B(n_184),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_264),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_277),
.B(n_294),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_279),
.A2(n_285),
.B(n_222),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_280),
.B(n_288),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_268),
.B(n_231),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_282),
.B(n_286),
.C(n_287),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_283),
.A2(n_284),
.B1(n_252),
.B2(n_253),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_270),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_266),
.A2(n_246),
.B1(n_242),
.B2(n_248),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_231),
.C(n_225),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_269),
.B(n_226),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_263),
.B(n_258),
.C(n_276),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_290),
.C(n_291),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_258),
.B(n_228),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_227),
.C(n_234),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_234),
.C(n_233),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_292),
.B(n_275),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_254),
.Y(n_294)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_296),
.Y(n_301)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_298),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_295),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_299),
.B(n_307),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_262),
.Y(n_304)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_304),
.Y(n_330)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_298),
.Y(n_305)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_305),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_308),
.B1(n_296),
.B2(n_289),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_297),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_283),
.A2(n_270),
.B1(n_260),
.B2(n_256),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_309),
.B(n_316),
.Y(n_320)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_310),
.B(n_282),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_279),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_311),
.B(n_315),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_236),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_312),
.B(n_232),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_287),
.B(n_221),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_303),
.B(n_297),
.C(n_286),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_317),
.B(n_322),
.C(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_319),
.Y(n_339)
);

NOR2x1_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_291),
.Y(n_321)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_321),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_302),
.B(n_292),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_323),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_301),
.A2(n_284),
.B1(n_257),
.B2(n_221),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_324),
.A2(n_318),
.B1(n_314),
.B2(n_325),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_303),
.B(n_285),
.C(n_256),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_302),
.B(n_278),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_327),
.B(n_328),
.C(n_312),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_281),
.C(n_267),
.Y(n_328)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_329),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_330),
.A2(n_308),
.B1(n_306),
.B2(n_301),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_332),
.B(n_333),
.Y(n_345)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_320),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_331),
.A2(n_305),
.B1(n_309),
.B2(n_313),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_335),
.A2(n_340),
.B1(n_244),
.B2(n_232),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_343),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_326),
.A2(n_311),
.B1(n_261),
.B2(n_307),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_320),
.B(n_281),
.Y(n_341)
);

OAI21x1_ASAP7_75t_L g348 ( 
.A1(n_341),
.A2(n_321),
.B(n_244),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_334),
.B(n_327),
.C(n_317),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_344),
.B(n_347),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_342),
.B(n_322),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_349),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_337),
.B(n_328),
.C(n_300),
.Y(n_347)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_348),
.Y(n_353)
);

OAI21xp5_ASAP7_75t_SL g349 ( 
.A1(n_341),
.A2(n_329),
.B(n_255),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_350),
.B(n_338),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g352 ( 
.A(n_351),
.B(n_340),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_352),
.B(n_355),
.Y(n_360)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_345),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_356),
.B(n_350),
.Y(n_358)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_358),
.Y(n_362)
);

AOI322xp5_ASAP7_75t_L g359 ( 
.A1(n_353),
.A2(n_335),
.A3(n_339),
.B1(n_332),
.B2(n_354),
.C1(n_352),
.C2(n_346),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_361),
.C(n_356),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_357),
.B(n_339),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_SL g363 ( 
.A1(n_360),
.A2(n_337),
.B(n_343),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_363),
.B(n_364),
.Y(n_365)
);

AOI321xp33_ASAP7_75t_SL g366 ( 
.A1(n_362),
.A2(n_244),
.A3(n_274),
.B1(n_243),
.B2(n_197),
.C(n_191),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_274),
.B(n_191),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_243),
.C(n_244),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_368),
.A2(n_365),
.B(n_212),
.Y(n_369)
);

BUFx24_ASAP7_75t_SL g370 ( 
.A(n_369),
.Y(n_370)
);


endmodule