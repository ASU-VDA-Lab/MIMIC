module real_aes_8816_n_270 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_270);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_270;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_673;
wire n_386;
wire n_792;
wire n_518;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_857;
wire n_461;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_660;
wire n_814;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_626;
wire n_400;
wire n_539;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_352;
wire n_824;
wire n_875;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_748;
wire n_781;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_296;
wire n_702;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_720;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_481;
wire n_691;
wire n_498;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_290;
wire n_365;
wire n_637;
wire n_526;
wire n_692;
wire n_544;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_679;
wire n_520;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_721;
wire n_446;
wire n_681;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_639;
wire n_587;
wire n_546;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_687;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_SL g843 ( .A1(n_0), .A2(n_166), .B1(n_594), .B2(n_844), .Y(n_843) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_1), .A2(n_45), .B1(n_362), .B2(n_364), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_2), .A2(n_256), .B1(n_665), .B2(n_833), .Y(n_832) );
AOI22xp33_ASAP7_75t_SL g716 ( .A1(n_3), .A2(n_200), .B1(n_511), .B2(n_717), .Y(n_716) );
CKINVDCx20_ASAP7_75t_R g876 ( .A(n_4), .Y(n_876) );
CKINVDCx20_ASAP7_75t_R g288 ( .A(n_5), .Y(n_288) );
AOI22xp33_ASAP7_75t_SL g354 ( .A1(n_6), .A2(n_263), .B1(n_355), .B2(n_358), .Y(n_354) );
AOI222xp33_ASAP7_75t_L g500 ( .A1(n_7), .A2(n_31), .B1(n_120), .B2(n_328), .C1(n_405), .C2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_SL g570 ( .A1(n_8), .A2(n_35), .B1(n_512), .B2(n_571), .Y(n_570) );
CKINVDCx20_ASAP7_75t_R g770 ( .A(n_9), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g609 ( .A1(n_10), .A2(n_129), .B1(n_375), .B2(n_590), .Y(n_609) );
AOI22xp33_ASAP7_75t_L g744 ( .A1(n_11), .A2(n_205), .B1(n_745), .B2(n_747), .Y(n_744) );
CKINVDCx20_ASAP7_75t_R g488 ( .A(n_12), .Y(n_488) );
AOI22xp33_ASAP7_75t_SL g865 ( .A1(n_13), .A2(n_60), .B1(n_558), .B2(n_866), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_14), .A2(n_218), .B1(n_346), .B2(n_592), .Y(n_591) );
CKINVDCx20_ASAP7_75t_R g676 ( .A(n_15), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g304 ( .A(n_16), .Y(n_304) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_17), .A2(n_142), .B1(n_411), .B2(n_451), .Y(n_450) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_18), .Y(n_614) );
AOI221xp5_ASAP7_75t_L g489 ( .A1(n_19), .A2(n_44), .B1(n_490), .B2(n_492), .C(n_493), .Y(n_489) );
AOI221xp5_ASAP7_75t_L g471 ( .A1(n_20), .A2(n_214), .B1(n_472), .B2(n_474), .C(n_475), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_21), .B(n_633), .Y(n_632) );
CKINVDCx20_ASAP7_75t_R g674 ( .A(n_22), .Y(n_674) );
CKINVDCx20_ASAP7_75t_R g680 ( .A(n_23), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_24), .A2(n_204), .B1(n_341), .B2(n_684), .Y(n_683) );
CKINVDCx20_ASAP7_75t_R g774 ( .A(n_25), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_26), .A2(n_264), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g374 ( .A1(n_27), .A2(n_48), .B1(n_375), .B2(n_377), .Y(n_374) );
AO22x2_ASAP7_75t_L g293 ( .A1(n_28), .A2(n_87), .B1(n_294), .B2(n_295), .Y(n_293) );
INVx1_ASAP7_75t_L g824 ( .A(n_28), .Y(n_824) );
CKINVDCx20_ASAP7_75t_R g595 ( .A(n_29), .Y(n_595) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_30), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_32), .A2(n_234), .B1(n_362), .B2(n_364), .Y(n_580) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_33), .A2(n_73), .B1(n_482), .B2(n_485), .C(n_486), .Y(n_481) );
CKINVDCx20_ASAP7_75t_R g401 ( .A(n_34), .Y(n_401) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_36), .A2(n_188), .B1(n_385), .B2(n_515), .Y(n_514) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_37), .A2(n_149), .B1(n_743), .B2(n_779), .Y(n_778) );
AOI22xp33_ASAP7_75t_L g806 ( .A1(n_38), .A2(n_131), .B1(n_382), .B2(n_807), .Y(n_806) );
AOI22xp33_ASAP7_75t_SL g563 ( .A1(n_39), .A2(n_190), .B1(n_564), .B2(n_565), .Y(n_563) );
CKINVDCx20_ASAP7_75t_R g582 ( .A(n_40), .Y(n_582) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_41), .Y(n_785) );
AOI22xp33_ASAP7_75t_SL g863 ( .A1(n_42), .A2(n_182), .B1(n_706), .B2(n_864), .Y(n_863) );
CKINVDCx20_ASAP7_75t_R g877 ( .A(n_43), .Y(n_877) );
AO22x2_ASAP7_75t_L g297 ( .A1(n_46), .A2(n_89), .B1(n_294), .B2(n_298), .Y(n_297) );
INVx1_ASAP7_75t_L g825 ( .A(n_46), .Y(n_825) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_47), .A2(n_97), .B1(n_362), .B2(n_568), .Y(n_567) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_49), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_50), .A2(n_246), .B1(n_568), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g659 ( .A1(n_51), .A2(n_191), .B1(n_341), .B2(n_346), .Y(n_659) );
CKINVDCx20_ASAP7_75t_R g767 ( .A(n_52), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_53), .B(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g510 ( .A1(n_54), .A2(n_235), .B1(n_511), .B2(n_512), .Y(n_510) );
AOI22xp5_ASAP7_75t_L g338 ( .A1(n_55), .A2(n_84), .B1(n_339), .B2(n_341), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_56), .A2(n_90), .B1(n_395), .B2(n_396), .Y(n_394) );
CKINVDCx20_ASAP7_75t_R g772 ( .A(n_57), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_58), .A2(n_109), .B1(n_376), .B2(n_803), .Y(n_802) );
AOI222xp33_ASAP7_75t_L g845 ( .A1(n_59), .A2(n_147), .B1(n_155), .B2(n_311), .C1(n_411), .C2(n_650), .Y(n_845) );
AOI22xp33_ASAP7_75t_SL g869 ( .A1(n_61), .A2(n_68), .B1(n_719), .B2(n_870), .Y(n_869) );
CKINVDCx20_ASAP7_75t_R g626 ( .A(n_62), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_63), .A2(n_226), .B1(n_536), .B2(n_594), .Y(n_793) );
AOI22xp33_ASAP7_75t_SL g805 ( .A1(n_64), .A2(n_229), .B1(n_355), .B2(n_358), .Y(n_805) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_65), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g333 ( .A(n_66), .Y(n_333) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_67), .A2(n_85), .B1(n_536), .B2(n_736), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_69), .Y(n_625) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_70), .Y(n_648) );
AOI22xp33_ASAP7_75t_SL g718 ( .A1(n_71), .A2(n_127), .B1(n_719), .B2(n_720), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g437 ( .A(n_72), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_74), .B(n_535), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_75), .A2(n_93), .B1(n_355), .B2(n_519), .Y(n_518) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_76), .A2(n_154), .B1(n_163), .B2(n_405), .C1(n_501), .C2(n_594), .Y(n_593) );
CKINVDCx20_ASAP7_75t_R g635 ( .A(n_77), .Y(n_635) );
AOI22xp33_ASAP7_75t_SL g871 ( .A1(n_78), .A2(n_105), .B1(n_592), .B2(n_872), .Y(n_871) );
AOI22xp33_ASAP7_75t_SL g703 ( .A1(n_79), .A2(n_222), .B1(n_536), .B2(n_650), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g777 ( .A1(n_80), .A2(n_86), .B1(n_341), .B2(n_750), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g345 ( .A1(n_81), .A2(n_186), .B1(n_346), .B2(n_349), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_82), .A2(n_145), .B1(n_388), .B2(n_391), .Y(n_387) );
AOI22xp33_ASAP7_75t_SL g707 ( .A1(n_83), .A2(n_136), .B1(n_491), .B2(n_708), .Y(n_707) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_88), .Y(n_739) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_91), .A2(n_470), .B1(n_503), .B2(n_504), .Y(n_469) );
INVx1_ASAP7_75t_L g503 ( .A(n_91), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_92), .A2(n_254), .B1(n_408), .B2(n_561), .Y(n_560) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_94), .Y(n_764) );
INVx1_ASAP7_75t_L g278 ( .A(n_95), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_96), .A2(n_189), .B1(n_432), .B2(n_434), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g781 ( .A1(n_98), .A2(n_250), .B1(n_564), .B2(n_782), .Y(n_781) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_99), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g574 ( .A(n_100), .Y(n_574) );
AOI22xp5_ASAP7_75t_L g605 ( .A1(n_101), .A2(n_606), .B1(n_638), .B2(n_639), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g638 ( .A(n_101), .Y(n_638) );
INVx1_ASAP7_75t_L g274 ( .A(n_102), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_103), .A2(n_170), .B1(n_341), .B2(n_590), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g837 ( .A1(n_104), .A2(n_236), .B1(n_429), .B2(n_838), .Y(n_837) );
CKINVDCx20_ASAP7_75t_R g879 ( .A(n_106), .Y(n_879) );
CKINVDCx20_ASAP7_75t_R g527 ( .A(n_107), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_108), .A2(n_130), .B1(n_317), .B2(n_561), .Y(n_677) );
CKINVDCx20_ASAP7_75t_R g441 ( .A(n_110), .Y(n_441) );
AOI22xp5_ASAP7_75t_L g316 ( .A1(n_111), .A2(n_259), .B1(n_317), .B2(n_321), .Y(n_316) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_112), .A2(n_187), .B1(n_429), .B2(n_430), .Y(n_428) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_113), .A2(n_237), .B1(n_463), .B2(n_466), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g525 ( .A(n_114), .Y(n_525) );
AOI211xp5_ASAP7_75t_L g873 ( .A1(n_115), .A2(n_874), .B(n_875), .C(n_878), .Y(n_873) );
CKINVDCx20_ASAP7_75t_R g487 ( .A(n_116), .Y(n_487) );
AOI22xp33_ASAP7_75t_SL g656 ( .A1(n_117), .A2(n_119), .B1(n_321), .B2(n_587), .Y(n_656) );
OA22x2_ASAP7_75t_L g641 ( .A1(n_118), .A2(n_642), .B1(n_643), .B2(n_667), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_118), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_121), .B(n_492), .Y(n_796) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_122), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_123), .B(n_559), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_124), .A2(n_128), .B1(n_565), .B2(n_579), .Y(n_578) );
OA22x2_ASAP7_75t_L g668 ( .A1(n_125), .A2(n_669), .B1(n_670), .B2(n_691), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_125), .Y(n_669) );
CKINVDCx20_ASAP7_75t_R g406 ( .A(n_126), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_132), .A2(n_251), .B1(n_395), .B2(n_434), .Y(n_839) );
CKINVDCx20_ASAP7_75t_R g636 ( .A(n_133), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_134), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_135), .B(n_556), .Y(n_555) );
XNOR2x2_ASAP7_75t_L g424 ( .A(n_137), .B(n_425), .Y(n_424) );
AND2x2_ASAP7_75t_L g277 ( .A(n_138), .B(n_278), .Y(n_277) );
CKINVDCx20_ASAP7_75t_R g497 ( .A(n_139), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_140), .A2(n_169), .B1(n_432), .B2(n_522), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_141), .Y(n_442) );
CKINVDCx20_ASAP7_75t_R g621 ( .A(n_143), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g834 ( .A1(n_144), .A2(n_150), .B1(n_803), .B2(n_835), .Y(n_834) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_146), .B(n_653), .Y(n_652) );
CKINVDCx20_ASAP7_75t_R g416 ( .A(n_148), .Y(n_416) );
CKINVDCx20_ASAP7_75t_R g859 ( .A(n_151), .Y(n_859) );
AND2x6_ASAP7_75t_L g273 ( .A(n_152), .B(n_274), .Y(n_273) );
HB1xp67_ASAP7_75t_L g818 ( .A(n_152), .Y(n_818) );
AO22x2_ASAP7_75t_L g303 ( .A1(n_153), .A2(n_216), .B1(n_294), .B2(n_298), .Y(n_303) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_156), .A2(n_185), .B1(n_485), .B2(n_750), .Y(n_749) );
AOI22xp33_ASAP7_75t_SL g710 ( .A1(n_157), .A2(n_225), .B1(n_592), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g860 ( .A(n_158), .Y(n_860) );
AOI22xp33_ASAP7_75t_SL g454 ( .A1(n_159), .A2(n_230), .B1(n_455), .B2(n_459), .Y(n_454) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_160), .A2(n_248), .B1(n_346), .B2(n_689), .Y(n_688) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_161), .Y(n_792) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_162), .A2(n_260), .B1(n_396), .B2(n_714), .Y(n_713) );
AOI211xp5_ASAP7_75t_L g270 ( .A1(n_164), .A2(n_271), .B(n_279), .C(n_826), .Y(n_270) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_165), .A2(n_203), .B1(n_532), .B2(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g752 ( .A(n_167), .Y(n_752) );
AOI22xp33_ASAP7_75t_SL g705 ( .A1(n_168), .A2(n_223), .B1(n_322), .B2(n_706), .Y(n_705) );
AOI22xp33_ASAP7_75t_SL g666 ( .A1(n_171), .A2(n_255), .B1(n_349), .B2(n_363), .Y(n_666) );
CKINVDCx20_ASAP7_75t_R g728 ( .A(n_172), .Y(n_728) );
CKINVDCx20_ASAP7_75t_R g436 ( .A(n_173), .Y(n_436) );
AOI22xp33_ASAP7_75t_L g797 ( .A1(n_174), .A2(n_184), .B1(n_457), .B2(n_650), .Y(n_797) );
CKINVDCx20_ASAP7_75t_R g494 ( .A(n_175), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_176), .B(n_459), .Y(n_765) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_177), .A2(n_242), .B1(n_664), .B2(n_665), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_178), .A2(n_179), .B1(n_393), .B2(n_801), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g610 ( .A1(n_180), .A2(n_211), .B1(n_434), .B2(n_611), .Y(n_610) );
AO22x2_ASAP7_75t_L g301 ( .A1(n_181), .A2(n_239), .B1(n_294), .B2(n_295), .Y(n_301) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_183), .Y(n_738) );
AOI22xp33_ASAP7_75t_SL g660 ( .A1(n_192), .A2(n_219), .B1(n_433), .B2(n_661), .Y(n_660) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_193), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_194), .Y(n_479) );
AOI22xp33_ASAP7_75t_SL g572 ( .A1(n_195), .A2(n_231), .B1(n_430), .B2(n_573), .Y(n_572) );
CKINVDCx20_ASAP7_75t_R g530 ( .A(n_196), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g649 ( .A1(n_197), .A2(n_241), .B1(n_502), .B2(n_650), .Y(n_649) );
CKINVDCx20_ASAP7_75t_R g679 ( .A(n_198), .Y(n_679) );
CKINVDCx20_ASAP7_75t_R g631 ( .A(n_199), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g506 ( .A1(n_201), .A2(n_507), .B1(n_544), .B2(n_545), .Y(n_506) );
CKINVDCx20_ASAP7_75t_R g544 ( .A(n_201), .Y(n_544) );
CKINVDCx20_ASAP7_75t_R g619 ( .A(n_202), .Y(n_619) );
INVx1_ASAP7_75t_L g841 ( .A(n_206), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_207), .A2(n_247), .B1(n_573), .B2(n_743), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_208), .B(n_584), .Y(n_795) );
AOI22xp33_ASAP7_75t_SL g553 ( .A1(n_209), .A2(n_252), .B1(n_321), .B2(n_536), .Y(n_553) );
NAND2xp5_ASAP7_75t_SL g557 ( .A(n_210), .B(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_212), .B(n_411), .Y(n_410) );
XOR2xp5_ASAP7_75t_L g827 ( .A(n_213), .B(n_828), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g538 ( .A(n_215), .Y(n_538) );
NOR2xp33_ASAP7_75t_L g822 ( .A(n_216), .B(n_823), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g414 ( .A(n_217), .Y(n_414) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_220), .Y(n_673) );
OA22x2_ASAP7_75t_L g697 ( .A1(n_221), .A2(n_698), .B1(n_699), .B2(n_721), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_221), .Y(n_698) );
CKINVDCx20_ASAP7_75t_R g629 ( .A(n_224), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_227), .B(n_559), .Y(n_842) );
INVx1_ASAP7_75t_L g368 ( .A(n_228), .Y(n_368) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_232), .Y(n_808) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_233), .Y(n_476) );
INVxp67_ASAP7_75t_L g853 ( .A(n_238), .Y(n_853) );
XNOR2xp5_ASAP7_75t_L g855 ( .A(n_238), .B(n_856), .Y(n_855) );
INVx1_ASAP7_75t_L g821 ( .A(n_239), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g552 ( .A(n_240), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g690 ( .A1(n_243), .A2(n_249), .B1(n_362), .B2(n_592), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g751 ( .A1(n_244), .A2(n_258), .B1(n_341), .B2(n_686), .Y(n_751) );
CKINVDCx20_ASAP7_75t_R g399 ( .A(n_245), .Y(n_399) );
AOI22xp5_ASAP7_75t_L g370 ( .A1(n_253), .A2(n_371), .B1(n_421), .B2(n_422), .Y(n_370) );
INVx1_ASAP7_75t_L g421 ( .A(n_253), .Y(n_421) );
INVx1_ASAP7_75t_L g294 ( .A(n_257), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_257), .Y(n_296) );
CKINVDCx20_ASAP7_75t_R g729 ( .A(n_261), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g409 ( .A(n_262), .Y(n_409) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_265), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g381 ( .A1(n_266), .A2(n_269), .B1(n_382), .B2(n_384), .Y(n_381) );
CKINVDCx20_ASAP7_75t_R g326 ( .A(n_267), .Y(n_326) );
CKINVDCx20_ASAP7_75t_R g861 ( .A(n_268), .Y(n_861) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_275), .Y(n_272) );
HB1xp67_ASAP7_75t_L g817 ( .A(n_274), .Y(n_817) );
OAI21xp5_ASAP7_75t_L g851 ( .A1(n_275), .A2(n_816), .B(n_852), .Y(n_851) );
CKINVDCx20_ASAP7_75t_R g275 ( .A(n_276), .Y(n_275) );
INVxp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AOI221xp5_ASAP7_75t_L g279 ( .A1(n_280), .A2(n_602), .B1(n_811), .B2(n_812), .C(n_813), .Y(n_279) );
INVxp67_ASAP7_75t_L g811 ( .A(n_280), .Y(n_811) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_282), .B1(n_423), .B2(n_601), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI22xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_284), .B1(n_369), .B2(n_370), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
XNOR2xp5_ASAP7_75t_L g723 ( .A(n_284), .B(n_724), .Y(n_723) );
XOR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_368), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_286), .B(n_336), .Y(n_285) );
NOR3xp33_ASAP7_75t_L g286 ( .A(n_287), .B(n_309), .C(n_325), .Y(n_286) );
OAI22xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B1(n_304), .B2(n_305), .Y(n_287) );
OAI22xp5_ASAP7_75t_L g672 ( .A1(n_289), .A2(n_402), .B1(n_673), .B2(n_674), .Y(n_672) );
BUFx3_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_290), .Y(n_400) );
INVx2_ASAP7_75t_L g540 ( .A(n_290), .Y(n_540) );
OR2x2_ASAP7_75t_L g290 ( .A(n_291), .B(n_299), .Y(n_290) );
INVx2_ASAP7_75t_L g340 ( .A(n_291), .Y(n_340) );
OR2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_297), .Y(n_291) );
AND2x2_ASAP7_75t_L g308 ( .A(n_292), .B(n_297), .Y(n_308) );
AND2x2_ASAP7_75t_L g344 ( .A(n_292), .B(n_332), .Y(n_344) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g312 ( .A(n_293), .B(n_297), .Y(n_312) );
AND2x2_ASAP7_75t_L g320 ( .A(n_293), .B(n_303), .Y(n_320) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g298 ( .A(n_296), .Y(n_298) );
INVx2_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
INVx1_ASAP7_75t_L g367 ( .A(n_297), .Y(n_367) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
NAND2x1p5_ASAP7_75t_L g307 ( .A(n_300), .B(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g363 ( .A(n_300), .B(n_344), .Y(n_363) );
AND2x4_ASAP7_75t_L g465 ( .A(n_300), .B(n_340), .Y(n_465) );
AND2x6_ASAP7_75t_L g467 ( .A(n_300), .B(n_308), .Y(n_467) );
AND2x2_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g314 ( .A(n_301), .Y(n_314) );
INVx1_ASAP7_75t_L g319 ( .A(n_301), .Y(n_319) );
INVx1_ASAP7_75t_L g324 ( .A(n_301), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_301), .B(n_303), .Y(n_352) );
AND2x2_ASAP7_75t_L g313 ( .A(n_302), .B(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g343 ( .A(n_303), .B(n_324), .Y(n_343) );
OA211x2_ASAP7_75t_L g840 ( .A1(n_305), .A2(n_841), .B(n_842), .C(n_843), .Y(n_840) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g402 ( .A(n_306), .Y(n_402) );
INVx2_ASAP7_75t_L g637 ( .A(n_306), .Y(n_637) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g543 ( .A(n_307), .Y(n_543) );
AND2x4_ASAP7_75t_L g357 ( .A(n_308), .B(n_313), .Y(n_357) );
AND2x2_ASAP7_75t_L g360 ( .A(n_308), .B(n_343), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_308), .B(n_343), .Y(n_478) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_315), .B(n_316), .Y(n_309) );
INVx4_ASAP7_75t_L g405 ( .A(n_310), .Y(n_405) );
BUFx2_ASAP7_75t_L g734 ( .A(n_310), .Y(n_734) );
INVx4_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g448 ( .A(n_311), .Y(n_448) );
INVx2_ASAP7_75t_L g529 ( .A(n_311), .Y(n_529) );
BUFx3_ASAP7_75t_L g647 ( .A(n_311), .Y(n_647) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_311), .Y(n_684) );
AND2x6_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
AND2x4_ASAP7_75t_L g322 ( .A(n_312), .B(n_323), .Y(n_322) );
INVx1_ASAP7_75t_L g419 ( .A(n_312), .Y(n_419) );
AND2x6_ASAP7_75t_L g339 ( .A(n_313), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g348 ( .A(n_313), .B(n_344), .Y(n_348) );
BUFx6f_ASAP7_75t_L g412 ( .A(n_317), .Y(n_412) );
BUFx12f_ASAP7_75t_L g502 ( .A(n_317), .Y(n_502) );
BUFx6f_ASAP7_75t_L g536 ( .A(n_317), .Y(n_536) );
AND2x4_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g331 ( .A(n_319), .B(n_332), .Y(n_331) );
AND2x4_ASAP7_75t_L g330 ( .A(n_320), .B(n_331), .Y(n_330) );
NAND2x1p5_ASAP7_75t_L g334 ( .A(n_320), .B(n_335), .Y(n_334) );
AND2x4_ASAP7_75t_L g457 ( .A(n_320), .B(n_458), .Y(n_457) );
BUFx2_ASAP7_75t_SL g321 ( .A(n_322), .Y(n_321) );
BUFx6f_ASAP7_75t_L g461 ( .A(n_322), .Y(n_461) );
BUFx2_ASAP7_75t_SL g594 ( .A(n_322), .Y(n_594) );
BUFx3_ASAP7_75t_L g864 ( .A(n_322), .Y(n_864) );
INVx1_ASAP7_75t_L g420 ( .A(n_323), .Y(n_420) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_327), .B1(n_333), .B2(n_334), .Y(n_325) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_SL g630 ( .A(n_328), .Y(n_630) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g773 ( .A(n_329), .Y(n_773) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_330), .Y(n_408) );
BUFx2_ASAP7_75t_L g532 ( .A(n_330), .Y(n_532) );
BUFx6f_ASAP7_75t_L g586 ( .A(n_330), .Y(n_586) );
BUFx4f_ASAP7_75t_SL g650 ( .A(n_330), .Y(n_650) );
INVx1_ASAP7_75t_L g335 ( .A(n_332), .Y(n_335) );
BUFx3_ASAP7_75t_L g415 ( .A(n_334), .Y(n_415) );
INVx4_ASAP7_75t_L g496 ( .A(n_334), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g624 ( .A1(n_334), .A2(n_625), .B1(n_626), .B2(n_627), .Y(n_624) );
AND2x2_ASAP7_75t_L g807 ( .A(n_335), .B(n_351), .Y(n_807) );
NOR2xp33_ASAP7_75t_L g336 ( .A(n_337), .B(n_353), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_338), .B(n_345), .Y(n_337) );
INVx11_ASAP7_75t_L g380 ( .A(n_339), .Y(n_380) );
INVx11_ASAP7_75t_L g513 ( .A(n_339), .Y(n_513) );
INVx1_ASAP7_75t_L g520 ( .A(n_341), .Y(n_520) );
BUFx2_ASAP7_75t_L g870 ( .A(n_341), .Y(n_870) );
BUFx3_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
BUFx3_ASAP7_75t_L g393 ( .A(n_342), .Y(n_393) );
BUFx3_ASAP7_75t_L g571 ( .A(n_342), .Y(n_571) );
BUFx3_ASAP7_75t_L g838 ( .A(n_342), .Y(n_838) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_343), .B(n_344), .Y(n_445) );
AND2x4_ASAP7_75t_L g350 ( .A(n_344), .B(n_351), .Y(n_350) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_L g779 ( .A(n_347), .Y(n_779) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_348), .Y(n_376) );
BUFx2_ASAP7_75t_SL g573 ( .A(n_348), .Y(n_573) );
BUFx2_ASAP7_75t_SL g874 ( .A(n_348), .Y(n_874) );
BUFx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
BUFx3_ASAP7_75t_L g385 ( .A(n_350), .Y(n_385) );
BUFx2_ASAP7_75t_SL g430 ( .A(n_350), .Y(n_430) );
BUFx3_ASAP7_75t_L g474 ( .A(n_350), .Y(n_474) );
BUFx3_ASAP7_75t_L g592 ( .A(n_350), .Y(n_592) );
BUFx2_ASAP7_75t_SL g743 ( .A(n_350), .Y(n_743) );
BUFx3_ASAP7_75t_L g803 ( .A(n_350), .Y(n_803) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x6_ASAP7_75t_L g366 ( .A(n_352), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_361), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g440 ( .A1(n_356), .A2(n_441), .B1(n_442), .B2(n_443), .Y(n_440) );
INVx2_ASAP7_75t_L g564 ( .A(n_356), .Y(n_564) );
INVx2_ASAP7_75t_L g579 ( .A(n_356), .Y(n_579) );
INVx3_ASAP7_75t_L g665 ( .A(n_356), .Y(n_665) );
INVx6_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx3_ASAP7_75t_L g390 ( .A(n_357), .Y(n_390) );
BUFx3_ASAP7_75t_L g686 ( .A(n_357), .Y(n_686) );
BUFx3_ASAP7_75t_L g719 ( .A(n_357), .Y(n_719) );
INVx3_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g395 ( .A(n_359), .Y(n_395) );
INVx4_ASAP7_75t_L g433 ( .A(n_359), .Y(n_433) );
BUFx3_ASAP7_75t_L g566 ( .A(n_359), .Y(n_566) );
INVx1_ASAP7_75t_L g612 ( .A(n_359), .Y(n_612) );
INVx5_ASAP7_75t_L g689 ( .A(n_359), .Y(n_689) );
INVx8_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g872 ( .A(n_362), .Y(n_872) );
BUFx3_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
INVx2_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_363), .Y(n_439) );
BUFx3_ASAP7_75t_L g516 ( .A(n_363), .Y(n_516) );
BUFx3_ASAP7_75t_L g784 ( .A(n_363), .Y(n_784) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
BUFx2_ASAP7_75t_L g396 ( .A(n_365), .Y(n_396) );
BUFx2_ASAP7_75t_L g434 ( .A(n_365), .Y(n_434) );
BUFx4f_ASAP7_75t_SL g522 ( .A(n_365), .Y(n_522) );
BUFx2_ASAP7_75t_L g568 ( .A(n_365), .Y(n_568) );
INVx6_ASAP7_75t_SL g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g661 ( .A(n_366), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_366), .A2(n_418), .B1(n_679), .B2(n_680), .Y(n_678) );
INVx1_ASAP7_75t_L g747 ( .A(n_366), .Y(n_747) );
INVx1_ASAP7_75t_L g458 ( .A(n_367), .Y(n_458) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx2_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_372), .B(n_397), .Y(n_371) );
NOR2xp33_ASAP7_75t_L g372 ( .A(n_373), .B(n_386), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_381), .Y(n_373) );
BUFx3_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
INVx3_ASAP7_75t_L g473 ( .A(n_376), .Y(n_473) );
BUFx3_ASAP7_75t_L g511 ( .A(n_376), .Y(n_511) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_378), .A2(n_436), .B1(n_437), .B2(n_438), .Y(n_435) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx5_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_SL g484 ( .A(n_380), .Y(n_484) );
INVx1_ASAP7_75t_L g590 ( .A(n_380), .Y(n_590) );
HB1xp67_ASAP7_75t_L g712 ( .A(n_380), .Y(n_712) );
INVx4_ASAP7_75t_L g801 ( .A(n_380), .Y(n_801) );
INVx2_ASAP7_75t_L g833 ( .A(n_380), .Y(n_833) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
BUFx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_387), .B(n_394), .Y(n_386) );
INVx2_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g486 ( .A1(n_389), .A2(n_443), .B1(n_487), .B2(n_488), .Y(n_486) );
INVx3_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
HB1xp67_ASAP7_75t_L g714 ( .A(n_395), .Y(n_714) );
NOR3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_403), .C(n_413), .Y(n_397) );
OAI22xp5_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_401), .B2(n_402), .Y(n_398) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_400), .A2(n_635), .B1(n_636), .B2(n_637), .Y(n_634) );
INVx1_ASAP7_75t_L g769 ( .A(n_400), .Y(n_769) );
OA211x2_ASAP7_75t_L g581 ( .A1(n_402), .A2(n_582), .B(n_583), .C(n_585), .Y(n_581) );
OAI221xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_406), .B1(n_407), .B2(n_409), .C(n_410), .Y(n_403) );
OAI221xp5_ASAP7_75t_L g628 ( .A1(n_404), .A2(n_629), .B1(n_630), .B2(n_631), .C(n_632), .Y(n_628) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx4_ASAP7_75t_L g452 ( .A(n_408), .Y(n_452) );
BUFx2_ASAP7_75t_L g736 ( .A(n_408), .Y(n_736) );
BUFx4f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g763 ( .A(n_412), .Y(n_763) );
OAI22xp5_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_415), .B1(n_416), .B2(n_417), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_415), .A2(n_772), .B1(n_773), .B2(n_774), .Y(n_771) );
BUFx2_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_418), .Y(n_499) );
OR2x6_ASAP7_75t_L g418 ( .A(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_L g601 ( .A(n_423), .Y(n_601) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_468), .B1(n_599), .B2(n_600), .Y(n_423) );
INVx2_ASAP7_75t_L g600 ( .A(n_424), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g425 ( .A(n_426), .B(n_446), .Y(n_425) );
NOR3xp33_ASAP7_75t_L g426 ( .A(n_427), .B(n_435), .C(n_440), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_428), .B(n_431), .Y(n_427) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g746 ( .A(n_433), .Y(n_746) );
INVx1_ASAP7_75t_L g480 ( .A(n_434), .Y(n_480) );
INVx4_ASAP7_75t_L g485 ( .A(n_438), .Y(n_485) );
INVx3_ASAP7_75t_L g835 ( .A(n_438), .Y(n_835) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx1_ASAP7_75t_L g617 ( .A(n_444), .Y(n_617) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
NOR2xp33_ASAP7_75t_L g446 ( .A(n_447), .B(n_453), .Y(n_446) );
OAI21xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B(n_450), .Y(n_447) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_448), .A2(n_702), .B(n_703), .Y(n_701) );
INVx3_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_454), .B(n_462), .Y(n_453) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g844 ( .A(n_456), .Y(n_844) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
BUFx2_ASAP7_75t_L g561 ( .A(n_457), .Y(n_561) );
BUFx3_ASAP7_75t_L g587 ( .A(n_457), .Y(n_587) );
BUFx2_ASAP7_75t_L g706 ( .A(n_457), .Y(n_706) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g491 ( .A(n_464), .Y(n_491) );
INVx5_ASAP7_75t_L g559 ( .A(n_464), .Y(n_559) );
INVx2_ASAP7_75t_L g584 ( .A(n_464), .Y(n_584) );
INVx4_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
BUFx4f_ASAP7_75t_L g492 ( .A(n_467), .Y(n_492) );
BUFx2_ASAP7_75t_L g556 ( .A(n_467), .Y(n_556) );
INVx1_ASAP7_75t_SL g654 ( .A(n_467), .Y(n_654) );
INVx1_ASAP7_75t_L g599 ( .A(n_468), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_469), .A2(n_505), .B1(n_597), .B2(n_598), .Y(n_468) );
INVx1_ASAP7_75t_L g597 ( .A(n_469), .Y(n_597) );
INVx1_ASAP7_75t_L g504 ( .A(n_470), .Y(n_504) );
AND4x1_ASAP7_75t_L g470 ( .A(n_471), .B(n_481), .C(n_489), .D(n_500), .Y(n_470) );
INVx2_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B1(n_479), .B2(n_480), .Y(n_475) );
OAI22xp5_ASAP7_75t_SL g875 ( .A1(n_477), .A2(n_480), .B1(n_876), .B2(n_877), .Y(n_875) );
BUFx2_ASAP7_75t_R g477 ( .A(n_478), .Y(n_477) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx1_ASAP7_75t_L g867 ( .A(n_492), .Y(n_867) );
OAI22xp5_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_495), .B1(n_497), .B2(n_498), .Y(n_493) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx3_ASAP7_75t_SL g526 ( .A(n_496), .Y(n_526) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_498), .A2(n_525), .B1(n_526), .B2(n_527), .Y(n_524) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_L g627 ( .A(n_499), .Y(n_627) );
BUFx4f_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g598 ( .A(n_505), .Y(n_598) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_546), .B1(n_547), .B2(n_596), .Y(n_505) );
INVx1_ASAP7_75t_L g596 ( .A(n_506), .Y(n_596) );
INVx1_ASAP7_75t_SL g545 ( .A(n_507), .Y(n_545) );
AND2x2_ASAP7_75t_SL g507 ( .A(n_508), .B(n_523), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_514), .Y(n_509) );
INVx1_ASAP7_75t_L g880 ( .A(n_512), .Y(n_880) );
INVx4_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx4_ASAP7_75t_L g664 ( .A(n_513), .Y(n_664) );
OAI21xp33_ASAP7_75t_SL g675 ( .A1(n_513), .A2(n_676), .B(n_677), .Y(n_675) );
INVx2_ASAP7_75t_SL g750 ( .A(n_513), .Y(n_750) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g620 ( .A(n_516), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_521), .Y(n_517) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
NOR3xp33_ASAP7_75t_SL g523 ( .A(n_524), .B(n_528), .C(n_537), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_526), .A2(n_627), .B1(n_738), .B2(n_739), .Y(n_737) );
OAI221xp5_ASAP7_75t_SL g528 ( .A1(n_529), .A2(n_530), .B1(n_531), .B2(n_533), .C(n_534), .Y(n_528) );
OAI21xp5_ASAP7_75t_SL g551 ( .A1(n_529), .A2(n_552), .B(n_553), .Y(n_551) );
OAI222xp33_ASAP7_75t_L g858 ( .A1(n_529), .A2(n_630), .B1(n_763), .B2(n_859), .C1(n_860), .C2(n_861), .Y(n_858) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx3_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
BUFx2_ASAP7_75t_L g633 ( .A(n_536), .Y(n_633) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_538), .A2(n_539), .B1(n_541), .B2(n_542), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_539), .A2(n_728), .B1(n_729), .B2(n_730), .Y(n_727) );
INVx1_ASAP7_75t_SL g539 ( .A(n_540), .Y(n_539) );
BUFx3_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g731 ( .A(n_543), .Y(n_731) );
INVx2_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
XNOR2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_575), .Y(n_547) );
XOR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_574), .Y(n_548) );
NAND3x1_ASAP7_75t_L g549 ( .A(n_550), .B(n_562), .C(n_569), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_554), .Y(n_550) );
NAND3xp33_ASAP7_75t_L g554 ( .A(n_555), .B(n_557), .C(n_560), .Y(n_554) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_567), .Y(n_562) );
INVx2_ASAP7_75t_L g615 ( .A(n_564), .Y(n_615) );
INVx3_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
BUFx3_ASAP7_75t_L g720 ( .A(n_571), .Y(n_720) );
XOR2x2_ASAP7_75t_L g575 ( .A(n_576), .B(n_595), .Y(n_575) );
NAND4xp75_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .C(n_588), .D(n_593), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
AND2x2_ASAP7_75t_L g588 ( .A(n_589), .B(n_591), .Y(n_588) );
INVxp67_ASAP7_75t_L g622 ( .A(n_592), .Y(n_622) );
INVx1_ASAP7_75t_L g812 ( .A(n_602), .Y(n_812) );
AOI22xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B1(n_694), .B2(n_810), .Y(n_602) );
INVx2_ASAP7_75t_SL g603 ( .A(n_604), .Y(n_603) );
OA22x2_ASAP7_75t_L g604 ( .A1(n_605), .A2(n_640), .B1(n_692), .B2(n_693), .Y(n_604) );
INVx1_ASAP7_75t_L g692 ( .A(n_605), .Y(n_692) );
INVx1_ASAP7_75t_L g639 ( .A(n_606), .Y(n_639) );
AND2x2_ASAP7_75t_SL g606 ( .A(n_607), .B(n_623), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g607 ( .A(n_608), .B(n_613), .C(n_618), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_615), .B1(n_616), .B2(n_617), .Y(n_613) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_620), .B1(n_621), .B2(n_622), .Y(n_618) );
INVx1_ASAP7_75t_L g717 ( .A(n_620), .Y(n_717) );
NOR3xp33_ASAP7_75t_SL g623 ( .A(n_624), .B(n_628), .C(n_634), .Y(n_623) );
INVx1_ASAP7_75t_L g693 ( .A(n_640), .Y(n_693) );
XOR2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_668), .Y(n_640) );
INVx1_ASAP7_75t_L g667 ( .A(n_643), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_644), .B(n_657), .Y(n_643) );
NOR2xp67_ASAP7_75t_L g644 ( .A(n_645), .B(n_651), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_646), .A2(n_648), .B(n_649), .Y(n_645) );
INVx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_655), .C(n_656), .Y(n_651) );
INVx1_ASAP7_75t_SL g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_SL g708 ( .A(n_654), .Y(n_708) );
NOR2x1_ASAP7_75t_L g657 ( .A(n_658), .B(n_662), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_663), .B(n_666), .Y(n_662) );
INVx2_ASAP7_75t_L g691 ( .A(n_670), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_671), .B(n_681), .Y(n_670) );
NOR3xp33_ASAP7_75t_L g671 ( .A(n_672), .B(n_675), .C(n_678), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_687), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx2_ASAP7_75t_L g761 ( .A(n_684), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_689), .Y(n_782) );
INVx1_ASAP7_75t_L g810 ( .A(n_694), .Y(n_810) );
AOI22xp5_ASAP7_75t_SL g694 ( .A1(n_695), .A2(n_753), .B1(n_754), .B2(n_809), .Y(n_694) );
INVx1_ASAP7_75t_L g809 ( .A(n_695), .Y(n_809) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_696), .A2(n_697), .B1(n_722), .B2(n_723), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g721 ( .A(n_699), .Y(n_721) );
NAND3x1_ASAP7_75t_L g699 ( .A(n_700), .B(n_709), .C(n_715), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_704), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_707), .Y(n_704) );
AND2x2_ASAP7_75t_L g709 ( .A(n_710), .B(n_713), .Y(n_709) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
AND2x2_ASAP7_75t_L g715 ( .A(n_716), .B(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
XOR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_752), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_726), .B(n_740), .Y(n_725) );
NOR3xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_732), .C(n_737), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_730), .A2(n_767), .B1(n_768), .B2(n_770), .Y(n_766) );
INVx2_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
OAI21xp33_ASAP7_75t_L g732 ( .A1(n_733), .A2(n_734), .B(n_735), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_748), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_742), .B(n_744), .Y(n_741) );
INVx3_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
XOR2xp5_ASAP7_75t_L g754 ( .A(n_755), .B(n_786), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
XOR2x2_ASAP7_75t_L g757 ( .A(n_758), .B(n_785), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_775), .Y(n_758) );
NOR3xp33_ASAP7_75t_L g759 ( .A(n_760), .B(n_766), .C(n_771), .Y(n_759) );
OAI221xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .C(n_765), .Y(n_760) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_761), .A2(n_792), .B(n_793), .Y(n_791) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_776), .B(n_780), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_783), .Y(n_780) );
INVx2_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
XOR2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_808), .Y(n_788) );
NAND2xp5_ASAP7_75t_SL g789 ( .A(n_790), .B(n_798), .Y(n_789) );
NOR2xp33_ASAP7_75t_L g790 ( .A(n_791), .B(n_794), .Y(n_790) );
NAND3xp33_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .C(n_797), .Y(n_794) );
NOR2x1_ASAP7_75t_L g798 ( .A(n_799), .B(n_804), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_802), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_805), .B(n_806), .Y(n_804) );
INVx1_ASAP7_75t_SL g813 ( .A(n_814), .Y(n_813) );
NOR2x1_ASAP7_75t_L g814 ( .A(n_815), .B(n_819), .Y(n_814) );
OR2x2_ASAP7_75t_SL g881 ( .A(n_815), .B(n_820), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_817), .Y(n_816) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_817), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_817), .B(n_849), .Y(n_852) );
CKINVDCx16_ASAP7_75t_R g849 ( .A(n_818), .Y(n_849) );
CKINVDCx20_ASAP7_75t_R g819 ( .A(n_820), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_821), .B(n_822), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_824), .B(n_825), .Y(n_823) );
OAI322xp33_ASAP7_75t_L g826 ( .A1(n_827), .A2(n_846), .A3(n_847), .B1(n_850), .B2(n_853), .C1(n_854), .C2(n_881), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g828 ( .A(n_829), .Y(n_828) );
HB1xp67_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
NAND4xp75_ASAP7_75t_L g830 ( .A(n_831), .B(n_836), .C(n_840), .D(n_845), .Y(n_830) );
AND2x2_ASAP7_75t_L g831 ( .A(n_832), .B(n_834), .Y(n_831) );
AND2x2_ASAP7_75t_L g836 ( .A(n_837), .B(n_839), .Y(n_836) );
HB1xp67_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
CKINVDCx20_ASAP7_75t_R g850 ( .A(n_851), .Y(n_850) );
HB1xp67_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NAND3x1_ASAP7_75t_L g856 ( .A(n_857), .B(n_868), .C(n_873), .Y(n_856) );
NOR2xp33_ASAP7_75t_L g857 ( .A(n_858), .B(n_862), .Y(n_857) );
NAND2xp5_ASAP7_75t_L g862 ( .A(n_863), .B(n_865), .Y(n_862) );
INVx1_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
AND2x2_ASAP7_75t_L g868 ( .A(n_869), .B(n_871), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_879), .B(n_880), .Y(n_878) );
endmodule