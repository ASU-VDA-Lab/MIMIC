module fake_jpeg_645_n_216 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_216);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_154;
wire n_127;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_25),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_28),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_15),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_1),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_27),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_34),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g63 ( 
.A(n_21),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_11),
.Y(n_64)
);

BUFx4f_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_13),
.Y(n_66)
);

BUFx16f_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_49),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_5),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_1),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_14),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_79),
.Y(n_97)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_71),
.Y(n_82)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_83),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_84),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_76),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g87 ( 
.A(n_56),
.Y(n_87)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_56),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_87),
.B(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_88),
.B(n_95),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_78),
.B1(n_73),
.B2(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_90),
.A2(n_92),
.B1(n_78),
.B2(n_67),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_66),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_100),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_82),
.A2(n_78),
.B1(n_73),
.B2(n_64),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_68),
.Y(n_95)
);

NAND2x1_ASAP7_75t_SL g121 ( 
.A(n_99),
.B(n_54),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_96),
.Y(n_104)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_104),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_98),
.A2(n_62),
.B1(n_53),
.B2(n_60),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_61),
.B1(n_65),
.B2(n_69),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g107 ( 
.A(n_93),
.Y(n_107)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_107),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_77),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_88),
.B(n_74),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_95),
.B(n_55),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_119),
.Y(n_133)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_98),
.Y(n_111)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_111),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_57),
.B1(n_58),
.B2(n_59),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_99),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_113),
.B(n_2),
.Y(n_136)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_101),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_115),
.B(n_116),
.Y(n_126)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_93),
.A2(n_65),
.B1(n_75),
.B2(n_70),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_118),
.A2(n_65),
.B1(n_97),
.B2(n_54),
.Y(n_125)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_67),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_120),
.B(n_94),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g140 ( 
.A(n_121),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_131),
.B1(n_144),
.B2(n_3),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_125),
.A2(n_141),
.B1(n_6),
.B2(n_7),
.Y(n_150)
);

AOI21x1_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_8),
.B(n_9),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_0),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_130),
.B(n_24),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_105),
.A2(n_117),
.B1(n_120),
.B2(n_119),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_107),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_132),
.B(n_138),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_2),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g152 ( 
.A(n_135),
.B(n_142),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_136),
.Y(n_168)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_137),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_103),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_104),
.A2(n_94),
.B1(n_4),
.B2(n_5),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_107),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_147),
.B(n_150),
.Y(n_176)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_122),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_149),
.B(n_153),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_23),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_157),
.C(n_166),
.Y(n_187)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_124),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_133),
.B(n_7),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_156),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_160),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_126),
.B(n_127),
.C(n_131),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_29),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_144),
.B(n_8),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_137),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_162),
.A2(n_164),
.B(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_129),
.B(n_10),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_134),
.A2(n_12),
.B(n_13),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_164),
.A2(n_17),
.B(n_18),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_14),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_165),
.B(n_167),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_134),
.B(n_32),
.C(n_47),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_145),
.B(n_15),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_16),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_16),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_170),
.B(n_31),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_172),
.B(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_125),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_180),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_151),
.B(n_19),
.C(n_20),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_146),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_185),
.Y(n_195)
);

OA21x2_ASAP7_75t_L g184 ( 
.A1(n_152),
.A2(n_22),
.B(n_30),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_184),
.A2(n_157),
.B1(n_169),
.B2(n_168),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_171),
.Y(n_189)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_189),
.Y(n_197)
);

HB1xp67_ASAP7_75t_L g202 ( 
.A(n_190),
.Y(n_202)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_173),
.Y(n_191)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_177),
.A2(n_168),
.B1(n_166),
.B2(n_39),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_193),
.A2(n_194),
.B1(n_184),
.B2(n_187),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_183),
.B1(n_175),
.B2(n_182),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_196),
.A2(n_175),
.B(n_184),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_199),
.A2(n_190),
.B(n_192),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_200),
.B(n_201),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_194),
.B(n_187),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_178),
.C(n_174),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_SL g207 ( 
.A(n_203),
.B(n_193),
.Y(n_207)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_198),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_205),
.B(n_207),
.C(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_206),
.B(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_208),
.B(n_209),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_210),
.B(n_188),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_SL g212 ( 
.A1(n_211),
.A2(n_204),
.B(n_176),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_212),
.A2(n_36),
.B(n_37),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_213),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_214),
.A2(n_40),
.B(n_44),
.Y(n_215)
);

XNOR2x2_ASAP7_75t_SL g216 ( 
.A(n_215),
.B(n_45),
.Y(n_216)
);


endmodule