module fake_netlist_5_1708_n_900 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_900);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_900;

wire n_676;
wire n_294;
wire n_431;
wire n_380;
wire n_419;
wire n_318;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_194;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_643;
wire n_620;
wire n_452;
wire n_885;
wire n_397;
wire n_493;
wire n_525;
wire n_880;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_501;
wire n_245;
wire n_284;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_629;
wire n_590;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_898;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_247;
wire n_368;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_516;
wire n_498;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_640;
wire n_275;
wire n_559;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_568;
wire n_509;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_186;
wire n_537;
wire n_191;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_878;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_883;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_449;
wire n_325;
wire n_862;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_896;
wire n_323;
wire n_569;
wire n_769;
wire n_195;
wire n_356;
wire n_227;
wire n_592;
wire n_894;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_886;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_192;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_750;
wire n_742;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_882;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_178;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_395;
wire n_432;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_888;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_184;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_772;
wire n_691;
wire n_881;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_402;
wire n_413;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_889;
wire n_277;
wire n_338;
wire n_571;
wire n_477;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_188;
wire n_190;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_892;
wire n_893;
wire n_891;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_632;
wire n_489;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_349;
wire n_585;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_884;
wire n_899;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_557;
wire n_182;
wire n_354;
wire n_575;
wire n_607;
wire n_647;
wire n_480;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_679;
wire n_710;
wire n_707;
wire n_832;
wire n_695;
wire n_795;
wire n_180;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_665;
wire n_602;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_879;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_179;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_895;
wire n_202;
wire n_266;
wire n_491;
wire n_272;
wire n_427;
wire n_791;
wire n_732;
wire n_193;
wire n_251;
wire n_352;
wire n_566;
wire n_565;
wire n_426;
wire n_520;
wire n_808;
wire n_409;
wire n_797;
wire n_887;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_890;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_187;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_103),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_69),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_94),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_70),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_30),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_55),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_117),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g189 ( 
.A(n_83),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_12),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_171),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_86),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_157),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_12),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_72),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_121),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_37),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_43),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_168),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_135),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_24),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_10),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_119),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_134),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_52),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g208 ( 
.A(n_131),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_62),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_99),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_38),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_104),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_44),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_41),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_35),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_174),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_77),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_32),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_153),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_7),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_112),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_84),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_116),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_36),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_5),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_128),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_97),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_154),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_100),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_66),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_9),
.Y(n_233)
);

BUFx10_ASAP7_75t_L g234 ( 
.A(n_74),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_136),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_166),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_46),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_61),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_63),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_161),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_120),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_173),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_82),
.Y(n_245)
);

BUFx10_ASAP7_75t_L g246 ( 
.A(n_75),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_114),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_160),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_106),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_48),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_147),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_177),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_167),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_80),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_73),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_90),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_102),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_42),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_18),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_15),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_165),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_26),
.Y(n_262)
);

BUFx10_ASAP7_75t_L g263 ( 
.A(n_59),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_76),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_105),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_85),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_212),
.B(n_0),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_179),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_203),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_0),
.Y(n_270)
);

INVx5_ASAP7_75t_L g271 ( 
.A(n_179),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_221),
.Y(n_273)
);

INVx5_ASAP7_75t_L g274 ( 
.A(n_179),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_221),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_208),
.B(n_1),
.Y(n_276)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_185),
.B(n_31),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_237),
.B(n_1),
.Y(n_278)
);

BUFx12f_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_221),
.B(n_2),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_185),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_2),
.Y(n_282)
);

AND2x4_ASAP7_75t_L g283 ( 
.A(n_235),
.B(n_3),
.Y(n_283)
);

BUFx8_ASAP7_75t_L g284 ( 
.A(n_221),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_180),
.Y(n_285)
);

INVx2_ASAP7_75t_SL g286 ( 
.A(n_259),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_235),
.Y(n_287)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_181),
.Y(n_288)
);

INVx5_ASAP7_75t_L g289 ( 
.A(n_234),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_189),
.B(n_3),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_202),
.Y(n_291)
);

AND2x4_ASAP7_75t_L g292 ( 
.A(n_186),
.B(n_187),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_188),
.B(n_4),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_241),
.B(n_4),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_200),
.B(n_5),
.Y(n_295)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_193),
.B(n_6),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_214),
.B(n_6),
.Y(n_298)
);

BUFx8_ASAP7_75t_SL g299 ( 
.A(n_238),
.Y(n_299)
);

INVx5_ASAP7_75t_L g300 ( 
.A(n_234),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_246),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_246),
.B(n_7),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_217),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_195),
.B(n_8),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_259),
.B(n_8),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_246),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_233),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_263),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_263),
.B(n_9),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_220),
.B(n_10),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_232),
.Y(n_311)
);

BUFx12f_ASAP7_75t_L g312 ( 
.A(n_263),
.Y(n_312)
);

INVx5_ASAP7_75t_L g313 ( 
.A(n_178),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_182),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_245),
.B(n_11),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_33),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_260),
.Y(n_318)
);

BUFx12f_ASAP7_75t_L g319 ( 
.A(n_184),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_190),
.B(n_13),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_194),
.B(n_13),
.Y(n_321)
);

BUFx8_ASAP7_75t_SL g322 ( 
.A(n_238),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_253),
.Y(n_323)
);

INVx5_ASAP7_75t_L g324 ( 
.A(n_183),
.Y(n_324)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_191),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_262),
.Y(n_327)
);

INVx2_ASAP7_75t_SL g328 ( 
.A(n_289),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_273),
.Y(n_329)
);

AOI22x1_ASAP7_75t_L g330 ( 
.A1(n_309),
.A2(n_227),
.B1(n_226),
.B2(n_225),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_302),
.A2(n_256),
.B1(n_257),
.B2(n_264),
.Y(n_331)
);

INVx8_ASAP7_75t_L g332 ( 
.A(n_312),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_275),
.Y(n_333)
);

OAI22xp33_ASAP7_75t_SL g334 ( 
.A1(n_267),
.A2(n_266),
.B1(n_192),
.B2(n_261),
.Y(n_334)
);

OAI22xp33_ASAP7_75t_L g335 ( 
.A1(n_301),
.A2(n_265),
.B1(n_258),
.B2(n_198),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_294),
.A2(n_223),
.B1(n_197),
.B2(n_255),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_268),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g338 ( 
.A1(n_305),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_338)
);

AO22x2_ASAP7_75t_L g339 ( 
.A1(n_305),
.A2(n_321),
.B1(n_283),
.B2(n_278),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_281),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_301),
.A2(n_265),
.B1(n_258),
.B2(n_204),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_281),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_314),
.B(n_196),
.Y(n_344)
);

OR2x6_ASAP7_75t_L g345 ( 
.A(n_279),
.B(n_218),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_281),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_290),
.A2(n_252),
.B1(n_251),
.B2(n_250),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_314),
.B(n_199),
.Y(n_348)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_289),
.B(n_201),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_321),
.A2(n_14),
.B1(n_16),
.B2(n_17),
.Y(n_350)
);

AO22x2_ASAP7_75t_L g351 ( 
.A1(n_283),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_222),
.B1(n_247),
.B2(n_243),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_SL g354 ( 
.A1(n_297),
.A2(n_248),
.B1(n_242),
.B2(n_240),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_268),
.Y(n_355)
);

AO22x2_ASAP7_75t_L g356 ( 
.A1(n_293),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.Y(n_356)
);

BUFx10_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_304),
.A2(n_319),
.B1(n_320),
.B2(n_279),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_287),
.Y(n_359)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_268),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_289),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_268),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_287),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_304),
.A2(n_215),
.B1(n_231),
.B2(n_230),
.Y(n_364)
);

BUFx6f_ASAP7_75t_SL g365 ( 
.A(n_306),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_287),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_SL g367 ( 
.A1(n_276),
.A2(n_236),
.B1(n_229),
.B2(n_228),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_312),
.B1(n_306),
.B2(n_316),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_288),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_289),
.B(n_296),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_296),
.B(n_205),
.Y(n_371)
);

AO22x2_ASAP7_75t_L g372 ( 
.A1(n_293),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_316),
.A2(n_211),
.B1(n_219),
.B2(n_216),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_316),
.A2(n_224),
.B1(n_213),
.B2(n_210),
.Y(n_374)
);

AND2x2_ASAP7_75t_SL g375 ( 
.A(n_270),
.B(n_22),
.Y(n_375)
);

OAI22xp33_ASAP7_75t_L g376 ( 
.A1(n_296),
.A2(n_209),
.B1(n_207),
.B2(n_206),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_295),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_377)
);

NOR2x1p5_ASAP7_75t_L g378 ( 
.A(n_282),
.B(n_25),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_L g379 ( 
.A1(n_296),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_288),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_300),
.B(n_34),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_288),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_382),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_370),
.B(n_300),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_332),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_340),
.Y(n_388)
);

INVxp33_ASAP7_75t_L g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_341),
.Y(n_390)
);

XOR2x2_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_299),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_358),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_300),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_343),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_346),
.Y(n_396)
);

AND2x6_ASAP7_75t_L g397 ( 
.A(n_381),
.B(n_277),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_357),
.B(n_300),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_355),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_347),
.B(n_308),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_360),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_332),
.Y(n_404)
);

AND2x6_ASAP7_75t_L g405 ( 
.A(n_377),
.B(n_295),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_363),
.Y(n_406)
);

OR2x6_ASAP7_75t_L g407 ( 
.A(n_351),
.B(n_285),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_352),
.B(n_308),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_366),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_333),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_329),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_373),
.A2(n_292),
.B(n_310),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_344),
.B(n_308),
.Y(n_415)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_339),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_360),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_378),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_349),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_308),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_339),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_330),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_351),
.Y(n_423)
);

NAND2x1p5_ASAP7_75t_L g424 ( 
.A(n_328),
.B(n_298),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_356),
.Y(n_425)
);

NAND2xp33_ASAP7_75t_R g426 ( 
.A(n_345),
.B(n_298),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_361),
.B(n_292),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_356),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_372),
.Y(n_429)
);

AND2x4_ASAP7_75t_L g430 ( 
.A(n_374),
.B(n_269),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_348),
.B(n_313),
.Y(n_431)
);

XOR2x2_ASAP7_75t_L g432 ( 
.A(n_368),
.B(n_299),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_345),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_371),
.B(n_313),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_331),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_338),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_336),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_338),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_334),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_350),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_350),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_354),
.B(n_292),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_379),
.Y(n_444)
);

AND2x2_ASAP7_75t_SL g445 ( 
.A(n_335),
.B(n_310),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_365),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_337),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_337),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_370),
.B(n_285),
.Y(n_450)
);

INVx8_ASAP7_75t_L g451 ( 
.A(n_332),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_393),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_399),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_448),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_387),
.Y(n_455)
);

INVx2_ASAP7_75t_SL g456 ( 
.A(n_419),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_419),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_450),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_414),
.B(n_313),
.Y(n_459)
);

AND2x2_ASAP7_75t_SL g460 ( 
.A(n_445),
.B(n_315),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_449),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_411),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_412),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_419),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_402),
.Y(n_465)
);

INVx2_ASAP7_75t_SL g466 ( 
.A(n_422),
.Y(n_466)
);

INVx2_ASAP7_75t_SL g467 ( 
.A(n_427),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_421),
.B(n_291),
.Y(n_468)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_436),
.A2(n_280),
.B(n_318),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_418),
.B(n_322),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_410),
.Y(n_471)
);

BUFx6f_ASAP7_75t_L g472 ( 
.A(n_438),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_416),
.B(n_291),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_402),
.Y(n_474)
);

OR2x2_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_327),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_414),
.B(n_288),
.Y(n_476)
);

AND2x4_ASAP7_75t_SL g477 ( 
.A(n_438),
.B(n_280),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_388),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

INVxp67_ASAP7_75t_SL g480 ( 
.A(n_383),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_397),
.B(n_303),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_443),
.A2(n_307),
.B(n_317),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_395),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_445),
.B(n_307),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_398),
.B(n_317),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_396),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_451),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_401),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_403),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_407),
.B(n_327),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_407),
.B(n_303),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_439),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_407),
.B(n_303),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_409),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_397),
.B(n_303),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_397),
.B(n_311),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_397),
.Y(n_499)
);

INVx3_ASAP7_75t_SL g500 ( 
.A(n_451),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_385),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_386),
.Y(n_502)
);

AND2x2_ASAP7_75t_SL g503 ( 
.A(n_440),
.B(n_311),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_394),
.B(n_313),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_420),
.B(n_311),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_430),
.B(n_311),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_430),
.B(n_326),
.Y(n_507)
);

INVx4_ASAP7_75t_L g508 ( 
.A(n_397),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_413),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_429),
.B(n_326),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_424),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_417),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_447),
.B(n_39),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_427),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_443),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_437),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_441),
.B(n_323),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_442),
.B(n_323),
.Y(n_518)
);

BUFx3_ASAP7_75t_L g519 ( 
.A(n_424),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_405),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_423),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_458),
.B(n_322),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_457),
.B(n_446),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_452),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_514),
.B(n_394),
.Y(n_525)
);

CKINVDCx8_ASAP7_75t_R g526 ( 
.A(n_455),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

CKINVDCx9p33_ASAP7_75t_R g528 ( 
.A(n_470),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_452),
.Y(n_529)
);

AND2x2_ASAP7_75t_L g530 ( 
.A(n_458),
.B(n_486),
.Y(n_530)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_475),
.B(n_444),
.Y(n_531)
);

NAND2x1p5_ASAP7_75t_L g532 ( 
.A(n_457),
.B(n_425),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_453),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_457),
.B(n_440),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_457),
.Y(n_535)
);

OR2x2_ASAP7_75t_L g536 ( 
.A(n_475),
.B(n_428),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_514),
.B(n_400),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_514),
.B(n_400),
.Y(n_538)
);

AND2x4_ASAP7_75t_L g539 ( 
.A(n_511),
.B(n_435),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_493),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_SL g541 ( 
.A(n_488),
.B(n_404),
.Y(n_541)
);

OR2x2_ASAP7_75t_L g542 ( 
.A(n_473),
.B(n_391),
.Y(n_542)
);

CKINVDCx16_ASAP7_75t_R g543 ( 
.A(n_492),
.Y(n_543)
);

BUFx2_ASAP7_75t_L g544 ( 
.A(n_485),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_511),
.B(n_405),
.Y(n_545)
);

INVx4_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

BUFx3_ASAP7_75t_L g547 ( 
.A(n_500),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_486),
.B(n_408),
.Y(n_548)
);

NOR2xp33_ASAP7_75t_L g549 ( 
.A(n_472),
.B(n_389),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_467),
.B(n_408),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_453),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_506),
.B(n_389),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_467),
.B(n_405),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_453),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_467),
.B(n_405),
.Y(n_555)
);

OR2x6_ASAP7_75t_L g556 ( 
.A(n_472),
.B(n_451),
.Y(n_556)
);

NOR2xp67_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_415),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_454),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_454),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_500),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g562 ( 
.A(n_500),
.B(n_392),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g563 ( 
.A(n_473),
.B(n_493),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_503),
.B(n_405),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_472),
.B(n_479),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_457),
.Y(n_566)
);

INVx6_ASAP7_75t_L g567 ( 
.A(n_491),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_503),
.B(n_415),
.Y(n_568)
);

INVx4_ASAP7_75t_L g569 ( 
.A(n_457),
.Y(n_569)
);

AND2x4_ASAP7_75t_L g570 ( 
.A(n_511),
.B(n_434),
.Y(n_570)
);

AND2x6_ASAP7_75t_L g571 ( 
.A(n_499),
.B(n_513),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_506),
.B(n_432),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_482),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_472),
.B(n_433),
.Y(n_574)
);

AND2x4_ASAP7_75t_L g575 ( 
.A(n_519),
.B(n_384),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_519),
.B(n_431),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_519),
.B(n_431),
.Y(n_577)
);

BUFx12f_ASAP7_75t_L g578 ( 
.A(n_491),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_482),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_503),
.B(n_324),
.Y(n_580)
);

NAND2x1p5_ASAP7_75t_L g581 ( 
.A(n_546),
.B(n_464),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_552),
.Y(n_582)
);

CKINVDCx6p67_ASAP7_75t_R g583 ( 
.A(n_547),
.Y(n_583)
);

BUFx4_ASAP7_75t_SL g584 ( 
.A(n_560),
.Y(n_584)
);

INVx1_ASAP7_75t_SL g585 ( 
.A(n_540),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_526),
.Y(n_586)
);

CKINVDCx12_ASAP7_75t_R g587 ( 
.A(n_556),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_546),
.B(n_464),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_573),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_535),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_573),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_578),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g593 ( 
.A(n_563),
.B(n_485),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

NOR2x1_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_520),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_579),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_535),
.Y(n_597)
);

BUFx2_ASAP7_75t_SL g598 ( 
.A(n_539),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_569),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_579),
.Y(n_600)
);

BUFx2_ASAP7_75t_L g601 ( 
.A(n_544),
.Y(n_601)
);

INVx6_ASAP7_75t_L g602 ( 
.A(n_535),
.Y(n_602)
);

INVx4_ASAP7_75t_L g603 ( 
.A(n_566),
.Y(n_603)
);

INVx2_ASAP7_75t_SL g604 ( 
.A(n_566),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_524),
.Y(n_605)
);

BUFx3_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_524),
.Y(n_607)
);

BUFx12f_ASAP7_75t_L g608 ( 
.A(n_531),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_525),
.B(n_472),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_527),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_539),
.Y(n_611)
);

INVx2_ASAP7_75t_SL g612 ( 
.A(n_566),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_542),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_571),
.Y(n_614)
);

INVx8_ASAP7_75t_L g615 ( 
.A(n_571),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_565),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_530),
.B(n_460),
.Y(n_617)
);

BUFx3_ASAP7_75t_L g618 ( 
.A(n_575),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_569),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_537),
.B(n_472),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_572),
.Y(n_621)
);

INVx1_ASAP7_75t_SL g622 ( 
.A(n_543),
.Y(n_622)
);

INVx3_ASAP7_75t_SL g623 ( 
.A(n_536),
.Y(n_623)
);

BUFx2_ASAP7_75t_SL g624 ( 
.A(n_570),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_541),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_571),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_575),
.Y(n_627)
);

BUFx3_ASAP7_75t_L g628 ( 
.A(n_523),
.Y(n_628)
);

BUFx12f_ASAP7_75t_L g629 ( 
.A(n_570),
.Y(n_629)
);

OAI22xp33_ASAP7_75t_L g630 ( 
.A1(n_593),
.A2(n_538),
.B1(n_550),
.B2(n_562),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_589),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_SL g632 ( 
.A1(n_608),
.A2(n_460),
.B1(n_549),
.B2(n_520),
.Y(n_632)
);

CKINVDCx8_ASAP7_75t_R g633 ( 
.A(n_592),
.Y(n_633)
);

AOI22xp33_ASAP7_75t_L g634 ( 
.A1(n_617),
.A2(n_460),
.B1(n_469),
.B2(n_548),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_586),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_596),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_SL g637 ( 
.A1(n_608),
.A2(n_520),
.B1(n_513),
.B2(n_564),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_591),
.Y(n_638)
);

BUFx4f_ASAP7_75t_SL g639 ( 
.A(n_629),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_626),
.B(n_619),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_593),
.B(n_617),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_585),
.Y(n_642)
);

BUFx2_ASAP7_75t_SL g643 ( 
.A(n_586),
.Y(n_643)
);

OAI22xp5_ASAP7_75t_L g644 ( 
.A1(n_616),
.A2(n_472),
.B1(n_479),
.B2(n_545),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_614),
.Y(n_645)
);

AOI22xp33_ASAP7_75t_L g646 ( 
.A1(n_582),
.A2(n_545),
.B1(n_534),
.B2(n_479),
.Y(n_646)
);

OAI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_613),
.A2(n_522),
.B(n_574),
.Y(n_647)
);

BUFx12f_ASAP7_75t_L g648 ( 
.A(n_592),
.Y(n_648)
);

OAI21xp33_ASAP7_75t_L g649 ( 
.A1(n_625),
.A2(n_477),
.B(n_507),
.Y(n_649)
);

INVx2_ASAP7_75t_SL g650 ( 
.A(n_584),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

BUFx2_ASAP7_75t_L g652 ( 
.A(n_623),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_621),
.Y(n_653)
);

BUFx2_ASAP7_75t_L g654 ( 
.A(n_623),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_605),
.Y(n_655)
);

NOR2x1_ASAP7_75t_L g656 ( 
.A(n_603),
.B(n_576),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_582),
.A2(n_479),
.B1(n_515),
.B2(n_477),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_582),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_607),
.Y(n_659)
);

AOI22xp33_ASAP7_75t_L g660 ( 
.A1(n_601),
.A2(n_479),
.B1(n_477),
.B2(n_494),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_601),
.A2(n_479),
.B1(n_492),
.B2(n_494),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_618),
.A2(n_479),
.B1(n_492),
.B2(n_494),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_594),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_591),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_611),
.Y(n_666)
);

OR2x2_ASAP7_75t_L g667 ( 
.A(n_622),
.B(n_507),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_611),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_629),
.Y(n_669)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_621),
.A2(n_426),
.B1(n_577),
.B2(n_576),
.Y(n_670)
);

AOI22xp33_ASAP7_75t_L g671 ( 
.A1(n_618),
.A2(n_491),
.B1(n_513),
.B2(n_459),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_594),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_631),
.Y(n_673)
);

BUFx8_ASAP7_75t_L g674 ( 
.A(n_672),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_647),
.B(n_606),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_649),
.A2(n_513),
.B1(n_577),
.B2(n_568),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_630),
.A2(n_557),
.B(n_580),
.Y(n_677)
);

OAI22xp5_ASAP7_75t_L g678 ( 
.A1(n_637),
.A2(n_598),
.B1(n_583),
.B2(n_555),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_637),
.A2(n_583),
.B1(n_553),
.B2(n_624),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_670),
.A2(n_532),
.B1(n_456),
.B2(n_627),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_632),
.A2(n_456),
.B1(n_471),
.B2(n_504),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_636),
.Y(n_682)
);

AOI22xp33_ASAP7_75t_L g683 ( 
.A1(n_632),
.A2(n_456),
.B1(n_471),
.B2(n_627),
.Y(n_683)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_630),
.A2(n_471),
.B1(n_469),
.B2(n_464),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_L g685 ( 
.A1(n_634),
.A2(n_464),
.B1(n_463),
.B2(n_505),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_651),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_641),
.B(n_606),
.Y(n_687)
);

AOI22xp33_ASAP7_75t_L g688 ( 
.A1(n_634),
.A2(n_464),
.B1(n_463),
.B2(n_505),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_638),
.Y(n_689)
);

OAI21xp5_ASAP7_75t_SL g690 ( 
.A1(n_657),
.A2(n_476),
.B(n_426),
.Y(n_690)
);

AOI222xp33_ASAP7_75t_L g691 ( 
.A1(n_642),
.A2(n_516),
.B1(n_468),
.B2(n_518),
.C1(n_517),
.C2(n_476),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_SL g692 ( 
.A1(n_646),
.A2(n_528),
.B(n_483),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_643),
.A2(n_571),
.B1(n_508),
.B2(n_499),
.Y(n_693)
);

AOI22xp33_ASAP7_75t_L g694 ( 
.A1(n_667),
.A2(n_464),
.B1(n_463),
.B2(n_483),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_665),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_635),
.A2(n_587),
.B1(n_480),
.B2(n_517),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_652),
.A2(n_464),
.B1(n_502),
.B2(n_501),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_640),
.Y(n_698)
);

AOI222xp33_ASAP7_75t_L g699 ( 
.A1(n_654),
.A2(n_516),
.B1(n_468),
.B2(n_518),
.C1(n_510),
.C2(n_521),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_660),
.A2(n_609),
.B1(n_620),
.B2(n_628),
.Y(n_700)
);

OAI22xp5_ASAP7_75t_L g701 ( 
.A1(n_671),
.A2(n_628),
.B1(n_480),
.B2(n_615),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_659),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_661),
.Y(n_704)
);

AOI22xp33_ASAP7_75t_L g705 ( 
.A1(n_663),
.A2(n_478),
.B1(n_502),
.B2(n_501),
.Y(n_705)
);

AOI22xp33_ASAP7_75t_L g706 ( 
.A1(n_662),
.A2(n_487),
.B1(n_478),
.B2(n_496),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_669),
.A2(n_496),
.B1(n_487),
.B2(n_466),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_666),
.B(n_510),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_640),
.Y(n_709)
);

AOI22xp5_ASAP7_75t_L g710 ( 
.A1(n_653),
.A2(n_587),
.B1(n_518),
.B2(n_595),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_658),
.A2(n_466),
.B1(n_508),
.B2(n_499),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_644),
.A2(n_615),
.B1(n_614),
.B2(n_626),
.Y(n_712)
);

BUFx6f_ASAP7_75t_L g713 ( 
.A(n_645),
.Y(n_713)
);

AOI22xp33_ASAP7_75t_L g714 ( 
.A1(n_669),
.A2(n_484),
.B1(n_489),
.B2(n_495),
.Y(n_714)
);

OAI222xp33_ASAP7_75t_L g715 ( 
.A1(n_656),
.A2(n_466),
.B1(n_527),
.B2(n_529),
.C1(n_554),
.C2(n_561),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_669),
.A2(n_668),
.B1(n_489),
.B2(n_484),
.Y(n_716)
);

OAI21xp5_ASAP7_75t_SL g717 ( 
.A1(n_650),
.A2(n_497),
.B(n_481),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_645),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_672),
.A2(n_462),
.B1(n_495),
.B2(n_490),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_664),
.B(n_521),
.Y(n_720)
);

OAI22xp33_ASAP7_75t_L g721 ( 
.A1(n_639),
.A2(n_508),
.B1(n_499),
.B2(n_614),
.Y(n_721)
);

NOR2x1_ASAP7_75t_L g722 ( 
.A(n_639),
.B(n_603),
.Y(n_722)
);

OAI21xp33_ASAP7_75t_L g723 ( 
.A1(n_633),
.A2(n_462),
.B(n_495),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_648),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_647),
.B(n_461),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_725),
.A2(n_489),
.B1(n_490),
.B2(n_484),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_687),
.B(n_482),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_675),
.A2(n_490),
.B1(n_499),
.B2(n_508),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_691),
.A2(n_499),
.B1(n_461),
.B2(n_498),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_699),
.A2(n_499),
.B1(n_497),
.B2(n_498),
.Y(n_730)
);

AOI22xp33_ASAP7_75t_SL g731 ( 
.A1(n_679),
.A2(n_614),
.B1(n_615),
.B2(n_626),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_696),
.A2(n_615),
.B1(n_481),
.B2(n_581),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_720),
.A2(n_512),
.B1(n_509),
.B2(n_284),
.Y(n_733)
);

AOI22xp33_ASAP7_75t_L g734 ( 
.A1(n_723),
.A2(n_676),
.B1(n_680),
.B2(n_678),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_701),
.A2(n_512),
.B1(n_509),
.B2(n_284),
.Y(n_735)
);

AOI221xp5_ASAP7_75t_L g736 ( 
.A1(n_690),
.A2(n_326),
.B1(n_323),
.B2(n_512),
.C(n_509),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_SL g737 ( 
.A1(n_674),
.A2(n_599),
.B1(n_619),
.B2(n_588),
.Y(n_737)
);

NAND3xp33_ASAP7_75t_L g738 ( 
.A(n_717),
.B(n_326),
.C(n_323),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_673),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_710),
.A2(n_588),
.B1(n_581),
.B2(n_599),
.Y(n_740)
);

AOI22xp33_ASAP7_75t_SL g741 ( 
.A1(n_674),
.A2(n_599),
.B1(n_619),
.B2(n_597),
.Y(n_741)
);

AOI22xp33_ASAP7_75t_L g742 ( 
.A1(n_677),
.A2(n_533),
.B1(n_551),
.B2(n_559),
.Y(n_742)
);

OAI22xp5_ASAP7_75t_L g743 ( 
.A1(n_719),
.A2(n_619),
.B1(n_602),
.B2(n_604),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_683),
.A2(n_554),
.B1(n_529),
.B2(n_558),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_682),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_692),
.A2(n_602),
.B1(n_619),
.B2(n_603),
.Y(n_746)
);

AOI22xp33_ASAP7_75t_SL g747 ( 
.A1(n_712),
.A2(n_597),
.B1(n_590),
.B2(n_602),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_689),
.B(n_558),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_719),
.A2(n_561),
.B1(n_465),
.B2(n_474),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_724),
.A2(n_681),
.B1(n_706),
.B2(n_705),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_SL g751 ( 
.A(n_707),
.B(n_597),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_695),
.Y(n_752)
);

OAI22xp5_ASAP7_75t_L g753 ( 
.A1(n_707),
.A2(n_602),
.B1(n_604),
.B2(n_612),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_711),
.A2(n_474),
.B1(n_465),
.B2(n_612),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_704),
.B(n_590),
.Y(n_755)
);

AOI22xp33_ASAP7_75t_L g756 ( 
.A1(n_711),
.A2(n_474),
.B1(n_465),
.B2(n_597),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_700),
.A2(n_474),
.B1(n_465),
.B2(n_597),
.Y(n_757)
);

AOI22xp33_ASAP7_75t_L g758 ( 
.A1(n_684),
.A2(n_590),
.B1(n_325),
.B2(n_324),
.Y(n_758)
);

OAI221xp5_ASAP7_75t_SL g759 ( 
.A1(n_697),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.C(n_30),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_716),
.A2(n_590),
.B1(n_325),
.B2(n_324),
.Y(n_760)
);

NAND3xp33_ASAP7_75t_L g761 ( 
.A(n_714),
.B(n_325),
.C(n_324),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_708),
.A2(n_685),
.B1(n_688),
.B2(n_718),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_709),
.A2(n_325),
.B1(n_272),
.B2(n_274),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_686),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_752),
.B(n_727),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_752),
.B(n_702),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_764),
.B(n_703),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_739),
.B(n_698),
.Y(n_768)
);

NAND3xp33_ASAP7_75t_L g769 ( 
.A(n_733),
.B(n_694),
.C(n_698),
.Y(n_769)
);

AND2x2_ASAP7_75t_SL g770 ( 
.A(n_734),
.B(n_698),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_739),
.B(n_698),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_737),
.B(n_713),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_745),
.B(n_713),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_745),
.B(n_713),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_764),
.B(n_713),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_755),
.B(n_693),
.Y(n_776)
);

AOI211xp5_ASAP7_75t_L g777 ( 
.A1(n_759),
.A2(n_721),
.B(n_715),
.C(n_29),
.Y(n_777)
);

NOR2x1p5_ASAP7_75t_L g778 ( 
.A(n_738),
.B(n_722),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_729),
.B(n_693),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_762),
.B(n_721),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_750),
.B(n_272),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_SL g782 ( 
.A1(n_732),
.A2(n_715),
.B1(n_272),
.B2(n_274),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_730),
.B(n_272),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_731),
.B(n_40),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_748),
.B(n_45),
.Y(n_785)
);

OA211x2_ASAP7_75t_L g786 ( 
.A1(n_736),
.A2(n_47),
.B(n_49),
.C(n_50),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_735),
.A2(n_274),
.B1(n_271),
.B2(n_54),
.Y(n_787)
);

NAND3xp33_ASAP7_75t_L g788 ( 
.A(n_726),
.B(n_274),
.C(n_271),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_751),
.A2(n_271),
.B1(n_53),
.B2(n_56),
.Y(n_789)
);

NAND3xp33_ASAP7_75t_L g790 ( 
.A(n_728),
.B(n_271),
.C(n_57),
.Y(n_790)
);

OAI22xp5_ASAP7_75t_L g791 ( 
.A1(n_746),
.A2(n_51),
.B1(n_58),
.B2(n_60),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_777),
.B(n_747),
.C(n_741),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_767),
.B(n_757),
.Y(n_793)
);

NAND4xp75_ASAP7_75t_L g794 ( 
.A(n_786),
.B(n_751),
.C(n_740),
.D(n_756),
.Y(n_794)
);

OAI211xp5_ASAP7_75t_SL g795 ( 
.A1(n_789),
.A2(n_772),
.B(n_787),
.C(n_768),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_767),
.B(n_761),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_765),
.B(n_758),
.Y(n_797)
);

NAND3xp33_ASAP7_75t_L g798 ( 
.A(n_769),
.B(n_763),
.C(n_760),
.Y(n_798)
);

AO21x2_ASAP7_75t_L g799 ( 
.A1(n_781),
.A2(n_743),
.B(n_753),
.Y(n_799)
);

AOI211xp5_ASAP7_75t_L g800 ( 
.A1(n_791),
.A2(n_64),
.B(n_65),
.C(n_67),
.Y(n_800)
);

NOR3xp33_ASAP7_75t_L g801 ( 
.A(n_785),
.B(n_744),
.C(n_754),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_770),
.A2(n_742),
.B1(n_749),
.B2(n_78),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_774),
.B(n_68),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_790),
.B(n_71),
.C(n_79),
.Y(n_804)
);

OR2x2_ASAP7_75t_L g805 ( 
.A(n_771),
.B(n_81),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_766),
.B(n_88),
.Y(n_806)
);

NOR3xp33_ASAP7_75t_L g807 ( 
.A(n_784),
.B(n_89),
.C(n_91),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_773),
.B(n_92),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_796),
.Y(n_809)
);

NAND4xp25_ASAP7_75t_L g810 ( 
.A(n_792),
.B(n_775),
.C(n_789),
.D(n_780),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_799),
.B(n_770),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_793),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_799),
.B(n_776),
.Y(n_813)
);

INVx1_ASAP7_75t_SL g814 ( 
.A(n_803),
.Y(n_814)
);

NAND4xp75_ASAP7_75t_L g815 ( 
.A(n_797),
.B(n_779),
.C(n_783),
.D(n_778),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_806),
.Y(n_816)
);

NAND4xp75_ASAP7_75t_SL g817 ( 
.A(n_794),
.B(n_782),
.C(n_788),
.D(n_96),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_805),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_809),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_813),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_818),
.Y(n_821)
);

XNOR2x1_ASAP7_75t_L g822 ( 
.A(n_814),
.B(n_798),
.Y(n_822)
);

XNOR2xp5_ASAP7_75t_L g823 ( 
.A(n_815),
.B(n_800),
.Y(n_823)
);

XOR2x2_ASAP7_75t_L g824 ( 
.A(n_817),
.B(n_807),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_823),
.B(n_811),
.Y(n_825)
);

OAI22xp5_ASAP7_75t_L g826 ( 
.A1(n_822),
.A2(n_811),
.B1(n_812),
.B2(n_813),
.Y(n_826)
);

INVx3_ASAP7_75t_L g827 ( 
.A(n_819),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_819),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_828),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_827),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_826),
.A2(n_824),
.B1(n_820),
.B2(n_810),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_827),
.Y(n_832)
);

AOI221xp5_ASAP7_75t_L g833 ( 
.A1(n_831),
.A2(n_825),
.B1(n_820),
.B2(n_821),
.C(n_816),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_829),
.Y(n_834)
);

OA22x2_ASAP7_75t_L g835 ( 
.A1(n_832),
.A2(n_816),
.B1(n_818),
.B2(n_808),
.Y(n_835)
);

AOI22x1_ASAP7_75t_L g836 ( 
.A1(n_834),
.A2(n_830),
.B1(n_795),
.B2(n_804),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_835),
.Y(n_837)
);

HB1xp67_ASAP7_75t_L g838 ( 
.A(n_833),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_834),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_839),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_838),
.B(n_830),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_838),
.B(n_782),
.Y(n_842)
);

NOR4xp25_ASAP7_75t_L g843 ( 
.A(n_837),
.B(n_802),
.C(n_95),
.D(n_98),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_836),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_839),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_838),
.A2(n_801),
.B1(n_101),
.B2(n_107),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_840),
.B(n_93),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_844),
.B(n_108),
.Y(n_848)
);

NOR3x1_ASAP7_75t_L g849 ( 
.A(n_841),
.B(n_109),
.C(n_110),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_845),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_842),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_843),
.B(n_113),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_846),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_844),
.B(n_115),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_841),
.Y(n_855)
);

AND3x1_ASAP7_75t_L g856 ( 
.A(n_853),
.B(n_118),
.C(n_122),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_855),
.Y(n_857)
);

AO22x2_ASAP7_75t_L g858 ( 
.A1(n_850),
.A2(n_123),
.B1(n_124),
.B2(n_125),
.Y(n_858)
);

INVx3_ASAP7_75t_L g859 ( 
.A(n_847),
.Y(n_859)
);

NAND4xp25_ASAP7_75t_L g860 ( 
.A(n_851),
.B(n_126),
.C(n_127),
.D(n_129),
.Y(n_860)
);

INVx4_ASAP7_75t_L g861 ( 
.A(n_849),
.Y(n_861)
);

INVxp67_ASAP7_75t_SL g862 ( 
.A(n_848),
.Y(n_862)
);

NAND5xp2_ASAP7_75t_L g863 ( 
.A(n_852),
.B(n_130),
.C(n_132),
.D(n_133),
.E(n_137),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_857),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_858),
.Y(n_865)
);

INVxp67_ASAP7_75t_SL g866 ( 
.A(n_862),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_859),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_856),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_858),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_861),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_863),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_860),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_857),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_866),
.Y(n_874)
);

HB1xp67_ASAP7_75t_L g875 ( 
.A(n_869),
.Y(n_875)
);

AOI22xp5_ASAP7_75t_L g876 ( 
.A1(n_870),
.A2(n_854),
.B1(n_139),
.B2(n_140),
.Y(n_876)
);

OAI22xp5_ASAP7_75t_SL g877 ( 
.A1(n_866),
.A2(n_868),
.B1(n_865),
.B2(n_871),
.Y(n_877)
);

HB1xp67_ASAP7_75t_L g878 ( 
.A(n_864),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_873),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_867),
.Y(n_880)
);

INVxp33_ASAP7_75t_SL g881 ( 
.A(n_871),
.Y(n_881)
);

AOI22xp33_ASAP7_75t_L g882 ( 
.A1(n_872),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_882)
);

AO22x2_ASAP7_75t_L g883 ( 
.A1(n_869),
.A2(n_176),
.B1(n_144),
.B2(n_145),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_875),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_874),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_877),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_878),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_879),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_880),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_886),
.A2(n_881),
.B1(n_876),
.B2(n_883),
.Y(n_890)
);

AOI22xp5_ASAP7_75t_L g891 ( 
.A1(n_884),
.A2(n_882),
.B1(n_146),
.B2(n_148),
.Y(n_891)
);

AOI22xp5_ASAP7_75t_L g892 ( 
.A1(n_887),
.A2(n_143),
.B1(n_149),
.B2(n_151),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_892),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_890),
.Y(n_894)
);

OAI22xp5_ASAP7_75t_L g895 ( 
.A1(n_894),
.A2(n_885),
.B1(n_889),
.B2(n_888),
.Y(n_895)
);

AOI22xp5_ASAP7_75t_L g896 ( 
.A1(n_893),
.A2(n_891),
.B1(n_888),
.B2(n_156),
.Y(n_896)
);

INVxp67_ASAP7_75t_L g897 ( 
.A(n_895),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_896),
.Y(n_898)
);

AOI221xp5_ASAP7_75t_L g899 ( 
.A1(n_897),
.A2(n_152),
.B1(n_155),
.B2(n_158),
.C(n_159),
.Y(n_899)
);

AOI211xp5_ASAP7_75t_L g900 ( 
.A1(n_899),
.A2(n_898),
.B(n_163),
.C(n_164),
.Y(n_900)
);


endmodule