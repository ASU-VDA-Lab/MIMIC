module fake_netlist_6_2974_n_1799 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_157, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1799);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_157;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1799;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g159 ( 
.A(n_1),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_80),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_41),
.Y(n_161)
);

INVx2_ASAP7_75t_SL g162 ( 
.A(n_114),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_89),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_126),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_44),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_1),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_34),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_17),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_71),
.Y(n_171)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_97),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_73),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_10),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_46),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_132),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_95),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_46),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_79),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_110),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_64),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_107),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_143),
.Y(n_184)
);

INVxp67_ASAP7_75t_SL g185 ( 
.A(n_54),
.Y(n_185)
);

BUFx8_ASAP7_75t_SL g186 ( 
.A(n_10),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_144),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_28),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_131),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_26),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_21),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_25),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_52),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_61),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_100),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_123),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_29),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g200 ( 
.A(n_32),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g202 ( 
.A(n_96),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_122),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_2),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_125),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_134),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_75),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_56),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_5),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_151),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_106),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_39),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_142),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_138),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_154),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_38),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g218 ( 
.A(n_33),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_141),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_41),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_91),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_137),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_42),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_128),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_30),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_87),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_155),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_36),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_127),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_22),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_27),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_84),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_156),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_60),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_76),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_111),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_81),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_2),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_47),
.Y(n_241)
);

INVx2_ASAP7_75t_SL g242 ( 
.A(n_129),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_109),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_0),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_55),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_13),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_33),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_59),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_108),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_157),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_29),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_83),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_69),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_30),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_119),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_16),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_23),
.Y(n_257)
);

INVx2_ASAP7_75t_SL g258 ( 
.A(n_82),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_105),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_90),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_31),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_45),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g263 ( 
.A(n_139),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_45),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_25),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_37),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_115),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_86),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_22),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_146),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_93),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_36),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_5),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_78),
.Y(n_275)
);

BUFx10_ASAP7_75t_L g276 ( 
.A(n_11),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_99),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_101),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_58),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_8),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_149),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_17),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_38),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_130),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_26),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_4),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_55),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_37),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_20),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_4),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_24),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_28),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_0),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_9),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_67),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_35),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_145),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_19),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_21),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_31),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_19),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_48),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_65),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_140),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_58),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_113),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_118),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_51),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_52),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_13),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_158),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_27),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_43),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_9),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_77),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_11),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_35),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_186),
.Y(n_318)
);

INVxp33_ASAP7_75t_SL g319 ( 
.A(n_241),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_262),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_262),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_162),
.B(n_3),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_196),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_285),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_292),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_192),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_163),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_292),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_210),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_302),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_302),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_213),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_162),
.B(n_3),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_164),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_182),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_308),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_308),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_159),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_168),
.Y(n_340)
);

INVxp67_ASAP7_75t_SL g341 ( 
.A(n_159),
.Y(n_341)
);

BUFx6f_ASAP7_75t_SL g342 ( 
.A(n_263),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_161),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_161),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_171),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_167),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_167),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_177),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_180),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_181),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_242),
.B(n_6),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_184),
.Y(n_352)
);

INVxp67_ASAP7_75t_SL g353 ( 
.A(n_188),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_194),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_192),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_197),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_188),
.Y(n_357)
);

CKINVDCx14_ASAP7_75t_R g358 ( 
.A(n_202),
.Y(n_358)
);

CKINVDCx16_ASAP7_75t_R g359 ( 
.A(n_218),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_189),
.Y(n_360)
);

INVxp67_ASAP7_75t_SL g361 ( 
.A(n_189),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_191),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_191),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_172),
.B(n_6),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_198),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_213),
.Y(n_366)
);

INVxp33_ASAP7_75t_SL g367 ( 
.A(n_165),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_195),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_203),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_206),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_218),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_195),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_208),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_211),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_208),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_L g376 ( 
.A(n_172),
.B(n_7),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_214),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_242),
.B(n_7),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_301),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_221),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_215),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_221),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_232),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_213),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_232),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_244),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_216),
.Y(n_387)
);

HB1xp67_ASAP7_75t_L g388 ( 
.A(n_301),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_276),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_222),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_244),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_223),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_251),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_333),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_322),
.B(n_258),
.Y(n_395)
);

OA21x2_ASAP7_75t_L g396 ( 
.A1(n_333),
.A2(n_166),
.B(n_160),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_333),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_355),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_364),
.B(n_276),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_366),
.Y(n_400)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_341),
.B(n_346),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

BUFx2_ASAP7_75t_L g403 ( 
.A(n_379),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_366),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_366),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_334),
.B(n_351),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_378),
.B(n_258),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_339),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_364),
.B(n_226),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_384),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_343),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_344),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_263),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_376),
.B(n_228),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_341),
.B(n_229),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

INVx3_ASAP7_75t_L g418 ( 
.A(n_384),
.Y(n_418)
);

BUFx2_ASAP7_75t_L g419 ( 
.A(n_388),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_384),
.B(n_172),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_346),
.B(n_172),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_347),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

AND2x4_ASAP7_75t_L g426 ( 
.A(n_353),
.B(n_190),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_320),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_321),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_319),
.B(n_160),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_353),
.B(n_190),
.Y(n_431)
);

INVx3_ASAP7_75t_L g432 ( 
.A(n_321),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_327),
.B(n_276),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_323),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_360),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_323),
.Y(n_437)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_325),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_325),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_362),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_326),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_326),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_361),
.B(n_235),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_329),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_361),
.B(n_237),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_329),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_362),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_331),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_386),
.B(n_205),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_368),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_331),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_332),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_380),
.Y(n_455)
);

BUFx6f_ASAP7_75t_L g456 ( 
.A(n_332),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_386),
.B(n_238),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_368),
.B(n_239),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_372),
.B(n_243),
.Y(n_459)
);

NAND2xp33_ASAP7_75t_SL g460 ( 
.A(n_375),
.B(n_199),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_337),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_372),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_327),
.B(n_276),
.Y(n_463)
);

AND2x4_ASAP7_75t_L g464 ( 
.A(n_382),
.B(n_205),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_337),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_439),
.Y(n_466)
);

BUFx6f_ASAP7_75t_SL g467 ( 
.A(n_426),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_429),
.B(n_328),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_404),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_409),
.B(n_415),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_420),
.Y(n_471)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_404),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_439),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_439),
.Y(n_474)
);

BUFx10_ASAP7_75t_L g475 ( 
.A(n_429),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_420),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_439),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_420),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_439),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_422),
.Y(n_480)
);

BUFx10_ASAP7_75t_L g481 ( 
.A(n_422),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_166),
.Y(n_482)
);

OR2x2_ASAP7_75t_L g483 ( 
.A(n_455),
.B(n_359),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_426),
.B(n_389),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_338),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_406),
.B(n_367),
.Y(n_487)
);

OAI22xp33_ASAP7_75t_SL g488 ( 
.A1(n_406),
.A2(n_173),
.B1(n_271),
.B2(n_272),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_409),
.B(n_415),
.Y(n_489)
);

INVx4_ASAP7_75t_L g490 ( 
.A(n_404),
.Y(n_490)
);

AND2x2_ASAP7_75t_SL g491 ( 
.A(n_396),
.B(n_252),
.Y(n_491)
);

AND2x2_ASAP7_75t_SL g492 ( 
.A(n_396),
.B(n_252),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_460),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_395),
.B(n_335),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_395),
.B(n_340),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_404),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_439),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_420),
.Y(n_498)
);

INVx6_ASAP7_75t_L g499 ( 
.A(n_422),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_422),
.B(n_173),
.Y(n_500)
);

INVx4_ASAP7_75t_L g501 ( 
.A(n_404),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_420),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_439),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_414),
.B(n_401),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_407),
.B(n_345),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g507 ( 
.A(n_460),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_397),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_396),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_426),
.B(n_338),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_397),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_407),
.B(n_348),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_426),
.A2(n_245),
.B1(n_268),
.B2(n_264),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_408),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_408),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

BUFx6f_ASAP7_75t_L g520 ( 
.A(n_404),
.Y(n_520)
);

NAND2x1p5_ASAP7_75t_L g521 ( 
.A(n_431),
.B(n_176),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_397),
.Y(n_522)
);

AOI22xp33_ASAP7_75t_L g523 ( 
.A1(n_431),
.A2(n_245),
.B1(n_268),
.B2(n_264),
.Y(n_523)
);

AOI22xp33_ASAP7_75t_L g524 ( 
.A1(n_431),
.A2(n_251),
.B1(n_254),
.B2(n_290),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_414),
.B(n_401),
.Y(n_525)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_455),
.B(n_359),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_414),
.B(n_349),
.Y(n_527)
);

AOI22xp33_ASAP7_75t_L g528 ( 
.A1(n_431),
.A2(n_254),
.B1(n_287),
.B2(n_288),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_405),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_401),
.B(n_350),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_411),
.Y(n_531)
);

AOI22xp33_ASAP7_75t_SL g532 ( 
.A1(n_403),
.A2(n_371),
.B1(n_293),
.B2(n_217),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_431),
.A2(n_273),
.B1(n_256),
.B2(n_290),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_404),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_405),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_405),
.Y(n_537)
);

BUFx2_ASAP7_75t_L g538 ( 
.A(n_403),
.Y(n_538)
);

BUFx8_ASAP7_75t_SL g539 ( 
.A(n_403),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_416),
.B(n_352),
.Y(n_540)
);

INVx2_ASAP7_75t_SL g541 ( 
.A(n_414),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

INVx4_ASAP7_75t_L g544 ( 
.A(n_410),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_427),
.Y(n_545)
);

BUFx10_ASAP7_75t_L g546 ( 
.A(n_451),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_414),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_427),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_451),
.Y(n_549)
);

AOI22xp33_ASAP7_75t_L g550 ( 
.A1(n_451),
.A2(n_256),
.B1(n_273),
.B2(n_309),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_412),
.Y(n_551)
);

INVx4_ASAP7_75t_L g552 ( 
.A(n_410),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_451),
.B(n_354),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_416),
.B(n_356),
.Y(n_554)
);

AOI22xp33_ASAP7_75t_L g555 ( 
.A1(n_451),
.A2(n_287),
.B1(n_286),
.B2(n_288),
.Y(n_555)
);

AND3x2_ASAP7_75t_L g556 ( 
.A(n_419),
.B(n_170),
.C(n_185),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_443),
.Y(n_557)
);

INVx1_ASAP7_75t_SL g558 ( 
.A(n_419),
.Y(n_558)
);

NOR2x1p5_ASAP7_75t_L g559 ( 
.A(n_443),
.B(n_318),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_427),
.Y(n_560)
);

OR2x2_ASAP7_75t_L g561 ( 
.A(n_445),
.B(n_371),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_413),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_413),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_427),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_464),
.A2(n_286),
.B1(n_309),
.B2(n_316),
.Y(n_565)
);

AOI22xp33_ASAP7_75t_L g566 ( 
.A1(n_464),
.A2(n_316),
.B1(n_380),
.B2(n_271),
.Y(n_566)
);

BUFx2_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx4_ASAP7_75t_SL g568 ( 
.A(n_410),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g569 ( 
.A(n_445),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_410),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_457),
.B(n_365),
.Y(n_571)
);

OR2x6_ASAP7_75t_L g572 ( 
.A(n_399),
.B(n_176),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_410),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_457),
.B(n_369),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_427),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_464),
.A2(n_281),
.B1(n_187),
.B2(n_207),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_410),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_458),
.B(n_370),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_SL g579 ( 
.A(n_433),
.B(n_374),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_458),
.B(n_377),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_417),
.Y(n_581)
);

AOI22xp33_ASAP7_75t_L g582 ( 
.A1(n_464),
.A2(n_231),
.B1(n_183),
.B2(n_187),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_459),
.B(n_392),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_417),
.Y(n_584)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_398),
.A2(n_336),
.B1(n_390),
.B2(n_387),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_398),
.B(n_459),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_433),
.B(n_381),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_423),
.B(n_382),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_423),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_427),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_424),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_424),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_399),
.B(n_358),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_427),
.Y(n_594)
);

AND2x6_ASAP7_75t_L g595 ( 
.A(n_464),
.B(n_213),
.Y(n_595)
);

INVx2_ASAP7_75t_SL g596 ( 
.A(n_463),
.Y(n_596)
);

AND2x6_ASAP7_75t_L g597 ( 
.A(n_410),
.B(n_213),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_425),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_425),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_437),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_463),
.B(n_213),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_430),
.A2(n_183),
.B1(n_207),
.B2(n_219),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_430),
.B(n_250),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_434),
.B(n_255),
.Y(n_604)
);

NAND2xp33_ASAP7_75t_R g605 ( 
.A(n_434),
.B(n_169),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_437),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_436),
.B(n_259),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_437),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_436),
.B(n_174),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_437),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_440),
.B(n_260),
.Y(n_611)
);

BUFx10_ASAP7_75t_L g612 ( 
.A(n_440),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_437),
.Y(n_613)
);

INVx1_ASAP7_75t_SL g614 ( 
.A(n_447),
.Y(n_614)
);

NOR2x1p5_ASAP7_75t_L g615 ( 
.A(n_447),
.B(n_175),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_394),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_480),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_480),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_471),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_557),
.B(n_428),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_509),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_557),
.B(n_428),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_487),
.A2(n_330),
.B1(n_324),
.B2(n_275),
.Y(n_623)
);

BUFx5_ASAP7_75t_L g624 ( 
.A(n_505),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_470),
.B(n_428),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_546),
.B(n_224),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_L g627 ( 
.A(n_489),
.B(n_267),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_494),
.B(n_428),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_471),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_495),
.B(n_428),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_506),
.B(n_432),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_514),
.B(n_432),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_476),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_569),
.B(n_586),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_554),
.B(n_432),
.Y(n_635)
);

AO22x2_ASAP7_75t_L g636 ( 
.A1(n_596),
.A2(n_248),
.B1(n_219),
.B2(n_231),
.Y(n_636)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_569),
.B(n_200),
.Y(n_637)
);

NAND2xp33_ASAP7_75t_L g638 ( 
.A(n_541),
.B(n_269),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_580),
.B(n_432),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_614),
.B(n_558),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_509),
.Y(n_641)
);

INVx2_ASAP7_75t_SL g642 ( 
.A(n_609),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_549),
.Y(n_643)
);

INVx8_ASAP7_75t_L g644 ( 
.A(n_467),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_504),
.B(n_432),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_546),
.B(n_224),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_525),
.B(n_438),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_491),
.A2(n_248),
.B1(n_234),
.B2(n_236),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_476),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_549),
.B(n_438),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_499),
.B(n_438),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_499),
.B(n_438),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_499),
.B(n_438),
.Y(n_653)
);

NOR2x1p5_ASAP7_75t_L g654 ( 
.A(n_483),
.B(n_178),
.Y(n_654)
);

OR2x6_ASAP7_75t_L g655 ( 
.A(n_538),
.B(n_373),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_478),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_499),
.B(n_437),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_546),
.B(n_224),
.Y(n_658)
);

NAND2xp33_ASAP7_75t_L g659 ( 
.A(n_541),
.B(n_277),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_486),
.B(n_437),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_478),
.Y(n_661)
);

AOI22xp5_ASAP7_75t_L g662 ( 
.A1(n_507),
.A2(n_467),
.B1(n_596),
.B2(n_530),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_486),
.B(n_437),
.Y(n_663)
);

O2A1O1Ixp33_ASAP7_75t_L g664 ( 
.A1(n_488),
.A2(n_462),
.B(n_448),
.C(n_452),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_546),
.B(n_481),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_586),
.B(n_373),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_498),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_481),
.B(n_547),
.Y(n_668)
);

OAI22xp5_ASAP7_75t_L g669 ( 
.A1(n_553),
.A2(n_234),
.B1(n_295),
.B2(n_303),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_512),
.B(n_446),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_574),
.B(n_270),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_498),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_481),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_512),
.B(n_446),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_578),
.B(n_446),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_502),
.Y(n_676)
);

BUFx5_ASAP7_75t_L g677 ( 
.A(n_505),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_502),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_588),
.Y(n_679)
);

NOR2xp67_ASAP7_75t_L g680 ( 
.A(n_585),
.B(n_448),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_513),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_481),
.B(n_224),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_513),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_583),
.B(n_446),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_522),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_547),
.B(n_446),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_588),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_574),
.B(n_224),
.Y(n_688)
);

OAI22xp5_ASAP7_75t_L g689 ( 
.A1(n_561),
.A2(n_303),
.B1(n_295),
.B2(n_306),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_491),
.B(n_224),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_609),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_L g692 ( 
.A(n_527),
.B(n_278),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_522),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_529),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g695 ( 
.A1(n_467),
.A2(n_315),
.B1(n_307),
.B2(n_304),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_538),
.Y(n_696)
);

BUFx5_ASAP7_75t_L g697 ( 
.A(n_508),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_482),
.B(n_446),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_491),
.B(n_284),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_598),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_561),
.B(n_179),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_L g703 ( 
.A(n_468),
.B(n_193),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_510),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_482),
.B(n_446),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_482),
.B(n_446),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_510),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_482),
.B(n_449),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_492),
.B(n_500),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_492),
.B(n_297),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_567),
.B(n_391),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_540),
.B(n_204),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_SL g713 ( 
.A(n_492),
.B(n_449),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_571),
.B(n_212),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_529),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_615),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_535),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_500),
.B(n_449),
.Y(n_718)
);

INVxp67_ASAP7_75t_SL g719 ( 
.A(n_616),
.Y(n_719)
);

AOI22xp5_ASAP7_75t_L g720 ( 
.A1(n_485),
.A2(n_342),
.B1(n_306),
.B2(n_249),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_511),
.Y(n_721)
);

NAND3xp33_ASAP7_75t_L g722 ( 
.A(n_605),
.B(n_601),
.C(n_566),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_500),
.B(n_449),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_500),
.B(n_449),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_511),
.B(n_449),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_516),
.B(n_449),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_567),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_516),
.B(n_449),
.Y(n_728)
);

O2A1O1Ixp33_ASAP7_75t_L g729 ( 
.A1(n_488),
.A2(n_518),
.B(n_519),
.C(n_517),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_517),
.B(n_453),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_518),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_598),
.B(n_453),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_531),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_531),
.B(n_453),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_542),
.B(n_453),
.Y(n_735)
);

NAND2xp5_ASAP7_75t_L g736 ( 
.A(n_542),
.B(n_453),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_551),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_551),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_SL g739 ( 
.A(n_598),
.B(n_612),
.Y(n_739)
);

CKINVDCx11_ASAP7_75t_R g740 ( 
.A(n_475),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_562),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_598),
.B(n_453),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_612),
.B(n_453),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_562),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_563),
.B(n_456),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_615),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_612),
.B(n_456),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_581),
.Y(n_748)
);

INVxp67_ASAP7_75t_SL g749 ( 
.A(n_616),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_612),
.B(n_456),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_581),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_SL g752 ( 
.A(n_483),
.B(n_201),
.Y(n_752)
);

INVxp33_ASAP7_75t_SL g753 ( 
.A(n_493),
.Y(n_753)
);

AOI22xp5_ASAP7_75t_L g754 ( 
.A1(n_485),
.A2(n_493),
.B1(n_579),
.B2(n_593),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_535),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_584),
.Y(n_756)
);

NOR3xp33_ASAP7_75t_L g757 ( 
.A(n_587),
.B(n_391),
.C(n_283),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_584),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_589),
.Y(n_759)
);

AND2x4_ASAP7_75t_L g760 ( 
.A(n_589),
.B(n_450),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_591),
.Y(n_761)
);

NOR3xp33_ASAP7_75t_L g762 ( 
.A(n_532),
.B(n_230),
.C(n_220),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_591),
.B(n_456),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_475),
.B(n_225),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_475),
.B(n_227),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_526),
.B(n_450),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_521),
.B(n_456),
.Y(n_767)
);

AO22x2_ASAP7_75t_L g768 ( 
.A1(n_526),
.A2(n_236),
.B1(n_249),
.B2(n_253),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_592),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_572),
.B(n_452),
.Y(n_770)
);

AOI22xp33_ASAP7_75t_L g771 ( 
.A1(n_602),
.A2(n_253),
.B1(n_311),
.B2(n_281),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_592),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_537),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_556),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_599),
.B(n_456),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_475),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_599),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_521),
.B(n_456),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_521),
.B(n_272),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_539),
.Y(n_780)
);

NOR2xp67_ASAP7_75t_L g781 ( 
.A(n_603),
.B(n_462),
.Y(n_781)
);

INVx2_ASAP7_75t_SL g782 ( 
.A(n_572),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_604),
.B(n_311),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_616),
.Y(n_784)
);

AOI221xp5_ASAP7_75t_L g785 ( 
.A1(n_524),
.A2(n_209),
.B1(n_299),
.B2(n_310),
.C(n_305),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_537),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_559),
.B(n_383),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_648),
.B(n_607),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_648),
.B(n_572),
.Y(n_789)
);

BUFx2_ASAP7_75t_L g790 ( 
.A(n_696),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_624),
.B(n_466),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_624),
.B(n_572),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_624),
.B(n_572),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_624),
.Y(n_794)
);

CKINVDCx11_ASAP7_75t_R g795 ( 
.A(n_740),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_624),
.B(n_528),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_679),
.B(n_559),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_619),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_634),
.B(n_611),
.Y(n_799)
);

AOI22xp5_ASAP7_75t_L g800 ( 
.A1(n_709),
.A2(n_573),
.B1(n_595),
.B2(n_515),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_619),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_634),
.B(n_533),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_633),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_671),
.B(n_550),
.C(n_555),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_671),
.B(n_523),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_713),
.A2(n_552),
.B(n_544),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_713),
.A2(n_552),
.B(n_544),
.Y(n_807)
);

A2O1A1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_729),
.A2(n_565),
.B(n_582),
.C(n_576),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_633),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_649),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_640),
.B(n_233),
.Y(n_811)
);

OAI22xp33_ASAP7_75t_L g812 ( 
.A1(n_687),
.A2(n_722),
.B1(n_752),
.B2(n_770),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_688),
.A2(n_479),
.B(n_466),
.C(n_473),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_661),
.Y(n_814)
);

BUFx8_ASAP7_75t_L g815 ( 
.A(n_774),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_677),
.B(n_469),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_661),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_643),
.Y(n_818)
);

OA21x2_ASAP7_75t_L g819 ( 
.A1(n_690),
.A2(n_497),
.B(n_479),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_677),
.Y(n_820)
);

AOI21xp5_ASAP7_75t_L g821 ( 
.A1(n_709),
.A2(n_684),
.B(n_675),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_677),
.B(n_469),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_677),
.B(n_484),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_677),
.B(n_473),
.Y(n_824)
);

BUFx4f_ASAP7_75t_L g825 ( 
.A(n_644),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_690),
.A2(n_503),
.B(n_497),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_SL g827 ( 
.A(n_753),
.B(n_342),
.Y(n_827)
);

AO21x1_ASAP7_75t_L g828 ( 
.A1(n_699),
.A2(n_503),
.B(n_477),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_668),
.A2(n_501),
.B(n_536),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_637),
.B(n_240),
.Y(n_830)
);

OAI22xp5_ASAP7_75t_L g831 ( 
.A1(n_639),
.A2(n_628),
.B1(n_631),
.B2(n_630),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_668),
.A2(n_501),
.B(n_536),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_632),
.A2(n_602),
.B1(n_474),
.B2(n_477),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_629),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_677),
.B(n_484),
.Y(n_835)
);

CKINVDCx20_ASAP7_75t_R g836 ( 
.A(n_780),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_656),
.Y(n_837)
);

AOI21xp5_ASAP7_75t_L g838 ( 
.A1(n_657),
.A2(n_536),
.B(n_544),
.Y(n_838)
);

AOI21xp5_ASAP7_75t_L g839 ( 
.A1(n_645),
.A2(n_501),
.B(n_552),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_635),
.A2(n_602),
.B1(n_474),
.B2(n_608),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_647),
.A2(n_490),
.B(n_496),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_666),
.B(n_602),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_697),
.B(n_484),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_660),
.A2(n_490),
.B(n_496),
.Y(n_844)
);

HB1xp67_ASAP7_75t_L g845 ( 
.A(n_727),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_667),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_663),
.A2(n_490),
.B(n_496),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_672),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_699),
.A2(n_595),
.B1(n_610),
.B2(n_608),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_697),
.B(n_534),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_697),
.B(n_534),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_655),
.Y(n_852)
);

AOI21xp5_ASAP7_75t_L g853 ( 
.A1(n_670),
.A2(n_496),
.B(n_520),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_676),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_674),
.A2(n_496),
.B(n_520),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_697),
.B(n_534),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_625),
.A2(n_520),
.B(n_570),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_665),
.A2(n_520),
.B(n_570),
.Y(n_858)
);

CKINVDCx8_ASAP7_75t_R g859 ( 
.A(n_655),
.Y(n_859)
);

BUFx4f_ASAP7_75t_L g860 ( 
.A(n_644),
.Y(n_860)
);

O2A1O1Ixp33_ASAP7_75t_L g861 ( 
.A1(n_688),
.A2(n_689),
.B(n_710),
.C(n_664),
.Y(n_861)
);

INVx3_ASAP7_75t_L g862 ( 
.A(n_643),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_623),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_665),
.A2(n_520),
.B(n_570),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_637),
.B(n_246),
.Y(n_865)
);

OAI21xp5_ASAP7_75t_L g866 ( 
.A1(n_710),
.A2(n_577),
.B(n_610),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_686),
.A2(n_705),
.B(n_698),
.Y(n_867)
);

BUFx3_ASAP7_75t_L g868 ( 
.A(n_644),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_697),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_697),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_678),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_702),
.B(n_247),
.Y(n_872)
);

AO21x1_ASAP7_75t_L g873 ( 
.A1(n_779),
.A2(n_613),
.B(n_606),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_721),
.B(n_577),
.Y(n_874)
);

AO21x1_ASAP7_75t_L g875 ( 
.A1(n_703),
.A2(n_613),
.B(n_606),
.Y(n_875)
);

OAI21x1_ASAP7_75t_L g876 ( 
.A1(n_706),
.A2(n_577),
.B(n_575),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_702),
.B(n_257),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_776),
.B(n_261),
.Y(n_878)
);

NOR2xp67_ASAP7_75t_L g879 ( 
.A(n_662),
.B(n_543),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_731),
.B(n_543),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_733),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_738),
.B(n_545),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_764),
.B(n_265),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_771),
.A2(n_595),
.B1(n_597),
.B2(n_266),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_741),
.B(n_545),
.Y(n_885)
);

OAI21xp33_ASAP7_75t_L g886 ( 
.A1(n_711),
.A2(n_274),
.B(n_279),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_744),
.B(n_548),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_748),
.B(n_548),
.Y(n_888)
);

INVx3_ASAP7_75t_L g889 ( 
.A(n_643),
.Y(n_889)
);

OAI21x1_ASAP7_75t_L g890 ( 
.A1(n_708),
.A2(n_600),
.B(n_560),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_733),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_718),
.A2(n_600),
.B(n_560),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_620),
.A2(n_594),
.B(n_590),
.Y(n_893)
);

AOI22xp33_ASAP7_75t_L g894 ( 
.A1(n_771),
.A2(n_595),
.B1(n_597),
.B2(n_280),
.Y(n_894)
);

INVx3_ASAP7_75t_L g895 ( 
.A(n_643),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_737),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_751),
.B(n_564),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_769),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_655),
.B(n_383),
.Y(n_899)
);

OAI21xp5_ASAP7_75t_L g900 ( 
.A1(n_622),
.A2(n_594),
.B(n_590),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_723),
.A2(n_564),
.B(n_575),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_756),
.B(n_595),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_769),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_651),
.A2(n_472),
.B(n_400),
.Y(n_904)
);

AOI21xp33_ASAP7_75t_L g905 ( 
.A1(n_703),
.A2(n_282),
.B(n_289),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_764),
.B(n_291),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_758),
.B(n_595),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_787),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_772),
.Y(n_909)
);

INVxp67_ASAP7_75t_L g910 ( 
.A(n_766),
.Y(n_910)
);

NOR2xp33_ASAP7_75t_L g911 ( 
.A(n_765),
.B(n_294),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_759),
.B(n_595),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_652),
.A2(n_472),
.B(n_394),
.Y(n_913)
);

HB1xp67_ASAP7_75t_L g914 ( 
.A(n_617),
.Y(n_914)
);

AOI22xp5_ASAP7_75t_L g915 ( 
.A1(n_781),
.A2(n_342),
.B1(n_597),
.B2(n_454),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_761),
.B(n_568),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_772),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_777),
.B(n_568),
.Y(n_918)
);

INVxp67_ASAP7_75t_SL g919 ( 
.A(n_673),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_653),
.A2(n_472),
.B(n_394),
.Y(n_920)
);

NOR2xp33_ASAP7_75t_L g921 ( 
.A(n_765),
.B(n_296),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_701),
.A2(n_707),
.B(n_704),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_701),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_704),
.B(n_568),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_760),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_707),
.Y(n_926)
);

BUFx2_ASAP7_75t_L g927 ( 
.A(n_636),
.Y(n_927)
);

A2O1A1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_712),
.A2(n_393),
.B(n_385),
.C(n_312),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_760),
.B(n_783),
.Y(n_929)
);

OAI321xp33_ASAP7_75t_L g930 ( 
.A1(n_669),
.A2(n_393),
.A3(n_385),
.B1(n_465),
.B2(n_441),
.C(n_461),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_650),
.A2(n_472),
.B(n_400),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_680),
.B(n_298),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_621),
.Y(n_933)
);

AOI22xp5_ASAP7_75t_L g934 ( 
.A1(n_618),
.A2(n_342),
.B1(n_597),
.B2(n_435),
.Y(n_934)
);

AOI21xp5_ASAP7_75t_L g935 ( 
.A1(n_724),
.A2(n_472),
.B(n_400),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_754),
.B(n_300),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_719),
.B(n_568),
.Y(n_937)
);

BUFx6f_ASAP7_75t_L g938 ( 
.A(n_673),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_724),
.A2(n_472),
.B(n_400),
.Y(n_939)
);

AOI22xp5_ASAP7_75t_L g940 ( 
.A1(n_627),
.A2(n_597),
.B1(n_465),
.B2(n_461),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_749),
.B(n_435),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_767),
.A2(n_400),
.B(n_418),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_767),
.A2(n_418),
.B(n_394),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_712),
.B(n_313),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_642),
.B(n_421),
.Y(n_945)
);

OAI22xp5_ASAP7_75t_L g946 ( 
.A1(n_782),
.A2(n_314),
.B1(n_317),
.B2(n_454),
.Y(n_946)
);

HB1xp67_ASAP7_75t_L g947 ( 
.A(n_700),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_673),
.B(n_441),
.Y(n_948)
);

AO21x2_ASAP7_75t_L g949 ( 
.A1(n_778),
.A2(n_442),
.B(n_461),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_714),
.B(n_441),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_778),
.A2(n_394),
.B(n_418),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_714),
.B(n_673),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_691),
.B(n_421),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_626),
.A2(n_418),
.B(n_454),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_700),
.B(n_739),
.Y(n_955)
);

AOI21x1_ASAP7_75t_L g956 ( 
.A1(n_732),
.A2(n_444),
.B(n_442),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_785),
.B(n_421),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_626),
.A2(n_418),
.B(n_444),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_739),
.B(n_8),
.Y(n_959)
);

OAI321xp33_ASAP7_75t_L g960 ( 
.A1(n_720),
.A2(n_435),
.A3(n_444),
.B1(n_15),
.B2(n_18),
.C(n_20),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_784),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_786),
.B(n_597),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_641),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_636),
.B(n_681),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_683),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_775),
.B(n_597),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_725),
.B(n_70),
.Y(n_967)
);

OAI21xp5_ASAP7_75t_L g968 ( 
.A1(n_682),
.A2(n_68),
.B(n_152),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_646),
.A2(n_66),
.B(n_150),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_646),
.A2(n_63),
.B(n_147),
.Y(n_970)
);

INVx3_ASAP7_75t_L g971 ( 
.A(n_685),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_658),
.A2(n_62),
.B(n_136),
.Y(n_972)
);

CKINVDCx10_ASAP7_75t_R g973 ( 
.A(n_654),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_693),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_762),
.A2(n_757),
.B(n_716),
.C(n_746),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_694),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_803),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_803),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_805),
.B(n_636),
.Y(n_979)
);

INVx3_ASAP7_75t_L g980 ( 
.A(n_938),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_872),
.Y(n_981)
);

AOI221x1_ASAP7_75t_L g982 ( 
.A1(n_928),
.A2(n_768),
.B1(n_734),
.B2(n_763),
.C(n_726),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_872),
.B(n_768),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_877),
.B(n_695),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_877),
.A2(n_692),
.B1(n_638),
.B2(n_659),
.Y(n_985)
);

BUFx3_ASAP7_75t_L g986 ( 
.A(n_790),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_821),
.A2(n_658),
.B(n_742),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_928),
.A2(n_682),
.B(n_728),
.C(n_730),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_836),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_SL g990 ( 
.A(n_799),
.B(n_743),
.Y(n_990)
);

BUFx6f_ASAP7_75t_L g991 ( 
.A(n_938),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_795),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_830),
.B(n_743),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_830),
.B(n_742),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_883),
.A2(n_750),
.B(n_747),
.C(n_735),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_865),
.B(n_750),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_865),
.B(n_747),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_883),
.B(n_736),
.Y(n_998)
);

NOR2xp33_ASAP7_75t_SL g999 ( 
.A(n_825),
.B(n_745),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_799),
.B(n_773),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_906),
.B(n_715),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_868),
.Y(n_1002)
);

INVx2_ASAP7_75t_SL g1003 ( 
.A(n_845),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_798),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_906),
.B(n_768),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_794),
.A2(n_755),
.B(n_717),
.Y(n_1006)
);

OR2x6_ASAP7_75t_L g1007 ( 
.A(n_868),
.B(n_153),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_789),
.A2(n_135),
.B1(n_133),
.B2(n_124),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_911),
.B(n_12),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_911),
.B(n_12),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_921),
.A2(n_121),
.B1(n_120),
.B2(n_117),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_801),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_809),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_921),
.B(n_14),
.Y(n_1014)
);

NOR2xp33_ASAP7_75t_L g1015 ( 
.A(n_845),
.B(n_14),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_788),
.A2(n_796),
.B1(n_793),
.B2(n_792),
.Y(n_1016)
);

HB1xp67_ASAP7_75t_L g1017 ( 
.A(n_899),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_896),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_815),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_852),
.B(n_104),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_898),
.Y(n_1021)
);

BUFx12f_ASAP7_75t_L g1022 ( 
.A(n_815),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_973),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_810),
.Y(n_1024)
);

O2A1O1Ixp33_ASAP7_75t_L g1025 ( 
.A1(n_812),
.A2(n_15),
.B(n_23),
.C(n_24),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_816),
.A2(n_103),
.B(n_102),
.Y(n_1026)
);

AOI21xp33_ASAP7_75t_L g1027 ( 
.A1(n_936),
.A2(n_34),
.B(n_40),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_938),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_925),
.B(n_98),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_802),
.B(n_40),
.Y(n_1030)
);

A2O1A1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_802),
.A2(n_42),
.B(n_43),
.C(n_44),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_822),
.A2(n_94),
.B(n_92),
.Y(n_1032)
);

OAI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_861),
.A2(n_88),
.B(n_72),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_929),
.B(n_47),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_797),
.Y(n_1035)
);

BUFx2_ASAP7_75t_L g1036 ( 
.A(n_908),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_925),
.B(n_48),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_814),
.Y(n_1038)
);

BUFx12f_ASAP7_75t_L g1039 ( 
.A(n_797),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_823),
.A2(n_49),
.B(n_50),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_SL g1041 ( 
.A(n_812),
.B(n_49),
.Y(n_1041)
);

O2A1O1Ixp33_ASAP7_75t_L g1042 ( 
.A1(n_960),
.A2(n_50),
.B(n_51),
.C(n_53),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_835),
.A2(n_850),
.B(n_843),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_856),
.A2(n_53),
.B(n_54),
.Y(n_1044)
);

NOR2xp33_ASAP7_75t_L g1045 ( 
.A(n_863),
.B(n_57),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_817),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_820),
.A2(n_869),
.B1(n_870),
.B2(n_800),
.Y(n_1047)
);

OR2x6_ASAP7_75t_L g1048 ( 
.A(n_938),
.B(n_57),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_944),
.B(n_957),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_903),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_818),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_905),
.A2(n_964),
.B(n_959),
.C(n_975),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_825),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_841),
.A2(n_839),
.B(n_831),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_820),
.A2(n_869),
.B1(n_870),
.B2(n_804),
.Y(n_1055)
);

AOI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_806),
.A2(n_807),
.B(n_867),
.Y(n_1056)
);

CKINVDCx8_ASAP7_75t_R g1057 ( 
.A(n_945),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_903),
.Y(n_1058)
);

O2A1O1Ixp5_ASAP7_75t_L g1059 ( 
.A1(n_875),
.A2(n_873),
.B(n_828),
.C(n_826),
.Y(n_1059)
);

INVx2_ASAP7_75t_SL g1060 ( 
.A(n_945),
.Y(n_1060)
);

AOI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_936),
.A2(n_932),
.B1(n_811),
.B2(n_910),
.Y(n_1061)
);

AOI21xp5_ASAP7_75t_L g1062 ( 
.A1(n_844),
.A2(n_847),
.B(n_829),
.Y(n_1062)
);

A2O1A1Ixp33_ASAP7_75t_L g1063 ( 
.A1(n_959),
.A2(n_811),
.B(n_808),
.C(n_848),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_975),
.A2(n_833),
.B(n_840),
.C(n_950),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_818),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_860),
.Y(n_1066)
);

CKINVDCx20_ASAP7_75t_R g1067 ( 
.A(n_860),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_808),
.A2(n_837),
.B(n_846),
.C(n_854),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_834),
.A2(n_871),
.B1(n_955),
.B2(n_919),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_842),
.B(n_917),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_832),
.A2(n_851),
.B(n_922),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_851),
.A2(n_853),
.B(n_855),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_923),
.A2(n_926),
.B1(n_881),
.B2(n_909),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_SL g1074 ( 
.A(n_947),
.B(n_878),
.Y(n_1074)
);

NAND3xp33_ASAP7_75t_L g1075 ( 
.A(n_878),
.B(n_886),
.C(n_946),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_838),
.A2(n_791),
.B(n_824),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_914),
.B(n_927),
.Y(n_1077)
);

O2A1O1Ixp5_ASAP7_75t_L g1078 ( 
.A1(n_967),
.A2(n_866),
.B(n_948),
.C(n_900),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_862),
.Y(n_1079)
);

INVx2_ASAP7_75t_SL g1080 ( 
.A(n_953),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_914),
.B(n_947),
.Y(n_1081)
);

AND2x2_ASAP7_75t_L g1082 ( 
.A(n_953),
.B(n_859),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_862),
.Y(n_1083)
);

NAND2x1_ASAP7_75t_L g1084 ( 
.A(n_923),
.B(n_926),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_L g1085 ( 
.A(n_891),
.B(n_889),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_827),
.B(n_961),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_879),
.B(n_889),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_895),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_967),
.A2(n_885),
.B(n_897),
.C(n_880),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_895),
.A2(n_974),
.B1(n_963),
.B2(n_965),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_933),
.Y(n_1091)
);

OAI21xp33_ASAP7_75t_L g1092 ( 
.A1(n_884),
.A2(n_894),
.B(n_968),
.Y(n_1092)
);

BUFx2_ASAP7_75t_L g1093 ( 
.A(n_971),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_971),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_941),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_791),
.A2(n_824),
.B(n_857),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_L g1097 ( 
.A(n_976),
.B(n_888),
.Y(n_1097)
);

INVx4_ASAP7_75t_L g1098 ( 
.A(n_976),
.Y(n_1098)
);

AND2x4_ASAP7_75t_L g1099 ( 
.A(n_948),
.B(n_887),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_SL g1100 ( 
.A(n_969),
.B(n_972),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_882),
.A2(n_930),
.B(n_874),
.C(n_912),
.Y(n_1101)
);

NOR3xp33_ASAP7_75t_SL g1102 ( 
.A(n_902),
.B(n_907),
.C(n_918),
.Y(n_1102)
);

NOR3xp33_ASAP7_75t_SL g1103 ( 
.A(n_916),
.B(n_966),
.C(n_970),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_937),
.A2(n_924),
.B(n_864),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_SL g1105 ( 
.A(n_884),
.B(n_894),
.Y(n_1105)
);

AND2x2_ASAP7_75t_L g1106 ( 
.A(n_819),
.B(n_949),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_915),
.B(n_849),
.Y(n_1107)
);

O2A1O1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_966),
.A2(n_813),
.B(n_893),
.C(n_962),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_819),
.B(n_956),
.Y(n_1109)
);

NAND2xp5_ASAP7_75t_L g1110 ( 
.A(n_892),
.B(n_901),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_949),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_819),
.B(n_858),
.Y(n_1112)
);

AND2x2_ASAP7_75t_L g1113 ( 
.A(n_940),
.B(n_934),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_890),
.Y(n_1114)
);

AND2x2_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_951),
.Y(n_1115)
);

O2A1O1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_954),
.A2(n_958),
.B(n_943),
.C(n_931),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_904),
.A2(n_913),
.B(n_920),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_876),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_935),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_939),
.Y(n_1120)
);

A2O1A1Ixp33_ASAP7_75t_L g1121 ( 
.A1(n_805),
.A2(n_872),
.B(n_877),
.C(n_883),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_805),
.A2(n_928),
.B(n_812),
.C(n_406),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1104),
.A2(n_1062),
.B(n_1072),
.Y(n_1123)
);

CKINVDCx5p33_ASAP7_75t_R g1124 ( 
.A(n_989),
.Y(n_1124)
);

AO21x1_ASAP7_75t_L g1125 ( 
.A1(n_981),
.A2(n_994),
.B(n_993),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_SL g1126 ( 
.A1(n_1121),
.A2(n_1092),
.B(n_1105),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1071),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_977),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1004),
.Y(n_1129)
);

BUFx3_ASAP7_75t_L g1130 ( 
.A(n_986),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_993),
.B(n_994),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1066),
.B(n_1053),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_1012),
.Y(n_1133)
);

CKINVDCx8_ASAP7_75t_R g1134 ( 
.A(n_1023),
.Y(n_1134)
);

OAI21x1_ASAP7_75t_L g1135 ( 
.A1(n_1096),
.A2(n_1076),
.B(n_1117),
.Y(n_1135)
);

HB1xp67_ASAP7_75t_L g1136 ( 
.A(n_1003),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_1118),
.A2(n_1033),
.B(n_1112),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_992),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1063),
.A2(n_1122),
.B(n_1064),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_996),
.B(n_997),
.Y(n_1140)
);

O2A1O1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1009),
.A2(n_1010),
.B(n_1014),
.C(n_1030),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_978),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_996),
.B(n_997),
.Y(n_1143)
);

CKINVDCx5p33_ASAP7_75t_R g1144 ( 
.A(n_1022),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1013),
.Y(n_1145)
);

OR2x6_ASAP7_75t_L g1146 ( 
.A(n_1007),
.B(n_1066),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1043),
.A2(n_1116),
.B(n_987),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1095),
.A2(n_1107),
.B(n_1110),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1116),
.A2(n_1114),
.B(n_1055),
.Y(n_1149)
);

NOR2xp67_ASAP7_75t_SL g1150 ( 
.A(n_1057),
.B(n_1019),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1041),
.A2(n_990),
.B(n_984),
.C(n_1122),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1095),
.A2(n_1089),
.B(n_998),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1002),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_1017),
.B(n_1030),
.Y(n_1154)
);

O2A1O1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_984),
.A2(n_1049),
.B(n_1027),
.C(n_1005),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1089),
.A2(n_998),
.B(n_1016),
.Y(n_1156)
);

AOI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_995),
.A2(n_1100),
.B(n_985),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1001),
.A2(n_1078),
.B(n_1108),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_982),
.A2(n_1109),
.A3(n_1111),
.B(n_1047),
.Y(n_1159)
);

CKINVDCx11_ASAP7_75t_R g1160 ( 
.A(n_1067),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1001),
.A2(n_1078),
.B(n_1108),
.Y(n_1161)
);

AOI21xp5_ASAP7_75t_L g1162 ( 
.A1(n_1064),
.A2(n_1101),
.B(n_988),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1073),
.A2(n_1069),
.A3(n_979),
.B(n_983),
.Y(n_1163)
);

AND2x4_ASAP7_75t_L g1164 ( 
.A(n_1060),
.B(n_1080),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1031),
.A2(n_1045),
.B(n_1025),
.C(n_1052),
.Y(n_1165)
);

BUFx4f_ASAP7_75t_L g1166 ( 
.A(n_1035),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1024),
.Y(n_1167)
);

OAI22xp5_ASAP7_75t_L g1168 ( 
.A1(n_1042),
.A2(n_1061),
.B1(n_1048),
.B2(n_1075),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1059),
.A2(n_1106),
.B(n_1120),
.Y(n_1169)
);

OA21x2_ASAP7_75t_L g1170 ( 
.A1(n_1119),
.A2(n_1006),
.B(n_1102),
.Y(n_1170)
);

NOR2xp33_ASAP7_75t_SL g1171 ( 
.A(n_1042),
.B(n_1048),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_1025),
.A2(n_1052),
.B(n_1074),
.C(n_1037),
.Y(n_1172)
);

NAND3x1_ASAP7_75t_L g1173 ( 
.A(n_1082),
.B(n_1086),
.C(n_1015),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1101),
.A2(n_988),
.B(n_1097),
.Y(n_1174)
);

AOI21x1_ASAP7_75t_L g1175 ( 
.A1(n_1000),
.A2(n_1087),
.B(n_1113),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1070),
.B(n_1068),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1008),
.A2(n_1098),
.A3(n_1040),
.B(n_1044),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1115),
.A2(n_1068),
.B(n_1099),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1099),
.A2(n_999),
.B(n_1084),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1085),
.A2(n_1029),
.B(n_1034),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_1058),
.B(n_1018),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1103),
.A2(n_1102),
.B(n_1032),
.Y(n_1182)
);

AOI21xp33_ASAP7_75t_L g1183 ( 
.A1(n_1077),
.A2(n_1017),
.B(n_1046),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1021),
.B(n_1050),
.Y(n_1184)
);

AO32x2_ASAP7_75t_L g1185 ( 
.A1(n_1098),
.A2(n_1079),
.A3(n_1028),
.B1(n_1103),
.B2(n_1077),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_1039),
.Y(n_1186)
);

BUFx10_ASAP7_75t_L g1187 ( 
.A(n_1081),
.Y(n_1187)
);

AOI21xp33_ASAP7_75t_L g1188 ( 
.A1(n_1038),
.A2(n_1011),
.B(n_1048),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1026),
.A2(n_1051),
.B(n_1065),
.Y(n_1189)
);

OAI22xp5_ASAP7_75t_L g1190 ( 
.A1(n_1007),
.A2(n_1020),
.B1(n_1090),
.B2(n_1088),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_1091),
.A2(n_1094),
.B(n_1093),
.C(n_1083),
.Y(n_1191)
);

INVx2_ASAP7_75t_L g1192 ( 
.A(n_1083),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1051),
.A2(n_1065),
.B(n_1079),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_980),
.A2(n_1007),
.B(n_1028),
.Y(n_1194)
);

INVx2_ASAP7_75t_SL g1195 ( 
.A(n_1036),
.Y(n_1195)
);

INVx6_ASAP7_75t_SL g1196 ( 
.A(n_1020),
.Y(n_1196)
);

AO31x2_ASAP7_75t_L g1197 ( 
.A1(n_980),
.A2(n_991),
.A3(n_1020),
.B(n_1065),
.Y(n_1197)
);

INVx3_ASAP7_75t_L g1198 ( 
.A(n_1065),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_991),
.B(n_981),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_991),
.A2(n_1121),
.B(n_981),
.C(n_906),
.Y(n_1200)
);

INVx2_ASAP7_75t_SL g1201 ( 
.A(n_991),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_986),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1203)
);

AOI21x1_ASAP7_75t_SL g1204 ( 
.A1(n_1009),
.A2(n_1014),
.B(n_1010),
.Y(n_1204)
);

BUFx10_ASAP7_75t_L g1205 ( 
.A(n_1015),
.Y(n_1205)
);

O2A1O1Ixp33_ASAP7_75t_SL g1206 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1105),
.C(n_1063),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1208)
);

BUFx6f_ASAP7_75t_L g1209 ( 
.A(n_991),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1210)
);

OAI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_SL g1212 ( 
.A1(n_1121),
.A2(n_1092),
.B(n_673),
.Y(n_1212)
);

OR2x6_ASAP7_75t_L g1213 ( 
.A(n_1007),
.B(n_644),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1121),
.A2(n_984),
.B(n_981),
.C(n_993),
.Y(n_1214)
);

OAI22x1_ASAP7_75t_L g1215 ( 
.A1(n_1030),
.A2(n_984),
.B1(n_1061),
.B2(n_1041),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_986),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1121),
.B(n_1061),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1121),
.A2(n_1054),
.B(n_1056),
.Y(n_1219)
);

AOI21x1_ASAP7_75t_L g1220 ( 
.A1(n_1107),
.A2(n_952),
.B(n_990),
.Y(n_1220)
);

BUFx12f_ASAP7_75t_L g1221 ( 
.A(n_992),
.Y(n_1221)
);

OAI21x1_ASAP7_75t_L g1222 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1224)
);

INVx4_ASAP7_75t_SL g1225 ( 
.A(n_991),
.Y(n_1225)
);

OAI22x1_ASAP7_75t_L g1226 ( 
.A1(n_1030),
.A2(n_984),
.B1(n_1061),
.B2(n_1041),
.Y(n_1226)
);

NOR4xp25_ASAP7_75t_L g1227 ( 
.A(n_1121),
.B(n_981),
.C(n_1025),
.D(n_1122),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1228)
);

INVx2_ASAP7_75t_SL g1229 ( 
.A(n_986),
.Y(n_1229)
);

OAI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1063),
.Y(n_1230)
);

AND2x2_ASAP7_75t_L g1231 ( 
.A(n_1017),
.B(n_640),
.Y(n_1231)
);

BUFx10_ASAP7_75t_L g1232 ( 
.A(n_1015),
.Y(n_1232)
);

OA21x2_ASAP7_75t_L g1233 ( 
.A1(n_1059),
.A2(n_1078),
.B(n_875),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_986),
.Y(n_1234)
);

O2A1O1Ixp33_ASAP7_75t_SL g1235 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1105),
.C(n_1063),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_977),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1059),
.A2(n_1078),
.B(n_875),
.Y(n_1237)
);

AO22x2_ASAP7_75t_L g1238 ( 
.A1(n_981),
.A2(n_1041),
.B1(n_982),
.B2(n_1105),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_1121),
.A2(n_1054),
.B(n_1056),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1056),
.A2(n_952),
.B(n_1054),
.Y(n_1241)
);

INVx1_ASAP7_75t_SL g1242 ( 
.A(n_986),
.Y(n_1242)
);

NOR2x1_ASAP7_75t_L g1243 ( 
.A(n_989),
.B(n_1066),
.Y(n_1243)
);

O2A1O1Ixp33_ASAP7_75t_L g1244 ( 
.A1(n_1121),
.A2(n_981),
.B(n_906),
.C(n_911),
.Y(n_1244)
);

BUFx8_ASAP7_75t_SL g1245 ( 
.A(n_989),
.Y(n_1245)
);

BUFx6f_ASAP7_75t_L g1246 ( 
.A(n_991),
.Y(n_1246)
);

INVx4_ASAP7_75t_L g1247 ( 
.A(n_1065),
.Y(n_1247)
);

A2O1A1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1121),
.A2(n_984),
.B(n_981),
.C(n_993),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1121),
.A2(n_981),
.B(n_906),
.C(n_911),
.Y(n_1249)
);

OA21x2_ASAP7_75t_L g1250 ( 
.A1(n_1059),
.A2(n_1078),
.B(n_875),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_981),
.B(n_1121),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_982),
.A2(n_875),
.A3(n_873),
.B(n_828),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1105),
.C(n_1063),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1007),
.B(n_644),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1004),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_986),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1121),
.A2(n_981),
.B(n_906),
.C(n_911),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1004),
.Y(n_1258)
);

AO31x2_ASAP7_75t_L g1259 ( 
.A1(n_982),
.A2(n_875),
.A3(n_873),
.B(n_828),
.Y(n_1259)
);

OAI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1063),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1261)
);

BUFx2_ASAP7_75t_L g1262 ( 
.A(n_986),
.Y(n_1262)
);

AOI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1107),
.A2(n_952),
.B(n_990),
.Y(n_1263)
);

AO32x2_ASAP7_75t_L g1264 ( 
.A1(n_1016),
.A2(n_1069),
.A3(n_1055),
.B1(n_1047),
.B2(n_833),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1121),
.A2(n_1092),
.B(n_673),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1104),
.A2(n_890),
.B(n_876),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1121),
.A2(n_984),
.B(n_981),
.C(n_993),
.Y(n_1267)
);

AO31x2_ASAP7_75t_L g1268 ( 
.A1(n_982),
.A2(n_875),
.A3(n_873),
.B(n_828),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1121),
.A2(n_981),
.B(n_1063),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_992),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1214),
.A2(n_1248),
.B1(n_1267),
.B2(n_1140),
.Y(n_1271)
);

INVx6_ASAP7_75t_L g1272 ( 
.A(n_1247),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_1217),
.B2(n_1168),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1168),
.A2(n_1171),
.B1(n_1131),
.B2(n_1140),
.Y(n_1274)
);

BUFx4f_ASAP7_75t_SL g1275 ( 
.A(n_1221),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1129),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1133),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1171),
.A2(n_1131),
.B1(n_1143),
.B2(n_1269),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1130),
.Y(n_1279)
);

BUFx2_ASAP7_75t_L g1280 ( 
.A(n_1202),
.Y(n_1280)
);

BUFx8_ASAP7_75t_SL g1281 ( 
.A(n_1245),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1160),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1143),
.A2(n_1269),
.B1(n_1230),
.B2(n_1260),
.Y(n_1283)
);

BUFx4f_ASAP7_75t_SL g1284 ( 
.A(n_1270),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1145),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1230),
.A2(n_1260),
.B1(n_1251),
.B2(n_1139),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1251),
.A2(n_1139),
.B1(n_1125),
.B2(n_1238),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1167),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1238),
.A2(n_1188),
.B1(n_1154),
.B2(n_1190),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1244),
.A2(n_1249),
.B1(n_1257),
.B2(n_1173),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1247),
.Y(n_1291)
);

BUFx2_ASAP7_75t_SL g1292 ( 
.A(n_1153),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1188),
.A2(n_1190),
.B1(n_1157),
.B2(n_1232),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1205),
.A2(n_1232),
.B1(n_1199),
.B2(n_1146),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_SL g1295 ( 
.A1(n_1205),
.A2(n_1187),
.B1(n_1254),
.B2(n_1213),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1146),
.A2(n_1231),
.B1(n_1196),
.B2(n_1183),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1155),
.B(n_1141),
.Y(n_1297)
);

AND2x2_ASAP7_75t_L g1298 ( 
.A(n_1227),
.B(n_1142),
.Y(n_1298)
);

CKINVDCx6p67_ASAP7_75t_R g1299 ( 
.A(n_1213),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_SL g1300 ( 
.A1(n_1187),
.A2(n_1254),
.B1(n_1213),
.B2(n_1146),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1227),
.B(n_1195),
.Y(n_1301)
);

CKINVDCx11_ASAP7_75t_R g1302 ( 
.A(n_1134),
.Y(n_1302)
);

AOI22x1_ASAP7_75t_L g1303 ( 
.A1(n_1156),
.A2(n_1174),
.B1(n_1152),
.B2(n_1162),
.Y(n_1303)
);

OAI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1254),
.A2(n_1196),
.B1(n_1242),
.B2(n_1234),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_SL g1305 ( 
.A1(n_1182),
.A2(n_1194),
.B1(n_1165),
.B2(n_1166),
.Y(n_1305)
);

BUFx12f_ASAP7_75t_L g1306 ( 
.A(n_1138),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1183),
.A2(n_1243),
.B1(n_1182),
.B2(n_1164),
.Y(n_1307)
);

BUFx12f_ASAP7_75t_L g1308 ( 
.A(n_1124),
.Y(n_1308)
);

INVx6_ASAP7_75t_L g1309 ( 
.A(n_1225),
.Y(n_1309)
);

INVx1_ASAP7_75t_L g1310 ( 
.A(n_1255),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1151),
.B(n_1200),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1164),
.A2(n_1178),
.B1(n_1176),
.B2(n_1194),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1144),
.Y(n_1313)
);

CKINVDCx11_ASAP7_75t_R g1314 ( 
.A(n_1234),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1258),
.Y(n_1315)
);

BUFx8_ASAP7_75t_L g1316 ( 
.A(n_1216),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1209),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1186),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1176),
.A2(n_1158),
.B1(n_1161),
.B2(n_1262),
.Y(n_1319)
);

BUFx8_ASAP7_75t_L g1320 ( 
.A(n_1132),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_1166),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1136),
.A2(n_1180),
.B1(n_1150),
.B2(n_1242),
.Y(n_1322)
);

OAI21xp5_ASAP7_75t_L g1323 ( 
.A1(n_1126),
.A2(n_1148),
.B(n_1172),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1209),
.Y(n_1324)
);

CKINVDCx20_ASAP7_75t_R g1325 ( 
.A(n_1256),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1256),
.A2(n_1137),
.B1(n_1239),
.B2(n_1219),
.Y(n_1326)
);

AOI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1132),
.A2(n_1235),
.B1(n_1206),
.B2(n_1253),
.Y(n_1327)
);

AOI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1137),
.A2(n_1219),
.B1(n_1239),
.B2(n_1179),
.Y(n_1328)
);

INVx4_ASAP7_75t_L g1329 ( 
.A(n_1225),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1229),
.A2(n_1265),
.B1(n_1212),
.B2(n_1198),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1236),
.A2(n_1192),
.B1(n_1170),
.B2(n_1169),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1170),
.A2(n_1169),
.B1(n_1181),
.B2(n_1198),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1225),
.Y(n_1333)
);

BUFx8_ASAP7_75t_L g1334 ( 
.A(n_1209),
.Y(n_1334)
);

BUFx10_ASAP7_75t_L g1335 ( 
.A(n_1246),
.Y(n_1335)
);

AOI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1181),
.A2(n_1233),
.B1(n_1237),
.B2(n_1250),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1233),
.A2(n_1237),
.B1(n_1250),
.B2(n_1184),
.Y(n_1337)
);

AOI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1191),
.A2(n_1189),
.B1(n_1201),
.B2(n_1184),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1175),
.A2(n_1220),
.B1(n_1263),
.B2(n_1193),
.Y(n_1339)
);

BUFx2_ASAP7_75t_SL g1340 ( 
.A(n_1246),
.Y(n_1340)
);

BUFx10_ASAP7_75t_L g1341 ( 
.A(n_1204),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1197),
.Y(n_1342)
);

INVxp67_ASAP7_75t_SL g1343 ( 
.A(n_1149),
.Y(n_1343)
);

INVx3_ASAP7_75t_L g1344 ( 
.A(n_1197),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1203),
.A2(n_1241),
.B1(n_1208),
.B2(n_1228),
.Y(n_1345)
);

AOI22xp33_ASAP7_75t_L g1346 ( 
.A1(n_1207),
.A2(n_1240),
.B1(n_1147),
.B2(n_1127),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1135),
.A2(n_1123),
.B1(n_1222),
.B2(n_1223),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1210),
.A2(n_1224),
.B1(n_1261),
.B2(n_1266),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1185),
.Y(n_1349)
);

INVx1_ASAP7_75t_SL g1350 ( 
.A(n_1185),
.Y(n_1350)
);

CKINVDCx6p67_ASAP7_75t_R g1351 ( 
.A(n_1177),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1163),
.Y(n_1352)
);

AOI22xp33_ASAP7_75t_SL g1353 ( 
.A1(n_1264),
.A2(n_1177),
.B1(n_1218),
.B2(n_1211),
.Y(n_1353)
);

BUFx4_ASAP7_75t_SL g1354 ( 
.A(n_1163),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1177),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1264),
.A2(n_1159),
.B1(n_1252),
.B2(n_1259),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_1159),
.Y(n_1357)
);

CKINVDCx5p33_ASAP7_75t_R g1358 ( 
.A(n_1264),
.Y(n_1358)
);

AOI22xp5_ASAP7_75t_L g1359 ( 
.A1(n_1252),
.A2(n_984),
.B1(n_981),
.B2(n_872),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1252),
.A2(n_1215),
.B1(n_1226),
.B2(n_984),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1259),
.A2(n_1215),
.B1(n_1226),
.B2(n_984),
.Y(n_1361)
);

BUFx12f_ASAP7_75t_L g1362 ( 
.A(n_1259),
.Y(n_1362)
);

BUFx3_ASAP7_75t_L g1363 ( 
.A(n_1268),
.Y(n_1363)
);

OAI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1268),
.A2(n_1121),
.B(n_981),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1268),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1129),
.Y(n_1366)
);

AND2x2_ASAP7_75t_L g1367 ( 
.A(n_1154),
.B(n_1214),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1129),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1128),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1131),
.B(n_981),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1372)
);

CKINVDCx20_ASAP7_75t_R g1373 ( 
.A(n_1245),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1129),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_SL g1375 ( 
.A1(n_1171),
.A2(n_984),
.B1(n_981),
.B2(n_752),
.Y(n_1375)
);

INVx6_ASAP7_75t_L g1376 ( 
.A(n_1247),
.Y(n_1376)
);

BUFx6f_ASAP7_75t_L g1377 ( 
.A(n_1209),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_L g1378 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1171),
.A2(n_981),
.B1(n_752),
.B2(n_863),
.Y(n_1379)
);

AOI22xp33_ASAP7_75t_L g1380 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1225),
.Y(n_1381)
);

BUFx12f_ASAP7_75t_L g1382 ( 
.A(n_1160),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1130),
.Y(n_1384)
);

BUFx3_ASAP7_75t_L g1385 ( 
.A(n_1130),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1131),
.B(n_981),
.Y(n_1386)
);

BUFx8_ASAP7_75t_L g1387 ( 
.A(n_1221),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1129),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_SL g1389 ( 
.A1(n_1171),
.A2(n_984),
.B1(n_981),
.B2(n_752),
.Y(n_1389)
);

BUFx6f_ASAP7_75t_L g1390 ( 
.A(n_1209),
.Y(n_1390)
);

INVx1_ASAP7_75t_SL g1391 ( 
.A(n_1234),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_1146),
.Y(n_1392)
);

INVx6_ASAP7_75t_L g1393 ( 
.A(n_1247),
.Y(n_1393)
);

INVx3_ASAP7_75t_SL g1394 ( 
.A(n_1124),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1234),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1129),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1245),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1215),
.A2(n_1226),
.B1(n_984),
.B2(n_981),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_1202),
.Y(n_1400)
);

OA21x2_ASAP7_75t_L g1401 ( 
.A1(n_1303),
.A2(n_1323),
.B(n_1364),
.Y(n_1401)
);

INVxp67_ASAP7_75t_L g1402 ( 
.A(n_1280),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1365),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1370),
.B(n_1386),
.Y(n_1404)
);

INVxp67_ASAP7_75t_L g1405 ( 
.A(n_1400),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1375),
.B(n_1389),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_SL g1407 ( 
.A1(n_1290),
.A2(n_1271),
.B1(n_1358),
.B2(n_1297),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1363),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1392),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1363),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1362),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1362),
.Y(n_1412)
);

OAI211xp5_ASAP7_75t_L g1413 ( 
.A1(n_1371),
.A2(n_1399),
.B(n_1372),
.C(n_1395),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1298),
.B(n_1367),
.Y(n_1414)
);

HB1xp67_ASAP7_75t_L g1415 ( 
.A(n_1276),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_1344),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1344),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1352),
.Y(n_1418)
);

OAI21x1_ASAP7_75t_L g1419 ( 
.A1(n_1348),
.A2(n_1347),
.B(n_1346),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1344),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1367),
.B(n_1378),
.Y(n_1421)
);

INVxp33_ASAP7_75t_L g1422 ( 
.A(n_1314),
.Y(n_1422)
);

INVx2_ASAP7_75t_L g1423 ( 
.A(n_1342),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1357),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1287),
.B(n_1358),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1357),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1351),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1301),
.B(n_1350),
.Y(n_1428)
);

INVxp67_ASAP7_75t_SL g1429 ( 
.A(n_1311),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1360),
.B(n_1361),
.Y(n_1430)
);

NAND2xp33_ASAP7_75t_R g1431 ( 
.A(n_1321),
.B(n_1313),
.Y(n_1431)
);

BUFx4f_ASAP7_75t_SL g1432 ( 
.A(n_1382),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1277),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1345),
.A2(n_1328),
.B(n_1339),
.Y(n_1434)
);

CKINVDCx12_ASAP7_75t_R g1435 ( 
.A(n_1302),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1326),
.A2(n_1343),
.B(n_1331),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1355),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1354),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1285),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1288),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1310),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1315),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1379),
.B(n_1325),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1366),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1349),
.Y(n_1445)
);

INVx2_ASAP7_75t_L g1446 ( 
.A(n_1368),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1374),
.Y(n_1447)
);

INVx1_ASAP7_75t_SL g1448 ( 
.A(n_1391),
.Y(n_1448)
);

INVx2_ASAP7_75t_SL g1449 ( 
.A(n_1392),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1388),
.Y(n_1450)
);

INVx4_ASAP7_75t_L g1451 ( 
.A(n_1329),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1337),
.A2(n_1332),
.B(n_1336),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1359),
.A2(n_1327),
.B1(n_1299),
.B2(n_1396),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1397),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1356),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1380),
.B(n_1383),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1319),
.B(n_1283),
.Y(n_1457)
);

INVxp33_ASAP7_75t_L g1458 ( 
.A(n_1314),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1312),
.B(n_1369),
.Y(n_1459)
);

AOI22xp33_ASAP7_75t_SL g1460 ( 
.A1(n_1349),
.A2(n_1325),
.B1(n_1316),
.B2(n_1382),
.Y(n_1460)
);

AOI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1273),
.A2(n_1305),
.B1(n_1274),
.B2(n_1286),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1341),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1281),
.Y(n_1463)
);

OR2x6_ASAP7_75t_L g1464 ( 
.A(n_1329),
.B(n_1381),
.Y(n_1464)
);

INVx6_ASAP7_75t_L g1465 ( 
.A(n_1320),
.Y(n_1465)
);

INVx4_ASAP7_75t_L g1466 ( 
.A(n_1381),
.Y(n_1466)
);

BUFx3_ASAP7_75t_L g1467 ( 
.A(n_1320),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1338),
.A2(n_1293),
.B(n_1278),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1289),
.A2(n_1296),
.B1(n_1307),
.B2(n_1322),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1330),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1317),
.B(n_1324),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1300),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1294),
.B(n_1304),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1295),
.A2(n_1334),
.B(n_1309),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1414),
.B(n_1394),
.Y(n_1476)
);

OR2x2_ASAP7_75t_L g1477 ( 
.A(n_1428),
.B(n_1394),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1429),
.B(n_1390),
.Y(n_1478)
);

AND2x4_ASAP7_75t_L g1479 ( 
.A(n_1411),
.B(n_1384),
.Y(n_1479)
);

OR2x2_ASAP7_75t_L g1480 ( 
.A(n_1445),
.B(n_1415),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1445),
.B(n_1385),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1433),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1447),
.B(n_1292),
.Y(n_1483)
);

AND2x4_ASAP7_75t_L g1484 ( 
.A(n_1412),
.B(n_1279),
.Y(n_1484)
);

OA21x2_ASAP7_75t_L g1485 ( 
.A1(n_1434),
.A2(n_1321),
.B(n_1335),
.Y(n_1485)
);

AO32x2_ASAP7_75t_L g1486 ( 
.A1(n_1449),
.A2(n_1390),
.A3(n_1377),
.B1(n_1335),
.B2(n_1340),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1473),
.B(n_1385),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1473),
.B(n_1384),
.Y(n_1488)
);

NOR2x1_ASAP7_75t_SL g1489 ( 
.A(n_1464),
.B(n_1308),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1441),
.B(n_1272),
.Y(n_1490)
);

AND2x4_ASAP7_75t_L g1491 ( 
.A(n_1409),
.B(n_1279),
.Y(n_1491)
);

OA21x2_ASAP7_75t_L g1492 ( 
.A1(n_1434),
.A2(n_1335),
.B(n_1313),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_1463),
.Y(n_1493)
);

O2A1O1Ixp33_ASAP7_75t_SL g1494 ( 
.A1(n_1453),
.A2(n_1398),
.B(n_1373),
.C(n_1282),
.Y(n_1494)
);

AOI221xp5_ASAP7_75t_L g1495 ( 
.A1(n_1461),
.A2(n_1282),
.B1(n_1373),
.B2(n_1398),
.C(n_1318),
.Y(n_1495)
);

A2O1A1Ixp33_ASAP7_75t_L g1496 ( 
.A1(n_1468),
.A2(n_1443),
.B(n_1413),
.C(n_1407),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1406),
.A2(n_1469),
.B1(n_1460),
.B2(n_1456),
.Y(n_1497)
);

OR2x2_ASAP7_75t_L g1498 ( 
.A(n_1441),
.B(n_1308),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1475),
.B(n_1309),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1425),
.B(n_1474),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_L g1501 ( 
.A(n_1474),
.B(n_1318),
.Y(n_1501)
);

A2O1A1Ixp33_ASAP7_75t_SL g1502 ( 
.A1(n_1462),
.A2(n_1393),
.B(n_1291),
.C(n_1376),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1439),
.Y(n_1503)
);

AOI22xp5_ASAP7_75t_L g1504 ( 
.A1(n_1457),
.A2(n_1387),
.B1(n_1302),
.B2(n_1284),
.Y(n_1504)
);

BUFx6f_ASAP7_75t_L g1505 ( 
.A(n_1467),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1446),
.B(n_1281),
.Y(n_1506)
);

NOR2xp33_ASAP7_75t_L g1507 ( 
.A(n_1421),
.B(n_1291),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1446),
.B(n_1306),
.Y(n_1508)
);

AOI22xp33_ASAP7_75t_L g1509 ( 
.A1(n_1457),
.A2(n_1387),
.B1(n_1306),
.B2(n_1275),
.Y(n_1509)
);

INVx4_ASAP7_75t_SL g1510 ( 
.A(n_1465),
.Y(n_1510)
);

A2O1A1Ixp33_ASAP7_75t_L g1511 ( 
.A1(n_1468),
.A2(n_1333),
.B(n_1471),
.C(n_1430),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1439),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1401),
.A2(n_1471),
.B(n_1436),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1450),
.B(n_1454),
.Y(n_1514)
);

NAND3xp33_ASAP7_75t_L g1515 ( 
.A(n_1401),
.B(n_1404),
.C(n_1402),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1405),
.B(n_1459),
.Y(n_1516)
);

OAI21x1_ASAP7_75t_L g1517 ( 
.A1(n_1419),
.A2(n_1436),
.B(n_1452),
.Y(n_1517)
);

A2O1A1Ixp33_ASAP7_75t_L g1518 ( 
.A1(n_1475),
.A2(n_1467),
.B(n_1438),
.C(n_1470),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1472),
.B(n_1454),
.Y(n_1519)
);

OR2x2_ASAP7_75t_L g1520 ( 
.A(n_1454),
.B(n_1440),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1467),
.A2(n_1438),
.B(n_1470),
.C(n_1452),
.Y(n_1521)
);

AOI22xp5_ASAP7_75t_L g1522 ( 
.A1(n_1459),
.A2(n_1401),
.B1(n_1448),
.B2(n_1435),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1435),
.A2(n_1422),
.B1(n_1458),
.B2(n_1432),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1503),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1512),
.Y(n_1525)
);

AND2x4_ASAP7_75t_SL g1526 ( 
.A(n_1499),
.B(n_1464),
.Y(n_1526)
);

AOI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1497),
.A2(n_1401),
.B1(n_1459),
.B2(n_1465),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1514),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1493),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1513),
.B(n_1517),
.Y(n_1530)
);

INVx6_ASAP7_75t_L g1531 ( 
.A(n_1510),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1482),
.B(n_1455),
.Y(n_1532)
);

OAI22xp5_ASAP7_75t_L g1533 ( 
.A1(n_1496),
.A2(n_1465),
.B1(n_1464),
.B2(n_1459),
.Y(n_1533)
);

INVxp67_ASAP7_75t_L g1534 ( 
.A(n_1515),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1519),
.B(n_1423),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1513),
.B(n_1424),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1515),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1520),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1480),
.B(n_1418),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1490),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1522),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1522),
.B(n_1417),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1490),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1485),
.B(n_1416),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1477),
.B(n_1418),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1499),
.B(n_1427),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1485),
.B(n_1417),
.Y(n_1547)
);

AND2x2_ASAP7_75t_L g1548 ( 
.A(n_1492),
.B(n_1417),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1497),
.A2(n_1465),
.B1(n_1464),
.B2(n_1442),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1516),
.B(n_1442),
.Y(n_1550)
);

INVx2_ASAP7_75t_L g1551 ( 
.A(n_1486),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1500),
.B(n_1444),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1478),
.Y(n_1553)
);

BUFx12f_ASAP7_75t_L g1554 ( 
.A(n_1505),
.Y(n_1554)
);

OR2x2_ASAP7_75t_L g1555 ( 
.A(n_1551),
.B(n_1521),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1553),
.B(n_1437),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1544),
.Y(n_1557)
);

OR2x2_ASAP7_75t_L g1558 ( 
.A(n_1551),
.B(n_1426),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1536),
.B(n_1408),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1546),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1524),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1534),
.B(n_1537),
.Y(n_1562)
);

INVx3_ASAP7_75t_L g1563 ( 
.A(n_1547),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1547),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_SL g1565 ( 
.A(n_1533),
.B(n_1511),
.Y(n_1565)
);

NAND4xp25_ASAP7_75t_SL g1566 ( 
.A(n_1527),
.B(n_1495),
.C(n_1504),
.D(n_1509),
.Y(n_1566)
);

AND2x2_ASAP7_75t_SL g1567 ( 
.A(n_1526),
.B(n_1501),
.Y(n_1567)
);

INVx3_ASAP7_75t_L g1568 ( 
.A(n_1547),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1534),
.B(n_1403),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1537),
.B(n_1403),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1410),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1541),
.B(n_1437),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1527),
.A2(n_1495),
.B(n_1504),
.Y(n_1573)
);

OR2x2_ASAP7_75t_L g1574 ( 
.A(n_1541),
.B(n_1410),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1548),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1524),
.Y(n_1576)
);

INVx4_ASAP7_75t_L g1577 ( 
.A(n_1531),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1530),
.B(n_1420),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1525),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1533),
.A2(n_1518),
.B(n_1494),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1542),
.B(n_1535),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1528),
.Y(n_1582)
);

OR2x6_ASAP7_75t_L g1583 ( 
.A(n_1549),
.B(n_1499),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1525),
.Y(n_1584)
);

BUFx3_ASAP7_75t_L g1585 ( 
.A(n_1531),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1542),
.B(n_1486),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1564),
.B(n_1542),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1561),
.Y(n_1588)
);

AOI22xp33_ASAP7_75t_L g1589 ( 
.A1(n_1566),
.A2(n_1549),
.B1(n_1507),
.B2(n_1523),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1540),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1557),
.Y(n_1591)
);

NAND4xp25_ASAP7_75t_L g1592 ( 
.A(n_1562),
.B(n_1509),
.C(n_1507),
.D(n_1487),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1561),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1562),
.B(n_1553),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1574),
.Y(n_1595)
);

INVx1_ASAP7_75t_SL g1596 ( 
.A(n_1555),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1561),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1576),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1576),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1576),
.Y(n_1600)
);

INVxp67_ASAP7_75t_SL g1601 ( 
.A(n_1562),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1555),
.B(n_1574),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1579),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1555),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1575),
.B(n_1540),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1575),
.B(n_1538),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1560),
.B(n_1526),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1575),
.B(n_1538),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1579),
.Y(n_1609)
);

OR2x2_ASAP7_75t_L g1610 ( 
.A(n_1555),
.B(n_1574),
.Y(n_1610)
);

OR2x2_ASAP7_75t_L g1611 ( 
.A(n_1574),
.B(n_1539),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1582),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1579),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1584),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1586),
.B(n_1538),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1569),
.B(n_1543),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1557),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1569),
.B(n_1543),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1580),
.B(n_1479),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1572),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1586),
.B(n_1535),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1586),
.B(n_1535),
.Y(n_1622)
);

INVx1_ASAP7_75t_L g1623 ( 
.A(n_1584),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1601),
.B(n_1594),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1621),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1596),
.B(n_1569),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1588),
.Y(n_1627)
);

AND2x2_ASAP7_75t_SL g1628 ( 
.A(n_1589),
.B(n_1565),
.Y(n_1628)
);

INVx1_ASAP7_75t_L g1629 ( 
.A(n_1588),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1593),
.Y(n_1630)
);

INVx4_ASAP7_75t_L g1631 ( 
.A(n_1607),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1601),
.B(n_1581),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1621),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1596),
.B(n_1570),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1593),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1607),
.B(n_1560),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1597),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

AO22x1_ASAP7_75t_L g1639 ( 
.A1(n_1604),
.A2(n_1580),
.B1(n_1577),
.B2(n_1585),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1607),
.B(n_1560),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_SL g1641 ( 
.A(n_1619),
.B(n_1565),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1621),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1594),
.B(n_1581),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1592),
.B(n_1581),
.Y(n_1644)
);

INVxp33_ASAP7_75t_L g1645 ( 
.A(n_1592),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1602),
.B(n_1570),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1616),
.B(n_1581),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1616),
.B(n_1559),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1607),
.B(n_1560),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1622),
.Y(n_1651)
);

OAI33xp33_ASAP7_75t_L g1652 ( 
.A1(n_1602),
.A2(n_1610),
.A3(n_1570),
.B1(n_1618),
.B2(n_1613),
.B3(n_1599),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1598),
.Y(n_1653)
);

OR2x2_ASAP7_75t_L g1654 ( 
.A(n_1610),
.B(n_1572),
.Y(n_1654)
);

AND2x4_ASAP7_75t_L g1655 ( 
.A(n_1607),
.B(n_1577),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1598),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_SL g1657 ( 
.A(n_1620),
.B(n_1565),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1599),
.Y(n_1658)
);

NAND2x1_ASAP7_75t_L g1659 ( 
.A(n_1587),
.B(n_1586),
.Y(n_1659)
);

OAI33xp33_ASAP7_75t_L g1660 ( 
.A1(n_1618),
.A2(n_1556),
.A3(n_1558),
.B1(n_1572),
.B2(n_1532),
.B3(n_1545),
.Y(n_1660)
);

OR2x2_ASAP7_75t_L g1661 ( 
.A(n_1611),
.B(n_1620),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1611),
.B(n_1572),
.Y(n_1662)
);

INVx2_ASAP7_75t_L g1663 ( 
.A(n_1622),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1622),
.B(n_1559),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1600),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1587),
.B(n_1559),
.Y(n_1666)
);

NAND3xp33_ASAP7_75t_L g1667 ( 
.A(n_1657),
.B(n_1573),
.C(n_1580),
.Y(n_1667)
);

OA211x2_ASAP7_75t_L g1668 ( 
.A1(n_1657),
.A2(n_1566),
.B(n_1556),
.C(n_1532),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1645),
.B(n_1587),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1645),
.B(n_1571),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1644),
.B(n_1552),
.Y(n_1671)
);

OR2x2_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1595),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1628),
.B(n_1571),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1646),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1552),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1631),
.B(n_1655),
.Y(n_1676)
);

NAND4xp75_ASAP7_75t_SL g1677 ( 
.A(n_1636),
.B(n_1571),
.C(n_1608),
.D(n_1606),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1628),
.B(n_1641),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1627),
.Y(n_1679)
);

NOR2xp33_ASAP7_75t_L g1680 ( 
.A(n_1641),
.B(n_1523),
.Y(n_1680)
);

NAND3xp33_ASAP7_75t_L g1681 ( 
.A(n_1639),
.B(n_1573),
.C(n_1612),
.Y(n_1681)
);

NAND2xp33_ASAP7_75t_L g1682 ( 
.A(n_1624),
.B(n_1529),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.B(n_1615),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1631),
.B(n_1615),
.Y(n_1684)
);

AND2x4_ASAP7_75t_L g1685 ( 
.A(n_1655),
.B(n_1577),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1629),
.Y(n_1686)
);

INVxp67_ASAP7_75t_L g1687 ( 
.A(n_1626),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1655),
.B(n_1615),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1647),
.B(n_1571),
.Y(n_1689)
);

AOI22xp33_ASAP7_75t_L g1690 ( 
.A1(n_1652),
.A2(n_1583),
.B1(n_1567),
.B2(n_1577),
.Y(n_1690)
);

OA21x2_ASAP7_75t_L g1691 ( 
.A1(n_1630),
.A2(n_1617),
.B(n_1591),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1635),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1647),
.B(n_1634),
.Y(n_1693)
);

INVx1_ASAP7_75t_SL g1694 ( 
.A(n_1636),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1643),
.B(n_1545),
.Y(n_1695)
);

INVx1_ASAP7_75t_SL g1696 ( 
.A(n_1640),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1640),
.B(n_1590),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1660),
.B(n_1506),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1637),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1634),
.B(n_1578),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1638),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1653),
.Y(n_1702)
);

AOI332xp33_ASAP7_75t_L g1703 ( 
.A1(n_1674),
.A2(n_1656),
.A3(n_1665),
.B1(n_1658),
.B2(n_1663),
.B3(n_1625),
.C1(n_1651),
.C2(n_1633),
.Y(n_1703)
);

OR2x2_ASAP7_75t_L g1704 ( 
.A(n_1669),
.B(n_1648),
.Y(n_1704)
);

OAI322xp33_ASAP7_75t_L g1705 ( 
.A1(n_1678),
.A2(n_1659),
.A3(n_1661),
.B1(n_1654),
.B2(n_1662),
.C1(n_1666),
.C2(n_1651),
.Y(n_1705)
);

OAI22xp5_ASAP7_75t_L g1706 ( 
.A1(n_1667),
.A2(n_1573),
.B1(n_1659),
.B2(n_1583),
.Y(n_1706)
);

OR2x2_ASAP7_75t_L g1707 ( 
.A(n_1673),
.B(n_1664),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1676),
.B(n_1650),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1678),
.B(n_1625),
.Y(n_1709)
);

INVxp67_ASAP7_75t_L g1710 ( 
.A(n_1680),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1676),
.B(n_1650),
.Y(n_1711)
);

AOI22xp33_ASAP7_75t_L g1712 ( 
.A1(n_1680),
.A2(n_1583),
.B1(n_1642),
.B2(n_1633),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1679),
.Y(n_1713)
);

AOI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1681),
.A2(n_1583),
.B1(n_1642),
.B2(n_1663),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1685),
.B(n_1585),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1690),
.A2(n_1661),
.B1(n_1654),
.B2(n_1585),
.C(n_1577),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1686),
.Y(n_1717)
);

OR2x2_ASAP7_75t_L g1718 ( 
.A(n_1670),
.B(n_1649),
.Y(n_1718)
);

OAI22xp33_ASAP7_75t_L g1719 ( 
.A1(n_1698),
.A2(n_1583),
.B1(n_1577),
.B2(n_1585),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1692),
.Y(n_1720)
);

AOI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1682),
.A2(n_1612),
.B(n_1489),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1699),
.Y(n_1722)
);

O2A1O1Ixp33_ASAP7_75t_L g1723 ( 
.A1(n_1682),
.A2(n_1502),
.B(n_1662),
.C(n_1508),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1701),
.Y(n_1724)
);

OAI322xp33_ASAP7_75t_L g1725 ( 
.A1(n_1698),
.A2(n_1591),
.A3(n_1617),
.B1(n_1558),
.B2(n_1613),
.C1(n_1609),
.C2(n_1600),
.Y(n_1725)
);

OR2x2_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1550),
.Y(n_1726)
);

AOI22xp5_ASAP7_75t_L g1727 ( 
.A1(n_1668),
.A2(n_1583),
.B1(n_1567),
.B2(n_1546),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1702),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1708),
.B(n_1685),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1713),
.Y(n_1730)
);

AND2x2_ASAP7_75t_L g1731 ( 
.A(n_1708),
.B(n_1685),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1711),
.B(n_1715),
.Y(n_1732)
);

OA21x2_ASAP7_75t_SL g1733 ( 
.A1(n_1703),
.A2(n_1696),
.B(n_1694),
.Y(n_1733)
);

NAND2x1_ASAP7_75t_SL g1734 ( 
.A(n_1717),
.B(n_1683),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1710),
.B(n_1687),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1720),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1714),
.B(n_1688),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1714),
.A2(n_1693),
.B1(n_1675),
.B2(n_1688),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1722),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1724),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1728),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1709),
.Y(n_1742)
);

INVxp67_ASAP7_75t_L g1743 ( 
.A(n_1710),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1704),
.Y(n_1744)
);

OAI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1712),
.A2(n_1716),
.B(n_1706),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1719),
.B(n_1683),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1729),
.B(n_1684),
.Y(n_1748)
);

OR2x2_ASAP7_75t_L g1749 ( 
.A(n_1735),
.B(n_1707),
.Y(n_1749)
);

AND2x2_ASAP7_75t_SL g1750 ( 
.A(n_1742),
.B(n_1431),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1743),
.B(n_1719),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1737),
.B(n_1732),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1741),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1741),
.Y(n_1754)
);

INVx2_ASAP7_75t_SL g1755 ( 
.A(n_1734),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1734),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1730),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1744),
.B(n_1705),
.Y(n_1758)
);

INVx1_ASAP7_75t_SL g1759 ( 
.A(n_1750),
.Y(n_1759)
);

NAND4xp75_ASAP7_75t_L g1760 ( 
.A(n_1755),
.B(n_1747),
.C(n_1737),
.D(n_1733),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1748),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_L g1762 ( 
.A(n_1758),
.B(n_1745),
.C(n_1746),
.D(n_1732),
.Y(n_1762)
);

NOR3xp33_ASAP7_75t_L g1763 ( 
.A(n_1751),
.B(n_1738),
.C(n_1736),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1750),
.B(n_1729),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_L g1765 ( 
.A(n_1758),
.B(n_1747),
.Y(n_1765)
);

AOI221xp5_ASAP7_75t_L g1766 ( 
.A1(n_1756),
.A2(n_1725),
.B1(n_1753),
.B2(n_1752),
.C(n_1757),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1749),
.B(n_1739),
.Y(n_1767)
);

AOI21xp33_ASAP7_75t_SL g1768 ( 
.A1(n_1765),
.A2(n_1753),
.B(n_1740),
.Y(n_1768)
);

OAI22xp5_ASAP7_75t_L g1769 ( 
.A1(n_1760),
.A2(n_1727),
.B1(n_1721),
.B2(n_1731),
.Y(n_1769)
);

AOI211xp5_ASAP7_75t_L g1770 ( 
.A1(n_1762),
.A2(n_1754),
.B(n_1731),
.C(n_1723),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1761),
.B(n_1759),
.Y(n_1771)
);

OAI222xp33_ASAP7_75t_L g1772 ( 
.A1(n_1764),
.A2(n_1672),
.B1(n_1718),
.B2(n_1697),
.C1(n_1700),
.C2(n_1726),
.Y(n_1772)
);

AOI32xp33_ASAP7_75t_L g1773 ( 
.A1(n_1769),
.A2(n_1763),
.A3(n_1766),
.B1(n_1767),
.B2(n_1697),
.Y(n_1773)
);

OAI311xp33_ASAP7_75t_L g1774 ( 
.A1(n_1771),
.A2(n_1770),
.A3(n_1768),
.B1(n_1772),
.C1(n_1672),
.Y(n_1774)
);

OAI22xp5_ASAP7_75t_L g1775 ( 
.A1(n_1769),
.A2(n_1689),
.B1(n_1695),
.B2(n_1531),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1768),
.B(n_1691),
.C(n_1488),
.Y(n_1776)
);

AOI21xp5_ASAP7_75t_L g1777 ( 
.A1(n_1769),
.A2(n_1691),
.B(n_1484),
.Y(n_1777)
);

AOI222xp33_ASAP7_75t_L g1778 ( 
.A1(n_1769),
.A2(n_1476),
.B1(n_1481),
.B2(n_1567),
.C1(n_1677),
.C2(n_1479),
.Y(n_1778)
);

NOR3xp33_ASAP7_75t_L g1779 ( 
.A(n_1773),
.B(n_1484),
.C(n_1498),
.Y(n_1779)
);

XOR2xp5_ASAP7_75t_L g1780 ( 
.A(n_1775),
.B(n_1505),
.Y(n_1780)
);

NOR4xp75_ASAP7_75t_L g1781 ( 
.A(n_1774),
.B(n_1563),
.C(n_1568),
.D(n_1606),
.Y(n_1781)
);

INVx1_ASAP7_75t_SL g1782 ( 
.A(n_1777),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_SL g1783 ( 
.A(n_1776),
.B(n_1505),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1782),
.A2(n_1778),
.B(n_1691),
.Y(n_1784)
);

NAND3x1_ASAP7_75t_L g1785 ( 
.A(n_1781),
.B(n_1568),
.C(n_1563),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_L g1786 ( 
.A(n_1779),
.B(n_1483),
.C(n_1466),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_SL g1787 ( 
.A1(n_1784),
.A2(n_1780),
.B1(n_1785),
.B2(n_1786),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1787),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1788),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1788),
.B(n_1783),
.Y(n_1790)
);

AOI22xp33_ASAP7_75t_L g1791 ( 
.A1(n_1789),
.A2(n_1554),
.B1(n_1617),
.B2(n_1591),
.Y(n_1791)
);

INVx1_ASAP7_75t_SL g1792 ( 
.A(n_1790),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1792),
.Y(n_1793)
);

AOI21x1_ASAP7_75t_L g1794 ( 
.A1(n_1791),
.A2(n_1623),
.B(n_1614),
.Y(n_1794)
);

NOR2x1p5_ASAP7_75t_L g1795 ( 
.A(n_1793),
.B(n_1451),
.Y(n_1795)
);

NOR2xp33_ASAP7_75t_L g1796 ( 
.A(n_1795),
.B(n_1794),
.Y(n_1796)
);

OAI22xp33_ASAP7_75t_L g1797 ( 
.A1(n_1796),
.A2(n_1623),
.B1(n_1614),
.B2(n_1609),
.Y(n_1797)
);

AOI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1797),
.A2(n_1603),
.B1(n_1568),
.B2(n_1563),
.C(n_1605),
.Y(n_1798)
);

AOI211xp5_ASAP7_75t_L g1799 ( 
.A1(n_1798),
.A2(n_1502),
.B(n_1491),
.C(n_1603),
.Y(n_1799)
);


endmodule