module fake_netlist_6_3881_n_1843 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1843);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1843;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_170;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_738;
wire n_189;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_527;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1775;
wire n_1773;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_1810;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_14),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_155),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_15),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_67),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_103),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_23),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_33),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g170 ( 
.A(n_39),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_64),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_27),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_18),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_140),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_73),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_100),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_36),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_26),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_153),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_61),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_59),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_60),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_18),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_90),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_84),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_54),
.Y(n_189)
);

INVx1_ASAP7_75t_SL g190 ( 
.A(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_62),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_16),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_15),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_109),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_127),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_97),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_56),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_12),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g200 ( 
.A(n_28),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_42),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_7),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_160),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_7),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_42),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_5),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_132),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

BUFx10_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_8),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_137),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_24),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_23),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_89),
.Y(n_215)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_145),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_88),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_71),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_83),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_117),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_111),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_27),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_11),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_151),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_134),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_6),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_65),
.Y(n_228)
);

BUFx8_ASAP7_75t_SL g229 ( 
.A(n_33),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_25),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_75),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_60),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_26),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_120),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_28),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_51),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_116),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_66),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_76),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_86),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_24),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_45),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_131),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_125),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_61),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_104),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g249 ( 
.A(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_154),
.Y(n_251)
);

INVxp67_ASAP7_75t_SL g252 ( 
.A(n_159),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_14),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_56),
.Y(n_254)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_130),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_152),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_114),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_22),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_148),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_53),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_85),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_95),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_133),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_2),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_135),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_105),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_118),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_74),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_79),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_59),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_30),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_6),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_139),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_150),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_41),
.Y(n_277)
);

BUFx10_ASAP7_75t_L g278 ( 
.A(n_62),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_77),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_46),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_91),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_47),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_41),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_136),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_107),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_80),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_10),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_0),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_82),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_110),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_50),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_146),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_19),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_93),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_34),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_115),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_53),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_144),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_63),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_124),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_113),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_141),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_149),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_99),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_162),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_147),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_21),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_98),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_13),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_32),
.Y(n_313)
);

BUFx10_ASAP7_75t_L g314 ( 
.A(n_161),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_30),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_57),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_101),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_72),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_35),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_20),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_87),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_39),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_12),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_40),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_157),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_17),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_11),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_106),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_32),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_229),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_200),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_200),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_249),
.B(n_1),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_221),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_208),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_212),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_215),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_311),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_217),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_220),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_225),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_226),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_228),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_200),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_255),
.B(n_266),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_200),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_237),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_200),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_200),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_200),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_251),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_200),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_168),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_163),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_168),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_216),
.Y(n_356)
);

INVxp67_ASAP7_75t_SL g357 ( 
.A(n_185),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_185),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_234),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_239),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_186),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_227),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_255),
.B(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_227),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_269),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_240),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_245),
.Y(n_367)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_186),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

INVxp67_ASAP7_75t_SL g370 ( 
.A(n_315),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_256),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_257),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_316),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_316),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_211),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_210),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_178),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_263),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_211),
.B(n_3),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_178),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_184),
.Y(n_381)
);

INVxp67_ASAP7_75t_SL g382 ( 
.A(n_165),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_184),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_264),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_267),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_L g386 ( 
.A(n_294),
.B(n_3),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_169),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_214),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_164),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_222),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_216),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_182),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_230),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_216),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_232),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_286),
.B(n_4),
.Y(n_396)
);

CKINVDCx16_ASAP7_75t_R g397 ( 
.A(n_210),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_233),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_191),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_192),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g401 ( 
.A(n_294),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_193),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_167),
.B(n_4),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_243),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_210),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_164),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_167),
.B(n_5),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_216),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_174),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_331),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_350),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_361),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g413 ( 
.A(n_333),
.B(n_194),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_331),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

INVx3_ASAP7_75t_L g416 ( 
.A(n_350),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_332),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_332),
.B(n_308),
.Y(n_418)
);

OA21x2_ASAP7_75t_L g419 ( 
.A1(n_407),
.A2(n_213),
.B(n_207),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_384),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_346),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_346),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

CKINVDCx6p67_ASAP7_75t_R g426 ( 
.A(n_338),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_348),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_349),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_349),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_377),
.B(n_308),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_345),
.B(n_363),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_377),
.B(n_194),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_352),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_356),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_356),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_356),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_391),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g440 ( 
.A(n_391),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

BUFx6f_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_387),
.Y(n_445)
);

BUFx3_ASAP7_75t_L g446 ( 
.A(n_407),
.Y(n_446)
);

AND2x6_ASAP7_75t_L g447 ( 
.A(n_333),
.B(n_219),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_408),
.Y(n_448)
);

INVx3_ASAP7_75t_L g449 ( 
.A(n_408),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_392),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_385),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_380),
.B(n_381),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_386),
.B(n_268),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_355),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_408),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_399),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_353),
.Y(n_459)
);

INVx4_ASAP7_75t_L g460 ( 
.A(n_335),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_355),
.B(n_219),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_380),
.B(n_241),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_400),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_353),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_354),
.B(n_190),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_358),
.Y(n_466)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_403),
.B(n_241),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_381),
.B(n_260),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_402),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_402),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_386),
.B(n_268),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_358),
.Y(n_473)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_362),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_396),
.B(n_260),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_362),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_364),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_364),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_369),
.Y(n_479)
);

OA21x2_ASAP7_75t_L g480 ( 
.A1(n_369),
.A2(n_236),
.B(n_235),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_376),
.B(n_268),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_373),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_373),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_357),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_379),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_421),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_415),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_439),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_415),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g490 ( 
.A(n_465),
.B(n_338),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_446),
.B(n_336),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_410),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g493 ( 
.A1(n_431),
.A2(n_204),
.B1(n_223),
.B2(n_179),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_415),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_415),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_431),
.B(n_337),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_465),
.B(n_339),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_446),
.B(n_357),
.Y(n_498)
);

BUFx3_ASAP7_75t_L g499 ( 
.A(n_418),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_421),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_411),
.Y(n_501)
);

BUFx8_ASAP7_75t_SL g502 ( 
.A(n_451),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_411),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_410),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_414),
.Y(n_505)
);

INVxp67_ASAP7_75t_SL g506 ( 
.A(n_484),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_411),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_412),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_439),
.Y(n_509)
);

BUFx2_ASAP7_75t_L g510 ( 
.A(n_412),
.Y(n_510)
);

INVx5_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_414),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_417),
.Y(n_513)
);

AND2x2_ASAP7_75t_SL g514 ( 
.A(n_485),
.B(n_270),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_446),
.B(n_340),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_417),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_418),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_446),
.A2(n_475),
.B1(n_485),
.B2(n_467),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_411),
.Y(n_519)
);

BUFx8_ASAP7_75t_SL g520 ( 
.A(n_451),
.Y(n_520)
);

AND2x6_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_270),
.Y(n_521)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_439),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_L g523 ( 
.A(n_475),
.B(n_341),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_411),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_475),
.A2(n_379),
.B1(n_382),
.B2(n_247),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_342),
.Y(n_526)
);

BUFx6f_ASAP7_75t_L g527 ( 
.A(n_439),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_420),
.Y(n_528)
);

INVx3_ASAP7_75t_L g529 ( 
.A(n_439),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_485),
.B(n_343),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_485),
.B(n_376),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_485),
.B(n_397),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_416),
.Y(n_533)
);

OAI22xp33_ASAP7_75t_L g534 ( 
.A1(n_456),
.A2(n_405),
.B1(n_397),
.B2(n_170),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_416),
.Y(n_535)
);

INVxp33_ASAP7_75t_L g536 ( 
.A(n_430),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_416),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_484),
.B(n_359),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_481),
.A2(n_261),
.B1(n_320),
.B2(n_258),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_416),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_416),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_435),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_435),
.Y(n_543)
);

XNOR2x1_ASAP7_75t_L g544 ( 
.A(n_467),
.B(n_163),
.Y(n_544)
);

AND2x4_ASAP7_75t_L g545 ( 
.A(n_418),
.B(n_461),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_435),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_419),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_460),
.B(n_405),
.Y(n_549)
);

CKINVDCx6p67_ASAP7_75t_R g550 ( 
.A(n_426),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_460),
.B(n_456),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g552 ( 
.A(n_419),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_484),
.B(n_360),
.Y(n_553)
);

CKINVDCx6p67_ASAP7_75t_R g554 ( 
.A(n_426),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_418),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_422),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g557 ( 
.A(n_430),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_475),
.B(n_366),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_460),
.B(n_367),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_435),
.Y(n_561)
);

OAI22x1_ASAP7_75t_L g562 ( 
.A1(n_481),
.A2(n_287),
.B1(n_283),
.B2(n_301),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_436),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_436),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_475),
.A2(n_447),
.B1(n_413),
.B2(n_461),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_426),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_423),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_460),
.B(n_371),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_436),
.Y(n_569)
);

AND2x6_ASAP7_75t_L g570 ( 
.A(n_418),
.B(n_325),
.Y(n_570)
);

INVxp67_ASAP7_75t_SL g571 ( 
.A(n_439),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_423),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_436),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_460),
.B(n_372),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_475),
.B(n_378),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_424),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_419),
.Y(n_577)
);

HB1xp67_ASAP7_75t_L g578 ( 
.A(n_430),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_424),
.Y(n_579)
);

INVx4_ASAP7_75t_L g580 ( 
.A(n_439),
.Y(n_580)
);

AO21x2_ASAP7_75t_L g581 ( 
.A1(n_427),
.A2(n_171),
.B(n_166),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_419),
.Y(n_582)
);

BUFx10_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_427),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_453),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_425),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_428),
.Y(n_587)
);

OAI22xp33_ASAP7_75t_L g588 ( 
.A1(n_472),
.A2(n_254),
.B1(n_253),
.B2(n_173),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_472),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_475),
.B(n_388),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_425),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_428),
.Y(n_592)
);

NAND2x1p5_ASAP7_75t_L g593 ( 
.A(n_419),
.B(n_175),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_461),
.B(n_390),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_439),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_475),
.A2(n_296),
.B1(n_271),
.B2(n_273),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_429),
.Y(n_597)
);

INVx1_ASAP7_75t_SL g598 ( 
.A(n_452),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_429),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_433),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_475),
.B(n_393),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_433),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_433),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_434),
.Y(n_604)
);

INVxp33_ASAP7_75t_SL g605 ( 
.A(n_452),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_475),
.B(n_395),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_461),
.B(n_398),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_434),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_434),
.Y(n_609)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_432),
.B(n_370),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_461),
.B(n_404),
.Y(n_611)
);

INVx4_ASAP7_75t_L g612 ( 
.A(n_440),
.Y(n_612)
);

INVx1_ASAP7_75t_SL g613 ( 
.A(n_452),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_425),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_432),
.B(n_389),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_425),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_449),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_440),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_480),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_419),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_480),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_449),
.Y(n_622)
);

INVx6_ASAP7_75t_L g623 ( 
.A(n_440),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_480),
.B(n_361),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_449),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_449),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_413),
.B(n_252),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_440),
.Y(n_628)
);

INVx4_ASAP7_75t_L g629 ( 
.A(n_440),
.Y(n_629)
);

AND2x6_ASAP7_75t_L g630 ( 
.A(n_432),
.B(n_325),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_444),
.B(n_406),
.Y(n_631)
);

INVx2_ASAP7_75t_SL g632 ( 
.A(n_480),
.Y(n_632)
);

INVx1_ASAP7_75t_SL g633 ( 
.A(n_462),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_449),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_SL g635 ( 
.A(n_462),
.B(n_409),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_457),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_496),
.B(n_413),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_538),
.B(n_413),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_545),
.Y(n_639)
);

NAND2x1p5_ASAP7_75t_L g640 ( 
.A(n_545),
.B(n_480),
.Y(n_640)
);

BUFx5_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_514),
.B(n_440),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_514),
.B(n_413),
.Y(n_643)
);

NOR3xp33_ASAP7_75t_L g644 ( 
.A(n_615),
.B(n_188),
.C(n_180),
.Y(n_644)
);

NAND2x1_ASAP7_75t_L g645 ( 
.A(n_545),
.B(n_413),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_545),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_514),
.B(n_413),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_557),
.B(n_375),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_498),
.B(n_447),
.Y(n_649)
);

OR2x6_ASAP7_75t_L g650 ( 
.A(n_508),
.B(n_383),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_536),
.B(n_375),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_524),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_498),
.B(n_447),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_518),
.B(n_440),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_553),
.B(n_174),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_506),
.B(n_447),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_499),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_499),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_551),
.A2(n_447),
.B1(n_334),
.B2(n_347),
.Y(n_659)
);

A2O1A1Ixp33_ASAP7_75t_L g660 ( 
.A1(n_624),
.A2(n_462),
.B(n_468),
.C(n_368),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_499),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_502),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_491),
.B(n_176),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_633),
.B(n_526),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_517),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_SL g666 ( 
.A(n_566),
.B(n_351),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_517),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_524),
.Y(n_668)
);

O2A1O1Ixp33_ASAP7_75t_L g669 ( 
.A1(n_624),
.A2(n_619),
.B(n_552),
.C(n_548),
.Y(n_669)
);

HB1xp67_ASAP7_75t_L g670 ( 
.A(n_578),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_565),
.B(n_530),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_520),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_517),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_515),
.B(n_447),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_555),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_544),
.A2(n_305),
.B1(n_250),
.B2(n_265),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_607),
.B(n_447),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_524),
.Y(n_678)
);

NOR2x1p5_ASAP7_75t_L g679 ( 
.A(n_550),
.B(n_330),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_492),
.B(n_447),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_585),
.B(n_440),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_492),
.B(n_447),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_590),
.B(n_442),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_555),
.B(n_444),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_601),
.B(n_442),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_504),
.B(n_480),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_504),
.B(n_505),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_605),
.B(n_176),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_505),
.B(n_442),
.Y(n_689)
);

BUFx3_ASAP7_75t_L g690 ( 
.A(n_555),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_497),
.B(n_177),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_535),
.Y(n_692)
);

AND2x2_ASAP7_75t_SL g693 ( 
.A(n_525),
.B(n_195),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_535),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_512),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_512),
.B(n_442),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_508),
.B(n_401),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_510),
.B(n_401),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_513),
.B(n_516),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_516),
.B(n_442),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_510),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_528),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_537),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_537),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_606),
.B(n_442),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_528),
.B(n_442),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_547),
.Y(n_707)
);

INVxp33_ASAP7_75t_L g708 ( 
.A(n_539),
.Y(n_708)
);

OAI22xp5_ASAP7_75t_L g709 ( 
.A1(n_551),
.A2(n_365),
.B1(n_281),
.B2(n_303),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_589),
.B(n_177),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_547),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_556),
.B(n_448),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_544),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_551),
.A2(n_468),
.B1(n_279),
.B2(n_289),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_556),
.B(n_448),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_560),
.B(n_448),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_537),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_560),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_511),
.B(n_448),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_511),
.B(n_448),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_567),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_567),
.B(n_448),
.Y(n_722)
);

INVx4_ASAP7_75t_L g723 ( 
.A(n_511),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_630),
.B(n_216),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_SL g725 ( 
.A(n_511),
.B(n_448),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_572),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_630),
.B(n_216),
.Y(n_727)
);

OAI21xp5_ASAP7_75t_L g728 ( 
.A1(n_621),
.A2(n_438),
.B(n_437),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_598),
.B(n_187),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_576),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_631),
.Y(n_731)
);

INVx4_ASAP7_75t_SL g732 ( 
.A(n_570),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_511),
.B(n_216),
.Y(n_733)
);

AND2x4_ASAP7_75t_L g734 ( 
.A(n_610),
.B(n_445),
.Y(n_734)
);

BUFx5_ASAP7_75t_L g735 ( 
.A(n_582),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_613),
.B(n_187),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_576),
.Y(n_737)
);

A2O1A1Ixp33_ASAP7_75t_L g738 ( 
.A1(n_582),
.A2(n_468),
.B(n_368),
.C(n_288),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_577),
.A2(n_298),
.B1(n_274),
.B2(n_272),
.Y(n_739)
);

AO221x1_ASAP7_75t_L g740 ( 
.A1(n_562),
.A2(n_312),
.B1(n_277),
.B2(n_280),
.C(n_282),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_540),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_511),
.B(n_216),
.Y(n_742)
);

AO22x2_ASAP7_75t_L g743 ( 
.A1(n_548),
.A2(n_324),
.B1(n_291),
.B2(n_313),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_579),
.B(n_457),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_579),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_SL g746 ( 
.A(n_577),
.B(n_203),
.Y(n_746)
);

OR2x6_ASAP7_75t_L g747 ( 
.A(n_635),
.B(n_531),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_584),
.B(n_457),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_584),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_587),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_532),
.B(n_197),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_587),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_594),
.B(n_611),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_540),
.Y(n_754)
);

NAND2xp33_ASAP7_75t_L g755 ( 
.A(n_630),
.B(n_197),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_592),
.B(n_457),
.Y(n_756)
);

NAND3xp33_ASAP7_75t_L g757 ( 
.A(n_596),
.B(n_383),
.C(n_276),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_592),
.B(n_474),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_550),
.Y(n_759)
);

AOI22xp33_ASAP7_75t_L g760 ( 
.A1(n_552),
.A2(n_327),
.B1(n_370),
.B2(n_374),
.Y(n_760)
);

NOR2xp67_ASAP7_75t_SL g761 ( 
.A(n_619),
.B(n_209),
.Y(n_761)
);

AND2x6_ASAP7_75t_L g762 ( 
.A(n_558),
.B(n_218),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_540),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_490),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_620),
.A2(n_632),
.B1(n_621),
.B2(n_593),
.Y(n_765)
);

AND2x4_ASAP7_75t_L g766 ( 
.A(n_597),
.B(n_445),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_597),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_575),
.B(n_620),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_599),
.B(n_474),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_599),
.B(n_474),
.Y(n_770)
);

INVx3_ASAP7_75t_L g771 ( 
.A(n_623),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_551),
.B(n_206),
.Y(n_772)
);

OAI22xp5_ASAP7_75t_L g773 ( 
.A1(n_632),
.A2(n_302),
.B1(n_275),
.B2(n_262),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_600),
.B(n_602),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_583),
.B(n_224),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_541),
.Y(n_776)
);

INVx2_ASAP7_75t_SL g777 ( 
.A(n_562),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_593),
.A2(n_238),
.B1(n_231),
.B2(n_244),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_541),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_523),
.A2(n_549),
.B1(n_559),
.B2(n_568),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_493),
.B(n_450),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_574),
.A2(n_630),
.B1(n_627),
.B2(n_570),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_600),
.B(n_602),
.Y(n_783)
);

BUFx2_ASAP7_75t_L g784 ( 
.A(n_486),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_493),
.B(n_450),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_630),
.B(n_206),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_603),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_603),
.B(n_474),
.Y(n_788)
);

BUFx6f_ASAP7_75t_L g789 ( 
.A(n_583),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_604),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_604),
.B(n_474),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_608),
.B(n_437),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_608),
.B(n_437),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_539),
.B(n_454),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_609),
.B(n_571),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_541),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_609),
.B(n_438),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_630),
.B(n_438),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_630),
.B(n_441),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_L g800 ( 
.A1(n_593),
.A2(n_246),
.B1(n_248),
.B2(n_285),
.Y(n_800)
);

OAI22xp5_ASAP7_75t_L g801 ( 
.A1(n_596),
.A2(n_317),
.B1(n_318),
.B2(n_328),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_667),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_641),
.B(n_735),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_728),
.A2(n_612),
.B(n_580),
.Y(n_804)
);

AOI21xp5_ASAP7_75t_L g805 ( 
.A1(n_768),
.A2(n_612),
.B(n_580),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_768),
.A2(n_612),
.B(n_580),
.Y(n_806)
);

OAI21xp5_ASAP7_75t_L g807 ( 
.A1(n_669),
.A2(n_614),
.B(n_591),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_787),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_731),
.B(n_534),
.Y(n_809)
);

NAND2xp33_ASAP7_75t_SL g810 ( 
.A(n_708),
.B(n_554),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_691),
.B(n_588),
.Y(n_811)
);

AOI21xp33_ASAP7_75t_L g812 ( 
.A1(n_691),
.A2(n_500),
.B(n_581),
.Y(n_812)
);

O2A1O1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_660),
.A2(n_614),
.B(n_581),
.C(n_591),
.Y(n_813)
);

BUFx6f_ASAP7_75t_L g814 ( 
.A(n_667),
.Y(n_814)
);

AOI21xp5_ASAP7_75t_L g815 ( 
.A1(n_654),
.A2(n_612),
.B(n_580),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_639),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_664),
.B(n_554),
.Y(n_817)
);

NAND2xp33_ASAP7_75t_SL g818 ( 
.A(n_781),
.B(n_276),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_654),
.A2(n_629),
.B(n_595),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_648),
.B(n_581),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_790),
.Y(n_821)
);

AOI222xp33_ASAP7_75t_L g822 ( 
.A1(n_713),
.A2(n_273),
.B1(n_271),
.B2(n_292),
.C1(n_300),
.C2(n_205),
.Y(n_822)
);

AOI21xp5_ASAP7_75t_L g823 ( 
.A1(n_683),
.A2(n_629),
.B(n_595),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_695),
.Y(n_824)
);

O2A1O1Ixp5_ASAP7_75t_L g825 ( 
.A1(n_761),
.A2(n_529),
.B(n_522),
.C(n_509),
.Y(n_825)
);

INVx2_ASAP7_75t_SL g826 ( 
.A(n_701),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_683),
.A2(n_705),
.B(n_685),
.Y(n_827)
);

NOR2x1_ASAP7_75t_L g828 ( 
.A(n_679),
.B(n_290),
.Y(n_828)
);

NOR3xp33_ASAP7_75t_L g829 ( 
.A(n_753),
.B(n_455),
.C(n_454),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_698),
.Y(n_830)
);

AOI21xp5_ASAP7_75t_L g831 ( 
.A1(n_685),
.A2(n_629),
.B(n_595),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_702),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_662),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_651),
.B(n_455),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_646),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_764),
.B(n_488),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_670),
.B(n_488),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_655),
.B(n_509),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_L g839 ( 
.A1(n_671),
.A2(n_616),
.B(n_586),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_667),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_729),
.B(n_458),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_705),
.A2(n_642),
.B(n_671),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_655),
.B(n_663),
.Y(n_843)
);

AND2x2_ASAP7_75t_L g844 ( 
.A(n_729),
.B(n_458),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_789),
.A2(n_629),
.B(n_595),
.Y(n_845)
);

OR2x2_ASAP7_75t_L g846 ( 
.A(n_697),
.B(n_463),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_663),
.B(n_509),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_734),
.B(n_509),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_734),
.B(n_522),
.Y(n_849)
);

AOI21x1_ASAP7_75t_L g850 ( 
.A1(n_719),
.A2(n_725),
.B(n_720),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_667),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_789),
.A2(n_595),
.B(n_527),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_670),
.B(n_522),
.Y(n_853)
);

INVx2_ASAP7_75t_L g854 ( 
.A(n_707),
.Y(n_854)
);

BUFx12f_ASAP7_75t_L g855 ( 
.A(n_759),
.Y(n_855)
);

O2A1O1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_660),
.A2(n_471),
.B(n_463),
.C(n_469),
.Y(n_856)
);

AOI22xp33_ASAP7_75t_L g857 ( 
.A1(n_693),
.A2(n_521),
.B1(n_570),
.B2(n_259),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_711),
.B(n_718),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_736),
.B(n_753),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_721),
.B(n_522),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_789),
.A2(n_595),
.B(n_527),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_726),
.B(n_529),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_730),
.B(n_529),
.Y(n_863)
);

AOI22xp5_ASAP7_75t_L g864 ( 
.A1(n_780),
.A2(n_570),
.B1(n_521),
.B2(n_583),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_684),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_650),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_736),
.B(n_469),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_737),
.B(n_529),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_784),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_688),
.B(n_618),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_650),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_789),
.A2(n_628),
.B(n_527),
.Y(n_872)
);

A2O1A1Ixp33_ASAP7_75t_L g873 ( 
.A1(n_739),
.A2(n_470),
.B(n_471),
.C(n_183),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_745),
.B(n_618),
.Y(n_874)
);

INVx3_ASAP7_75t_L g875 ( 
.A(n_690),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_649),
.A2(n_628),
.B(n_527),
.Y(n_876)
);

A2O1A1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_739),
.A2(n_470),
.B(n_202),
.C(n_205),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_653),
.A2(n_628),
.B(n_527),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_795),
.A2(n_723),
.B(n_647),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_723),
.A2(n_628),
.B(n_527),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_L g881 ( 
.A(n_641),
.B(n_570),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_641),
.B(n_583),
.Y(n_882)
);

O2A1O1Ixp5_ASAP7_75t_L g883 ( 
.A1(n_773),
.A2(n_618),
.B(n_495),
.C(n_564),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_641),
.B(n_628),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_749),
.B(n_618),
.Y(n_885)
);

OAI22x1_ASAP7_75t_L g886 ( 
.A1(n_777),
.A2(n_296),
.B1(n_173),
.B2(n_181),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_750),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_766),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_SL g889 ( 
.A1(n_738),
.A2(n_617),
.B(n_634),
.C(n_626),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_766),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_752),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_643),
.A2(n_628),
.B(n_636),
.Y(n_892)
);

OAI21xp33_ASAP7_75t_L g893 ( 
.A1(n_688),
.A2(n_301),
.B(n_181),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_767),
.B(n_570),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_746),
.A2(n_570),
.B(n_521),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_640),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_641),
.B(n_501),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_657),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_687),
.B(n_521),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_640),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_674),
.A2(n_656),
.B(n_765),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_710),
.B(n_623),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_699),
.B(n_521),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_765),
.B(n_778),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_658),
.Y(n_905)
);

INVx3_ASAP7_75t_L g906 ( 
.A(n_690),
.Y(n_906)
);

INVx4_ASAP7_75t_L g907 ( 
.A(n_732),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_746),
.A2(n_521),
.B(n_495),
.Y(n_908)
);

AOI21xp33_ASAP7_75t_L g909 ( 
.A1(n_751),
.A2(n_172),
.B(n_183),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_650),
.B(n_476),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_641),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_735),
.B(n_501),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_710),
.B(n_623),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_798),
.A2(n_533),
.B(n_519),
.Y(n_914)
);

AOI21x1_ASAP7_75t_L g915 ( 
.A1(n_719),
.A2(n_569),
.B(n_563),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_799),
.A2(n_519),
.B(n_507),
.Y(n_916)
);

OAI21xp5_ASAP7_75t_L g917 ( 
.A1(n_686),
.A2(n_521),
.B(n_563),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_747),
.Y(n_918)
);

O2A1O1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_801),
.A2(n_561),
.B(n_489),
.C(n_542),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_735),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_661),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_637),
.A2(n_503),
.B(n_507),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_785),
.B(n_242),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_735),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_735),
.Y(n_925)
);

OAI21xp5_ASAP7_75t_L g926 ( 
.A1(n_638),
.A2(n_564),
.B(n_569),
.Y(n_926)
);

BUFx6f_ASAP7_75t_L g927 ( 
.A(n_645),
.Y(n_927)
);

AND2x4_ASAP7_75t_L g928 ( 
.A(n_665),
.B(n_476),
.Y(n_928)
);

OAI21xp33_ASAP7_75t_L g929 ( 
.A1(n_794),
.A2(n_199),
.B(n_172),
.Y(n_929)
);

AOI22xp33_ASAP7_75t_L g930 ( 
.A1(n_693),
.A2(n_242),
.B1(n_259),
.B2(n_278),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_672),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_677),
.A2(n_503),
.B(n_626),
.Y(n_932)
);

OR2x6_ASAP7_75t_SL g933 ( 
.A(n_709),
.B(n_189),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_673),
.Y(n_934)
);

BUFx2_ASAP7_75t_L g935 ( 
.A(n_747),
.Y(n_935)
);

OAI321xp33_ASAP7_75t_L g936 ( 
.A1(n_751),
.A2(n_482),
.A3(n_478),
.B1(n_242),
.B2(n_278),
.C(n_259),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_738),
.A2(n_494),
.B(n_487),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_800),
.B(n_494),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_675),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_775),
.A2(n_634),
.B(n_626),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_778),
.B(n_487),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_771),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_775),
.A2(n_634),
.B(n_625),
.Y(n_943)
);

NOR2x1p5_ASAP7_75t_L g944 ( 
.A(n_757),
.B(n_189),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_800),
.A2(n_196),
.B(n_198),
.C(n_199),
.Y(n_945)
);

INVx1_ASAP7_75t_SL g946 ( 
.A(n_666),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_774),
.B(n_487),
.Y(n_947)
);

OAI21xp5_ASAP7_75t_L g948 ( 
.A1(n_680),
.A2(n_546),
.B(n_489),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_783),
.B(n_489),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_772),
.A2(n_196),
.B(n_198),
.C(n_201),
.Y(n_950)
);

BUFx3_ASAP7_75t_L g951 ( 
.A(n_771),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_758),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_681),
.A2(n_625),
.B1(n_622),
.B2(n_617),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_676),
.B(n_278),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_735),
.B(n_542),
.Y(n_955)
);

AOI22xp33_ASAP7_75t_L g956 ( 
.A1(n_743),
.A2(n_322),
.B1(n_202),
.B2(n_283),
.Y(n_956)
);

OAI21xp5_ASAP7_75t_L g957 ( 
.A1(n_682),
.A2(n_542),
.B(n_543),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_772),
.A2(n_323),
.B(n_287),
.C(n_292),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_681),
.A2(n_696),
.B(n_689),
.Y(n_959)
);

OAI22xp5_ASAP7_75t_L g960 ( 
.A1(n_659),
.A2(n_289),
.B1(n_309),
.B2(n_307),
.Y(n_960)
);

OAI21xp33_ASAP7_75t_L g961 ( 
.A1(n_644),
.A2(n_326),
.B(n_300),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_760),
.B(n_543),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_700),
.A2(n_625),
.B(n_622),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_706),
.A2(n_622),
.B(n_617),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_712),
.A2(n_443),
.B(n_441),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_714),
.B(n_201),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_676),
.B(n_644),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_769),
.B(n_770),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_715),
.A2(n_441),
.B(n_443),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_676),
.B(n_478),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_716),
.A2(n_443),
.B(n_561),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_740),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_788),
.A2(n_573),
.B(n_561),
.C(n_546),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_744),
.B(n_546),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_720),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_722),
.A2(n_573),
.B(n_477),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_782),
.B(n_573),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_748),
.B(n_279),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_791),
.A2(n_482),
.B(n_479),
.C(n_477),
.Y(n_979)
);

NOR2x1_ASAP7_75t_L g980 ( 
.A(n_755),
.B(n_459),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_756),
.B(n_284),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_786),
.A2(n_479),
.B(n_477),
.C(n_459),
.Y(n_982)
);

BUFx2_ASAP7_75t_L g983 ( 
.A(n_743),
.Y(n_983)
);

INVxp67_ASAP7_75t_L g984 ( 
.A(n_743),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_824),
.Y(n_985)
);

OR2x6_ASAP7_75t_SL g986 ( 
.A(n_843),
.B(n_310),
.Y(n_986)
);

AOI22x1_ASAP7_75t_L g987 ( 
.A1(n_952),
.A2(n_668),
.B1(n_796),
.B2(n_652),
.Y(n_987)
);

INVx1_ASAP7_75t_SL g988 ( 
.A(n_869),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_881),
.A2(n_727),
.B(n_724),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_808),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_859),
.B(n_792),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_802),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_859),
.B(n_793),
.Y(n_993)
);

INVxp33_ASAP7_75t_L g994 ( 
.A(n_923),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_820),
.B(n_797),
.Y(n_995)
);

O2A1O1Ixp33_ASAP7_75t_L g996 ( 
.A1(n_811),
.A2(n_733),
.B(n_742),
.C(n_763),
.Y(n_996)
);

OAI22xp5_ASAP7_75t_L g997 ( 
.A1(n_811),
.A2(n_329),
.B1(n_326),
.B2(n_319),
.Y(n_997)
);

BUFx3_ASAP7_75t_L g998 ( 
.A(n_931),
.Y(n_998)
);

AOI21x1_ASAP7_75t_L g999 ( 
.A1(n_977),
.A2(n_779),
.B(n_776),
.Y(n_999)
);

INVx3_ASAP7_75t_L g1000 ( 
.A(n_802),
.Y(n_1000)
);

O2A1O1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_909),
.A2(n_733),
.B(n_742),
.C(n_754),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_804),
.A2(n_725),
.B(n_732),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_824),
.Y(n_1003)
);

OA21x2_ASAP7_75t_L g1004 ( 
.A1(n_827),
.A2(n_703),
.B(n_741),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_809),
.A2(n_694),
.B(n_717),
.C(n_704),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_802),
.Y(n_1006)
);

NOR2xp33_ASAP7_75t_L g1007 ( 
.A(n_809),
.B(n_678),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_841),
.B(n_692),
.Y(n_1008)
);

CKINVDCx16_ASAP7_75t_R g1009 ( 
.A(n_855),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_844),
.B(n_867),
.Y(n_1010)
);

O2A1O1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_950),
.A2(n_479),
.B(n_459),
.C(n_293),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_802),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_882),
.A2(n_762),
.B(n_309),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_814),
.Y(n_1014)
);

OAI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_904),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_830),
.B(n_293),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_817),
.B(n_284),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_834),
.B(n_832),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_SL g1019 ( 
.A(n_966),
.B(n_329),
.C(n_295),
.Y(n_1019)
);

A2O1A1Ixp33_ASAP7_75t_SL g1020 ( 
.A1(n_902),
.A2(n_459),
.B(n_762),
.C(n_293),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_803),
.A2(n_762),
.B(n_295),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_846),
.B(n_314),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_832),
.B(n_854),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

AOI22xp5_ASAP7_75t_L g1025 ( 
.A1(n_935),
.A2(n_762),
.B1(n_297),
.B2(n_307),
.Y(n_1025)
);

INVx3_ASAP7_75t_SL g1026 ( 
.A(n_833),
.Y(n_1026)
);

BUFx3_ASAP7_75t_L g1027 ( 
.A(n_931),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_817),
.B(n_321),
.Y(n_1028)
);

INVx2_ASAP7_75t_SL g1029 ( 
.A(n_826),
.Y(n_1029)
);

A2O1A1Ixp33_ASAP7_75t_L g1030 ( 
.A1(n_966),
.A2(n_321),
.B(n_299),
.C(n_304),
.Y(n_1030)
);

NOR2xp67_ASAP7_75t_SL g1031 ( 
.A(n_907),
.B(n_297),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_814),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_808),
.B(n_762),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_SL g1034 ( 
.A(n_812),
.B(n_299),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_893),
.B(n_306),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_814),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_821),
.B(n_483),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_821),
.B(n_483),
.Y(n_1038)
);

NOR2xp33_ASAP7_75t_L g1039 ( 
.A(n_946),
.B(n_306),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_887),
.B(n_483),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_803),
.A2(n_304),
.B(n_473),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_891),
.B(n_483),
.Y(n_1042)
);

BUFx2_ASAP7_75t_L g1043 ( 
.A(n_871),
.Y(n_1043)
);

A2O1A1Ixp33_ASAP7_75t_L g1044 ( 
.A1(n_842),
.A2(n_483),
.B(n_473),
.C(n_466),
.Y(n_1044)
);

NOR2xp67_ASAP7_75t_SL g1045 ( 
.A(n_907),
.B(n_855),
.Y(n_1045)
);

HB1xp67_ASAP7_75t_L g1046 ( 
.A(n_918),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_891),
.B(n_870),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_816),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_858),
.B(n_483),
.Y(n_1049)
);

OAI22xp5_ASAP7_75t_L g1050 ( 
.A1(n_873),
.A2(n_473),
.B1(n_466),
.B2(n_464),
.Y(n_1050)
);

INVxp67_ASAP7_75t_L g1051 ( 
.A(n_970),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_870),
.B(n_483),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_933),
.B(n_314),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_902),
.B(n_483),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_950),
.A2(n_314),
.B(n_10),
.C(n_13),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_836),
.B(n_473),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_835),
.Y(n_1057)
);

O2A1O1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_958),
.A2(n_936),
.B(n_877),
.C(n_945),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_814),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_898),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_928),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_873),
.A2(n_473),
.B(n_466),
.C(n_464),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_901),
.A2(n_473),
.B(n_466),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_958),
.A2(n_9),
.B(n_17),
.C(n_19),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_879),
.A2(n_464),
.B(n_466),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_836),
.B(n_466),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_954),
.B(n_888),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_SL g1068 ( 
.A(n_890),
.B(n_464),
.Y(n_1068)
);

BUFx3_ASAP7_75t_L g1069 ( 
.A(n_866),
.Y(n_1069)
);

O2A1O1Ixp5_ASAP7_75t_L g1070 ( 
.A1(n_913),
.A2(n_108),
.B(n_129),
.C(n_128),
.Y(n_1070)
);

OR2x2_ASAP7_75t_SL g1071 ( 
.A(n_910),
.B(n_20),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_913),
.B(n_464),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_928),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_959),
.A2(n_464),
.B(n_126),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_905),
.Y(n_1075)
);

BUFx6f_ASAP7_75t_L g1076 ( 
.A(n_840),
.Y(n_1076)
);

NOR3xp33_ASAP7_75t_SL g1077 ( 
.A(n_818),
.B(n_21),
.C(n_22),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_884),
.A2(n_123),
.B(n_122),
.Y(n_1078)
);

INVx4_ASAP7_75t_L g1079 ( 
.A(n_840),
.Y(n_1079)
);

BUFx3_ASAP7_75t_L g1080 ( 
.A(n_951),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_R g1081 ( 
.A(n_810),
.B(n_851),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_921),
.Y(n_1082)
);

NOR3xp33_ASAP7_75t_L g1083 ( 
.A(n_929),
.B(n_29),
.C(n_31),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_968),
.B(n_121),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_884),
.A2(n_955),
.B(n_845),
.Y(n_1085)
);

AOI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_847),
.A2(n_838),
.B(n_852),
.Y(n_1086)
);

AND2x4_ASAP7_75t_L g1087 ( 
.A(n_865),
.B(n_875),
.Y(n_1087)
);

AOI21xp33_ASAP7_75t_L g1088 ( 
.A1(n_856),
.A2(n_29),
.B(n_31),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_861),
.A2(n_872),
.B(n_977),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_877),
.A2(n_945),
.B(n_829),
.C(n_895),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_875),
.B(n_78),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_837),
.B(n_34),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_934),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_815),
.A2(n_102),
.B(n_96),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_928),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_837),
.B(n_853),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_972),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_853),
.B(n_35),
.Y(n_1098)
);

O2A1O1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_960),
.A2(n_36),
.B(n_37),
.C(n_38),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_956),
.A2(n_37),
.B1(n_40),
.B2(n_43),
.Y(n_1100)
);

NOR2xp33_ASAP7_75t_L g1101 ( 
.A(n_967),
.B(n_43),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_899),
.A2(n_94),
.B(n_81),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_903),
.A2(n_70),
.B(n_69),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_911),
.A2(n_68),
.B(n_45),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_911),
.A2(n_63),
.B(n_46),
.Y(n_1105)
);

AO31x2_ASAP7_75t_L g1106 ( 
.A1(n_983),
.A2(n_44),
.A3(n_47),
.B(n_48),
.Y(n_1106)
);

NOR2xp67_ASAP7_75t_L g1107 ( 
.A(n_886),
.B(n_48),
.Y(n_1107)
);

NAND2x1p5_ASAP7_75t_L g1108 ( 
.A(n_840),
.B(n_49),
.Y(n_1108)
);

OR2x2_ASAP7_75t_L g1109 ( 
.A(n_939),
.B(n_49),
.Y(n_1109)
);

HB1xp67_ASAP7_75t_L g1110 ( 
.A(n_984),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_947),
.B(n_50),
.Y(n_1111)
);

NOR3xp33_ASAP7_75t_SL g1112 ( 
.A(n_961),
.B(n_52),
.C(n_55),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_906),
.B(n_58),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_SL g1114 ( 
.A(n_972),
.B(n_52),
.C(n_57),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_906),
.B(n_58),
.Y(n_1115)
);

BUFx4f_ASAP7_75t_SL g1116 ( 
.A(n_840),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_949),
.B(n_848),
.Y(n_1117)
);

AO21x1_ASAP7_75t_L g1118 ( 
.A1(n_813),
.A2(n_979),
.B(n_937),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_920),
.A2(n_924),
.B(n_925),
.Y(n_1119)
);

OAI22xp5_ASAP7_75t_SL g1120 ( 
.A1(n_930),
.A2(n_956),
.B1(n_857),
.B2(n_822),
.Y(n_1120)
);

OAI21xp33_ASAP7_75t_L g1121 ( 
.A1(n_930),
.A2(n_857),
.B(n_978),
.Y(n_1121)
);

O2A1O1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_981),
.A2(n_889),
.B(n_944),
.C(n_849),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_L g1123 ( 
.A(n_951),
.Y(n_1123)
);

A2O1A1Ixp33_ASAP7_75t_L g1124 ( 
.A1(n_864),
.A2(n_894),
.B(n_908),
.C(n_892),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_825),
.A2(n_941),
.B(n_916),
.C(n_914),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_920),
.A2(n_924),
.B(n_925),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_942),
.Y(n_1127)
);

NAND2xp5_ASAP7_75t_L g1128 ( 
.A(n_896),
.B(n_900),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_975),
.B(n_896),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_975),
.Y(n_1130)
);

NOR2xp33_ASAP7_75t_L g1131 ( 
.A(n_900),
.B(n_975),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_889),
.A2(n_868),
.B(n_874),
.C(n_863),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_860),
.Y(n_1133)
);

BUFx4f_ASAP7_75t_L g1134 ( 
.A(n_975),
.Y(n_1134)
);

INVx2_ASAP7_75t_L g1135 ( 
.A(n_990),
.Y(n_1135)
);

O2A1O1Ixp5_ASAP7_75t_SL g1136 ( 
.A1(n_1088),
.A2(n_807),
.B(n_839),
.C(n_897),
.Y(n_1136)
);

AOI221x1_ASAP7_75t_L g1137 ( 
.A1(n_1088),
.A2(n_876),
.B1(n_878),
.B2(n_819),
.C(n_823),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1057),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_989),
.A2(n_805),
.B(n_806),
.Y(n_1139)
);

INVx2_ASAP7_75t_SL g1140 ( 
.A(n_998),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_993),
.B(n_962),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1086),
.A2(n_938),
.B(n_831),
.Y(n_1142)
);

AND2x2_ASAP7_75t_L g1143 ( 
.A(n_1051),
.B(n_828),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_985),
.Y(n_1144)
);

NAND3xp33_ASAP7_75t_SL g1145 ( 
.A(n_1083),
.B(n_922),
.C(n_932),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1003),
.Y(n_1146)
);

OAI22xp5_ASAP7_75t_L g1147 ( 
.A1(n_1120),
.A2(n_862),
.B1(n_885),
.B2(n_927),
.Y(n_1147)
);

BUFx3_ASAP7_75t_L g1148 ( 
.A(n_1027),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_1121),
.A2(n_980),
.B(n_919),
.C(n_963),
.Y(n_1149)
);

AOI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_1054),
.A2(n_917),
.B(n_897),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_991),
.B(n_927),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1074),
.A2(n_912),
.B(n_926),
.Y(n_1152)
);

AND2x4_ASAP7_75t_L g1153 ( 
.A(n_1080),
.B(n_1123),
.Y(n_1153)
);

NOR2xp33_ASAP7_75t_L g1154 ( 
.A(n_1010),
.B(n_850),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_1072),
.A2(n_912),
.B(n_974),
.Y(n_1155)
);

NOR2x1_ASAP7_75t_SL g1156 ( 
.A(n_1047),
.B(n_927),
.Y(n_1156)
);

INVx8_ASAP7_75t_L g1157 ( 
.A(n_1006),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1035),
.A2(n_943),
.B1(n_940),
.B2(n_953),
.Y(n_1158)
);

NOR2xp33_ASAP7_75t_L g1159 ( 
.A(n_994),
.B(n_988),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1072),
.A2(n_880),
.B(n_957),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1084),
.A2(n_948),
.B(n_964),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_991),
.B(n_965),
.Y(n_1162)
);

O2A1O1Ixp5_ASAP7_75t_L g1163 ( 
.A1(n_1017),
.A2(n_883),
.B(n_976),
.C(n_915),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_1026),
.Y(n_1164)
);

AOI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_1084),
.A2(n_982),
.B(n_973),
.Y(n_1165)
);

OA21x2_ASAP7_75t_L g1166 ( 
.A1(n_1044),
.A2(n_971),
.B(n_969),
.Y(n_1166)
);

AOI31xp67_ASAP7_75t_L g1167 ( 
.A1(n_1034),
.A2(n_1052),
.A3(n_1066),
.B(n_1056),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_995),
.B(n_1007),
.Y(n_1169)
);

AO31x2_ASAP7_75t_L g1170 ( 
.A1(n_1062),
.A2(n_1125),
.A3(n_1050),
.B(n_1124),
.Y(n_1170)
);

AND2x2_ASAP7_75t_L g1171 ( 
.A(n_1022),
.B(n_1067),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1039),
.B(n_1018),
.Y(n_1172)
);

AND2x6_ASAP7_75t_SL g1173 ( 
.A(n_1053),
.B(n_1101),
.Y(n_1173)
);

INVx5_ASAP7_75t_L g1174 ( 
.A(n_1006),
.Y(n_1174)
);

AOI221xp5_ASAP7_75t_L g1175 ( 
.A1(n_997),
.A2(n_1015),
.B1(n_1100),
.B2(n_1058),
.C(n_1099),
.Y(n_1175)
);

NAND2x1p5_ASAP7_75t_L g1176 ( 
.A(n_1134),
.B(n_992),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1085),
.A2(n_1119),
.B(n_1126),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1043),
.Y(n_1178)
);

INVx2_ASAP7_75t_L g1179 ( 
.A(n_1024),
.Y(n_1179)
);

AOI22xp5_ASAP7_75t_L g1180 ( 
.A1(n_1028),
.A2(n_1073),
.B1(n_1095),
.B2(n_1061),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_995),
.B(n_1047),
.Y(n_1181)
);

AOI211x1_ASAP7_75t_L g1182 ( 
.A1(n_1100),
.A2(n_1015),
.B(n_1093),
.C(n_1075),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1002),
.A2(n_1117),
.B(n_1052),
.Y(n_1183)
);

A2O1A1Ixp33_ASAP7_75t_L g1184 ( 
.A1(n_1122),
.A2(n_1090),
.B(n_1030),
.C(n_1011),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1117),
.A2(n_1132),
.B(n_1008),
.Y(n_1185)
);

AOI21xp33_ASAP7_75t_L g1186 ( 
.A1(n_1092),
.A2(n_1098),
.B(n_1055),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1096),
.B(n_1133),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1016),
.B(n_1110),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_987),
.A2(n_1063),
.B(n_1038),
.Y(n_1189)
);

OAI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_1056),
.A2(n_1066),
.B(n_996),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1049),
.A2(n_1005),
.B(n_1001),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1006),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1070),
.A2(n_1033),
.B(n_1050),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_997),
.A2(n_1048),
.B1(n_1087),
.B2(n_1115),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1060),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1019),
.B(n_1046),
.Y(n_1196)
);

AO32x2_ASAP7_75t_L g1197 ( 
.A1(n_992),
.A2(n_1079),
.A3(n_1012),
.B1(n_1020),
.B2(n_1106),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1128),
.A2(n_1129),
.B(n_1023),
.Y(n_1198)
);

OAI21x1_ASAP7_75t_L g1199 ( 
.A1(n_1037),
.A2(n_1038),
.B(n_1040),
.Y(n_1199)
);

BUFx6f_ASAP7_75t_L g1200 ( 
.A(n_1123),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1033),
.A2(n_1111),
.B(n_1094),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1037),
.A2(n_1040),
.B(n_1042),
.Y(n_1202)
);

OAI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1042),
.A2(n_1103),
.B(n_1102),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1131),
.B(n_1128),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1013),
.A2(n_1021),
.B(n_1041),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1087),
.A2(n_1091),
.B1(n_1082),
.B2(n_1107),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1112),
.B(n_1114),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1064),
.A2(n_1077),
.B(n_1113),
.C(n_1109),
.Y(n_1208)
);

O2A1O1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1105),
.A2(n_1108),
.B(n_1104),
.C(n_1068),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1134),
.A2(n_1004),
.B(n_1078),
.Y(n_1210)
);

BUFx4f_ASAP7_75t_SL g1211 ( 
.A(n_1069),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1127),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1091),
.A2(n_1130),
.B(n_1079),
.Y(n_1213)
);

AO32x2_ASAP7_75t_L g1214 ( 
.A1(n_1012),
.A2(n_1106),
.A3(n_986),
.B1(n_1071),
.B2(n_1029),
.Y(n_1214)
);

OA21x2_ASAP7_75t_L g1215 ( 
.A1(n_1025),
.A2(n_1106),
.B(n_1108),
.Y(n_1215)
);

O2A1O1Ixp33_ASAP7_75t_SL g1216 ( 
.A1(n_1000),
.A2(n_1032),
.B(n_1081),
.C(n_1031),
.Y(n_1216)
);

NAND2x1p5_ASAP7_75t_L g1217 ( 
.A(n_1014),
.B(n_1076),
.Y(n_1217)
);

AOI22xp5_ASAP7_75t_L g1218 ( 
.A1(n_1097),
.A2(n_1009),
.B1(n_1045),
.B2(n_1123),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1116),
.A2(n_1014),
.B1(n_1036),
.B2(n_1059),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1036),
.A2(n_811),
.B(n_859),
.C(n_843),
.Y(n_1220)
);

OR2x6_ASAP7_75t_L g1221 ( 
.A(n_1059),
.B(n_1076),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1059),
.A2(n_989),
.B(n_881),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1076),
.A2(n_989),
.B(n_881),
.Y(n_1223)
);

OAI21x1_ASAP7_75t_L g1224 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1224)
);

AO31x2_ASAP7_75t_L g1225 ( 
.A1(n_1118),
.A2(n_1062),
.A3(n_1044),
.B(n_1125),
.Y(n_1225)
);

O2A1O1Ixp5_ASAP7_75t_L g1226 ( 
.A1(n_1074),
.A2(n_843),
.B(n_811),
.C(n_691),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1010),
.B(n_731),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1229)
);

A2O1A1Ixp33_ASAP7_75t_L g1230 ( 
.A1(n_1121),
.A2(n_811),
.B(n_859),
.C(n_843),
.Y(n_1230)
);

OAI22x1_ASAP7_75t_L g1231 ( 
.A1(n_1101),
.A2(n_811),
.B1(n_859),
.B2(n_539),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1051),
.B(n_923),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_988),
.Y(n_1234)
);

BUFx3_ASAP7_75t_L g1235 ( 
.A(n_998),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_993),
.B(n_991),
.Y(n_1236)
);

OA21x2_ASAP7_75t_L g1237 ( 
.A1(n_1074),
.A2(n_1118),
.B(n_1044),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1010),
.B(n_731),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1239)
);

NOR2xp33_ASAP7_75t_SL g1240 ( 
.A(n_1120),
.B(n_811),
.Y(n_1240)
);

INVx2_ASAP7_75t_L g1241 ( 
.A(n_990),
.Y(n_1241)
);

OAI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_1124),
.A2(n_811),
.B(n_843),
.Y(n_1242)
);

AOI21xp5_ASAP7_75t_L g1243 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1243)
);

NOR2xp33_ASAP7_75t_L g1244 ( 
.A(n_1010),
.B(n_731),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1010),
.B(n_859),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1118),
.A2(n_1062),
.A3(n_1044),
.B(n_1125),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1057),
.Y(n_1247)
);

OR2x2_ASAP7_75t_L g1248 ( 
.A(n_988),
.B(n_713),
.Y(n_1248)
);

OR2x2_ASAP7_75t_L g1249 ( 
.A(n_988),
.B(n_713),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1121),
.A2(n_811),
.B(n_859),
.C(n_843),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1010),
.B(n_859),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1057),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1080),
.B(n_1123),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1124),
.A2(n_811),
.B(n_843),
.Y(n_1257)
);

NAND2x1p5_ASAP7_75t_L g1258 ( 
.A(n_1134),
.B(n_802),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1057),
.Y(n_1259)
);

O2A1O1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1030),
.A2(n_811),
.B(n_843),
.C(n_731),
.Y(n_1260)
);

NOR2xp33_ASAP7_75t_L g1261 ( 
.A(n_1010),
.B(n_731),
.Y(n_1261)
);

OR2x6_ASAP7_75t_L g1262 ( 
.A(n_998),
.B(n_1027),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1264)
);

BUFx2_ASAP7_75t_L g1265 ( 
.A(n_988),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1057),
.Y(n_1266)
);

OR2x2_ASAP7_75t_L g1267 ( 
.A(n_988),
.B(n_713),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_SL g1268 ( 
.A(n_1010),
.B(n_859),
.Y(n_1268)
);

OAI21x1_ASAP7_75t_L g1269 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_988),
.B(n_713),
.Y(n_1270)
);

O2A1O1Ixp5_ASAP7_75t_L g1271 ( 
.A1(n_1074),
.A2(n_843),
.B(n_811),
.C(n_691),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1057),
.Y(n_1272)
);

NAND3xp33_ASAP7_75t_L g1273 ( 
.A(n_1083),
.B(n_811),
.C(n_843),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1010),
.B(n_859),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1275)
);

AO31x2_ASAP7_75t_L g1276 ( 
.A1(n_1118),
.A2(n_1062),
.A3(n_1044),
.B(n_1125),
.Y(n_1276)
);

OAI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1101),
.A2(n_811),
.B1(n_859),
.B2(n_539),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_990),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1281)
);

OAI21x1_ASAP7_75t_L g1282 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1283)
);

O2A1O1Ixp5_ASAP7_75t_L g1284 ( 
.A1(n_1074),
.A2(n_843),
.B(n_811),
.C(n_691),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_999),
.A2(n_1089),
.B(n_1065),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_989),
.A2(n_881),
.B(n_728),
.Y(n_1286)
);

BUFx10_ASAP7_75t_L g1287 ( 
.A(n_1039),
.Y(n_1287)
);

AOI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1052),
.A2(n_1072),
.B(n_1054),
.Y(n_1288)
);

BUFx3_ASAP7_75t_L g1289 ( 
.A(n_998),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1010),
.B(n_859),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1174),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1240),
.A2(n_1277),
.B1(n_1231),
.B2(n_1273),
.Y(n_1292)
);

OAI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1240),
.A2(n_1273),
.B1(n_1253),
.B2(n_1245),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_SL g1295 ( 
.A(n_1230),
.B(n_1252),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_L g1296 ( 
.A1(n_1175),
.A2(n_1257),
.B1(n_1242),
.B2(n_1274),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1138),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1195),
.Y(n_1298)
);

INVxp67_ASAP7_75t_SL g1299 ( 
.A(n_1151),
.Y(n_1299)
);

CKINVDCx11_ASAP7_75t_R g1300 ( 
.A(n_1287),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1236),
.A2(n_1169),
.B1(n_1172),
.B2(n_1257),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1242),
.A2(n_1290),
.B1(n_1268),
.B2(n_1186),
.Y(n_1302)
);

BUFx6f_ASAP7_75t_L g1303 ( 
.A(n_1174),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1247),
.Y(n_1304)
);

INVx6_ASAP7_75t_L g1305 ( 
.A(n_1192),
.Y(n_1305)
);

AO22x1_ASAP7_75t_L g1306 ( 
.A1(n_1244),
.A2(n_1261),
.B1(n_1207),
.B2(n_1171),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1186),
.A2(n_1236),
.B1(n_1169),
.B2(n_1287),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1144),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1255),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1141),
.A2(n_1187),
.B1(n_1181),
.B2(n_1233),
.Y(n_1310)
);

CKINVDCx6p67_ASAP7_75t_R g1311 ( 
.A(n_1148),
.Y(n_1311)
);

INVx1_ASAP7_75t_SL g1312 ( 
.A(n_1265),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_L g1313 ( 
.A1(n_1141),
.A2(n_1187),
.B1(n_1181),
.B2(n_1194),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1196),
.A2(n_1145),
.B1(n_1188),
.B2(n_1143),
.Y(n_1314)
);

CKINVDCx11_ASAP7_75t_R g1315 ( 
.A(n_1173),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1259),
.Y(n_1316)
);

INVx5_ASAP7_75t_L g1317 ( 
.A(n_1221),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1146),
.Y(n_1318)
);

INVx2_ASAP7_75t_SL g1319 ( 
.A(n_1235),
.Y(n_1319)
);

CKINVDCx20_ASAP7_75t_R g1320 ( 
.A(n_1164),
.Y(n_1320)
);

INVx1_ASAP7_75t_SL g1321 ( 
.A(n_1248),
.Y(n_1321)
);

HB1xp67_ASAP7_75t_SL g1322 ( 
.A(n_1289),
.Y(n_1322)
);

NAND2x1p5_ASAP7_75t_L g1323 ( 
.A(n_1192),
.B(n_1200),
.Y(n_1323)
);

INVx3_ASAP7_75t_SL g1324 ( 
.A(n_1262),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1154),
.A2(n_1162),
.B1(n_1206),
.B2(n_1215),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1220),
.A2(n_1178),
.B1(n_1260),
.B2(n_1151),
.Y(n_1326)
);

INVx3_ASAP7_75t_L g1327 ( 
.A(n_1258),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_1153),
.Y(n_1328)
);

OAI21xp33_ASAP7_75t_L g1329 ( 
.A1(n_1184),
.A2(n_1208),
.B(n_1159),
.Y(n_1329)
);

BUFx4f_ASAP7_75t_SL g1330 ( 
.A(n_1153),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_1249),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1266),
.Y(n_1332)
);

OAI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1178),
.A2(n_1213),
.B1(n_1267),
.B2(n_1270),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1262),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1272),
.Y(n_1335)
);

INVx3_ASAP7_75t_SL g1336 ( 
.A(n_1262),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_SL g1337 ( 
.A1(n_1173),
.A2(n_1215),
.B1(n_1156),
.B2(n_1211),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1204),
.A2(n_1180),
.B1(n_1182),
.B2(n_1147),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1204),
.A2(n_1237),
.B1(n_1147),
.B2(n_1185),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1218),
.A2(n_1140),
.B1(n_1219),
.B2(n_1176),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_L g1341 ( 
.A1(n_1237),
.A2(n_1135),
.B1(n_1278),
.B2(n_1241),
.Y(n_1341)
);

INVx6_ASAP7_75t_L g1342 ( 
.A(n_1192),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1190),
.A2(n_1152),
.B1(n_1193),
.B2(n_1212),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1256),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1256),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1176),
.A2(n_1258),
.B1(n_1158),
.B2(n_1210),
.Y(n_1346)
);

AOI22xp33_ASAP7_75t_L g1347 ( 
.A1(n_1190),
.A2(n_1193),
.B1(n_1198),
.B2(n_1271),
.Y(n_1347)
);

BUFx10_ASAP7_75t_L g1348 ( 
.A(n_1200),
.Y(n_1348)
);

OAI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1201),
.A2(n_1284),
.B1(n_1226),
.B2(n_1191),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_SL g1350 ( 
.A1(n_1205),
.A2(n_1203),
.B1(n_1201),
.B2(n_1214),
.Y(n_1350)
);

OAI22xp5_ASAP7_75t_L g1351 ( 
.A1(n_1229),
.A2(n_1264),
.B1(n_1286),
.B2(n_1251),
.Y(n_1351)
);

CKINVDCx14_ASAP7_75t_R g1352 ( 
.A(n_1221),
.Y(n_1352)
);

BUFx10_ASAP7_75t_L g1353 ( 
.A(n_1221),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1232),
.A2(n_1243),
.B1(n_1281),
.B2(n_1279),
.Y(n_1354)
);

OAI22xp33_ASAP7_75t_L g1355 ( 
.A1(n_1205),
.A2(n_1137),
.B1(n_1183),
.B2(n_1203),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1157),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1217),
.Y(n_1357)
);

BUFx12f_ASAP7_75t_L g1358 ( 
.A(n_1217),
.Y(n_1358)
);

INVx8_ASAP7_75t_L g1359 ( 
.A(n_1157),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1157),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1202),
.A2(n_1165),
.B1(n_1150),
.B2(n_1161),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1166),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1202),
.A2(n_1254),
.B1(n_1250),
.B2(n_1275),
.Y(n_1363)
);

INVx6_ASAP7_75t_L g1364 ( 
.A(n_1216),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1197),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1197),
.Y(n_1366)
);

INVx6_ASAP7_75t_L g1367 ( 
.A(n_1197),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1155),
.A2(n_1199),
.B1(n_1142),
.B2(n_1160),
.Y(n_1368)
);

OAI22xp5_ASAP7_75t_L g1369 ( 
.A1(n_1222),
.A2(n_1223),
.B1(n_1209),
.B2(n_1149),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1214),
.Y(n_1370)
);

BUFx3_ASAP7_75t_L g1371 ( 
.A(n_1177),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_1168),
.Y(n_1372)
);

AOI22xp33_ASAP7_75t_L g1373 ( 
.A1(n_1166),
.A2(n_1139),
.B1(n_1189),
.B2(n_1285),
.Y(n_1373)
);

BUFx5_ASAP7_75t_L g1374 ( 
.A(n_1224),
.Y(n_1374)
);

OAI22xp5_ASAP7_75t_L g1375 ( 
.A1(n_1288),
.A2(n_1167),
.B1(n_1136),
.B2(n_1170),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1225),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1163),
.Y(n_1377)
);

HB1xp67_ASAP7_75t_L g1378 ( 
.A(n_1246),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1246),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1276),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1227),
.A2(n_1239),
.B1(n_1263),
.B2(n_1269),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1280),
.A2(n_1282),
.B1(n_1283),
.B2(n_1276),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1383)
);

AOI22xp5_ASAP7_75t_L g1384 ( 
.A1(n_1240),
.A2(n_811),
.B1(n_1277),
.B2(n_1231),
.Y(n_1384)
);

INVx6_ASAP7_75t_L g1385 ( 
.A(n_1174),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1138),
.Y(n_1386)
);

CKINVDCx6p67_ASAP7_75t_R g1387 ( 
.A(n_1148),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1164),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1174),
.Y(n_1389)
);

BUFx8_ASAP7_75t_L g1390 ( 
.A(n_1234),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1164),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_1234),
.Y(n_1392)
);

INVx1_ASAP7_75t_SL g1393 ( 
.A(n_1234),
.Y(n_1393)
);

BUFx2_ASAP7_75t_SL g1394 ( 
.A(n_1148),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1179),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1138),
.Y(n_1397)
);

BUFx3_ASAP7_75t_L g1398 ( 
.A(n_1148),
.Y(n_1398)
);

CKINVDCx16_ASAP7_75t_R g1399 ( 
.A(n_1148),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_L g1400 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1400)
);

INVx6_ASAP7_75t_L g1401 ( 
.A(n_1174),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_811),
.B2(n_859),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1240),
.A2(n_843),
.B1(n_1277),
.B2(n_1231),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1240),
.A2(n_811),
.B1(n_1277),
.B2(n_1231),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1406)
);

AND2x2_ASAP7_75t_L g1407 ( 
.A(n_1228),
.B(n_1238),
.Y(n_1407)
);

BUFx4f_ASAP7_75t_SL g1408 ( 
.A(n_1148),
.Y(n_1408)
);

INVx3_ASAP7_75t_L g1409 ( 
.A(n_1258),
.Y(n_1409)
);

BUFx3_ASAP7_75t_L g1410 ( 
.A(n_1148),
.Y(n_1410)
);

BUFx4f_ASAP7_75t_L g1411 ( 
.A(n_1262),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1412)
);

INVx6_ASAP7_75t_L g1413 ( 
.A(n_1174),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1164),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_L g1415 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1415)
);

AOI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1240),
.A2(n_1120),
.B1(n_1277),
.B2(n_1231),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1321),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1294),
.B(n_1407),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1376),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1379),
.Y(n_1420)
);

INVx2_ASAP7_75t_SL g1421 ( 
.A(n_1411),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1380),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1378),
.Y(n_1423)
);

INVx2_ASAP7_75t_SL g1424 ( 
.A(n_1411),
.Y(n_1424)
);

AO21x2_ASAP7_75t_L g1425 ( 
.A1(n_1355),
.A2(n_1349),
.B(n_1375),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1291),
.Y(n_1426)
);

BUFx3_ASAP7_75t_L g1427 ( 
.A(n_1324),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1299),
.B(n_1308),
.Y(n_1428)
);

BUFx2_ASAP7_75t_L g1429 ( 
.A(n_1377),
.Y(n_1429)
);

BUFx3_ASAP7_75t_L g1430 ( 
.A(n_1324),
.Y(n_1430)
);

AOI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1369),
.A2(n_1295),
.B(n_1351),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1388),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1367),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1308),
.B(n_1318),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1370),
.Y(n_1435)
);

AO21x2_ASAP7_75t_L g1436 ( 
.A1(n_1354),
.A2(n_1295),
.B(n_1365),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1373),
.A2(n_1381),
.B(n_1368),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1317),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1366),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1301),
.B(n_1310),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1318),
.Y(n_1441)
);

OAI21x1_ASAP7_75t_L g1442 ( 
.A1(n_1373),
.A2(n_1368),
.B(n_1381),
.Y(n_1442)
);

INVx2_ASAP7_75t_L g1443 ( 
.A(n_1362),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1310),
.B(n_1313),
.Y(n_1444)
);

HB1xp67_ASAP7_75t_L g1445 ( 
.A(n_1333),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_SL g1446 ( 
.A1(n_1402),
.A2(n_1326),
.B1(n_1364),
.B2(n_1338),
.Y(n_1446)
);

INVxp33_ASAP7_75t_L g1447 ( 
.A(n_1322),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1346),
.B(n_1371),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1384),
.B(n_1404),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1374),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_L g1451 ( 
.A(n_1313),
.B(n_1307),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1367),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1367),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1297),
.Y(n_1454)
);

INVx2_ASAP7_75t_L g1455 ( 
.A(n_1374),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1298),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1304),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1372),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1309),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1363),
.A2(n_1361),
.B(n_1347),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1363),
.A2(n_1361),
.B(n_1347),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1331),
.B(n_1329),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1316),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1332),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1335),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1386),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1397),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1383),
.A2(n_1416),
.B1(n_1406),
.B2(n_1415),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1350),
.A2(n_1339),
.B(n_1296),
.Y(n_1469)
);

OAI21x1_ASAP7_75t_L g1470 ( 
.A1(n_1343),
.A2(n_1339),
.B(n_1341),
.Y(n_1470)
);

OR2x2_ASAP7_75t_L g1471 ( 
.A(n_1292),
.B(n_1314),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1395),
.B(n_1400),
.Y(n_1472)
);

AO21x2_ASAP7_75t_L g1473 ( 
.A1(n_1403),
.A2(n_1293),
.B(n_1396),
.Y(n_1473)
);

BUFx3_ASAP7_75t_L g1474 ( 
.A(n_1336),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1395),
.A2(n_1406),
.B1(n_1412),
.B2(n_1405),
.Y(n_1475)
);

AO21x1_ASAP7_75t_SL g1476 ( 
.A1(n_1400),
.A2(n_1412),
.B(n_1405),
.Y(n_1476)
);

OA21x2_ASAP7_75t_L g1477 ( 
.A1(n_1343),
.A2(n_1325),
.B(n_1341),
.Y(n_1477)
);

BUFx2_ASAP7_75t_L g1478 ( 
.A(n_1334),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1292),
.A2(n_1315),
.B1(n_1296),
.B2(n_1314),
.Y(n_1479)
);

BUFx3_ASAP7_75t_L g1480 ( 
.A(n_1336),
.Y(n_1480)
);

OAI22xp5_ASAP7_75t_L g1481 ( 
.A1(n_1307),
.A2(n_1302),
.B1(n_1352),
.B2(n_1337),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1325),
.B(n_1306),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1382),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1364),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1312),
.A2(n_1393),
.B1(n_1392),
.B2(n_1364),
.Y(n_1485)
);

OAI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1340),
.A2(n_1357),
.B(n_1327),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1317),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1353),
.Y(n_1488)
);

INVx2_ASAP7_75t_L g1489 ( 
.A(n_1353),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1327),
.Y(n_1490)
);

OAI21xp5_ASAP7_75t_L g1491 ( 
.A1(n_1446),
.A2(n_1345),
.B(n_1319),
.Y(n_1491)
);

AND2x2_ASAP7_75t_L g1492 ( 
.A(n_1449),
.B(n_1328),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1445),
.B(n_1328),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1468),
.B(n_1398),
.C(n_1410),
.D(n_1315),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1417),
.B(n_1390),
.Y(n_1495)
);

OR2x6_ASAP7_75t_L g1496 ( 
.A(n_1469),
.B(n_1394),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_L g1497 ( 
.A1(n_1479),
.A2(n_1409),
.B(n_1323),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1449),
.B(n_1390),
.Y(n_1498)
);

AND2x2_ASAP7_75t_L g1499 ( 
.A(n_1478),
.B(n_1344),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_SL g1500 ( 
.A(n_1485),
.B(n_1399),
.Y(n_1500)
);

INVx5_ASAP7_75t_L g1501 ( 
.A(n_1458),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1454),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1475),
.A2(n_1352),
.B1(n_1330),
.B2(n_1311),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1442),
.A2(n_1391),
.B(n_1413),
.Y(n_1504)
);

A2O1A1Ixp33_ASAP7_75t_L g1505 ( 
.A1(n_1462),
.A2(n_1398),
.B(n_1410),
.C(n_1360),
.Y(n_1505)
);

INVx11_ASAP7_75t_L g1506 ( 
.A(n_1447),
.Y(n_1506)
);

OR2x2_ASAP7_75t_L g1507 ( 
.A(n_1428),
.B(n_1454),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1418),
.B(n_1320),
.Y(n_1508)
);

OAI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1451),
.A2(n_1356),
.B(n_1360),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1456),
.Y(n_1510)
);

CKINVDCx8_ASAP7_75t_R g1511 ( 
.A(n_1432),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1429),
.B(n_1348),
.Y(n_1512)
);

NOR2x1_ASAP7_75t_R g1513 ( 
.A(n_1427),
.B(n_1414),
.Y(n_1513)
);

OAI21xp5_ASAP7_75t_L g1514 ( 
.A1(n_1451),
.A2(n_1356),
.B(n_1300),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1472),
.A2(n_1387),
.B1(n_1408),
.B2(n_1305),
.Y(n_1515)
);

AOI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1472),
.A2(n_1481),
.B1(n_1471),
.B2(n_1444),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1428),
.B(n_1414),
.Y(n_1517)
);

BUFx12f_ASAP7_75t_L g1518 ( 
.A(n_1421),
.Y(n_1518)
);

AOI22xp5_ASAP7_75t_L g1519 ( 
.A1(n_1481),
.A2(n_1358),
.B1(n_1413),
.B2(n_1305),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1482),
.A2(n_1291),
.B(n_1401),
.Y(n_1520)
);

AOI22xp5_ASAP7_75t_L g1521 ( 
.A1(n_1471),
.A2(n_1358),
.B1(n_1305),
.B2(n_1342),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1442),
.A2(n_1342),
.B(n_1385),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1456),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1457),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1444),
.A2(n_1303),
.B(n_1389),
.C(n_1359),
.Y(n_1525)
);

AO21x2_ASAP7_75t_L g1526 ( 
.A1(n_1437),
.A2(n_1342),
.B(n_1385),
.Y(n_1526)
);

NOR2x1_ASAP7_75t_SL g1527 ( 
.A(n_1473),
.B(n_1389),
.Y(n_1527)
);

O2A1O1Ixp33_ASAP7_75t_SL g1528 ( 
.A1(n_1484),
.A2(n_1401),
.B(n_1413),
.C(n_1359),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1434),
.B(n_1427),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1428),
.B(n_1434),
.Y(n_1530)
);

NOR2x1_ASAP7_75t_SL g1531 ( 
.A(n_1473),
.B(n_1389),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1440),
.A2(n_1359),
.B(n_1461),
.C(n_1460),
.Y(n_1532)
);

AO32x1_ASAP7_75t_L g1533 ( 
.A1(n_1483),
.A2(n_1422),
.A3(n_1420),
.B1(n_1419),
.B2(n_1423),
.Y(n_1533)
);

O2A1O1Ixp33_ASAP7_75t_L g1534 ( 
.A1(n_1440),
.A2(n_1486),
.B(n_1421),
.C(n_1424),
.Y(n_1534)
);

O2A1O1Ixp33_ASAP7_75t_L g1535 ( 
.A1(n_1486),
.A2(n_1424),
.B(n_1484),
.C(n_1488),
.Y(n_1535)
);

AOI221xp5_ASAP7_75t_L g1536 ( 
.A1(n_1425),
.A2(n_1483),
.B1(n_1473),
.B2(n_1428),
.C(n_1436),
.Y(n_1536)
);

NOR2x1_ASAP7_75t_SL g1537 ( 
.A(n_1473),
.B(n_1431),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_L g1538 ( 
.A1(n_1460),
.A2(n_1461),
.B(n_1470),
.Y(n_1538)
);

AOI221xp5_ASAP7_75t_L g1539 ( 
.A1(n_1425),
.A2(n_1436),
.B1(n_1466),
.B2(n_1459),
.C(n_1464),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1427),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1470),
.A2(n_1477),
.B(n_1442),
.Y(n_1541)
);

CKINVDCx16_ASAP7_75t_R g1542 ( 
.A(n_1430),
.Y(n_1542)
);

OR2x6_ASAP7_75t_L g1543 ( 
.A(n_1448),
.B(n_1438),
.Y(n_1543)
);

AND2x4_ASAP7_75t_L g1544 ( 
.A(n_1430),
.B(n_1474),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1430),
.B(n_1474),
.Y(n_1545)
);

OR2x2_ASAP7_75t_L g1546 ( 
.A(n_1459),
.B(n_1463),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1488),
.B(n_1489),
.Y(n_1547)
);

AO21x1_ASAP7_75t_L g1548 ( 
.A1(n_1490),
.A2(n_1423),
.B(n_1465),
.Y(n_1548)
);

AO32x2_ASAP7_75t_L g1549 ( 
.A1(n_1438),
.A2(n_1426),
.A3(n_1435),
.B1(n_1436),
.B2(n_1425),
.Y(n_1549)
);

HB1xp67_ASAP7_75t_L g1550 ( 
.A(n_1441),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1489),
.B(n_1474),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1502),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1510),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1523),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1524),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1541),
.B(n_1436),
.Y(n_1556)
);

INVxp67_ASAP7_75t_SL g1557 ( 
.A(n_1548),
.Y(n_1557)
);

AND2x4_ASAP7_75t_SL g1558 ( 
.A(n_1543),
.B(n_1496),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1541),
.B(n_1538),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1538),
.B(n_1425),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1522),
.Y(n_1561)
);

AOI221x1_ASAP7_75t_SL g1562 ( 
.A1(n_1494),
.A2(n_1476),
.B1(n_1467),
.B2(n_1465),
.C(n_1466),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1546),
.Y(n_1563)
);

INVx4_ASAP7_75t_L g1564 ( 
.A(n_1496),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1522),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1494),
.A2(n_1476),
.B1(n_1477),
.B2(n_1448),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1507),
.B(n_1530),
.Y(n_1567)
);

INVx1_ASAP7_75t_SL g1568 ( 
.A(n_1547),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1550),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1549),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1549),
.B(n_1439),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_1504),
.Y(n_1572)
);

OAI21xp5_ASAP7_75t_SL g1573 ( 
.A1(n_1519),
.A2(n_1433),
.B(n_1487),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1549),
.B(n_1439),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1533),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1533),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1526),
.Y(n_1577)
);

BUFx2_ASAP7_75t_SL g1578 ( 
.A(n_1501),
.Y(n_1578)
);

AOI21xp5_ASAP7_75t_R g1579 ( 
.A1(n_1503),
.A2(n_1480),
.B(n_1426),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1504),
.B(n_1543),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1496),
.A2(n_1477),
.B1(n_1480),
.B2(n_1448),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1537),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1527),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1531),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1529),
.Y(n_1585)
);

OAI221xp5_ASAP7_75t_SL g1586 ( 
.A1(n_1566),
.A2(n_1516),
.B1(n_1534),
.B2(n_1539),
.C(n_1519),
.Y(n_1586)
);

BUFx3_ASAP7_75t_L g1587 ( 
.A(n_1558),
.Y(n_1587)
);

NAND3xp33_ASAP7_75t_L g1588 ( 
.A(n_1557),
.B(n_1500),
.C(n_1516),
.Y(n_1588)
);

OR2x2_ASAP7_75t_L g1589 ( 
.A(n_1570),
.B(n_1452),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1561),
.Y(n_1590)
);

NAND3xp33_ASAP7_75t_SL g1591 ( 
.A(n_1566),
.B(n_1535),
.C(n_1514),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1553),
.Y(n_1592)
);

INVx2_ASAP7_75t_SL g1593 ( 
.A(n_1553),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1559),
.B(n_1536),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1559),
.B(n_1433),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1559),
.B(n_1452),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1552),
.Y(n_1597)
);

NAND2xp5_ASAP7_75t_L g1598 ( 
.A(n_1569),
.B(n_1532),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1570),
.B(n_1453),
.Y(n_1599)
);

INVx1_ASAP7_75t_SL g1600 ( 
.A(n_1568),
.Y(n_1600)
);

AOI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1581),
.A2(n_1497),
.B1(n_1514),
.B2(n_1515),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1571),
.B(n_1448),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1557),
.Y(n_1603)
);

AND2x4_ASAP7_75t_SL g1604 ( 
.A(n_1564),
.B(n_1544),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1552),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1568),
.Y(n_1606)
);

INVx4_ASAP7_75t_L g1607 ( 
.A(n_1564),
.Y(n_1607)
);

NOR2x1_ASAP7_75t_L g1608 ( 
.A(n_1564),
.B(n_1545),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1581),
.A2(n_1497),
.B1(n_1491),
.B2(n_1492),
.Y(n_1609)
);

AO21x2_ASAP7_75t_L g1610 ( 
.A1(n_1570),
.A2(n_1437),
.B(n_1422),
.Y(n_1610)
);

INVx1_ASAP7_75t_SL g1611 ( 
.A(n_1577),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1554),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1571),
.B(n_1448),
.Y(n_1613)
);

NOR2xp33_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1498),
.Y(n_1614)
);

BUFx2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1574),
.Y(n_1616)
);

BUFx2_ASAP7_75t_L g1617 ( 
.A(n_1582),
.Y(n_1617)
);

AO21x2_ASAP7_75t_L g1618 ( 
.A1(n_1570),
.A2(n_1450),
.B(n_1455),
.Y(n_1618)
);

INVx3_ASAP7_75t_L g1619 ( 
.A(n_1561),
.Y(n_1619)
);

INVxp67_ASAP7_75t_SL g1620 ( 
.A(n_1561),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1554),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1555),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1556),
.B(n_1443),
.Y(n_1623)
);

HB1xp67_ASAP7_75t_L g1624 ( 
.A(n_1593),
.Y(n_1624)
);

BUFx2_ASAP7_75t_L g1625 ( 
.A(n_1608),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1616),
.B(n_1556),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1616),
.B(n_1556),
.Y(n_1627)
);

OR2x2_ASAP7_75t_L g1628 ( 
.A(n_1589),
.B(n_1575),
.Y(n_1628)
);

NOR2xp67_ASAP7_75t_L g1629 ( 
.A(n_1603),
.B(n_1564),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1592),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1608),
.B(n_1561),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1616),
.B(n_1602),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1602),
.B(n_1560),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1597),
.Y(n_1635)
);

CKINVDCx5p33_ASAP7_75t_R g1636 ( 
.A(n_1614),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1589),
.B(n_1575),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1597),
.Y(n_1638)
);

INVxp67_ASAP7_75t_SL g1639 ( 
.A(n_1603),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1605),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1594),
.B(n_1563),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1605),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1589),
.B(n_1576),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1618),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1612),
.Y(n_1645)
);

INVx5_ASAP7_75t_SL g1646 ( 
.A(n_1610),
.Y(n_1646)
);

INVx2_ASAP7_75t_L g1647 ( 
.A(n_1618),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1612),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1613),
.B(n_1560),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1621),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

NAND2x1p5_ASAP7_75t_L g1652 ( 
.A(n_1607),
.B(n_1564),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1621),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1622),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1618),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1613),
.B(n_1594),
.Y(n_1656)
);

OR2x2_ASAP7_75t_L g1657 ( 
.A(n_1599),
.B(n_1576),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1622),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1613),
.B(n_1565),
.Y(n_1659)
);

INVx2_ASAP7_75t_SL g1660 ( 
.A(n_1593),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1594),
.B(n_1565),
.Y(n_1661)
);

AND2x2_ASAP7_75t_L g1662 ( 
.A(n_1615),
.B(n_1565),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1641),
.B(n_1656),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1636),
.B(n_1588),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1641),
.B(n_1598),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1656),
.B(n_1604),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1635),
.Y(n_1667)
);

AOI322xp5_ASAP7_75t_L g1668 ( 
.A1(n_1639),
.A2(n_1591),
.A3(n_1609),
.B1(n_1601),
.B2(n_1598),
.C1(n_1595),
.C2(n_1611),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1635),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1567),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1639),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1636),
.B(n_1588),
.Y(n_1672)
);

NOR2x1_ASAP7_75t_L g1673 ( 
.A(n_1625),
.B(n_1591),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1625),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1638),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1661),
.B(n_1596),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1638),
.Y(n_1677)
);

INVxp67_ASAP7_75t_L g1678 ( 
.A(n_1625),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1640),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1661),
.B(n_1567),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1661),
.B(n_1596),
.Y(n_1681)
);

OR2x2_ASAP7_75t_L g1682 ( 
.A(n_1632),
.B(n_1567),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1652),
.A2(n_1586),
.B1(n_1601),
.B2(n_1609),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1640),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1629),
.B(n_1600),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1633),
.B(n_1587),
.Y(n_1686)
);

OR2x2_ASAP7_75t_L g1687 ( 
.A(n_1632),
.B(n_1600),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1632),
.B(n_1606),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1633),
.B(n_1604),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1633),
.B(n_1606),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1642),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1642),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1645),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1634),
.B(n_1596),
.Y(n_1694)
);

INVxp67_ASAP7_75t_L g1695 ( 
.A(n_1645),
.Y(n_1695)
);

NOR2xp67_ASAP7_75t_L g1696 ( 
.A(n_1629),
.B(n_1607),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1648),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1648),
.Y(n_1698)
);

AOI22xp5_ASAP7_75t_L g1699 ( 
.A1(n_1652),
.A2(n_1558),
.B1(n_1573),
.B2(n_1580),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1634),
.B(n_1587),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1650),
.Y(n_1701)
);

NOR2x1p5_ASAP7_75t_L g1702 ( 
.A(n_1634),
.B(n_1587),
.Y(n_1702)
);

AND2x4_ASAP7_75t_L g1703 ( 
.A(n_1631),
.B(n_1607),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1660),
.Y(n_1704)
);

INVx2_ASAP7_75t_L g1705 ( 
.A(n_1660),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1664),
.B(n_1649),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1697),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1697),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1667),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1669),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_R g1711 ( 
.A(n_1664),
.B(n_1511),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1675),
.Y(n_1712)
);

NAND2x1_ASAP7_75t_SL g1713 ( 
.A(n_1673),
.B(n_1631),
.Y(n_1713)
);

OR2x2_ASAP7_75t_L g1714 ( 
.A(n_1663),
.B(n_1628),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1677),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1679),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1670),
.B(n_1649),
.Y(n_1717)
);

INVx4_ASAP7_75t_L g1718 ( 
.A(n_1685),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1702),
.B(n_1649),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1684),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1614),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1665),
.B(n_1623),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1691),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1696),
.B(n_1631),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1692),
.Y(n_1725)
);

INVx1_ASAP7_75t_SL g1726 ( 
.A(n_1672),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1683),
.B(n_1586),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1671),
.B(n_1623),
.Y(n_1728)
);

OR2x2_ASAP7_75t_L g1729 ( 
.A(n_1671),
.B(n_1628),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1676),
.B(n_1623),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1681),
.B(n_1666),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1693),
.Y(n_1732)
);

AND2x2_ASAP7_75t_SL g1733 ( 
.A(n_1703),
.B(n_1542),
.Y(n_1733)
);

OAI322xp33_ASAP7_75t_L g1734 ( 
.A1(n_1674),
.A2(n_1643),
.A3(n_1637),
.B1(n_1628),
.B2(n_1657),
.C1(n_1652),
.C2(n_1611),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1698),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1686),
.B(n_1562),
.Y(n_1736)
);

OAI22xp5_ASAP7_75t_L g1737 ( 
.A1(n_1699),
.A2(n_1579),
.B1(n_1505),
.B2(n_1587),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1686),
.B(n_1652),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1685),
.A2(n_1513),
.B(n_1495),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1700),
.B(n_1690),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1700),
.B(n_1659),
.Y(n_1741)
);

OAI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1727),
.A2(n_1678),
.B1(n_1674),
.B2(n_1562),
.C(n_1695),
.Y(n_1742)
);

CKINVDCx14_ASAP7_75t_R g1743 ( 
.A(n_1711),
.Y(n_1743)
);

AOI32xp33_ASAP7_75t_L g1744 ( 
.A1(n_1721),
.A2(n_1703),
.A3(n_1631),
.B1(n_1689),
.B2(n_1659),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_SL g1745 ( 
.A1(n_1726),
.A2(n_1678),
.B(n_1573),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1707),
.Y(n_1746)
);

AOI31xp33_ASAP7_75t_SL g1747 ( 
.A1(n_1736),
.A2(n_1695),
.A3(n_1687),
.B(n_1688),
.Y(n_1747)
);

NAND3xp33_ASAP7_75t_L g1748 ( 
.A(n_1718),
.B(n_1705),
.C(n_1704),
.Y(n_1748)
);

OAI22xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1733),
.A2(n_1508),
.B1(n_1518),
.B2(n_1703),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1733),
.B(n_1680),
.Y(n_1750)
);

AOI21xp5_ASAP7_75t_L g1751 ( 
.A1(n_1739),
.A2(n_1701),
.B(n_1631),
.Y(n_1751)
);

AND2x4_ASAP7_75t_L g1752 ( 
.A(n_1718),
.B(n_1704),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1706),
.B(n_1694),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1713),
.A2(n_1607),
.B1(n_1705),
.B2(n_1682),
.C(n_1520),
.Y(n_1754)
);

OAI22xp5_ASAP7_75t_L g1755 ( 
.A1(n_1737),
.A2(n_1579),
.B1(n_1607),
.B2(n_1572),
.Y(n_1755)
);

AOI22xp5_ASAP7_75t_L g1756 ( 
.A1(n_1719),
.A2(n_1580),
.B1(n_1558),
.B2(n_1572),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1718),
.A2(n_1620),
.B(n_1525),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1740),
.B(n_1650),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1708),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_L g1760 ( 
.A(n_1711),
.B(n_1572),
.Y(n_1760)
);

AOI22xp33_ASAP7_75t_L g1761 ( 
.A1(n_1738),
.A2(n_1558),
.B1(n_1580),
.B2(n_1572),
.Y(n_1761)
);

INVx1_ASAP7_75t_SL g1762 ( 
.A(n_1738),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1719),
.A2(n_1572),
.B1(n_1646),
.B2(n_1584),
.Y(n_1763)
);

OR2x2_ASAP7_75t_L g1764 ( 
.A(n_1731),
.B(n_1637),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1717),
.B(n_1722),
.Y(n_1765)
);

OAI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1729),
.A2(n_1620),
.B(n_1551),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1728),
.B(n_1506),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1762),
.B(n_1709),
.Y(n_1768)
);

AOI221xp5_ASAP7_75t_L g1769 ( 
.A1(n_1745),
.A2(n_1742),
.B1(n_1734),
.B2(n_1744),
.C(n_1746),
.Y(n_1769)
);

OAI22xp5_ASAP7_75t_L g1770 ( 
.A1(n_1745),
.A2(n_1724),
.B1(n_1729),
.B2(n_1741),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1759),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1743),
.B(n_1710),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1749),
.A2(n_1750),
.B1(n_1755),
.B2(n_1760),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1767),
.B(n_1712),
.Y(n_1774)
);

NOR2xp67_ASAP7_75t_L g1775 ( 
.A(n_1748),
.B(n_1724),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1758),
.Y(n_1776)
);

AO21x1_ASAP7_75t_SL g1777 ( 
.A1(n_1757),
.A2(n_1716),
.B(n_1715),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_SL g1778 ( 
.A(n_1754),
.B(n_1724),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1752),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1764),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1752),
.A2(n_1741),
.B1(n_1735),
.B2(n_1732),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1753),
.B(n_1720),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1747),
.A2(n_1646),
.B1(n_1572),
.B2(n_1714),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1751),
.B(n_1723),
.Y(n_1784)
);

INVxp67_ASAP7_75t_L g1785 ( 
.A(n_1765),
.Y(n_1785)
);

INVx1_ASAP7_75t_SL g1786 ( 
.A(n_1766),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1756),
.Y(n_1787)
);

OAI32xp33_ASAP7_75t_L g1788 ( 
.A1(n_1783),
.A2(n_1763),
.A3(n_1714),
.B1(n_1725),
.B2(n_1761),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1779),
.B(n_1730),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1785),
.B(n_1659),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1768),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1780),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1772),
.Y(n_1793)
);

NOR2x1_ASAP7_75t_L g1794 ( 
.A(n_1775),
.B(n_1637),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1771),
.Y(n_1795)
);

AOI211x1_ASAP7_75t_SL g1796 ( 
.A1(n_1770),
.A2(n_1644),
.B(n_1655),
.C(n_1647),
.Y(n_1796)
);

NAND4xp25_ASAP7_75t_SL g1797 ( 
.A(n_1769),
.B(n_1662),
.C(n_1521),
.D(n_1626),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1781),
.B(n_1615),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1776),
.B(n_1653),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1792),
.Y(n_1800)
);

NOR4xp25_ASAP7_75t_L g1801 ( 
.A(n_1797),
.B(n_1783),
.C(n_1784),
.D(n_1786),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1790),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1793),
.B(n_1777),
.Y(n_1803)
);

NAND3xp33_ASAP7_75t_SL g1804 ( 
.A(n_1791),
.B(n_1778),
.C(n_1773),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_SL g1805 ( 
.A(n_1794),
.B(n_1782),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1795),
.B(n_1787),
.C(n_1774),
.Y(n_1806)
);

NOR3xp33_ASAP7_75t_L g1807 ( 
.A(n_1788),
.B(n_1789),
.C(n_1798),
.Y(n_1807)
);

AOI222xp33_ASAP7_75t_L g1808 ( 
.A1(n_1799),
.A2(n_1646),
.B1(n_1644),
.B2(n_1655),
.C1(n_1651),
.C2(n_1647),
.Y(n_1808)
);

AOI21x1_ASAP7_75t_L g1809 ( 
.A1(n_1799),
.A2(n_1624),
.B(n_1662),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1796),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_SL g1811 ( 
.A1(n_1794),
.A2(n_1660),
.B(n_1662),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_SL g1812 ( 
.A1(n_1801),
.A2(n_1521),
.B1(n_1499),
.B2(n_1643),
.C(n_1657),
.Y(n_1812)
);

AOI221xp5_ASAP7_75t_L g1813 ( 
.A1(n_1804),
.A2(n_1655),
.B1(n_1644),
.B2(n_1647),
.C(n_1651),
.Y(n_1813)
);

AOI22xp5_ASAP7_75t_L g1814 ( 
.A1(n_1804),
.A2(n_1512),
.B1(n_1545),
.B2(n_1604),
.Y(n_1814)
);

NOR4xp25_ASAP7_75t_SL g1815 ( 
.A(n_1805),
.B(n_1617),
.C(n_1615),
.D(n_1528),
.Y(n_1815)
);

NOR3xp33_ASAP7_75t_L g1816 ( 
.A(n_1806),
.B(n_1517),
.C(n_1480),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1816),
.B(n_1803),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1814),
.B(n_1807),
.Y(n_1818)
);

OR2x2_ASAP7_75t_L g1819 ( 
.A(n_1812),
.B(n_1802),
.Y(n_1819)
);

NAND2xp5_ASAP7_75t_L g1820 ( 
.A(n_1815),
.B(n_1800),
.Y(n_1820)
);

OAI221xp5_ASAP7_75t_L g1821 ( 
.A1(n_1813),
.A2(n_1811),
.B1(n_1810),
.B2(n_1809),
.C(n_1808),
.Y(n_1821)
);

INVx2_ASAP7_75t_L g1822 ( 
.A(n_1814),
.Y(n_1822)
);

NOR2x1_ASAP7_75t_L g1823 ( 
.A(n_1820),
.B(n_1643),
.Y(n_1823)
);

OAI221xp5_ASAP7_75t_L g1824 ( 
.A1(n_1821),
.A2(n_1617),
.B1(n_1657),
.B2(n_1590),
.C(n_1619),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1822),
.Y(n_1825)
);

NAND4xp75_ASAP7_75t_L g1826 ( 
.A(n_1818),
.B(n_1626),
.C(n_1627),
.D(n_1583),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1817),
.B(n_1626),
.Y(n_1827)
);

AOI21xp5_ASAP7_75t_L g1828 ( 
.A1(n_1824),
.A2(n_1819),
.B(n_1624),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1823),
.B(n_1653),
.Y(n_1829)
);

NOR3xp33_ASAP7_75t_L g1830 ( 
.A(n_1825),
.B(n_1509),
.C(n_1493),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1829),
.Y(n_1831)
);

BUFx3_ASAP7_75t_L g1832 ( 
.A(n_1831),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1832),
.Y(n_1833)
);

NOR2x1_ASAP7_75t_SL g1834 ( 
.A(n_1832),
.B(n_1826),
.Y(n_1834)
);

AOI22x1_ASAP7_75t_L g1835 ( 
.A1(n_1833),
.A2(n_1828),
.B1(n_1827),
.B2(n_1834),
.Y(n_1835)
);

OAI22xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1833),
.A2(n_1830),
.B1(n_1540),
.B2(n_1578),
.Y(n_1836)
);

AOI21xp33_ASAP7_75t_SL g1837 ( 
.A1(n_1835),
.A2(n_1658),
.B(n_1654),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1836),
.B(n_1654),
.Y(n_1838)
);

OAI22xp5_ASAP7_75t_SL g1839 ( 
.A1(n_1838),
.A2(n_1578),
.B1(n_1540),
.B2(n_1617),
.Y(n_1839)
);

AOI211x1_ASAP7_75t_L g1840 ( 
.A1(n_1839),
.A2(n_1837),
.B(n_1658),
.C(n_1630),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_L g1841 ( 
.A1(n_1840),
.A2(n_1646),
.B1(n_1590),
.B2(n_1619),
.Y(n_1841)
);

AOI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1841),
.A2(n_1627),
.B1(n_1646),
.B2(n_1619),
.Y(n_1842)
);

AOI211xp5_ASAP7_75t_L g1843 ( 
.A1(n_1842),
.A2(n_1540),
.B(n_1651),
.C(n_1647),
.Y(n_1843)
);


endmodule