module fake_aes_5872_n_556 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_556);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_556;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_29), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_57), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_59), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_35), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_41), .Y(n_82) );
CKINVDCx16_ASAP7_75t_R g83 ( .A(n_63), .Y(n_83) );
INVxp33_ASAP7_75t_L g84 ( .A(n_69), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_47), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_21), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_33), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_30), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_61), .Y(n_89) );
CKINVDCx20_ASAP7_75t_R g90 ( .A(n_26), .Y(n_90) );
CKINVDCx14_ASAP7_75t_R g91 ( .A(n_5), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_5), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_19), .Y(n_93) );
INVx2_ASAP7_75t_L g94 ( .A(n_7), .Y(n_94) );
CKINVDCx20_ASAP7_75t_R g95 ( .A(n_72), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_50), .Y(n_96) );
CKINVDCx20_ASAP7_75t_R g97 ( .A(n_27), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_18), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_0), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_34), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_53), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_44), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_13), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_77), .Y(n_104) );
CKINVDCx16_ASAP7_75t_R g105 ( .A(n_64), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_43), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_39), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_7), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_8), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_71), .Y(n_112) );
HB1xp67_ASAP7_75t_L g113 ( .A(n_111), .Y(n_113) );
AND2x2_ASAP7_75t_SL g114 ( .A(n_102), .B(n_36), .Y(n_114) );
AND2x4_ASAP7_75t_L g115 ( .A(n_102), .B(n_0), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_91), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_85), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_90), .Y(n_118) );
AND2x2_ASAP7_75t_L g119 ( .A(n_84), .B(n_1), .Y(n_119) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_83), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_85), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_86), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_86), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_87), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_87), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_88), .Y(n_126) );
BUFx3_ASAP7_75t_L g127 ( .A(n_88), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_89), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_89), .Y(n_129) );
AO21x2_ASAP7_75t_L g130 ( .A1(n_98), .A2(n_2), .B(n_3), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_98), .Y(n_131) );
HB1xp67_ASAP7_75t_L g132 ( .A(n_103), .Y(n_132) );
BUFx6f_ASAP7_75t_L g133 ( .A(n_112), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_112), .Y(n_134) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_94), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_80), .Y(n_137) );
NOR2xp33_ASAP7_75t_SL g138 ( .A(n_114), .B(n_116), .Y(n_138) );
NOR2xp33_ASAP7_75t_L g139 ( .A(n_116), .B(n_104), .Y(n_139) );
OAI22xp5_ASAP7_75t_SL g140 ( .A1(n_120), .A2(n_110), .B1(n_103), .B2(n_97), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_133), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_133), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_133), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_127), .B(n_101), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_113), .B(n_105), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_133), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_132), .B(n_109), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_133), .Y(n_149) );
NAND2x1p5_ASAP7_75t_L g150 ( .A(n_114), .B(n_108), .Y(n_150) );
INVx4_ASAP7_75t_L g151 ( .A(n_115), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_133), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_135), .Y(n_153) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_114), .B(n_78), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
AND2x2_ASAP7_75t_L g156 ( .A(n_115), .B(n_94), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_135), .Y(n_157) );
AND2x4_ASAP7_75t_L g158 ( .A(n_115), .B(n_92), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_135), .Y(n_159) );
BUFx10_ASAP7_75t_L g160 ( .A(n_118), .Y(n_160) );
INVx4_ASAP7_75t_L g161 ( .A(n_127), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
AOI22xp5_ASAP7_75t_L g163 ( .A1(n_119), .A2(n_95), .B1(n_106), .B2(n_99), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_117), .B(n_107), .Y(n_164) );
AOI22xp5_ASAP7_75t_L g165 ( .A1(n_119), .A2(n_107), .B1(n_100), .B2(n_78), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_143), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_143), .B(n_100), .Y(n_167) );
BUFx3_ASAP7_75t_L g168 ( .A(n_158), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_143), .B(n_122), .Y(n_169) );
INVx1_ASAP7_75t_SL g170 ( .A(n_146), .Y(n_170) );
NAND2xp33_ASAP7_75t_L g171 ( .A(n_150), .B(n_129), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_146), .B(n_122), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_151), .B(n_124), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_158), .Y(n_174) );
INVx3_ASAP7_75t_L g175 ( .A(n_151), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_161), .Y(n_177) );
NAND2xp33_ASAP7_75t_SL g178 ( .A(n_154), .B(n_124), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_139), .B(n_126), .Y(n_179) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_160), .Y(n_180) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_150), .A2(n_130), .B1(n_117), .B2(n_121), .Y(n_181) );
AND2x2_ASAP7_75t_L g182 ( .A(n_165), .B(n_126), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_156), .Y(n_183) );
INVx2_ASAP7_75t_SL g184 ( .A(n_161), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_138), .A2(n_130), .B1(n_121), .B2(n_129), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_142), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_145), .B(n_128), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_156), .Y(n_188) );
INVx2_ASAP7_75t_SL g189 ( .A(n_161), .Y(n_189) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_164), .A2(n_128), .B(n_134), .Y(n_190) );
AND2x2_ASAP7_75t_L g191 ( .A(n_165), .B(n_131), .Y(n_191) );
BUFx3_ASAP7_75t_L g192 ( .A(n_158), .Y(n_192) );
INVx2_ASAP7_75t_SL g193 ( .A(n_158), .Y(n_193) );
INVx4_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_163), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g196 ( .A(n_148), .B(n_131), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_153), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_142), .Y(n_199) );
AOI22xp5_ASAP7_75t_L g200 ( .A1(n_140), .A2(n_130), .B1(n_134), .B2(n_137), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g201 ( .A(n_163), .B(n_137), .Y(n_201) );
AND2x2_ASAP7_75t_L g202 ( .A(n_182), .B(n_160), .Y(n_202) );
OAI22xp5_ASAP7_75t_L g203 ( .A1(n_193), .A2(n_123), .B1(n_125), .B2(n_136), .Y(n_203) );
AOI22xp5_ASAP7_75t_L g204 ( .A1(n_201), .A2(n_160), .B1(n_125), .B2(n_123), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_179), .B(n_136), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_175), .Y(n_206) );
BUFx2_ASAP7_75t_L g207 ( .A(n_168), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_168), .Y(n_208) );
BUFx12f_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
NOR2xp67_ASAP7_75t_SL g210 ( .A(n_193), .B(n_81), .Y(n_210) );
INVx4_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_187), .A2(n_135), .B(n_93), .C(n_96), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_172), .Y(n_213) );
NOR2x1_ASAP7_75t_L g214 ( .A(n_172), .B(n_82), .Y(n_214) );
BUFx2_ASAP7_75t_L g215 ( .A(n_174), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_196), .B(n_4), .Y(n_216) );
AND2x2_ASAP7_75t_L g217 ( .A(n_182), .B(n_4), .Y(n_217) );
AOI22xp5_ASAP7_75t_L g218 ( .A1(n_170), .A2(n_152), .B1(n_144), .B2(n_147), .Y(n_218) );
A2O1A1Ixp33_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_162), .B(n_155), .C(n_152), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_166), .Y(n_220) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_174), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_175), .Y(n_222) );
BUFx3_ASAP7_75t_L g223 ( .A(n_174), .Y(n_223) );
INVx3_ASAP7_75t_L g224 ( .A(n_175), .Y(n_224) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_170), .A2(n_149), .B1(n_144), .B2(n_147), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_166), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_192), .Y(n_227) );
CKINVDCx20_ASAP7_75t_R g228 ( .A(n_191), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_175), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_191), .Y(n_230) );
INVx2_ASAP7_75t_SL g231 ( .A(n_192), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_176), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_196), .B(n_6), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_183), .B(n_6), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_169), .A2(n_149), .B(n_141), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_194), .Y(n_236) );
NAND2x1p5_ASAP7_75t_L g237 ( .A(n_221), .B(n_194), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_213), .B(n_195), .Y(n_238) );
BUFx8_ASAP7_75t_L g239 ( .A(n_209), .Y(n_239) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_219), .A2(n_185), .B(n_181), .Y(n_240) );
AO31x2_ASAP7_75t_L g241 ( .A1(n_212), .A2(n_190), .A3(n_162), .B(n_157), .Y(n_241) );
OAI21x1_ASAP7_75t_L g242 ( .A1(n_235), .A2(n_185), .B(n_173), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_217), .B(n_183), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_220), .A2(n_193), .B(n_169), .Y(n_244) );
OAI21x1_ASAP7_75t_L g245 ( .A1(n_234), .A2(n_173), .B(n_197), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_221), .Y(n_246) );
NAND2x1p5_ASAP7_75t_L g247 ( .A(n_221), .B(n_194), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_236), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_220), .Y(n_249) );
INVx8_ASAP7_75t_L g250 ( .A(n_236), .Y(n_250) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_216), .A2(n_141), .B(n_153), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_202), .B(n_194), .Y(n_252) );
BUFx6f_ASAP7_75t_L g253 ( .A(n_221), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_233), .A2(n_197), .B(n_199), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_226), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_217), .B(n_188), .Y(n_256) );
OR2x6_ASAP7_75t_L g257 ( .A(n_207), .B(n_192), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_226), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_232), .Y(n_259) );
INVx6_ASAP7_75t_L g260 ( .A(n_221), .Y(n_260) );
BUFx2_ASAP7_75t_L g261 ( .A(n_207), .Y(n_261) );
OA21x2_ASAP7_75t_L g262 ( .A1(n_205), .A2(n_157), .B(n_159), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_232), .Y(n_263) );
BUFx8_ASAP7_75t_L g264 ( .A(n_209), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_252), .A2(n_230), .B1(n_228), .B2(n_200), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_256), .B(n_249), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_254), .A2(n_171), .B(n_178), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_238), .A2(n_202), .B1(n_230), .B2(n_228), .Y(n_268) );
OAI211xp5_ASAP7_75t_L g269 ( .A1(n_243), .A2(n_200), .B(n_204), .C(n_214), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_249), .Y(n_270) );
OAI221xp5_ASAP7_75t_L g271 ( .A1(n_238), .A2(n_188), .B1(n_215), .B2(n_227), .C(n_203), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_261), .Y(n_272) );
AOI221xp5_ASAP7_75t_L g273 ( .A1(n_256), .A2(n_255), .B1(n_258), .B2(n_259), .C(n_263), .Y(n_273) );
INVx3_ASAP7_75t_L g274 ( .A(n_237), .Y(n_274) );
OAI22xp5_ASAP7_75t_L g275 ( .A1(n_257), .A2(n_215), .B1(n_208), .B2(n_211), .Y(n_275) );
AOI21xp5_ASAP7_75t_L g276 ( .A1(n_254), .A2(n_206), .B(n_229), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_263), .B(n_206), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_248), .B(n_211), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_244), .B(n_211), .Y(n_279) );
OAI22xp5_ASAP7_75t_L g280 ( .A1(n_257), .A2(n_208), .B1(n_231), .B2(n_223), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_248), .B(n_208), .Y(n_281) );
AOI22xp33_ASAP7_75t_SL g282 ( .A1(n_250), .A2(n_223), .B1(n_231), .B2(n_224), .Y(n_282) );
CKINVDCx5p33_ASAP7_75t_R g283 ( .A(n_239), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_245), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_253), .Y(n_285) );
INVx3_ASAP7_75t_L g286 ( .A(n_237), .Y(n_286) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_284), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_266), .B(n_240), .Y(n_288) );
INVx2_ASAP7_75t_L g289 ( .A(n_284), .Y(n_289) );
INVx3_ASAP7_75t_L g290 ( .A(n_274), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_266), .B(n_261), .Y(n_291) );
AND2x2_ASAP7_75t_L g292 ( .A(n_270), .B(n_240), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_270), .B(n_240), .Y(n_293) );
AND2x4_ASAP7_75t_L g294 ( .A(n_274), .B(n_253), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_273), .B(n_240), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
AND2x2_ASAP7_75t_SL g297 ( .A(n_265), .B(n_279), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_285), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_277), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_279), .Y(n_300) );
OAI22xp5_ASAP7_75t_L g301 ( .A1(n_265), .A2(n_250), .B1(n_257), .B2(n_247), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_286), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_286), .Y(n_304) );
AND2x2_ASAP7_75t_SL g305 ( .A(n_278), .B(n_250), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_274), .B(n_237), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_269), .B(n_241), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_274), .B(n_241), .Y(n_308) );
AOI22xp33_ASAP7_75t_L g309 ( .A1(n_268), .A2(n_250), .B1(n_257), .B2(n_264), .Y(n_309) );
OR2x2_ASAP7_75t_L g310 ( .A(n_300), .B(n_272), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_291), .Y(n_311) );
AND2x4_ASAP7_75t_L g312 ( .A(n_300), .B(n_286), .Y(n_312) );
OAI221xp5_ASAP7_75t_L g313 ( .A1(n_309), .A2(n_271), .B1(n_282), .B2(n_281), .C(n_275), .Y(n_313) );
OR2x2_ASAP7_75t_L g314 ( .A(n_288), .B(n_286), .Y(n_314) );
NOR2x1_ASAP7_75t_L g315 ( .A(n_301), .B(n_280), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_305), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_294), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_288), .B(n_280), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_291), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_301), .B(n_283), .C(n_275), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_289), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_289), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_296), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_293), .B(n_285), .Y(n_324) );
AOI33xp33_ASAP7_75t_L g325 ( .A1(n_296), .A2(n_281), .A3(n_278), .B1(n_10), .B2(n_11), .B3(n_12), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_299), .Y(n_326) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g328 ( .A1(n_307), .A2(n_278), .B1(n_267), .B2(n_167), .C(n_276), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_293), .B(n_241), .Y(n_329) );
OAI211xp5_ASAP7_75t_SL g330 ( .A1(n_307), .A2(n_159), .B(n_239), .C(n_264), .Y(n_330) );
CKINVDCx20_ASAP7_75t_R g331 ( .A(n_306), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_297), .B(n_278), .Y(n_332) );
NOR2xp33_ASAP7_75t_L g333 ( .A(n_297), .B(n_239), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_289), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_305), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_293), .B(n_246), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_287), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_292), .B(n_241), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_287), .Y(n_339) );
OR2x2_ASAP7_75t_L g340 ( .A(n_308), .B(n_241), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_303), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_314), .B(n_308), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_321), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_329), .B(n_292), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_311), .B(n_297), .Y(n_345) );
AND2x2_ASAP7_75t_L g346 ( .A(n_329), .B(n_298), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_319), .B(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_338), .B(n_298), .Y(n_349) );
AOI221x1_ASAP7_75t_L g350 ( .A1(n_330), .A2(n_320), .B1(n_333), .B2(n_337), .C(n_339), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_338), .B(n_298), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_326), .B(n_303), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_322), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_314), .B(n_295), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_322), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_324), .B(n_302), .Y(n_356) );
NAND3xp33_ASAP7_75t_L g357 ( .A(n_325), .B(n_304), .C(n_295), .Y(n_357) );
NAND2x1_ASAP7_75t_SL g358 ( .A(n_335), .B(n_290), .Y(n_358) );
INVxp67_ASAP7_75t_L g359 ( .A(n_327), .Y(n_359) );
NOR2x1_ASAP7_75t_L g360 ( .A(n_335), .B(n_290), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_324), .B(n_302), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_331), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_334), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_336), .B(n_302), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_334), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_341), .Y(n_366) );
AND2x2_ASAP7_75t_SL g367 ( .A(n_335), .B(n_305), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_340), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_336), .B(n_304), .Y(n_369) );
INVx6_ASAP7_75t_L g370 ( .A(n_312), .Y(n_370) );
BUFx3_ASAP7_75t_L g371 ( .A(n_331), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_336), .B(n_306), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_310), .B(n_290), .Y(n_374) );
OR2x2_ASAP7_75t_L g375 ( .A(n_318), .B(n_290), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_340), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_318), .B(n_317), .Y(n_377) );
OR2x2_ASAP7_75t_L g378 ( .A(n_317), .B(n_294), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_325), .B(n_294), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_312), .B(n_294), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_317), .B(n_262), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_312), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_315), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_332), .B(n_262), .Y(n_384) );
AND2x4_ASAP7_75t_L g385 ( .A(n_316), .B(n_253), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_316), .B(n_262), .Y(n_386) );
INVx3_ASAP7_75t_L g387 ( .A(n_328), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_313), .Y(n_388) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_359), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_372), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_344), .B(n_251), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_355), .Y(n_392) );
AOI22xp33_ASAP7_75t_L g393 ( .A1(n_388), .A2(n_246), .B1(n_260), .B2(n_264), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_368), .B(n_8), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_344), .B(n_251), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_366), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_342), .B(n_9), .Y(n_397) );
OR2x2_ASAP7_75t_L g398 ( .A(n_342), .B(n_9), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_377), .B(n_251), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_366), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_368), .B(n_10), .Y(n_401) );
AND2x4_ASAP7_75t_L g402 ( .A(n_377), .B(n_253), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_376), .B(n_11), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_347), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_346), .B(n_251), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_376), .B(n_12), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_383), .B(n_13), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_373), .B(n_14), .Y(n_408) );
OR2x2_ASAP7_75t_L g409 ( .A(n_346), .B(n_14), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_383), .B(n_15), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_352), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_371), .B(n_15), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_343), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_349), .B(n_16), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_343), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_348), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_371), .B(n_16), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_373), .B(n_17), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_349), .B(n_351), .Y(n_419) );
NAND2x1_ASAP7_75t_L g420 ( .A(n_360), .B(n_262), .Y(n_420) );
INVxp67_ASAP7_75t_L g421 ( .A(n_371), .Y(n_421) );
NAND2x1_ASAP7_75t_L g422 ( .A(n_360), .B(n_260), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_348), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_17), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_353), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_356), .B(n_245), .Y(n_426) );
AOI21xp5_ASAP7_75t_L g427 ( .A1(n_367), .A2(n_242), .B(n_253), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_353), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_356), .B(n_242), .Y(n_429) );
NAND2x1p5_ASAP7_75t_L g430 ( .A(n_367), .B(n_246), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_365), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_355), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_361), .B(n_247), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_365), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_361), .B(n_247), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_375), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_363), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_388), .B(n_260), .Y(n_438) );
OR2x2_ASAP7_75t_L g439 ( .A(n_354), .B(n_20), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_364), .B(n_22), .Y(n_440) );
OR2x2_ASAP7_75t_L g441 ( .A(n_354), .B(n_23), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_392), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_389), .Y(n_443) );
OAI22xp5_ASAP7_75t_L g444 ( .A1(n_430), .A2(n_367), .B1(n_362), .B2(n_388), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_389), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_396), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_419), .B(n_364), .Y(n_447) );
AOI32xp33_ASAP7_75t_L g448 ( .A1(n_408), .A2(n_387), .A3(n_379), .B1(n_386), .B2(n_345), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_419), .B(n_382), .Y(n_449) );
INVxp67_ASAP7_75t_L g450 ( .A(n_404), .Y(n_450) );
AOI221x1_ASAP7_75t_L g451 ( .A1(n_407), .A2(n_387), .B1(n_357), .B2(n_374), .C(n_382), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g452 ( .A1(n_430), .A2(n_370), .B1(n_387), .B2(n_357), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g453 ( .A1(n_409), .A2(n_387), .B1(n_370), .B2(n_375), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_435), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_390), .B(n_384), .Y(n_455) );
NOR2xp33_ASAP7_75t_L g456 ( .A(n_421), .B(n_370), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_411), .B(n_384), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_400), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_421), .Y(n_459) );
NAND2xp33_ASAP7_75t_L g460 ( .A(n_412), .B(n_386), .Y(n_460) );
INVxp67_ASAP7_75t_L g461 ( .A(n_417), .Y(n_461) );
AND2x2_ASAP7_75t_SL g462 ( .A(n_424), .B(n_381), .Y(n_462) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_438), .A2(n_369), .B1(n_370), .B2(n_382), .Y(n_463) );
INVxp67_ASAP7_75t_SL g464 ( .A(n_420), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_435), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_436), .B(n_369), .Y(n_466) );
OAI22xp5_ASAP7_75t_L g467 ( .A1(n_397), .A2(n_378), .B1(n_380), .B2(n_381), .Y(n_467) );
INVxp67_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_391), .B(n_350), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_413), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_391), .B(n_350), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g472 ( .A1(n_393), .A2(n_378), .B1(n_363), .B2(n_385), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_415), .Y(n_473) );
OAI21xp5_ASAP7_75t_L g474 ( .A1(n_398), .A2(n_358), .B(n_385), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_395), .B(n_358), .Y(n_475) );
AOI32xp33_ASAP7_75t_L g476 ( .A1(n_418), .A2(n_385), .A3(n_224), .B1(n_229), .B2(n_222), .Y(n_476) );
AOI222xp33_ASAP7_75t_L g477 ( .A1(n_393), .A2(n_385), .B1(n_210), .B2(n_260), .C1(n_222), .C2(n_224), .Y(n_477) );
AOI21xp5_ASAP7_75t_L g478 ( .A1(n_427), .A2(n_225), .B(n_218), .Y(n_478) );
AOI32xp33_ASAP7_75t_L g479 ( .A1(n_395), .A2(n_176), .A3(n_210), .B1(n_28), .B2(n_31), .Y(n_479) );
NOR3xp33_ASAP7_75t_SL g480 ( .A(n_414), .B(n_24), .C(n_25), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_416), .Y(n_481) );
O2A1O1Ixp33_ASAP7_75t_L g482 ( .A1(n_394), .A2(n_189), .B(n_184), .C(n_177), .Y(n_482) );
OR2x2_ASAP7_75t_L g483 ( .A(n_405), .B(n_32), .Y(n_483) );
XNOR2x1_ASAP7_75t_L g484 ( .A(n_406), .B(n_37), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_423), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_443), .B(n_428), .Y(n_486) );
AOI32xp33_ASAP7_75t_L g487 ( .A1(n_452), .A2(n_440), .A3(n_405), .B1(n_399), .B2(n_426), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_442), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_445), .Y(n_489) );
OAI221xp5_ASAP7_75t_SL g490 ( .A1(n_448), .A2(n_403), .B1(n_401), .B2(n_439), .C(n_441), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_444), .B(n_399), .Y(n_491) );
XNOR2xp5_ASAP7_75t_L g492 ( .A(n_484), .B(n_433), .Y(n_492) );
OAI321xp33_ASAP7_75t_L g493 ( .A1(n_444), .A2(n_440), .A3(n_438), .B1(n_426), .B2(n_429), .C(n_425), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_468), .A2(n_434), .B(n_431), .C(n_422), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_469), .B(n_429), .Y(n_495) );
INVx2_ASAP7_75t_SL g496 ( .A(n_454), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_462), .B(n_402), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_453), .A2(n_467), .B1(n_460), .B2(n_472), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_471), .B(n_437), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_485), .B(n_437), .Y(n_501) );
AOI21xp33_ASAP7_75t_L g502 ( .A1(n_482), .A2(n_432), .B(n_392), .Y(n_502) );
OAI221xp5_ASAP7_75t_L g503 ( .A1(n_474), .A2(n_432), .B1(n_402), .B2(n_189), .C(n_184), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_458), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_467), .A2(n_402), .B1(n_189), .B2(n_184), .C(n_177), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_464), .A2(n_177), .B(n_40), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_473), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_455), .B(n_38), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_450), .B(n_42), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_481), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_449), .B(n_45), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_461), .B(n_46), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_459), .B(n_48), .Y(n_514) );
AOI31xp33_ASAP7_75t_L g515 ( .A1(n_491), .A2(n_474), .A3(n_453), .B(n_477), .Y(n_515) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_500), .A2(n_475), .B(n_451), .Y(n_516) );
INVx2_ASAP7_75t_SL g517 ( .A(n_496), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_501), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_501), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_500), .B(n_457), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_499), .A2(n_456), .B1(n_463), .B2(n_465), .Y(n_521) );
INVxp67_ASAP7_75t_SL g522 ( .A(n_494), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_495), .B(n_447), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_493), .B(n_476), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_498), .A2(n_477), .B(n_479), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_503), .A2(n_466), .B1(n_483), .B2(n_478), .Y(n_526) );
AOI22xp5_ASAP7_75t_L g527 ( .A1(n_492), .A2(n_480), .B1(n_199), .B2(n_186), .Y(n_527) );
AOI221xp5_ASAP7_75t_L g528 ( .A1(n_490), .A2(n_199), .B1(n_186), .B2(n_198), .C(n_54), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g529 ( .A1(n_489), .A2(n_186), .B1(n_51), .B2(n_52), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_512), .A2(n_49), .B1(n_55), .B2(n_56), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_488), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_518), .Y(n_532) );
AOI211xp5_ASAP7_75t_L g533 ( .A1(n_524), .A2(n_502), .B(n_505), .C(n_513), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_525), .B(n_487), .C(n_507), .D(n_502), .Y(n_534) );
NAND3xp33_ASAP7_75t_SL g535 ( .A(n_528), .B(n_514), .C(n_510), .Y(n_535) );
NAND3xp33_ASAP7_75t_L g536 ( .A(n_515), .B(n_509), .C(n_511), .Y(n_536) );
OAI211xp5_ASAP7_75t_SL g537 ( .A1(n_522), .A2(n_508), .B(n_506), .C(n_504), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_519), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_526), .A2(n_497), .B1(n_486), .B2(n_198), .C(n_65), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_517), .A2(n_520), .B1(n_521), .B2(n_523), .C(n_531), .Y(n_540) );
INVxp67_ASAP7_75t_SL g541 ( .A(n_533), .Y(n_541) );
NOR3xp33_ASAP7_75t_SL g542 ( .A(n_534), .B(n_520), .C(n_523), .Y(n_542) );
OR5x1_ASAP7_75t_L g543 ( .A(n_537), .B(n_516), .C(n_527), .D(n_530), .E(n_529), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_540), .B(n_58), .Y(n_544) );
NOR3xp33_ASAP7_75t_SL g545 ( .A(n_536), .B(n_60), .C(n_62), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_541), .Y(n_546) );
NAND3x1_ASAP7_75t_L g547 ( .A(n_543), .B(n_539), .C(n_538), .Y(n_547) );
NOR3xp33_ASAP7_75t_L g548 ( .A(n_544), .B(n_535), .C(n_532), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_546), .B(n_542), .Y(n_549) );
INVx1_ASAP7_75t_L g550 ( .A(n_548), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_549), .Y(n_551) );
OAI22xp5_ASAP7_75t_L g552 ( .A1(n_550), .A2(n_547), .B1(n_545), .B2(n_198), .Y(n_552) );
AOI22x1_ASAP7_75t_L g553 ( .A1(n_551), .A2(n_67), .B1(n_68), .B2(n_70), .Y(n_553) );
OAI21xp5_ASAP7_75t_L g554 ( .A1(n_553), .A2(n_552), .B(n_75), .Y(n_554) );
AOI22x1_ASAP7_75t_L g555 ( .A1(n_554), .A2(n_73), .B1(n_76), .B2(n_198), .Y(n_555) );
AOI21xp5_ASAP7_75t_L g556 ( .A1(n_555), .A2(n_198), .B(n_549), .Y(n_556) );
endmodule