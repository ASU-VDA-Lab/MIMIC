module fake_ibex_1989_n_916 (n_151, n_147, n_85, n_167, n_128, n_84, n_64, n_3, n_73, n_152, n_171, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_161, n_29, n_143, n_106, n_177, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_164, n_38, n_124, n_37, n_110, n_47, n_169, n_108, n_10, n_82, n_21, n_27, n_165, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_175, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_173, n_120, n_93, n_168, n_155, n_162, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_172, n_49, n_40, n_66, n_17, n_74, n_90, n_176, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_166, n_163, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_170, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_159, n_158, n_132, n_174, n_157, n_160, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_916);

input n_151;
input n_147;
input n_85;
input n_167;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_171;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_161;
input n_29;
input n_143;
input n_106;
input n_177;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_164;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_169;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_165;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_175;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_173;
input n_120;
input n_93;
input n_168;
input n_155;
input n_162;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_172;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_176;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_166;
input n_163;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_170;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_159;
input n_158;
input n_132;
input n_174;
input n_157;
input n_160;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_916;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_707;
wire n_273;
wire n_309;
wire n_330;
wire n_328;
wire n_372;
wire n_293;
wire n_341;
wire n_418;
wire n_256;
wire n_193;
wire n_510;
wire n_845;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_873;
wire n_593;
wire n_862;
wire n_545;
wire n_909;
wire n_583;
wire n_887;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_872;
wire n_423;
wire n_608;
wire n_864;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_861;
wire n_449;
wire n_547;
wire n_727;
wire n_216;
wire n_915;
wire n_911;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_900;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_340;
wire n_375;
wire n_698;
wire n_901;
wire n_187;
wire n_667;
wire n_884;
wire n_682;
wire n_850;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_879;
wire n_723;
wire n_270;
wire n_383;
wire n_346;
wire n_886;
wire n_840;
wire n_561;
wire n_883;
wire n_417;
wire n_471;
wire n_846;
wire n_739;
wire n_755;
wire n_265;
wire n_853;
wire n_504;
wire n_859;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_875;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_671;
wire n_228;
wire n_711;
wire n_876;
wire n_552;
wire n_251;
wire n_384;
wire n_632;
wire n_373;
wire n_854;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_898;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_673;
wire n_732;
wire n_798;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_893;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_914;
wire n_835;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_694;
wire n_787;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_865;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_907;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_852;
wire n_789;
wire n_880;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_904;
wire n_842;
wire n_355;
wire n_767;
wire n_474;
wire n_878;
wire n_758;
wire n_594;
wire n_636;
wire n_710;
wire n_720;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_791;
wire n_715;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_849;
wire n_857;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_851;
wire n_689;
wire n_793;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_910;
wire n_635;
wire n_844;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_847;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_262;
wire n_299;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_696;
wire n_837;
wire n_796;
wire n_797;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_869;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_882;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_651;
wire n_365;
wire n_721;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_444;
wire n_200;
wire n_506;
wire n_564;
wire n_562;
wire n_868;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_905;
wire n_308;
wire n_675;
wire n_800;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_894;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_888;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_906;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_214;
wire n_238;
wire n_579;
wire n_843;
wire n_899;
wire n_902;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_817;
wire n_744;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_881;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_863;
wire n_415;
wire n_597;
wire n_288;
wire n_285;
wire n_320;
wire n_379;
wire n_247;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_858;
wire n_342;
wire n_233;
wire n_414;
wire n_385;
wire n_430;
wire n_729;
wire n_807;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_198;
wire n_264;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_820;
wire n_670;
wire n_805;
wire n_892;
wire n_390;
wire n_544;
wire n_891;
wire n_913;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_856;
wire n_668;
wire n_779;
wire n_871;
wire n_266;
wire n_294;
wire n_485;
wire n_870;
wire n_284;
wire n_811;
wire n_808;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_903;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_885;
wire n_513;
wire n_212;
wire n_588;
wire n_877;
wire n_693;
wire n_311;
wire n_860;
wire n_661;
wire n_848;
wire n_406;
wire n_606;
wire n_737;
wire n_896;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_867;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_889;
wire n_897;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_697;
wire n_816;
wire n_874;
wire n_890;
wire n_912;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_908;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_394;
wire n_364;
wire n_687;
wire n_895;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_855;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_866;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_100),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_147),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_29),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_146),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_113),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_158),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

NOR2xp67_ASAP7_75t_L g186 ( 
.A(n_123),
.B(n_115),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_55),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_140),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_145),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_166),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_120),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_75),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_60),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_54),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_152),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_133),
.B(n_79),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_42),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_37),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_71),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_84),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_80),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_168),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_174),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_82),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_51),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_58),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_38),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_19),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_33),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVxp33_ASAP7_75t_SL g218 ( 
.A(n_162),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_150),
.Y(n_219)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_44),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_144),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_131),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_83),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_85),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_175),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_65),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_141),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_47),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_154),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_32),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_3),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_114),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_46),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_41),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_136),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_77),
.Y(n_238)
);

INVxp67_ASAP7_75t_SL g239 ( 
.A(n_169),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_24),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_76),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_5),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_176),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_96),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_149),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_74),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_109),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_156),
.Y(n_248)
);

BUFx2_ASAP7_75t_SL g249 ( 
.A(n_29),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_18),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_40),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_56),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_129),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_86),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_24),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_49),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_128),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_23),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_67),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_119),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_11),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_62),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_110),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_7),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_137),
.Y(n_267)
);

NOR2xp67_ASAP7_75t_L g268 ( 
.A(n_8),
.B(n_95),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_78),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_151),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_43),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_177),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_121),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_139),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_66),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_142),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_173),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_171),
.Y(n_279)
);

HB1xp67_ASAP7_75t_L g280 ( 
.A(n_21),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_6),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_130),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_33),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_157),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_48),
.Y(n_285)
);

BUFx3_ASAP7_75t_L g286 ( 
.A(n_16),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_53),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_14),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_183),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_220),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_284),
.B(n_0),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_183),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_284),
.B(n_0),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_280),
.B(n_2),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_280),
.Y(n_295)
);

OAI21x1_ASAP7_75t_L g296 ( 
.A1(n_227),
.A2(n_81),
.B(n_170),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_203),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_287),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_265),
.B(n_2),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_286),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_182),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_180),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_185),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_258),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_181),
.B(n_7),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_180),
.Y(n_307)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

AOI22x1_ASAP7_75t_SL g309 ( 
.A1(n_201),
.A2(n_216),
.B1(n_232),
.B2(n_215),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_195),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_251),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_180),
.Y(n_312)
);

OA21x2_ASAP7_75t_L g313 ( 
.A1(n_178),
.A2(n_88),
.B(n_167),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_256),
.B(n_9),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_196),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_185),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_190),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g318 ( 
.A(n_195),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_196),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_10),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_281),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_196),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_233),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g324 ( 
.A(n_250),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_179),
.A2(n_89),
.B(n_165),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_266),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_233),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_196),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_205),
.Y(n_329)
);

INVx5_ASAP7_75t_L g330 ( 
.A(n_206),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_283),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_205),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_269),
.B(n_12),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_184),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_197),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_213),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g337 ( 
.A(n_262),
.Y(n_337)
);

INVx6_ASAP7_75t_L g338 ( 
.A(n_206),
.Y(n_338)
);

OA21x2_ASAP7_75t_L g339 ( 
.A1(n_192),
.A2(n_90),
.B(n_164),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_288),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_225),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_194),
.B(n_198),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_249),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_200),
.B(n_15),
.Y(n_344)
);

AND2x4_ASAP7_75t_L g345 ( 
.A(n_225),
.B(n_16),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_206),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_207),
.B(n_17),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_206),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_208),
.B(n_17),
.Y(n_349)
);

INVx3_ASAP7_75t_L g350 ( 
.A(n_233),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_254),
.Y(n_351)
);

INVx5_ASAP7_75t_L g352 ( 
.A(n_214),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_214),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_211),
.B(n_19),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_212),
.B(n_20),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_217),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_221),
.B(n_222),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_224),
.B(n_226),
.Y(n_358)
);

AOI22xp33_ASAP7_75t_SL g359 ( 
.A1(n_343),
.A2(n_246),
.B1(n_223),
.B2(n_253),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_345),
.B(n_228),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_299),
.Y(n_361)
);

CKINVDCx6p67_ASAP7_75t_R g362 ( 
.A(n_318),
.Y(n_362)
);

NAND3xp33_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_233),
.C(n_230),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_295),
.B(n_242),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_235),
.Y(n_365)
);

BUFx10_ASAP7_75t_L g366 ( 
.A(n_297),
.Y(n_366)
);

AND2x6_ASAP7_75t_L g367 ( 
.A(n_345),
.B(n_267),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_299),
.Y(n_368)
);

HB1xp67_ASAP7_75t_L g369 ( 
.A(n_324),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_300),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g371 ( 
.A(n_334),
.B(n_237),
.Y(n_371)
);

OR2x2_ASAP7_75t_L g372 ( 
.A(n_308),
.B(n_267),
.Y(n_372)
);

AOI22xp33_ASAP7_75t_L g373 ( 
.A1(n_289),
.A2(n_218),
.B1(n_255),
.B2(n_273),
.Y(n_373)
);

CKINVDCx6p67_ASAP7_75t_R g374 ( 
.A(n_318),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_301),
.Y(n_375)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_301),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_301),
.Y(n_377)
);

OR2x2_ASAP7_75t_L g378 ( 
.A(n_337),
.B(n_238),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_340),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_298),
.Y(n_380)
);

BUFx6f_ASAP7_75t_SL g381 ( 
.A(n_310),
.Y(n_381)
);

INVxp33_ASAP7_75t_L g382 ( 
.A(n_294),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_317),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_241),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_298),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_326),
.A2(n_264),
.B1(n_239),
.B2(n_244),
.Y(n_386)
);

OR2x6_ASAP7_75t_L g387 ( 
.A(n_305),
.B(n_268),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_289),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_307),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_307),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_342),
.B(n_252),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_292),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_R g393 ( 
.A(n_317),
.B(n_188),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_332),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_292),
.Y(n_395)
);

NAND2xp33_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_189),
.Y(n_396)
);

INVx4_ASAP7_75t_L g397 ( 
.A(n_304),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_304),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_307),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_331),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_335),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_302),
.B(n_257),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_191),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_351),
.B(n_193),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_302),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_316),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_312),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_291),
.Y(n_409)
);

AND3x2_ASAP7_75t_L g410 ( 
.A(n_293),
.B(n_199),
.C(n_261),
.Y(n_410)
);

BUFx6f_ASAP7_75t_SL g411 ( 
.A(n_309),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_316),
.B(n_276),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_329),
.B(n_341),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_358),
.B(n_277),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_312),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_312),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_329),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_312),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_341),
.B(n_278),
.Y(n_419)
);

BUFx3_ASAP7_75t_L g420 ( 
.A(n_303),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_306),
.Y(n_421)
);

NAND3xp33_ASAP7_75t_L g422 ( 
.A(n_333),
.B(n_279),
.C(n_285),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_315),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_354),
.A2(n_320),
.B1(n_314),
.B2(n_355),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_333),
.B(n_202),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_303),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_323),
.B(n_327),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_315),
.Y(n_428)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_344),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_315),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_347),
.B(n_282),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_349),
.B(n_214),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_319),
.Y(n_434)
);

CKINVDCx6p67_ASAP7_75t_R g435 ( 
.A(n_330),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_353),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_353),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_L g438 ( 
.A1(n_313),
.A2(n_260),
.B1(n_271),
.B2(n_282),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_336),
.B(n_204),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_323),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_330),
.Y(n_441)
);

BUFx8_ASAP7_75t_SL g442 ( 
.A(n_336),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_303),
.B(n_260),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_311),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_323),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_327),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_338),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_338),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_350),
.Y(n_449)
);

INVx4_ASAP7_75t_L g450 ( 
.A(n_330),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_303),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_296),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

NOR2xp33_ASAP7_75t_L g454 ( 
.A(n_409),
.B(n_187),
.Y(n_454)
);

NAND2xp33_ASAP7_75t_L g455 ( 
.A(n_367),
.B(n_209),
.Y(n_455)
);

AND2x4_ASAP7_75t_L g456 ( 
.A(n_429),
.B(n_296),
.Y(n_456)
);

A2O1A1Ixp33_ASAP7_75t_L g457 ( 
.A1(n_391),
.A2(n_186),
.B(n_350),
.C(n_263),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_424),
.B(n_210),
.Y(n_458)
);

O2A1O1Ixp33_ASAP7_75t_L g459 ( 
.A1(n_370),
.A2(n_350),
.B(n_325),
.C(n_339),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_444),
.A2(n_272),
.B1(n_229),
.B2(n_231),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_372),
.B(n_219),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_364),
.B(n_234),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_424),
.B(n_236),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_414),
.B(n_243),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_414),
.B(n_245),
.Y(n_465)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_382),
.A2(n_379),
.B1(n_361),
.B2(n_368),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_398),
.B(n_401),
.Y(n_467)
);

NAND2xp33_ASAP7_75t_L g468 ( 
.A(n_367),
.B(n_247),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_425),
.B(n_248),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_362),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_369),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_360),
.B(n_270),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_369),
.B(n_274),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_365),
.B(n_275),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_375),
.Y(n_475)
);

INVx2_ASAP7_75t_SL g476 ( 
.A(n_366),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_384),
.B(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_377),
.Y(n_478)
);

BUFx8_ASAP7_75t_L g479 ( 
.A(n_411),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_374),
.Y(n_480)
);

NAND3xp33_ASAP7_75t_L g481 ( 
.A(n_438),
.B(n_325),
.C(n_313),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_384),
.B(n_339),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g483 ( 
.A(n_397),
.B(n_260),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_404),
.B(n_303),
.Y(n_484)
);

NAND3xp33_ASAP7_75t_L g485 ( 
.A(n_438),
.B(n_373),
.C(n_371),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_380),
.Y(n_486)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_371),
.A2(n_352),
.B(n_338),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_431),
.A2(n_352),
.B(n_353),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_394),
.Y(n_489)
);

NOR2x1p5_ASAP7_75t_L g490 ( 
.A(n_439),
.B(n_442),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_373),
.B(n_422),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_383),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_405),
.B(n_396),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_385),
.B(n_352),
.Y(n_494)
);

NOR2xp67_ASAP7_75t_SL g495 ( 
.A(n_363),
.B(n_282),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_445),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_449),
.B(n_282),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_381),
.A2(n_353),
.B1(n_348),
.B2(n_346),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_447),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_448),
.Y(n_501)
);

AOI22xp33_ASAP7_75t_L g502 ( 
.A1(n_387),
.A2(n_348),
.B1(n_346),
.B2(n_328),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_388),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_392),
.Y(n_504)
);

INVxp67_ASAP7_75t_SL g505 ( 
.A(n_399),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_395),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_393),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_322),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_406),
.Y(n_509)
);

BUFx5_ASAP7_75t_L g510 ( 
.A(n_420),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_393),
.B(n_22),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_433),
.B(n_322),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_402),
.Y(n_514)
);

INVxp33_ASAP7_75t_L g515 ( 
.A(n_359),
.Y(n_515)
);

INVx3_ASAP7_75t_L g516 ( 
.A(n_417),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_413),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_403),
.B(n_322),
.Y(n_518)
);

AOI22xp33_ASAP7_75t_L g519 ( 
.A1(n_387),
.A2(n_348),
.B1(n_346),
.B2(n_328),
.Y(n_519)
);

NOR3xp33_ASAP7_75t_L g520 ( 
.A(n_386),
.B(n_22),
.C(n_23),
.Y(n_520)
);

OR2x2_ASAP7_75t_L g521 ( 
.A(n_387),
.B(n_25),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_403),
.B(n_412),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_412),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_419),
.B(n_36),
.Y(n_524)
);

AOI22xp33_ASAP7_75t_L g525 ( 
.A1(n_419),
.A2(n_443),
.B1(n_440),
.B2(n_446),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_411),
.A2(n_348),
.B1(n_346),
.B2(n_328),
.Y(n_526)
);

OAI221xp5_ASAP7_75t_L g527 ( 
.A1(n_427),
.A2(n_328),
.B1(n_27),
.B2(n_28),
.C(n_30),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_443),
.B(n_39),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_432),
.Y(n_529)
);

BUFx5_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_432),
.B(n_26),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_410),
.B(n_45),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_441),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_L g534 ( 
.A1(n_477),
.A2(n_450),
.B1(n_410),
.B2(n_451),
.Y(n_534)
);

OR2x6_ASAP7_75t_SL g535 ( 
.A(n_492),
.B(n_26),
.Y(n_535)
);

O2A1O1Ixp33_ASAP7_75t_L g536 ( 
.A1(n_491),
.A2(n_426),
.B(n_451),
.C(n_437),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_467),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_476),
.B(n_27),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_471),
.B(n_28),
.Y(n_539)
);

BUFx4f_ASAP7_75t_L g540 ( 
.A(n_499),
.Y(n_540)
);

BUFx2_ASAP7_75t_SL g541 ( 
.A(n_470),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_467),
.B(n_30),
.Y(n_542)
);

O2A1O1Ixp33_ASAP7_75t_L g543 ( 
.A1(n_458),
.A2(n_436),
.B(n_434),
.C(n_430),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_454),
.B(n_31),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_473),
.B(n_31),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_482),
.A2(n_456),
.B(n_493),
.Y(n_546)
);

AOI21x1_ASAP7_75t_L g547 ( 
.A1(n_456),
.A2(n_481),
.B(n_488),
.Y(n_547)
);

CKINVDCx10_ASAP7_75t_R g548 ( 
.A(n_479),
.Y(n_548)
);

OA21x2_ASAP7_75t_L g549 ( 
.A1(n_481),
.A2(n_428),
.B(n_423),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_461),
.B(n_34),
.Y(n_550)
);

CKINVDCx10_ASAP7_75t_R g551 ( 
.A(n_479),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_475),
.Y(n_552)
);

CKINVDCx10_ASAP7_75t_R g553 ( 
.A(n_480),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_L g554 ( 
.A1(n_466),
.A2(n_418),
.B1(n_416),
.B2(n_415),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_459),
.A2(n_416),
.B(n_415),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_514),
.B(n_34),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_499),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_462),
.B(n_35),
.Y(n_558)
);

BUFx12f_ASAP7_75t_L g559 ( 
.A(n_490),
.Y(n_559)
);

AOI21x1_ASAP7_75t_L g560 ( 
.A1(n_508),
.A2(n_408),
.B(n_400),
.Y(n_560)
);

OA22x2_ASAP7_75t_L g561 ( 
.A1(n_507),
.A2(n_35),
.B1(n_390),
.B2(n_389),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_464),
.B(n_50),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_465),
.B(n_52),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_515),
.B(n_163),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g565 ( 
.A(n_499),
.B(n_57),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_484),
.A2(n_59),
.B(n_61),
.Y(n_566)
);

O2A1O1Ixp5_ASAP7_75t_L g567 ( 
.A1(n_457),
.A2(n_63),
.B(n_64),
.C(n_68),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g568 ( 
.A1(n_505),
.A2(n_69),
.B(n_70),
.Y(n_568)
);

AOI21xp5_ASAP7_75t_L g569 ( 
.A1(n_455),
.A2(n_72),
.B(n_73),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_511),
.B(n_460),
.Y(n_570)
);

OAI21xp5_ASAP7_75t_L g571 ( 
.A1(n_485),
.A2(n_92),
.B(n_94),
.Y(n_571)
);

AOI21xp5_ASAP7_75t_L g572 ( 
.A1(n_468),
.A2(n_97),
.B(n_98),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g573 ( 
.A(n_527),
.B(n_99),
.C(n_101),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_516),
.B(n_161),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_486),
.B(n_102),
.Y(n_575)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_460),
.Y(n_576)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_522),
.A2(n_103),
.B(n_104),
.Y(n_577)
);

AO21x1_ASAP7_75t_L g578 ( 
.A1(n_513),
.A2(n_105),
.B(n_106),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_517),
.A2(n_107),
.B(n_108),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_503),
.A2(n_111),
.B1(n_112),
.B2(n_116),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_504),
.Y(n_581)
);

HB1xp67_ASAP7_75t_L g582 ( 
.A(n_506),
.Y(n_582)
);

INVxp67_ASAP7_75t_SL g583 ( 
.A(n_483),
.Y(n_583)
);

AND2x2_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_117),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_478),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_523),
.A2(n_118),
.B1(n_122),
.B2(n_124),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_472),
.A2(n_125),
.B(n_126),
.Y(n_587)
);

AOI21xp5_ASAP7_75t_L g588 ( 
.A1(n_474),
.A2(n_135),
.B(n_138),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_489),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_L g590 ( 
.A1(n_509),
.A2(n_512),
.B1(n_469),
.B2(n_453),
.Y(n_590)
);

OR2x6_ASAP7_75t_L g591 ( 
.A(n_526),
.B(n_153),
.Y(n_591)
);

AND2x4_ASAP7_75t_L g592 ( 
.A(n_529),
.B(n_533),
.Y(n_592)
);

NAND3xp33_ASAP7_75t_L g593 ( 
.A(n_502),
.B(n_519),
.C(n_532),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_500),
.Y(n_594)
);

AOI21xp5_ASAP7_75t_L g595 ( 
.A1(n_518),
.A2(n_496),
.B(n_494),
.Y(n_595)
);

OAI21x1_ASAP7_75t_L g596 ( 
.A1(n_487),
.A2(n_525),
.B(n_531),
.Y(n_596)
);

AOI21xp5_ASAP7_75t_L g597 ( 
.A1(n_487),
.A2(n_497),
.B(n_528),
.Y(n_597)
);

AO21x1_ASAP7_75t_L g598 ( 
.A1(n_524),
.A2(n_498),
.B(n_501),
.Y(n_598)
);

BUFx12f_ASAP7_75t_L g599 ( 
.A(n_510),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_495),
.A2(n_481),
.B(n_482),
.Y(n_600)
);

AND2x4_ASAP7_75t_L g601 ( 
.A(n_530),
.B(n_476),
.Y(n_601)
);

AOI21xp5_ASAP7_75t_L g602 ( 
.A1(n_530),
.A2(n_452),
.B(n_482),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_540),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_602),
.A2(n_546),
.B(n_600),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_537),
.B(n_570),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_576),
.A2(n_542),
.B1(n_582),
.B2(n_581),
.Y(n_606)
);

AO22x2_ASAP7_75t_L g607 ( 
.A1(n_538),
.A2(n_584),
.B1(n_590),
.B2(n_564),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_601),
.B(n_557),
.Y(n_608)
);

AO31x2_ASAP7_75t_L g609 ( 
.A1(n_598),
.A2(n_578),
.A3(n_555),
.B(n_569),
.Y(n_609)
);

BUFx5_ASAP7_75t_L g610 ( 
.A(n_599),
.Y(n_610)
);

INVx1_ASAP7_75t_SL g611 ( 
.A(n_538),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_540),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_547),
.A2(n_560),
.B(n_549),
.Y(n_613)
);

AO31x2_ASAP7_75t_L g614 ( 
.A1(n_572),
.A2(n_586),
.A3(n_568),
.B(n_587),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_556),
.B(n_545),
.Y(n_615)
);

A2O1A1Ixp33_ASAP7_75t_L g616 ( 
.A1(n_543),
.A2(n_550),
.B(n_585),
.C(n_552),
.Y(n_616)
);

OAI22xp5_ASAP7_75t_SL g617 ( 
.A1(n_559),
.A2(n_535),
.B1(n_551),
.B2(n_548),
.Y(n_617)
);

AO31x2_ASAP7_75t_L g618 ( 
.A1(n_588),
.A2(n_597),
.A3(n_580),
.B(n_579),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_539),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_596),
.A2(n_595),
.B(n_536),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_583),
.A2(n_562),
.B(n_563),
.Y(n_621)
);

AO31x2_ASAP7_75t_L g622 ( 
.A1(n_577),
.A2(n_566),
.A3(n_574),
.B(n_575),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_541),
.B(n_544),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_553),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_553),
.Y(n_625)
);

NAND3xp33_ASAP7_75t_L g626 ( 
.A(n_573),
.B(n_567),
.C(n_593),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_592),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_592),
.B(n_534),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_561),
.Y(n_629)
);

BUFx3_ASAP7_75t_L g630 ( 
.A(n_565),
.Y(n_630)
);

BUFx4f_ASAP7_75t_SL g631 ( 
.A(n_548),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_594),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_589),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_551),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_591),
.Y(n_635)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_591),
.A2(n_537),
.B1(n_576),
.B2(n_542),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_537),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_547),
.A2(n_602),
.B(n_600),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_537),
.B(n_471),
.Y(n_639)
);

OAI21x1_ASAP7_75t_L g640 ( 
.A1(n_547),
.A2(n_602),
.B(n_600),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_537),
.B(n_409),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_537),
.Y(n_642)
);

OR2x6_ASAP7_75t_L g643 ( 
.A(n_541),
.B(n_559),
.Y(n_643)
);

OAI21xp5_ASAP7_75t_L g644 ( 
.A1(n_546),
.A2(n_602),
.B(n_485),
.Y(n_644)
);

AO32x2_ASAP7_75t_L g645 ( 
.A1(n_534),
.A2(n_590),
.A3(n_586),
.B1(n_554),
.B2(n_526),
.Y(n_645)
);

OA21x2_ASAP7_75t_L g646 ( 
.A1(n_600),
.A2(n_481),
.B(n_571),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_537),
.B(n_409),
.Y(n_647)
);

INVx6_ASAP7_75t_SL g648 ( 
.A(n_538),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_537),
.B(n_409),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_537),
.Y(n_650)
);

O2A1O1Ixp33_ASAP7_75t_L g651 ( 
.A1(n_576),
.A2(n_491),
.B(n_477),
.C(n_457),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_537),
.B(n_409),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_537),
.B(n_409),
.Y(n_653)
);

NAND3x1_ASAP7_75t_L g654 ( 
.A(n_548),
.B(n_520),
.C(n_551),
.Y(n_654)
);

INVx4_ASAP7_75t_SL g655 ( 
.A(n_559),
.Y(n_655)
);

OR2x2_ASAP7_75t_L g656 ( 
.A(n_537),
.B(n_471),
.Y(n_656)
);

OA21x2_ASAP7_75t_L g657 ( 
.A1(n_600),
.A2(n_481),
.B(n_571),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_546),
.A2(n_602),
.B(n_485),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_537),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_537),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_537),
.B(n_409),
.Y(n_661)
);

NOR2xp33_ASAP7_75t_L g662 ( 
.A(n_576),
.B(n_514),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_537),
.B(n_471),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_537),
.B(n_409),
.Y(n_664)
);

BUFx2_ASAP7_75t_R g665 ( 
.A(n_535),
.Y(n_665)
);

AO31x2_ASAP7_75t_L g666 ( 
.A1(n_598),
.A2(n_578),
.A3(n_602),
.B(n_546),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_537),
.B(n_409),
.Y(n_667)
);

HB1xp67_ASAP7_75t_L g668 ( 
.A(n_537),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_537),
.B(n_409),
.Y(n_669)
);

OR2x6_ASAP7_75t_L g670 ( 
.A(n_541),
.B(n_559),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_537),
.B(n_409),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_537),
.B(n_471),
.Y(n_672)
);

AO31x2_ASAP7_75t_L g673 ( 
.A1(n_598),
.A2(n_578),
.A3(n_602),
.B(n_546),
.Y(n_673)
);

AND3x4_ASAP7_75t_L g674 ( 
.A(n_548),
.B(n_551),
.C(n_480),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_546),
.A2(n_602),
.B(n_485),
.Y(n_675)
);

AOI21xp5_ASAP7_75t_L g676 ( 
.A1(n_602),
.A2(n_546),
.B(n_452),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_537),
.B(n_601),
.Y(n_677)
);

BUFx2_ASAP7_75t_L g678 ( 
.A(n_537),
.Y(n_678)
);

AOI211x1_ASAP7_75t_L g679 ( 
.A1(n_537),
.A2(n_491),
.B(n_463),
.C(n_458),
.Y(n_679)
);

AOI21xp5_ASAP7_75t_L g680 ( 
.A1(n_602),
.A2(n_546),
.B(n_452),
.Y(n_680)
);

A2O1A1Ixp33_ASAP7_75t_L g681 ( 
.A1(n_537),
.A2(n_542),
.B(n_546),
.C(n_558),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_537),
.B(n_409),
.Y(n_682)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_537),
.B(n_471),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_546),
.A2(n_602),
.B(n_485),
.Y(n_684)
);

OA21x2_ASAP7_75t_L g685 ( 
.A1(n_600),
.A2(n_481),
.B(n_571),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_537),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_537),
.B(n_601),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_548),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_537),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_576),
.B(n_514),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_537),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_537),
.B(n_409),
.Y(n_692)
);

OAI21xp33_ASAP7_75t_L g693 ( 
.A1(n_537),
.A2(n_477),
.B(n_454),
.Y(n_693)
);

OA21x2_ASAP7_75t_L g694 ( 
.A1(n_613),
.A2(n_640),
.B(n_638),
.Y(n_694)
);

AO21x2_ASAP7_75t_L g695 ( 
.A1(n_620),
.A2(n_604),
.B(n_626),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_641),
.B(n_652),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_678),
.B(n_668),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_647),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_650),
.Y(n_699)
);

AO21x2_ASAP7_75t_L g700 ( 
.A1(n_644),
.A2(n_684),
.B(n_658),
.Y(n_700)
);

OR2x6_ASAP7_75t_L g701 ( 
.A(n_643),
.B(n_670),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_649),
.B(n_653),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_643),
.B(n_670),
.Y(n_703)
);

AND2x2_ASAP7_75t_L g704 ( 
.A(n_661),
.B(n_664),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_659),
.B(n_660),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_667),
.B(n_669),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_677),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_671),
.B(n_682),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_637),
.Y(n_709)
);

AND2x4_ASAP7_75t_L g710 ( 
.A(n_687),
.B(n_642),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_676),
.A2(n_680),
.B(n_675),
.Y(n_711)
);

BUFx2_ASAP7_75t_L g712 ( 
.A(n_648),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_692),
.Y(n_713)
);

AOI21xp5_ASAP7_75t_L g714 ( 
.A1(n_621),
.A2(n_681),
.B(n_636),
.Y(n_714)
);

CKINVDCx6p67_ASAP7_75t_R g715 ( 
.A(n_634),
.Y(n_715)
);

NAND3xp33_ASAP7_75t_L g716 ( 
.A(n_679),
.B(n_651),
.C(n_693),
.Y(n_716)
);

OAI21x1_ASAP7_75t_L g717 ( 
.A1(n_646),
.A2(n_685),
.B(n_657),
.Y(n_717)
);

OA21x2_ASAP7_75t_L g718 ( 
.A1(n_616),
.A2(n_628),
.B(n_629),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_605),
.B(n_672),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_SL g720 ( 
.A1(n_607),
.A2(n_606),
.B1(n_611),
.B2(n_617),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_686),
.B(n_691),
.Y(n_721)
);

INVx1_ASAP7_75t_SL g722 ( 
.A(n_648),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_689),
.Y(n_723)
);

AO21x2_ASAP7_75t_L g724 ( 
.A1(n_609),
.A2(n_673),
.B(n_666),
.Y(n_724)
);

OR2x6_ASAP7_75t_L g725 ( 
.A(n_687),
.B(n_683),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_631),
.Y(n_726)
);

AO21x1_ASAP7_75t_L g727 ( 
.A1(n_627),
.A2(n_619),
.B(n_662),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_656),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_630),
.B(n_615),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_633),
.Y(n_730)
);

INVx1_ASAP7_75t_SL g731 ( 
.A(n_610),
.Y(n_731)
);

AOI21xp5_ASAP7_75t_L g732 ( 
.A1(n_607),
.A2(n_639),
.B(n_663),
.Y(n_732)
);

OAI21x1_ASAP7_75t_L g733 ( 
.A1(n_666),
.A2(n_673),
.B(n_609),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_666),
.A2(n_673),
.B(n_618),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_632),
.Y(n_735)
);

AO31x2_ASAP7_75t_L g736 ( 
.A1(n_690),
.A2(n_618),
.A3(n_645),
.B(n_614),
.Y(n_736)
);

AO31x2_ASAP7_75t_L g737 ( 
.A1(n_618),
.A2(n_645),
.A3(n_614),
.B(n_622),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_622),
.A2(n_608),
.A3(n_623),
.B(n_654),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_608),
.Y(n_739)
);

AO21x2_ASAP7_75t_L g740 ( 
.A1(n_622),
.A2(n_612),
.B(n_665),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_603),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_674),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_655),
.Y(n_743)
);

INVx3_ASAP7_75t_L g744 ( 
.A(n_688),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_624),
.B(n_625),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_674),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_641),
.Y(n_747)
);

OAI22xp33_ASAP7_75t_L g748 ( 
.A1(n_635),
.A2(n_636),
.B1(n_537),
.B2(n_678),
.Y(n_748)
);

HB1xp67_ASAP7_75t_L g749 ( 
.A(n_668),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_650),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_641),
.B(n_652),
.Y(n_751)
);

NAND2x1p5_ASAP7_75t_L g752 ( 
.A(n_678),
.B(n_540),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

NAND3xp33_ASAP7_75t_SL g754 ( 
.A(n_635),
.B(n_335),
.C(n_317),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_641),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_641),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_641),
.B(n_652),
.Y(n_757)
);

OAI21xp5_ASAP7_75t_L g758 ( 
.A1(n_681),
.A2(n_485),
.B(n_693),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_641),
.Y(n_759)
);

NAND2x1p5_ASAP7_75t_L g760 ( 
.A(n_678),
.B(n_540),
.Y(n_760)
);

NAND2x1p5_ASAP7_75t_L g761 ( 
.A(n_678),
.B(n_540),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_641),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_641),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_641),
.Y(n_764)
);

INVx4_ASAP7_75t_SL g765 ( 
.A(n_701),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_699),
.B(n_750),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_699),
.B(n_750),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_747),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_749),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_749),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_709),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_697),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_694),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_696),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_755),
.Y(n_775)
);

AND2x4_ASAP7_75t_L g776 ( 
.A(n_738),
.B(n_710),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_756),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_705),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_759),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_704),
.B(n_708),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_762),
.Y(n_781)
);

OR2x6_ASAP7_75t_L g782 ( 
.A(n_701),
.B(n_703),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_763),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_764),
.Y(n_784)
);

AO21x2_ASAP7_75t_L g785 ( 
.A1(n_714),
.A2(n_711),
.B(n_758),
.Y(n_785)
);

OR2x6_ASAP7_75t_L g786 ( 
.A(n_701),
.B(n_703),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_723),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_718),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_698),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_713),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_720),
.A2(n_748),
.B1(n_751),
.B2(n_727),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_757),
.B(n_706),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_719),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_721),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_730),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_702),
.B(n_728),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_735),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_718),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_718),
.B(n_725),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_748),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_754),
.B(n_729),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_720),
.B(n_707),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_726),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_752),
.Y(n_804)
);

CKINVDCx20_ASAP7_75t_R g805 ( 
.A(n_726),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_736),
.Y(n_806)
);

OA21x2_ASAP7_75t_L g807 ( 
.A1(n_714),
.A2(n_734),
.B(n_733),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_766),
.B(n_767),
.Y(n_808)
);

AND2x2_ASAP7_75t_L g809 ( 
.A(n_766),
.B(n_724),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_767),
.B(n_724),
.Y(n_810)
);

AOI33xp33_ASAP7_75t_L g811 ( 
.A1(n_791),
.A2(n_722),
.A3(n_745),
.B1(n_743),
.B2(n_739),
.B3(n_731),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_771),
.B(n_700),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_769),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_773),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_770),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_765),
.B(n_746),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_800),
.A2(n_703),
.B1(n_716),
.B2(n_732),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_799),
.B(n_737),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_799),
.B(n_717),
.Y(n_819)
);

BUFx2_ASAP7_75t_L g820 ( 
.A(n_778),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_806),
.Y(n_821)
);

INVx5_ASAP7_75t_L g822 ( 
.A(n_782),
.Y(n_822)
);

HB1xp67_ASAP7_75t_L g823 ( 
.A(n_772),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_794),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_776),
.B(n_695),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_776),
.B(n_695),
.Y(n_826)
);

OR2x2_ASAP7_75t_L g827 ( 
.A(n_780),
.B(n_738),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_792),
.B(n_746),
.Y(n_828)
);

OAI211xp5_ASAP7_75t_L g829 ( 
.A1(n_801),
.A2(n_742),
.B(n_729),
.C(n_754),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_824),
.B(n_789),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_818),
.B(n_788),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_821),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_808),
.B(n_790),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_818),
.B(n_798),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_814),
.Y(n_835)
);

INVxp33_ASAP7_75t_L g836 ( 
.A(n_828),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_811),
.B(n_765),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_809),
.B(n_807),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_820),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_810),
.B(n_807),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_808),
.B(n_787),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_823),
.B(n_793),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_813),
.B(n_815),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_827),
.B(n_785),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_815),
.B(n_768),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_810),
.B(n_819),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_836),
.A2(n_802),
.B1(n_817),
.B2(n_822),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_846),
.B(n_825),
.Y(n_848)
);

NOR2xp67_ASAP7_75t_L g849 ( 
.A(n_837),
.B(n_742),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_835),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_832),
.Y(n_851)
);

NOR3xp33_ASAP7_75t_L g852 ( 
.A(n_843),
.B(n_829),
.C(n_796),
.Y(n_852)
);

INVxp67_ASAP7_75t_L g853 ( 
.A(n_839),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_830),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_831),
.B(n_826),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_833),
.B(n_841),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_831),
.B(n_826),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_845),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_842),
.B(n_827),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_832),
.Y(n_860)
);

OR2x2_ASAP7_75t_L g861 ( 
.A(n_844),
.B(n_812),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_834),
.B(n_819),
.Y(n_862)
);

OAI21xp5_ASAP7_75t_L g863 ( 
.A1(n_849),
.A2(n_829),
.B(n_817),
.Y(n_863)
);

OR2x2_ASAP7_75t_L g864 ( 
.A(n_861),
.B(n_844),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_858),
.B(n_838),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_854),
.B(n_838),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_851),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_853),
.Y(n_868)
);

INVxp67_ASAP7_75t_SL g869 ( 
.A(n_850),
.Y(n_869)
);

HB1xp67_ASAP7_75t_L g870 ( 
.A(n_861),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_851),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_862),
.B(n_840),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_860),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_870),
.Y(n_874)
);

AOI22xp5_ASAP7_75t_L g875 ( 
.A1(n_866),
.A2(n_852),
.B1(n_859),
.B2(n_847),
.Y(n_875)
);

OR2x2_ASAP7_75t_L g876 ( 
.A(n_864),
.B(n_862),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_872),
.B(n_855),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_872),
.B(n_855),
.Y(n_878)
);

INVxp67_ASAP7_75t_SL g879 ( 
.A(n_869),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_864),
.Y(n_880)
);

AND2x2_ASAP7_75t_L g881 ( 
.A(n_868),
.B(n_848),
.Y(n_881)
);

NAND2x1_ASAP7_75t_L g882 ( 
.A(n_863),
.B(n_839),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_873),
.B(n_857),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_873),
.B(n_857),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_875),
.B(n_865),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_883),
.Y(n_886)
);

AOI21x1_ASAP7_75t_L g887 ( 
.A1(n_882),
.A2(n_816),
.B(n_786),
.Y(n_887)
);

AOI221xp5_ASAP7_75t_L g888 ( 
.A1(n_874),
.A2(n_856),
.B1(n_774),
.B2(n_867),
.C(n_871),
.Y(n_888)
);

AOI211xp5_ASAP7_75t_L g889 ( 
.A1(n_885),
.A2(n_879),
.B(n_803),
.C(n_802),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_888),
.A2(n_883),
.B(n_884),
.Y(n_890)
);

OAI211xp5_ASAP7_75t_L g891 ( 
.A1(n_887),
.A2(n_803),
.B(n_805),
.C(n_744),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_891),
.B(n_744),
.C(n_889),
.Y(n_892)
);

NOR2xp33_ASAP7_75t_L g893 ( 
.A(n_890),
.B(n_886),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_893),
.Y(n_894)
);

NAND4xp25_ASAP7_75t_L g895 ( 
.A(n_892),
.B(n_753),
.C(n_712),
.D(n_715),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_R g896 ( 
.A(n_894),
.B(n_805),
.Y(n_896)
);

AOI221xp5_ASAP7_75t_L g897 ( 
.A1(n_895),
.A2(n_880),
.B1(n_795),
.B2(n_881),
.C(n_797),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_896),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_897),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_898),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_899),
.B(n_877),
.Y(n_901)
);

OAI21xp5_ASAP7_75t_L g902 ( 
.A1(n_900),
.A2(n_786),
.B(n_782),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_901),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_900),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_900),
.B(n_765),
.Y(n_905)
);

OAI22xp5_ASAP7_75t_L g906 ( 
.A1(n_904),
.A2(n_786),
.B1(n_782),
.B2(n_876),
.Y(n_906)
);

AOI22x1_ASAP7_75t_L g907 ( 
.A1(n_903),
.A2(n_760),
.B1(n_761),
.B2(n_741),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_SL g908 ( 
.A1(n_902),
.A2(n_761),
.B(n_741),
.Y(n_908)
);

AOI21xp33_ASAP7_75t_SL g909 ( 
.A1(n_905),
.A2(n_740),
.B(n_804),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_904),
.Y(n_910)
);

OAI21xp5_ASAP7_75t_L g911 ( 
.A1(n_910),
.A2(n_732),
.B(n_878),
.Y(n_911)
);

AOI222xp33_ASAP7_75t_L g912 ( 
.A1(n_906),
.A2(n_784),
.B1(n_783),
.B2(n_781),
.C1(n_779),
.C2(n_777),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_911),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_912),
.B(n_909),
.Y(n_914)
);

OA21x2_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_907),
.B(n_908),
.Y(n_915)
);

AOI21xp33_ASAP7_75t_SL g916 ( 
.A1(n_915),
.A2(n_913),
.B(n_775),
.Y(n_916)
);


endmodule