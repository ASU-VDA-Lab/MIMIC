module real_jpeg_16987_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

INVx1_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_0),
.Y(n_67)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_0),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_1),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_1),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_22),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_35),
.Y(n_34)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_2),
.B(n_42),
.Y(n_41)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_2),
.B(n_63),
.Y(n_62)
);

NAND2x1_ASAP7_75t_L g80 ( 
.A(n_2),
.B(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_2),
.B(n_90),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_2),
.B(n_131),
.Y(n_130)
);

NAND2x1_ASAP7_75t_L g179 ( 
.A(n_2),
.B(n_180),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_3),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_3),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_4),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_4),
.B(n_58),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_4),
.B(n_134),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_7),
.Y(n_171)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_7),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_8),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_8),
.B(n_32),
.Y(n_31)
);

AND2x4_ASAP7_75t_L g46 ( 
.A(n_8),
.B(n_47),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_8),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_8),
.B(n_120),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g168 ( 
.A(n_8),
.B(n_169),
.Y(n_168)
);

AND2x2_ASAP7_75t_SL g217 ( 
.A(n_8),
.B(n_180),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_9),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_9),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g122 ( 
.A(n_10),
.Y(n_122)
);

BUFx8_ASAP7_75t_L g180 ( 
.A(n_11),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_193),
.Y(n_12)
);

OAI21x1_ASAP7_75t_L g13 ( 
.A1(n_14),
.A2(n_156),
.B(n_192),
.Y(n_13)
);

AOI21x1_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_108),
.B(n_155),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_69),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_16),
.B(n_69),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_39),
.C(n_55),
.Y(n_16)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_17),
.B(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_30),
.Y(n_17)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_18),
.Y(n_146)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_19),
.A2(n_31),
.B(n_38),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_20),
.A2(n_21),
.B1(n_104),
.B2(n_107),
.Y(n_103)
);

INVx2_ASAP7_75t_SL g20 ( 
.A(n_21),
.Y(n_20)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_34),
.B(n_36),
.Y(n_33)
);

NAND2x1p5_ASAP7_75t_L g36 ( 
.A(n_21),
.B(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_24),
.Y(n_135)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_24),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_25),
.A2(n_133),
.B1(n_136),
.B2(n_137),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_25),
.Y(n_137)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_29),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

O2A1O1Ixp33_ASAP7_75t_R g129 ( 
.A1(n_31),
.A2(n_130),
.B(n_132),
.C(n_138),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_31),
.B(n_130),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_31),
.A2(n_37),
.B1(n_130),
.B2(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_34),
.A2(n_119),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_34),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_34),
.B(n_133),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_36),
.B(n_73),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_36),
.B(n_74),
.C(n_80),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_39),
.A2(n_55),
.B1(n_56),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_39),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.C(n_50),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_40),
.A2(n_41),
.B1(n_50),
.B2(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_41),
.B(n_206),
.Y(n_205)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_45),
.A2(n_46),
.B1(n_87),
.B2(n_97),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_45),
.A2(n_46),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_46),
.A2(n_89),
.B(n_91),
.C(n_138),
.Y(n_163)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_49),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g116 ( 
.A(n_50),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_50),
.A2(n_74),
.B1(n_82),
.B2(n_116),
.Y(n_202)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_105),
.Y(n_104)
);

OR2x2_ASAP7_75t_L g187 ( 
.A(n_51),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_68),
.Y(n_56)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_57),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_57),
.B(n_62),
.C(n_101),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_64),
.Y(n_189)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_65),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_65),
.A2(n_101),
.B1(n_167),
.B2(n_173),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_85),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_72),
.B1(n_83),
.B2(n_84),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_72),
.B(n_83),
.C(n_85),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_79),
.B1(n_80),
.B2(n_82),
.Y(n_73)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_98),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_86),
.B(n_99),
.C(n_103),
.Y(n_160)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_89),
.B1(n_91),
.B2(n_96),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_88),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_88),
.B(n_145),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_88),
.B(n_130),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_89),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g201 ( 
.A(n_89),
.B(n_130),
.C(n_179),
.Y(n_201)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_91),
.Y(n_96)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_99),
.A2(n_100),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_101),
.B(n_133),
.C(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_104),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_104),
.A2(n_107),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_107),
.B(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_107),
.A2(n_118),
.B(n_119),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_127),
.B(n_154),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_110),
.B(n_113),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_118),
.C(n_123),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_114),
.B(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_115),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_118),
.A2(n_123),
.B1(n_124),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_142),
.B(n_153),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_139),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_130),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_130),
.A2(n_151),
.B1(n_205),
.B2(n_210),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_132),
.B(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_133),
.A2(n_136),
.B1(n_168),
.B2(n_172),
.Y(n_167)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_149),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_148),
.B(n_152),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_146),
.B(n_147),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_158),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_160),
.B(n_161),
.C(n_174),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_166),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_163),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_164),
.B(n_166),
.C(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_167),
.Y(n_173)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_168),
.Y(n_172)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_191),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_182),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_176),
.B(n_182),
.C(n_191),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_176)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_177),
.Y(n_181)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_187),
.B(n_190),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_183),
.B(n_187),
.Y(n_190)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_190),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_223)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_228),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_195),
.B(n_196),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_213),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_211),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_227),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_223),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_218),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);


endmodule