module fake_aes_5788_n_33 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AND2x2_ASAP7_75t_SL g13 ( .A(n_6), .B(n_1), .Y(n_13) );
INVx5_ASAP7_75t_L g14 ( .A(n_2), .Y(n_14) );
AND2x4_ASAP7_75t_L g15 ( .A(n_3), .B(n_10), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_1), .Y(n_16) );
AOI22xp5_ASAP7_75t_L g17 ( .A1(n_2), .A2(n_8), .B1(n_11), .B2(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_14), .B(n_0), .Y(n_18) );
INVx1_ASAP7_75t_SL g19 ( .A(n_13), .Y(n_19) );
INVx3_ASAP7_75t_SL g20 ( .A(n_19), .Y(n_20) );
OAI22xp33_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_17), .B1(n_16), .B2(n_14), .Y(n_21) );
BUFx3_ASAP7_75t_L g22 ( .A(n_20), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
XOR2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
NOR2xp33_ASAP7_75t_L g25 ( .A(n_23), .B(n_22), .Y(n_25) );
OAI21xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_21), .B(n_17), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_24), .A2(n_15), .B1(n_18), .B2(n_14), .Y(n_27) );
NAND4xp25_ASAP7_75t_SL g28 ( .A(n_27), .B(n_12), .C(n_4), .D(n_3), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_26), .Y(n_29) );
OAI21xp5_ASAP7_75t_L g30 ( .A1(n_29), .A2(n_15), .B(n_4), .Y(n_30) );
BUFx6f_ASAP7_75t_L g31 ( .A(n_28), .Y(n_31) );
INVx1_ASAP7_75t_L g32 ( .A(n_31), .Y(n_32) );
AO221x2_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_30), .B1(n_31), .B2(n_7), .C(n_5), .Y(n_33) );
endmodule