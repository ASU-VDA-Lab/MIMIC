module real_jpeg_17001_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_332;
wire n_149;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_525;
wire n_288;
wire n_78;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_543;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_537;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_549;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_52),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_0),
.A2(n_66),
.B1(n_214),
.B2(n_218),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_0),
.A2(n_66),
.B1(n_272),
.B2(n_274),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_1),
.A2(n_71),
.B1(n_77),
.B2(n_81),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_1),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_1),
.A2(n_81),
.B1(n_182),
.B2(n_185),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_1),
.A2(n_81),
.B1(n_539),
.B2(n_542),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_2),
.Y(n_459)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_3),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_3),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_199),
.B1(n_203),
.B2(n_204),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_4),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_4),
.A2(n_204),
.B1(n_546),
.B2(n_551),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_5),
.Y(n_85)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_5),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g197 ( 
.A(n_5),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_5),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_6),
.A2(n_124),
.B1(n_127),
.B2(n_128),
.Y(n_123)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_6),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_6),
.A2(n_127),
.B1(n_242),
.B2(n_245),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_6),
.A2(n_127),
.B1(n_349),
.B2(n_352),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_6),
.A2(n_127),
.B1(n_315),
.B2(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_7),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_7),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_7),
.A2(n_117),
.B1(n_139),
.B2(n_210),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_7),
.A2(n_139),
.B1(n_325),
.B2(n_328),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_7),
.A2(n_139),
.B1(n_373),
.B2(n_378),
.Y(n_372)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_8),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_8),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g424 ( 
.A(n_8),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_9),
.B(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_9),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_9),
.A2(n_262),
.B(n_337),
.Y(n_336)
);

OAI32xp33_ASAP7_75t_L g356 ( 
.A1(n_9),
.A2(n_357),
.A3(n_360),
.B1(n_364),
.B2(n_369),
.Y(n_356)
);

OAI32xp33_ASAP7_75t_L g393 ( 
.A1(n_9),
.A2(n_357),
.A3(n_360),
.B1(n_364),
.B2(n_369),
.Y(n_393)
);

OAI32xp33_ASAP7_75t_L g395 ( 
.A1(n_9),
.A2(n_357),
.A3(n_360),
.B1(n_364),
.B2(n_369),
.Y(n_395)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_9),
.A2(n_320),
.B1(n_406),
.B2(n_409),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_9),
.B(n_249),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_9),
.A2(n_82),
.B1(n_384),
.B2(n_494),
.Y(n_493)
);

AOI22xp33_ASAP7_75t_SL g282 ( 
.A1(n_10),
.A2(n_283),
.B1(n_285),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_10),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_10),
.A2(n_287),
.B1(n_298),
.B2(n_303),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_10),
.A2(n_287),
.B1(n_421),
.B2(n_425),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_10),
.A2(n_287),
.B1(n_488),
.B2(n_495),
.Y(n_494)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_11),
.Y(n_103)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_11),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_11),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_11),
.Y(n_256)
);

OAI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_52),
.B1(n_57),
.B2(n_58),
.Y(n_51)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_12),
.A2(n_57),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_12),
.A2(n_57),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g559 ( 
.A1(n_12),
.A2(n_57),
.B1(n_263),
.B2(n_340),
.Y(n_559)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_13),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_14),
.A2(n_88),
.B1(n_90),
.B2(n_92),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_14),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_14),
.A2(n_92),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

BUFx4f_ASAP7_75t_L g377 ( 
.A(n_15),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_16),
.A2(n_117),
.B1(n_121),
.B2(n_122),
.Y(n_116)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_16),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_16),
.A2(n_121),
.B1(n_243),
.B2(n_307),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_16),
.A2(n_121),
.B1(n_398),
.B2(n_401),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g475 ( 
.A1(n_16),
.A2(n_121),
.B1(n_476),
.B2(n_480),
.Y(n_475)
);

BUFx8_ASAP7_75t_L g105 ( 
.A(n_17),
.Y(n_105)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_17),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_17),
.Y(n_126)
);

BUFx5_ASAP7_75t_L g129 ( 
.A(n_17),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_17),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_527),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_288),
.B(n_525),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_234),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_22),
.B(n_234),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_177),
.Y(n_22)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_23),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_98),
.C(n_131),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_25),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_69),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_26),
.A2(n_27),
.B1(n_69),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_51),
.B1(n_63),
.B2(n_65),
.Y(n_27)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_28),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_28),
.B(n_65),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_28),
.A2(n_63),
.B1(n_348),
.B2(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_28),
.A2(n_63),
.B1(n_397),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_28),
.A2(n_63),
.B1(n_420),
.B2(n_465),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_SL g543 ( 
.A1(n_28),
.A2(n_63),
.B1(n_544),
.B2(n_545),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

OAI22xp33_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_32),
.Y(n_164)
);

INVx6_ASAP7_75t_L g363 ( 
.A(n_32),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g426 ( 
.A(n_37),
.Y(n_426)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_38),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_38),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_38),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_43),
.B1(n_47),
.B2(n_49),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_41),
.Y(n_453)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_44),
.Y(n_275)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_45),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_46),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_48),
.Y(n_202)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_51),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_52),
.B(n_320),
.Y(n_454)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_56),
.Y(n_188)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_56),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_56),
.Y(n_468)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g552 ( 
.A(n_62),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_63),
.B(n_224),
.Y(n_223)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_64),
.A2(n_180),
.B1(n_181),
.B2(n_189),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_64),
.A2(n_180),
.B1(n_324),
.B2(n_332),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_64),
.A2(n_180),
.B1(n_324),
.B2(n_347),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_64),
.B(n_320),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_69),
.Y(n_517)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_82),
.B1(n_87),
.B2(n_93),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_70),
.A2(n_82),
.B1(n_270),
.B2(n_276),
.Y(n_269)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_76),
.Y(n_273)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_76),
.Y(n_431)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_77),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_82),
.A2(n_195),
.B(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_82),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g427 ( 
.A1(n_82),
.A2(n_428),
.B1(n_432),
.B2(n_436),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g497 ( 
.A1(n_82),
.A2(n_475),
.B1(n_494),
.B2(n_498),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_86),
.Y(n_82)
);

INVx5_ASAP7_75t_L g384 ( 
.A(n_83),
.Y(n_384)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_84),
.Y(n_230)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_85),
.Y(n_318)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_86),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_87),
.Y(n_227)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_89),
.Y(n_451)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_96),
.Y(n_435)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_96),
.Y(n_500)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_98),
.B(n_132),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_116),
.B1(n_123),
.B2(n_130),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_99),
.A2(n_123),
.B1(n_130),
.B2(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_99),
.A2(n_116),
.B1(n_130),
.B2(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_99),
.A2(n_130),
.B1(n_282),
.B2(n_336),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_99),
.A2(n_130),
.B1(n_209),
.B2(n_559),
.Y(n_558)
);

AO21x2_ASAP7_75t_L g99 ( 
.A1(n_100),
.A2(n_106),
.B(n_110),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_104),
.Y(n_100)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_106),
.A2(n_252),
.B1(n_261),
.B2(n_265),
.Y(n_251)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

AO22x2_ASAP7_75t_L g110 ( 
.A1(n_108),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_112),
.Y(n_176)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_112),
.Y(n_311)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_112),
.Y(n_359)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_113),
.Y(n_220)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_117),
.Y(n_122)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx5_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_126),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_126),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_129),
.Y(n_211)
);

NOR2x1_ASAP7_75t_R g319 ( 
.A(n_130),
.B(n_320),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_142),
.B1(n_168),
.B2(n_169),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_134),
.A2(n_143),
.B1(n_241),
.B2(n_249),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_137),
.Y(n_302)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_137),
.Y(n_414)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_138),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g248 ( 
.A(n_138),
.Y(n_248)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OAI22x1_ASAP7_75t_L g212 ( 
.A1(n_142),
.A2(n_168),
.B1(n_169),
.B2(n_213),
.Y(n_212)
);

OAI22xp33_ASAP7_75t_L g296 ( 
.A1(n_142),
.A2(n_168),
.B1(n_297),
.B2(n_306),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_142),
.A2(n_168),
.B1(n_306),
.B2(n_334),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_142),
.A2(n_168),
.B1(n_297),
.B2(n_405),
.Y(n_404)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_143),
.A2(n_249),
.B1(n_536),
.B2(n_537),
.Y(n_535)
);

OA21x2_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_152),
.B(n_158),
.Y(n_143)
);

INVxp33_ASAP7_75t_L g369 ( 
.A(n_144),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_149),
.Y(n_144)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_148),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_149),
.Y(n_542)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_151),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_151),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_156),
.Y(n_152)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g541 ( 
.A(n_156),
.Y(n_541)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g168 ( 
.A(n_158),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_162),
.B1(n_163),
.B2(n_165),
.Y(n_158)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_206),
.B1(n_232),
.B2(n_233),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_178),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_178),
.B(n_233),
.C(n_530),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_179),
.A2(n_193),
.B1(n_194),
.B2(n_205),
.Y(n_178)
);

INVxp33_ASAP7_75t_SL g205 ( 
.A(n_179),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_179),
.B(n_194),
.Y(n_560)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_181),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_183),
.Y(n_402)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_184),
.Y(n_353)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_188),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g544 ( 
.A(n_189),
.Y(n_544)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_193),
.A2(n_194),
.B1(n_557),
.B2(n_558),
.Y(n_556)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx12f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_198),
.Y(n_231)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_200),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_202),
.Y(n_381)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_206),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_221),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_208),
.B(n_212),
.C(n_221),
.Y(n_532)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx6_ASAP7_75t_L g340 ( 
.A(n_211),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g536 ( 
.A(n_213),
.Y(n_536)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_217),
.Y(n_305)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

HB1xp67_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_223),
.B(n_225),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_222),
.B(n_223),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_225),
.B(n_238),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_227),
.B1(n_228),
.B2(n_231),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_226),
.A2(n_271),
.B1(n_314),
.B2(n_318),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_226),
.A2(n_314),
.B1(n_372),
.B2(n_382),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_226),
.A2(n_382),
.B1(n_474),
.B2(n_482),
.Y(n_473)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx6_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_235),
.B(n_237),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g509 ( 
.A(n_239),
.B(n_510),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_250),
.C(n_280),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_240),
.A2(n_280),
.B1(n_281),
.B2(n_514),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_240),
.Y(n_514)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_248),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g512 ( 
.A(n_250),
.B(n_513),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_269),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_251),
.B(n_269),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g270 ( 
.A(n_271),
.Y(n_270)
);

INVx4_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_275),
.Y(n_317)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_508),
.B(n_523),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_385),
.B(n_507),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_341),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_292),
.B(n_341),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_321),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_294),
.B(n_295),
.C(n_321),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_312),
.C(n_319),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_296),
.B(n_344),
.Y(n_343)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_311),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_312),
.A2(n_313),
.B1(n_319),
.B2(n_345),
.Y(n_344)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_319),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_320),
.B(n_365),
.Y(n_364)
);

OAI21xp33_ASAP7_75t_SL g465 ( 
.A1(n_320),
.A2(n_454),
.B(n_466),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_320),
.B(n_490),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_335),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_333),
.Y(n_322)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_323),
.B(n_333),
.C(n_335),
.Y(n_518)
);

BUFx2_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_346),
.C(n_354),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_342),
.A2(n_343),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_346),
.A2(n_354),
.B1(n_355),
.B2(n_390),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_346),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_370),
.Y(n_355)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_363),
.Y(n_400)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_363),
.Y(n_448)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_363),
.Y(n_550)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_370),
.A2(n_371),
.B1(n_393),
.B2(n_394),
.Y(n_392)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_377),
.Y(n_481)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_381),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx3_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

OAI21x1_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_415),
.B(n_506),
.Y(n_385)
);

NOR2xp67_ASAP7_75t_SL g386 ( 
.A(n_387),
.B(n_391),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_391),
.Y(n_506)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_396),
.C(n_403),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_392),
.B(n_440),
.Y(n_439)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g440 ( 
.A1(n_396),
.A2(n_403),
.B1(n_404),
.B2(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_396),
.Y(n_441)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

BUFx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI21x1_ASAP7_75t_SL g415 ( 
.A1(n_416),
.A2(n_442),
.B(n_505),
.Y(n_415)
);

NAND2xp33_ASAP7_75t_SL g416 ( 
.A(n_417),
.B(n_439),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_417),
.B(n_439),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_427),
.C(n_437),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g470 ( 
.A1(n_418),
.A2(n_419),
.B1(n_437),
.B2(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_427),
.B(n_470),
.Y(n_469)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_428),
.Y(n_482)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx4_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx4_ASAP7_75t_SL g434 ( 
.A(n_435),
.Y(n_434)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g442 ( 
.A1(n_443),
.A2(n_471),
.B(n_504),
.Y(n_442)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_469),
.Y(n_443)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_444),
.B(n_469),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_463),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_445),
.A2(n_463),
.B1(n_464),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_445),
.Y(n_484)
);

OAI32xp33_ASAP7_75t_L g445 ( 
.A1(n_446),
.A2(n_449),
.A3(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_447),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_460),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

INVx3_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx8_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

INVx3_ASAP7_75t_L g461 ( 
.A(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_472),
.A2(n_485),
.B(n_503),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_483),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_473),
.B(n_483),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_476),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_478),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

OAI21xp5_ASAP7_75t_L g485 ( 
.A1(n_486),
.A2(n_496),
.B(n_502),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_493),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_489),
.Y(n_487)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_501),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_497),
.B(n_501),
.Y(n_502)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_499),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_511),
.B(n_519),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_509),
.B(n_511),
.C(n_524),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_515),
.C(n_518),
.Y(n_511)
);

XNOR2xp5_ASAP7_75t_SL g520 ( 
.A(n_512),
.B(n_521),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_516),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_518),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_520),
.B(n_522),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_520),
.B(n_522),
.Y(n_524)
);

INVxp67_ASAP7_75t_SL g525 ( 
.A(n_526),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_528),
.B(n_562),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_531),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_529),
.B(n_531),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_532),
.B(n_533),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_534),
.B(n_554),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g534 ( 
.A1(n_535),
.A2(n_543),
.B(n_553),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_535),
.B(n_543),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_547),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_550),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_552),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_555),
.A2(n_556),
.B1(n_560),
.B2(n_561),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_556),
.Y(n_555)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_560),
.Y(n_561)
);

INVxp33_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);


endmodule