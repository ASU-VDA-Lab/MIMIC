module fake_ariane_2304_n_87 (n_8, n_7, n_1, n_6, n_13, n_17, n_4, n_2, n_18, n_9, n_11, n_3, n_14, n_0, n_19, n_16, n_5, n_12, n_15, n_10, n_87);

input n_8;
input n_7;
input n_1;
input n_6;
input n_13;
input n_17;
input n_4;
input n_2;
input n_18;
input n_9;
input n_11;
input n_3;
input n_14;
input n_0;
input n_19;
input n_16;
input n_5;
input n_12;
input n_15;
input n_10;

output n_87;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_38;
wire n_47;
wire n_86;
wire n_75;
wire n_67;
wire n_34;
wire n_69;
wire n_74;
wire n_33;
wire n_40;
wire n_53;
wire n_21;
wire n_66;
wire n_71;
wire n_24;
wire n_49;
wire n_20;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_26;
wire n_46;
wire n_84;
wire n_36;
wire n_72;
wire n_44;
wire n_30;
wire n_82;
wire n_42;
wire n_31;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_32;
wire n_37;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_23;
wire n_61;
wire n_22;
wire n_43;
wire n_81;
wire n_27;
wire n_29;
wire n_41;
wire n_55;
wire n_28;
wire n_80;
wire n_68;
wire n_78;
wire n_39;
wire n_59;
wire n_63;
wire n_35;
wire n_54;
wire n_25;

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_10),
.A2(n_1),
.B(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_7),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_12),
.B(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_8),
.B(n_19),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22x1_ASAP7_75t_L g30 ( 
.A1(n_3),
.A2(n_2),
.B1(n_9),
.B2(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

OAI21x1_ASAP7_75t_L g32 ( 
.A1(n_4),
.A2(n_6),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_5),
.B(n_8),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g34 ( 
.A(n_11),
.B(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_21),
.B(n_16),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_30),
.A2(n_33),
.B1(n_26),
.B2(n_34),
.Y(n_38)
);

INVxp67_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_27),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_39),
.B(n_24),
.Y(n_41)
);

NOR2xp67_ASAP7_75t_L g42 ( 
.A(n_38),
.B(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_37),
.A2(n_33),
.B1(n_30),
.B2(n_34),
.Y(n_43)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_40),
.Y(n_44)
);

AOI221x1_ASAP7_75t_L g45 ( 
.A1(n_36),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.C(n_25),
.Y(n_45)
);

OAI21x1_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_32),
.B(n_28),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_29),
.Y(n_47)
);

AO21x2_ASAP7_75t_L g48 ( 
.A1(n_42),
.A2(n_32),
.B(n_25),
.Y(n_48)
);

AO21x2_ASAP7_75t_L g49 ( 
.A1(n_46),
.A2(n_32),
.B(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_29),
.Y(n_51)
);

AO21x1_ASAP7_75t_SL g52 ( 
.A1(n_43),
.A2(n_45),
.B(n_33),
.Y(n_52)
);

AO21x2_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_35),
.B(n_22),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_45),
.Y(n_54)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g56 ( 
.A(n_47),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_57),
.B(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_56),
.A2(n_51),
.B(n_48),
.Y(n_62)
);

HB1xp67_ASAP7_75t_L g63 ( 
.A(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_48),
.Y(n_66)
);

AOI221xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_52),
.B1(n_23),
.B2(n_31),
.C(n_48),
.Y(n_67)
);

OAI221xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_22),
.B1(n_31),
.B2(n_23),
.C(n_28),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_53),
.Y(n_69)
);

AOI211x1_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_61),
.B(n_65),
.C(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_53),
.Y(n_71)
);

XOR2x2_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_49),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_61),
.A2(n_31),
.B1(n_23),
.B2(n_22),
.Y(n_73)
);

NOR4xp25_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_35),
.C(n_66),
.D(n_22),
.Y(n_74)
);

A2O1A1Ixp33_ASAP7_75t_L g75 ( 
.A1(n_67),
.A2(n_23),
.B(n_31),
.C(n_20),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_53),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_71),
.A2(n_28),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_73),
.B(n_20),
.Y(n_78)
);

OAI21xp33_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_31),
.B(n_70),
.Y(n_79)
);

NAND4xp25_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_31),
.C(n_28),
.D(n_49),
.Y(n_80)
);

NOR3xp33_ASAP7_75t_SL g81 ( 
.A(n_75),
.B(n_49),
.C(n_20),
.Y(n_81)
);

NOR2xp67_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_20),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_81),
.A2(n_74),
.B1(n_77),
.B2(n_20),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_84),
.A2(n_80),
.B1(n_78),
.B2(n_20),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_75),
.B(n_49),
.Y(n_86)
);

OR2x6_ASAP7_75t_L g87 ( 
.A(n_86),
.B(n_85),
.Y(n_87)
);


endmodule