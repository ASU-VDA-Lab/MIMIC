module fake_netlist_5_2139_n_1668 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1668);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1668;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_226;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1580;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_171;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1598;
wire n_955;
wire n_163;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1623;
wire n_1565;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_284;
wire n_1128;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_254;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_314;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_259;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_168;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_261;
wire n_174;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_233;
wire n_572;
wire n_366;
wire n_815;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_280;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_774;
wire n_1628;
wire n_1514;
wire n_1335;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1440;
wire n_177;
wire n_421;
wire n_1356;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_198;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_209;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_481;
wire n_1554;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_167;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_276;
wire n_1225;
wire n_1520;
wire n_169;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_170;
wire n_161;
wire n_273;
wire n_585;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_166;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_4),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_45),
.Y(n_162)
);

BUFx8_ASAP7_75t_SL g163 ( 
.A(n_113),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_94),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_79),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_97),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_125),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_96),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_82),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_31),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_41),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_18),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_65),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_118),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_45),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_17),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_48),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_57),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_26),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_99),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_108),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_141),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_109),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_101),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_160),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g190 ( 
.A(n_138),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_127),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_19),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_92),
.Y(n_196)
);

BUFx8_ASAP7_75t_SL g197 ( 
.A(n_41),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_75),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_153),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_18),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_63),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_151),
.Y(n_203)
);

HB1xp67_ASAP7_75t_L g204 ( 
.A(n_107),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_147),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_126),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_156),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_100),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_43),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_103),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g211 ( 
.A(n_78),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_93),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

INVx2_ASAP7_75t_SL g214 ( 
.A(n_150),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_69),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_43),
.Y(n_216)
);

BUFx5_ASAP7_75t_L g217 ( 
.A(n_30),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_115),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_74),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_88),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_119),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_70),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_132),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_38),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_31),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_51),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_28),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g228 ( 
.A(n_30),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_8),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_51),
.Y(n_230)
);

INVx2_ASAP7_75t_SL g231 ( 
.A(n_28),
.Y(n_231)
);

BUFx10_ASAP7_75t_L g232 ( 
.A(n_116),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_110),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_10),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_71),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_59),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_72),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_112),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_17),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_22),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_77),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_124),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_111),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_25),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_15),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_34),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_20),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_11),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_140),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_105),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_9),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_46),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_142),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_146),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_58),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_145),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_35),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_81),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_29),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_5),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_46),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_13),
.Y(n_264)
);

BUFx10_ASAP7_75t_L g265 ( 
.A(n_39),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_5),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_48),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_135),
.Y(n_268)
);

BUFx10_ASAP7_75t_L g269 ( 
.A(n_76),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_102),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_73),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_89),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_90),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_39),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_67),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_47),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_114),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_47),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_117),
.Y(n_279)
);

BUFx2_ASAP7_75t_L g280 ( 
.A(n_84),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_144),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_0),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_50),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_61),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_19),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_134),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_4),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_0),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_120),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_87),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_25),
.Y(n_291)
);

BUFx5_ASAP7_75t_L g292 ( 
.A(n_54),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_6),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_9),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_123),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_52),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_33),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_26),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_128),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_33),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_50),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_23),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_23),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_34),
.Y(n_304)
);

INVx2_ASAP7_75t_SL g305 ( 
.A(n_6),
.Y(n_305)
);

BUFx10_ASAP7_75t_L g306 ( 
.A(n_55),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_24),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_95),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_149),
.Y(n_309)
);

BUFx5_ASAP7_75t_L g310 ( 
.A(n_104),
.Y(n_310)
);

BUFx5_ASAP7_75t_L g311 ( 
.A(n_159),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_14),
.Y(n_312)
);

INVx1_ASAP7_75t_SL g313 ( 
.A(n_12),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_11),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_49),
.Y(n_315)
);

BUFx8_ASAP7_75t_SL g316 ( 
.A(n_121),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_68),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_66),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_60),
.Y(n_319)
);

INVxp67_ASAP7_75t_SL g320 ( 
.A(n_164),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_217),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_217),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_197),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_217),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_176),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_216),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_176),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_195),
.B(n_280),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_217),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_217),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_197),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_165),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_204),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_166),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_212),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_167),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_217),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_168),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_212),
.Y(n_339)
);

NOR2xp67_ASAP7_75t_L g340 ( 
.A(n_230),
.B(n_1),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_217),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_232),
.Y(n_342)
);

NOR2xp67_ASAP7_75t_L g343 ( 
.A(n_231),
.B(n_1),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_169),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_170),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_261),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_234),
.B(n_2),
.Y(n_347)
);

BUFx2_ASAP7_75t_SL g348 ( 
.A(n_218),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_218),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_303),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_171),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_184),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_187),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_261),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_188),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_161),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_189),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_261),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_275),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_191),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_196),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_199),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_200),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_246),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_234),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_246),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_291),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_177),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_265),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_202),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_291),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_300),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_300),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_239),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_239),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_162),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_211),
.B(n_2),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_207),
.Y(n_379)
);

BUFx3_ASAP7_75t_L g380 ( 
.A(n_232),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_215),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_179),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_289),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_219),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_181),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_201),
.Y(n_386)
);

INVx1_ASAP7_75t_SL g387 ( 
.A(n_265),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_232),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_289),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_308),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_308),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_220),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_163),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_163),
.Y(n_394)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_347),
.B(n_366),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_321),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_325),
.A2(n_161),
.B1(n_174),
.B2(n_175),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_321),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_322),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_322),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_324),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_329),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_329),
.Y(n_404)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_330),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_330),
.Y(n_407)
);

INVx6_ASAP7_75t_L g408 ( 
.A(n_347),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_337),
.Y(n_409)
);

INVx3_ASAP7_75t_L g410 ( 
.A(n_337),
.Y(n_410)
);

AND2x2_ASAP7_75t_SL g411 ( 
.A(n_378),
.B(n_252),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_341),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_341),
.Y(n_413)
);

INVx3_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_346),
.B(n_211),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_348),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_352),
.B(n_214),
.Y(n_417)
);

OA21x2_ASAP7_75t_L g418 ( 
.A1(n_352),
.A2(n_226),
.B(n_209),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_355),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g420 ( 
.A(n_355),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_359),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_387),
.B(n_316),
.Y(n_422)
);

NAND2xp33_ASAP7_75t_L g423 ( 
.A(n_359),
.B(n_231),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_327),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_343),
.B(n_214),
.Y(n_427)
);

INVx3_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_375),
.B(n_173),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_367),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_368),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_335),
.A2(n_183),
.B1(n_314),
.B2(n_174),
.Y(n_432)
);

BUFx10_ASAP7_75t_L g433 ( 
.A(n_328),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_368),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_372),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_372),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_375),
.B(n_173),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_348),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_373),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_376),
.B(n_252),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_357),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_343),
.B(n_251),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_374),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_377),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_320),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_185),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_382),
.B(n_186),
.Y(n_450)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_382),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_385),
.Y(n_452)
);

OA21x2_ASAP7_75t_L g453 ( 
.A1(n_385),
.A2(n_262),
.B(n_248),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_386),
.B(n_251),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_386),
.B(n_305),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_342),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_342),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_340),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_333),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_326),
.B(n_305),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_380),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_332),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_350),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_334),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_336),
.B(n_193),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_338),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_465),
.B(n_344),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_456),
.B(n_345),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_351),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_433),
.B(n_369),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_395),
.B(n_388),
.Y(n_472)
);

AND3x2_ASAP7_75t_L g473 ( 
.A(n_422),
.B(n_278),
.C(n_198),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_396),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g477 ( 
.A1(n_411),
.A2(n_228),
.B1(n_245),
.B2(n_254),
.Y(n_477)
);

INVx3_ASAP7_75t_L g478 ( 
.A(n_407),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_416),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_398),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_396),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_398),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_433),
.B(n_369),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_456),
.B(n_395),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_401),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_398),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_401),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_401),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g489 ( 
.A(n_433),
.B(n_388),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_403),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_353),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_427),
.B(n_251),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_456),
.B(n_354),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_395),
.B(n_356),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g495 ( 
.A(n_395),
.B(n_358),
.Y(n_495)
);

AND2x6_ASAP7_75t_L g496 ( 
.A(n_427),
.B(n_251),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_399),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_403),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_456),
.B(n_361),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

BUFx2_ASAP7_75t_L g501 ( 
.A(n_405),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_427),
.B(n_362),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_433),
.B(n_363),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_407),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_433),
.B(n_364),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_438),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_399),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_416),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_465),
.B(n_371),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_399),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_400),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_407),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_411),
.A2(n_267),
.B1(n_294),
.B2(n_263),
.Y(n_513)
);

INVx3_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_404),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_404),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_397),
.B(n_323),
.Y(n_517)
);

NAND2xp33_ASAP7_75t_L g518 ( 
.A(n_459),
.B(n_379),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_400),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g520 ( 
.A(n_457),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_407),
.Y(n_521)
);

OR2x6_ASAP7_75t_L g522 ( 
.A(n_463),
.B(n_190),
.Y(n_522)
);

NAND2xp33_ASAP7_75t_SL g523 ( 
.A(n_405),
.B(n_331),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_404),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_433),
.B(n_381),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_400),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_447),
.B(n_384),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_406),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_427),
.B(n_392),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_427),
.B(n_221),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_413),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_448),
.B(n_315),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_406),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_427),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_407),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_406),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_411),
.B(n_223),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_411),
.B(n_233),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_408),
.B(n_235),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_447),
.B(n_339),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_409),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_438),
.B(n_269),
.Y(n_543)
);

INVx1_ASAP7_75t_SL g544 ( 
.A(n_405),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_407),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_457),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_408),
.B(n_236),
.Y(n_547)
);

OR2x2_ASAP7_75t_L g548 ( 
.A(n_442),
.B(n_288),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_408),
.A2(n_272),
.B1(n_271),
.B2(n_317),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_448),
.B(n_194),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_408),
.B(n_444),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_460),
.B(n_269),
.Y(n_552)
);

BUFx6f_ASAP7_75t_L g553 ( 
.A(n_407),
.Y(n_553)
);

OR2x2_ASAP7_75t_L g554 ( 
.A(n_442),
.B(n_293),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_407),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_408),
.A2(n_272),
.B1(n_271),
.B2(n_317),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_412),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_463),
.B(n_349),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_412),
.Y(n_559)
);

NAND2xp33_ASAP7_75t_SL g560 ( 
.A(n_464),
.B(n_393),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_412),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_463),
.B(n_460),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_448),
.B(n_269),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_413),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_408),
.B(n_238),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_408),
.B(n_242),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_463),
.B(n_360),
.Y(n_567)
);

INVx2_ASAP7_75t_SL g568 ( 
.A(n_466),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_444),
.B(n_244),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_444),
.B(n_255),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_460),
.B(n_306),
.Y(n_571)
);

AOI22xp33_ASAP7_75t_L g572 ( 
.A1(n_461),
.A2(n_453),
.B1(n_448),
.B2(n_450),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_409),
.Y(n_573)
);

INVx2_ASAP7_75t_SL g574 ( 
.A(n_466),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_409),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_466),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

AND2x2_ASAP7_75t_SL g578 ( 
.A(n_418),
.B(n_271),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_402),
.Y(n_579)
);

AND2x2_ASAP7_75t_L g580 ( 
.A(n_440),
.B(n_306),
.Y(n_580)
);

AND2x4_ASAP7_75t_L g581 ( 
.A(n_450),
.B(n_203),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_413),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_413),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_402),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_463),
.B(n_383),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_402),
.Y(n_586)
);

HB1xp67_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_459),
.B(n_389),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_421),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_412),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_440),
.B(n_306),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_421),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_440),
.B(n_313),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_412),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_412),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g596 ( 
.A1(n_397),
.A2(n_175),
.B1(n_314),
.B2(n_312),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_457),
.B(n_178),
.Y(n_597)
);

BUFx8_ASAP7_75t_SL g598 ( 
.A(n_425),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_402),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_402),
.Y(n_600)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_425),
.Y(n_601)
);

INVx2_ASAP7_75t_SL g602 ( 
.A(n_466),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_412),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_SL g604 ( 
.A(n_457),
.B(n_178),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_459),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_412),
.Y(n_606)
);

INVx4_ASAP7_75t_L g607 ( 
.A(n_412),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_402),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_421),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_462),
.B(n_390),
.Y(n_610)
);

INVx2_ASAP7_75t_SL g611 ( 
.A(n_462),
.Y(n_611)
);

BUFx3_ASAP7_75t_L g612 ( 
.A(n_457),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_410),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_568),
.B(n_457),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_513),
.A2(n_458),
.B1(n_444),
.B2(n_462),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_587),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_506),
.B(n_464),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_475),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_476),
.Y(n_619)
);

INVx2_ASAP7_75t_SL g620 ( 
.A(n_506),
.Y(n_620)
);

AND2x4_ASAP7_75t_L g621 ( 
.A(n_532),
.B(n_581),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_572),
.A2(n_458),
.B1(n_444),
.B2(n_462),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_562),
.B(n_444),
.Y(n_623)
);

NAND2xp33_ASAP7_75t_L g624 ( 
.A(n_538),
.B(n_457),
.Y(n_624)
);

INVx8_ASAP7_75t_L g625 ( 
.A(n_522),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_534),
.B(n_457),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_534),
.B(n_457),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g628 ( 
.A(n_479),
.B(n_458),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_537),
.B(n_429),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_568),
.B(n_429),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_574),
.B(n_437),
.Y(n_631)
);

INVx3_ASAP7_75t_L g632 ( 
.A(n_613),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_484),
.B(n_410),
.Y(n_633)
);

INVx3_ASAP7_75t_L g634 ( 
.A(n_613),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_472),
.B(n_577),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_472),
.B(n_394),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_476),
.Y(n_637)
);

A2O1A1Ixp33_ASAP7_75t_L g638 ( 
.A1(n_477),
.A2(n_410),
.B(n_449),
.C(n_450),
.Y(n_638)
);

OR2x2_ASAP7_75t_L g639 ( 
.A(n_544),
.B(n_397),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_481),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_598),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_576),
.B(n_410),
.Y(n_642)
);

NAND2x1p5_ASAP7_75t_L g643 ( 
.A(n_576),
.B(n_418),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_485),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_485),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_605),
.B(n_410),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_602),
.B(n_271),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_487),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_602),
.B(n_449),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_539),
.B(n_272),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_611),
.B(n_453),
.Y(n_651)
);

AOI22xp33_ASAP7_75t_L g652 ( 
.A1(n_578),
.A2(n_453),
.B1(n_418),
.B2(n_450),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_611),
.B(n_453),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_577),
.B(n_449),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_494),
.B(n_272),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_593),
.Y(n_656)
);

OAI22x1_ASAP7_75t_L g657 ( 
.A1(n_596),
.A2(n_477),
.B1(n_544),
.B2(n_501),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_527),
.B(n_453),
.Y(n_658)
);

AOI22xp5_ASAP7_75t_L g659 ( 
.A1(n_494),
.A2(n_391),
.B1(n_440),
.B2(n_281),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_495),
.B(n_467),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_613),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_495),
.B(n_455),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_578),
.A2(n_453),
.B1(n_418),
.B2(n_432),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_578),
.B(n_551),
.Y(n_664)
);

BUFx6f_ASAP7_75t_SL g665 ( 
.A(n_581),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_488),
.B(n_453),
.Y(n_666)
);

BUFx6f_ASAP7_75t_L g667 ( 
.A(n_520),
.Y(n_667)
);

AOI22xp5_ASAP7_75t_L g668 ( 
.A1(n_588),
.A2(n_277),
.B1(n_256),
.B2(n_284),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_490),
.B(n_418),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_468),
.B(n_422),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_532),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_509),
.B(n_449),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g673 ( 
.A1(n_610),
.A2(n_295),
.B1(n_258),
.B2(n_268),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_502),
.B(n_432),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_490),
.B(n_418),
.Y(n_675)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_548),
.B(n_432),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_498),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_529),
.B(n_317),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_501),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_L g680 ( 
.A(n_469),
.B(n_292),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_563),
.B(n_182),
.Y(n_681)
);

AND2x4_ASAP7_75t_SL g682 ( 
.A(n_522),
.B(n_265),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_498),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_515),
.B(n_420),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_L g685 ( 
.A1(n_548),
.A2(n_243),
.B1(n_237),
.B2(n_222),
.Y(n_685)
);

BUFx3_ASAP7_75t_L g686 ( 
.A(n_581),
.Y(n_686)
);

OR2x6_ASAP7_75t_L g687 ( 
.A(n_471),
.B(n_455),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_516),
.B(n_317),
.Y(n_688)
);

NOR2xp67_ASAP7_75t_SL g689 ( 
.A(n_520),
.B(n_205),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_516),
.B(n_420),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_524),
.B(n_420),
.Y(n_691)
);

AOI22xp33_ASAP7_75t_L g692 ( 
.A1(n_581),
.A2(n_446),
.B1(n_279),
.B2(n_206),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_524),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_540),
.A2(n_415),
.B(n_417),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_543),
.B(n_445),
.Y(n_695)
);

INVx1_ASAP7_75t_SL g696 ( 
.A(n_601),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_528),
.B(n_420),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_528),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_533),
.B(n_445),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_SL g700 ( 
.A1(n_596),
.A2(n_183),
.B1(n_180),
.B2(n_312),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_554),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_533),
.B(n_445),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_536),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_536),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_542),
.B(n_451),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_542),
.B(n_445),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_L g707 ( 
.A(n_470),
.B(n_292),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_573),
.B(n_445),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_550),
.A2(n_446),
.B1(n_318),
.B2(n_208),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_550),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_554),
.Y(n_711)
);

OAI22xp5_ASAP7_75t_L g712 ( 
.A1(n_522),
.A2(n_319),
.B1(n_210),
.B2(n_257),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_550),
.A2(n_290),
.B1(n_299),
.B2(n_260),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_552),
.B(n_445),
.Y(n_714)
);

OR2x2_ASAP7_75t_L g715 ( 
.A(n_541),
.B(n_180),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_575),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_580),
.B(n_430),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_522),
.A2(n_270),
.B1(n_286),
.B2(n_182),
.Y(n_718)
);

BUFx8_ASAP7_75t_L g719 ( 
.A(n_580),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_575),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_474),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_591),
.B(n_430),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_491),
.B(n_451),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_493),
.B(n_451),
.Y(n_724)
);

OAI22xp5_ASAP7_75t_SL g725 ( 
.A1(n_601),
.A2(n_229),
.B1(n_172),
.B2(n_192),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_579),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_571),
.B(n_213),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_503),
.B(n_224),
.Y(n_728)
);

CKINVDCx11_ASAP7_75t_R g729 ( 
.A(n_517),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_480),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_591),
.B(n_430),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_579),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_499),
.B(n_451),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_505),
.B(n_225),
.Y(n_734)
);

INVx1_ASAP7_75t_SL g735 ( 
.A(n_560),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_480),
.Y(n_736)
);

BUFx3_ASAP7_75t_L g737 ( 
.A(n_550),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_584),
.B(n_451),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_482),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_522),
.A2(n_273),
.B1(n_309),
.B2(n_415),
.Y(n_740)
);

NOR2xp67_ASAP7_75t_L g741 ( 
.A(n_479),
.B(n_417),
.Y(n_741)
);

AND2x2_ASAP7_75t_SL g742 ( 
.A(n_549),
.B(n_423),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_508),
.B(n_525),
.Y(n_743)
);

INVx2_ASAP7_75t_SL g744 ( 
.A(n_530),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_482),
.Y(n_745)
);

INVx2_ASAP7_75t_SL g746 ( 
.A(n_508),
.Y(n_746)
);

AO22x2_ASAP7_75t_L g747 ( 
.A1(n_489),
.A2(n_454),
.B1(n_441),
.B2(n_439),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_486),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_584),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_586),
.B(n_599),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_586),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_599),
.B(n_451),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_600),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_600),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_608),
.B(n_451),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_608),
.B(n_451),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_486),
.Y(n_757)
);

NOR3xp33_ASAP7_75t_L g758 ( 
.A(n_483),
.B(n_423),
.C(n_285),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_569),
.B(n_451),
.Y(n_759)
);

OR2x2_ASAP7_75t_L g760 ( 
.A(n_558),
.B(n_227),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_497),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_567),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_570),
.B(n_452),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_473),
.Y(n_764)
);

NOR2xp33_ASAP7_75t_L g765 ( 
.A(n_518),
.B(n_547),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_556),
.B(n_452),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_497),
.Y(n_767)
);

AOI22xp5_ASAP7_75t_L g768 ( 
.A1(n_597),
.A2(n_454),
.B1(n_310),
.B2(n_292),
.Y(n_768)
);

NOR2xp67_ASAP7_75t_L g769 ( 
.A(n_585),
.B(n_435),
.Y(n_769)
);

OAI22xp5_ASAP7_75t_L g770 ( 
.A1(n_672),
.A2(n_565),
.B1(n_566),
.B2(n_546),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_624),
.A2(n_612),
.B(n_520),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_660),
.B(n_620),
.Y(n_772)
);

AOI22xp5_ASAP7_75t_L g773 ( 
.A1(n_660),
.A2(n_674),
.B1(n_672),
.B2(n_630),
.Y(n_773)
);

NOR2x1_ASAP7_75t_L g774 ( 
.A(n_628),
.B(n_741),
.Y(n_774)
);

HB1xp67_ASAP7_75t_L g775 ( 
.A(n_679),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_641),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_630),
.B(n_504),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_623),
.A2(n_612),
.B(n_546),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_629),
.B(n_762),
.Y(n_779)
);

CKINVDCx5p33_ASAP7_75t_R g780 ( 
.A(n_729),
.Y(n_780)
);

AOI22xp5_ASAP7_75t_L g781 ( 
.A1(n_674),
.A2(n_604),
.B1(n_523),
.B2(n_492),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_631),
.B(n_504),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_631),
.A2(n_496),
.B1(n_492),
.B2(n_559),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_686),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_626),
.A2(n_612),
.B(n_546),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_626),
.A2(n_555),
.B(n_607),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_663),
.A2(n_492),
.B1(n_496),
.B2(n_311),
.Y(n_787)
);

INVx3_ASAP7_75t_L g788 ( 
.A(n_661),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_661),
.B(n_553),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_L g790 ( 
.A1(n_663),
.A2(n_535),
.B1(n_559),
.B2(n_545),
.Y(n_790)
);

A2O1A1Ixp33_ASAP7_75t_L g791 ( 
.A1(n_629),
.A2(n_535),
.B(n_504),
.C(n_545),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_661),
.B(n_553),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_627),
.A2(n_555),
.B(n_607),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_701),
.B(n_535),
.Y(n_794)
);

CKINVDCx8_ASAP7_75t_R g795 ( 
.A(n_687),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_686),
.Y(n_796)
);

O2A1O1Ixp33_ASAP7_75t_L g797 ( 
.A1(n_638),
.A2(n_656),
.B(n_671),
.C(n_658),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_627),
.A2(n_555),
.B(n_607),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_717),
.B(n_722),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_618),
.Y(n_800)
);

NAND2x1_ASAP7_75t_L g801 ( 
.A(n_720),
.B(n_478),
.Y(n_801)
);

BUFx3_ASAP7_75t_L g802 ( 
.A(n_719),
.Y(n_802)
);

AOI21xp5_ASAP7_75t_L g803 ( 
.A1(n_765),
.A2(n_555),
.B(n_607),
.Y(n_803)
);

AOI21xp5_ASAP7_75t_L g804 ( 
.A1(n_765),
.A2(n_521),
.B(n_557),
.Y(n_804)
);

BUFx6f_ASAP7_75t_L g805 ( 
.A(n_710),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_731),
.B(n_545),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_635),
.B(n_435),
.Y(n_807)
);

AOI21xp5_ASAP7_75t_L g808 ( 
.A1(n_733),
.A2(n_521),
.B(n_557),
.Y(n_808)
);

INVx3_ASAP7_75t_L g809 ( 
.A(n_661),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_662),
.B(n_769),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_759),
.A2(n_521),
.B(n_557),
.Y(n_811)
);

NOR2x1_ASAP7_75t_R g812 ( 
.A(n_711),
.B(n_517),
.Y(n_812)
);

HB1xp67_ASAP7_75t_L g813 ( 
.A(n_621),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_763),
.A2(n_553),
.B(n_557),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_676),
.B(n_559),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_664),
.A2(n_557),
.B(n_553),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_664),
.A2(n_553),
.B(n_590),
.Y(n_817)
);

INVx3_ASAP7_75t_L g818 ( 
.A(n_632),
.Y(n_818)
);

AOI21xp5_ASAP7_75t_L g819 ( 
.A1(n_723),
.A2(n_724),
.B(n_653),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_715),
.B(n_561),
.Y(n_820)
);

AND2x2_ASAP7_75t_SL g821 ( 
.A(n_682),
.B(n_454),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_728),
.A2(n_561),
.B(n_595),
.C(n_603),
.Y(n_822)
);

NAND3xp33_ASAP7_75t_L g823 ( 
.A(n_728),
.B(n_282),
.C(n_276),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_723),
.A2(n_590),
.B(n_561),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_649),
.A2(n_595),
.B1(n_606),
.B2(n_603),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_696),
.Y(n_826)
);

O2A1O1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_655),
.A2(n_511),
.B(n_526),
.C(n_500),
.Y(n_827)
);

AOI21xp5_ASAP7_75t_L g828 ( 
.A1(n_724),
.A2(n_651),
.B(n_633),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_649),
.B(n_595),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_654),
.B(n_478),
.Y(n_830)
);

BUFx2_ASAP7_75t_L g831 ( 
.A(n_719),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_694),
.A2(n_590),
.B(n_606),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_636),
.B(n_266),
.C(n_249),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_654),
.B(n_478),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_614),
.A2(n_666),
.B(n_642),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_621),
.B(n_478),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_640),
.Y(n_837)
);

BUFx12f_ASAP7_75t_L g838 ( 
.A(n_746),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_645),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_744),
.B(n_720),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_632),
.Y(n_841)
);

NOR2xp33_ASAP7_75t_L g842 ( 
.A(n_639),
.B(n_512),
.Y(n_842)
);

A2O1A1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_734),
.A2(n_512),
.B(n_606),
.C(n_603),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_SL g844 ( 
.A(n_735),
.B(n_734),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_648),
.Y(n_845)
);

AOI21xp5_ASAP7_75t_L g846 ( 
.A1(n_622),
.A2(n_590),
.B(n_603),
.Y(n_846)
);

AOI21x1_ASAP7_75t_L g847 ( 
.A1(n_750),
.A2(n_507),
.B(n_500),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_695),
.B(n_452),
.Y(n_848)
);

AOI21xp5_ASAP7_75t_L g849 ( 
.A1(n_699),
.A2(n_706),
.B(n_702),
.Y(n_849)
);

AOI22xp33_ASAP7_75t_L g850 ( 
.A1(n_742),
.A2(n_492),
.B1(n_496),
.B2(n_311),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_619),
.B(n_637),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_634),
.B(n_512),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_687),
.Y(n_853)
);

AOI21xp5_ASAP7_75t_L g854 ( 
.A1(n_708),
.A2(n_514),
.B(n_594),
.Y(n_854)
);

O2A1O1Ixp5_ASAP7_75t_L g855 ( 
.A1(n_650),
.A2(n_511),
.B(n_507),
.C(n_510),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_644),
.B(n_514),
.Y(n_856)
);

AOI21x1_ASAP7_75t_L g857 ( 
.A1(n_750),
.A2(n_564),
.B(n_519),
.Y(n_857)
);

INVx1_ASAP7_75t_SL g858 ( 
.A(n_760),
.Y(n_858)
);

BUFx4f_ASAP7_75t_L g859 ( 
.A(n_687),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_764),
.Y(n_860)
);

INVx2_ASAP7_75t_L g861 ( 
.A(n_677),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_695),
.B(n_514),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_677),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_669),
.A2(n_594),
.B(n_531),
.Y(n_864)
);

AOI22xp33_ASAP7_75t_L g865 ( 
.A1(n_742),
.A2(n_492),
.B1(n_496),
.B2(n_311),
.Y(n_865)
);

BUFx8_ASAP7_75t_L g866 ( 
.A(n_665),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_683),
.B(n_519),
.Y(n_867)
);

NOR2x1p5_ASAP7_75t_L g868 ( 
.A(n_616),
.B(n_240),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_675),
.A2(n_582),
.B(n_583),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_670),
.B(n_743),
.Y(n_870)
);

AND2x4_ASAP7_75t_L g871 ( 
.A(n_737),
.B(n_439),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_652),
.A2(n_582),
.B(n_531),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_698),
.B(n_703),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_657),
.Y(n_874)
);

O2A1O1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_647),
.A2(n_419),
.B(n_592),
.C(n_589),
.Y(n_875)
);

AO21x1_ASAP7_75t_L g876 ( 
.A1(n_650),
.A2(n_609),
.B(n_592),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_737),
.B(n_452),
.Y(n_877)
);

OAI321xp33_ASAP7_75t_L g878 ( 
.A1(n_700),
.A2(n_685),
.A3(n_725),
.B1(n_727),
.B2(n_718),
.C(n_659),
.Y(n_878)
);

AOI21xp5_ASAP7_75t_L g879 ( 
.A1(n_646),
.A2(n_667),
.B(n_766),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_681),
.B(n_439),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_667),
.A2(n_609),
.B(n_452),
.Y(n_881)
);

AOI21xp5_ASAP7_75t_L g882 ( 
.A1(n_667),
.A2(n_452),
.B(n_414),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_714),
.B(n_492),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_714),
.B(n_496),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_667),
.A2(n_452),
.B(n_414),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_680),
.A2(n_707),
.B(n_678),
.Y(n_886)
);

AOI21xp5_ASAP7_75t_L g887 ( 
.A1(n_678),
.A2(n_452),
.B(n_414),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_692),
.B(n_496),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_684),
.A2(n_452),
.B(n_414),
.Y(n_889)
);

BUFx4f_ASAP7_75t_L g890 ( 
.A(n_682),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_693),
.B(n_292),
.Y(n_891)
);

A2O1A1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_727),
.A2(n_434),
.B(n_428),
.C(n_436),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_SL g893 ( 
.A1(n_625),
.A2(n_274),
.B1(n_264),
.B2(n_259),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_726),
.B(n_316),
.Y(n_894)
);

OAI21xp33_ASAP7_75t_L g895 ( 
.A1(n_713),
.A2(n_304),
.B(n_247),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_732),
.B(n_241),
.Y(n_896)
);

OAI22xp33_ASAP7_75t_L g897 ( 
.A1(n_625),
.A2(n_716),
.B1(n_704),
.B2(n_615),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_690),
.A2(n_414),
.B(n_428),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_709),
.B(n_704),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_758),
.B(n_441),
.Y(n_900)
);

BUFx12f_ASAP7_75t_L g901 ( 
.A(n_643),
.Y(n_901)
);

AOI22xp5_ASAP7_75t_L g902 ( 
.A1(n_747),
.A2(n_419),
.B1(n_310),
.B2(n_311),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_L g903 ( 
.A(n_749),
.B(n_250),
.Y(n_903)
);

OAI22xp5_ASAP7_75t_L g904 ( 
.A1(n_643),
.A2(n_428),
.B1(n_436),
.B2(n_434),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_709),
.B(n_428),
.Y(n_905)
);

INVx2_ASAP7_75t_L g906 ( 
.A(n_721),
.Y(n_906)
);

A2O1A1Ixp33_ASAP7_75t_L g907 ( 
.A1(n_751),
.A2(n_753),
.B(n_754),
.C(n_713),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_691),
.A2(n_414),
.B(n_428),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_647),
.B(n_428),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_721),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_697),
.A2(n_436),
.B(n_434),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_738),
.A2(n_436),
.B(n_434),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_752),
.A2(n_436),
.B(n_434),
.Y(n_913)
);

OAI21xp33_ASAP7_75t_L g914 ( 
.A1(n_668),
.A2(n_673),
.B(n_283),
.Y(n_914)
);

NOR2xp33_ASAP7_75t_L g915 ( 
.A(n_665),
.B(n_253),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_730),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_755),
.A2(n_436),
.B(n_434),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_730),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_625),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_740),
.B(n_292),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_747),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_736),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_756),
.A2(n_443),
.B(n_426),
.Y(n_923)
);

INVxp67_ASAP7_75t_L g924 ( 
.A(n_747),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_736),
.B(n_419),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_739),
.B(n_443),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_705),
.A2(n_443),
.B(n_426),
.Y(n_927)
);

AO21x2_ASAP7_75t_L g928 ( 
.A1(n_712),
.A2(n_441),
.B(n_443),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_768),
.A2(n_302),
.B1(n_296),
.B2(n_297),
.Y(n_929)
);

AND2x4_ASAP7_75t_L g930 ( 
.A(n_745),
.B(n_767),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_745),
.A2(n_426),
.B(n_424),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_804),
.A2(n_803),
.B(n_849),
.Y(n_932)
);

AND2x4_ASAP7_75t_L g933 ( 
.A(n_813),
.B(n_761),
.Y(n_933)
);

BUFx6f_ASAP7_75t_L g934 ( 
.A(n_784),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_784),
.Y(n_935)
);

A2O1A1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_773),
.A2(n_761),
.B(n_757),
.C(n_748),
.Y(n_936)
);

BUFx2_ASAP7_75t_L g937 ( 
.A(n_775),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_813),
.B(n_757),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_828),
.A2(n_688),
.B(n_426),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_R g940 ( 
.A(n_776),
.B(n_287),
.Y(n_940)
);

OR2x6_ASAP7_75t_SL g941 ( 
.A(n_780),
.B(n_298),
.Y(n_941)
);

AOI21xp5_ASAP7_75t_L g942 ( 
.A1(n_829),
.A2(n_688),
.B(n_424),
.Y(n_942)
);

BUFx3_ASAP7_75t_L g943 ( 
.A(n_838),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_779),
.B(n_424),
.Y(n_944)
);

AND2x4_ASAP7_75t_L g945 ( 
.A(n_784),
.B(n_424),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_844),
.B(n_307),
.Y(n_946)
);

A2O1A1Ixp33_ASAP7_75t_L g947 ( 
.A1(n_878),
.A2(n_689),
.B(n_301),
.C(n_431),
.Y(n_947)
);

BUFx2_ASAP7_75t_L g948 ( 
.A(n_775),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_862),
.A2(n_431),
.B(n_130),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_874),
.A2(n_311),
.B1(n_310),
.B2(n_292),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_779),
.B(n_431),
.Y(n_951)
);

BUFx3_ASAP7_75t_L g952 ( 
.A(n_866),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_799),
.B(n_311),
.Y(n_953)
);

AND2x2_ASAP7_75t_L g954 ( 
.A(n_858),
.B(n_431),
.Y(n_954)
);

A2O1A1Ixp33_ASAP7_75t_SL g955 ( 
.A1(n_870),
.A2(n_310),
.B(n_106),
.C(n_158),
.Y(n_955)
);

A2O1A1Ixp33_ASAP7_75t_L g956 ( 
.A1(n_870),
.A2(n_431),
.B(n_310),
.C(n_10),
.Y(n_956)
);

XOR2xp5_ASAP7_75t_L g957 ( 
.A(n_831),
.B(n_154),
.Y(n_957)
);

NAND2x1p5_ASAP7_75t_L g958 ( 
.A(n_919),
.B(n_431),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_837),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_772),
.A2(n_3),
.B(n_7),
.C(n_12),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_842),
.B(n_431),
.Y(n_961)
);

INVxp67_ASAP7_75t_L g962 ( 
.A(n_826),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_839),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_930),
.Y(n_964)
);

O2A1O1Ixp5_ASAP7_75t_L g965 ( 
.A1(n_920),
.A2(n_310),
.B(n_152),
.C(n_148),
.Y(n_965)
);

AOI21x1_ASAP7_75t_L g966 ( 
.A1(n_862),
.A2(n_139),
.B(n_136),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_796),
.B(n_133),
.Y(n_967)
);

A2O1A1Ixp33_ASAP7_75t_L g968 ( 
.A1(n_797),
.A2(n_3),
.B(n_7),
.C(n_13),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_807),
.B(n_14),
.Y(n_969)
);

BUFx2_ASAP7_75t_L g970 ( 
.A(n_853),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_860),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_771),
.A2(n_808),
.B(n_811),
.Y(n_972)
);

A2O1A1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_815),
.A2(n_16),
.B(n_20),
.C(n_21),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_815),
.B(n_16),
.Y(n_974)
);

HB1xp67_ASAP7_75t_L g975 ( 
.A(n_840),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_866),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_930),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_819),
.A2(n_98),
.B(n_91),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_848),
.A2(n_86),
.B(n_83),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_770),
.A2(n_80),
.B(n_64),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_772),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_796),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_SL g983 ( 
.A(n_796),
.B(n_62),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_805),
.Y(n_984)
);

NOR2xp67_ASAP7_75t_SL g985 ( 
.A(n_795),
.B(n_21),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_880),
.B(n_22),
.Y(n_986)
);

O2A1O1Ixp33_ASAP7_75t_L g987 ( 
.A1(n_810),
.A2(n_24),
.B(n_27),
.C(n_29),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_851),
.B(n_27),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_L g989 ( 
.A(n_894),
.B(n_32),
.Y(n_989)
);

AND2x2_ASAP7_75t_L g990 ( 
.A(n_894),
.B(n_32),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_777),
.A2(n_56),
.B(n_53),
.Y(n_991)
);

AND2x2_ASAP7_75t_L g992 ( 
.A(n_896),
.B(n_35),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_873),
.B(n_820),
.Y(n_993)
);

AND2x4_ASAP7_75t_L g994 ( 
.A(n_805),
.B(n_36),
.Y(n_994)
);

AOI21xp5_ASAP7_75t_L g995 ( 
.A1(n_782),
.A2(n_36),
.B(n_37),
.Y(n_995)
);

OAI22xp5_ASAP7_75t_L g996 ( 
.A1(n_787),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_883),
.A2(n_42),
.B(n_44),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_805),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_802),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_787),
.A2(n_42),
.B1(n_44),
.B2(n_49),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_884),
.A2(n_52),
.B(n_879),
.Y(n_1001)
);

OAI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_899),
.A2(n_924),
.B1(n_921),
.B2(n_781),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_814),
.A2(n_846),
.B(n_834),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_924),
.A2(n_865),
.B1(n_850),
.B2(n_897),
.Y(n_1004)
);

NAND2xp33_ASAP7_75t_L g1005 ( 
.A(n_774),
.B(n_914),
.Y(n_1005)
);

A2O1A1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_823),
.A2(n_820),
.B(n_859),
.C(n_903),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_806),
.B(n_800),
.Y(n_1007)
);

BUFx8_ASAP7_75t_L g1008 ( 
.A(n_901),
.Y(n_1008)
);

A2O1A1Ixp33_ASAP7_75t_L g1009 ( 
.A1(n_859),
.A2(n_896),
.B(n_903),
.C(n_835),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_821),
.B(n_890),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_830),
.A2(n_778),
.B(n_897),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_872),
.A2(n_793),
.B(n_798),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_890),
.B(n_893),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_812),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_845),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_871),
.B(n_868),
.Y(n_1016)
);

O2A1O1Ixp33_ASAP7_75t_L g1017 ( 
.A1(n_929),
.A2(n_920),
.B(n_900),
.C(n_833),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_833),
.A2(n_871),
.B1(n_893),
.B2(n_836),
.Y(n_1018)
);

O2A1O1Ixp5_ASAP7_75t_L g1019 ( 
.A1(n_886),
.A2(n_876),
.B(n_791),
.C(n_822),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_915),
.B(n_794),
.Y(n_1020)
);

BUFx3_ASAP7_75t_L g1021 ( 
.A(n_919),
.Y(n_1021)
);

BUFx6f_ASAP7_75t_L g1022 ( 
.A(n_788),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_915),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_895),
.Y(n_1024)
);

BUFx4f_ASAP7_75t_L g1025 ( 
.A(n_788),
.Y(n_1025)
);

INVx2_ASAP7_75t_SL g1026 ( 
.A(n_809),
.Y(n_1026)
);

NAND2x1p5_ASAP7_75t_L g1027 ( 
.A(n_809),
.B(n_818),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_861),
.B(n_863),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_818),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_910),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_841),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_786),
.A2(n_832),
.B(n_785),
.Y(n_1032)
);

O2A1O1Ixp33_ASAP7_75t_SL g1033 ( 
.A1(n_843),
.A2(n_892),
.B(n_907),
.C(n_852),
.Y(n_1033)
);

INVxp67_ASAP7_75t_L g1034 ( 
.A(n_891),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_SL g1035 ( 
.A1(n_902),
.A2(n_850),
.B(n_865),
.C(n_827),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_906),
.Y(n_1036)
);

AND2x2_ASAP7_75t_L g1037 ( 
.A(n_916),
.B(n_922),
.Y(n_1037)
);

HB1xp67_ASAP7_75t_L g1038 ( 
.A(n_918),
.Y(n_1038)
);

CKINVDCx14_ASAP7_75t_R g1039 ( 
.A(n_888),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_867),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_790),
.A2(n_816),
.B(n_817),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_783),
.B(n_905),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_877),
.A2(n_856),
.B(n_852),
.C(n_825),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_789),
.A2(n_792),
.B1(n_925),
.B2(n_909),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_847),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_926),
.Y(n_1046)
);

BUFx2_ASAP7_75t_L g1047 ( 
.A(n_928),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_928),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_789),
.A2(n_792),
.B1(n_801),
.B2(n_904),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_923),
.Y(n_1050)
);

OR2x6_ASAP7_75t_L g1051 ( 
.A(n_854),
.B(n_824),
.Y(n_1051)
);

OAI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_864),
.A2(n_917),
.B(n_912),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_869),
.A2(n_911),
.B1(n_913),
.B2(n_908),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_881),
.B(n_882),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_875),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_857),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_927),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_898),
.B(n_889),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_931),
.Y(n_1059)
);

BUFx5_ASAP7_75t_L g1060 ( 
.A(n_855),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_L g1061 ( 
.A1(n_1009),
.A2(n_855),
.B(n_887),
.C(n_885),
.Y(n_1061)
);

NOR2xp33_ASAP7_75t_L g1062 ( 
.A(n_1020),
.B(n_962),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_1003),
.A2(n_1032),
.B(n_1011),
.Y(n_1064)
);

BUFx2_ASAP7_75t_R g1065 ( 
.A(n_952),
.Y(n_1065)
);

AOI21xp5_ASAP7_75t_L g1066 ( 
.A1(n_1005),
.A2(n_993),
.B(n_1041),
.Y(n_1066)
);

NOR2xp33_ASAP7_75t_L g1067 ( 
.A(n_1023),
.B(n_981),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_981),
.B(n_1040),
.Y(n_1068)
);

AO32x2_ASAP7_75t_L g1069 ( 
.A1(n_1002),
.A2(n_1004),
.A3(n_996),
.B1(n_1000),
.B2(n_1044),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_975),
.B(n_986),
.Y(n_1070)
);

NOR2xp67_ASAP7_75t_L g1071 ( 
.A(n_1018),
.B(n_964),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_939),
.A2(n_1053),
.B(n_1045),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_L g1073 ( 
.A1(n_1053),
.A2(n_1056),
.B(n_1019),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_992),
.B(n_969),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_1030),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1058),
.A2(n_1033),
.B(n_1006),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1024),
.B(n_954),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_959),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1046),
.B(n_1038),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_934),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_988),
.B(n_944),
.Y(n_1081)
);

INVxp67_ASAP7_75t_L g1082 ( 
.A(n_937),
.Y(n_1082)
);

AOI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_989),
.A2(n_1039),
.B1(n_1000),
.B2(n_996),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_973),
.A2(n_1013),
.B(n_968),
.C(n_956),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_990),
.B(n_970),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1007),
.B(n_933),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_SL g1087 ( 
.A(n_985),
.B(n_1021),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_1016),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_SL g1089 ( 
.A1(n_978),
.A2(n_955),
.B(n_983),
.C(n_967),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_961),
.A2(n_1051),
.B(n_1017),
.Y(n_1090)
);

AO31x2_ASAP7_75t_L g1091 ( 
.A1(n_1047),
.A2(n_1048),
.A3(n_1002),
.B(n_1001),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_963),
.Y(n_1092)
);

AND2x2_ASAP7_75t_SL g1093 ( 
.A(n_994),
.B(n_976),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_SL g1094 ( 
.A(n_1008),
.B(n_994),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_1051),
.A2(n_1042),
.B(n_1052),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_948),
.B(n_946),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_942),
.A2(n_1054),
.B(n_1049),
.Y(n_1097)
);

OAI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_974),
.A2(n_1004),
.B1(n_999),
.B2(n_943),
.Y(n_1098)
);

AOI221x1_ASAP7_75t_L g1099 ( 
.A1(n_980),
.A2(n_978),
.B1(n_997),
.B2(n_995),
.C(n_1049),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1043),
.A2(n_1007),
.B(n_1044),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_951),
.A2(n_936),
.B(n_1050),
.Y(n_1101)
);

INVx2_ASAP7_75t_L g1102 ( 
.A(n_1037),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_953),
.A2(n_949),
.B(n_1010),
.Y(n_1103)
);

CKINVDCx11_ASAP7_75t_R g1104 ( 
.A(n_941),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1028),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_940),
.Y(n_1106)
);

INVx3_ASAP7_75t_L g1107 ( 
.A(n_1031),
.Y(n_1107)
);

A2O1A1Ixp33_ASAP7_75t_L g1108 ( 
.A1(n_987),
.A2(n_1034),
.B(n_960),
.C(n_965),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1057),
.A2(n_966),
.B(n_1059),
.Y(n_1109)
);

AO31x2_ASAP7_75t_L g1110 ( 
.A1(n_1055),
.A2(n_947),
.A3(n_991),
.B(n_979),
.Y(n_1110)
);

AND2x2_ASAP7_75t_L g1111 ( 
.A(n_1016),
.B(n_1029),
.Y(n_1111)
);

AO32x2_ASAP7_75t_L g1112 ( 
.A1(n_984),
.A2(n_1026),
.A3(n_1060),
.B1(n_950),
.B2(n_1015),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_977),
.A2(n_1036),
.B(n_1025),
.C(n_938),
.Y(n_1113)
);

AOI221xp5_ASAP7_75t_L g1114 ( 
.A1(n_1014),
.A2(n_971),
.B1(n_957),
.B2(n_933),
.C(n_938),
.Y(n_1114)
);

OAI22x1_ASAP7_75t_L g1115 ( 
.A1(n_1027),
.A2(n_984),
.B1(n_945),
.B2(n_958),
.Y(n_1115)
);

AOI22xp5_ASAP7_75t_L g1116 ( 
.A1(n_1008),
.A2(n_1031),
.B1(n_935),
.B2(n_982),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1022),
.Y(n_1117)
);

OAI22xp33_ASAP7_75t_L g1118 ( 
.A1(n_934),
.A2(n_935),
.B1(n_982),
.B2(n_998),
.Y(n_1118)
);

O2A1O1Ixp33_ASAP7_75t_SL g1119 ( 
.A1(n_1060),
.A2(n_958),
.B(n_1022),
.C(n_934),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_935),
.A2(n_982),
.B(n_998),
.Y(n_1120)
);

OA21x2_ASAP7_75t_L g1121 ( 
.A1(n_1060),
.A2(n_1022),
.B(n_998),
.Y(n_1121)
);

BUFx12f_ASAP7_75t_L g1122 ( 
.A(n_1060),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1060),
.B(n_1021),
.Y(n_1123)
);

OR2x2_ASAP7_75t_L g1124 ( 
.A(n_962),
.B(n_506),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_937),
.Y(n_1126)
);

AOI221x1_ASAP7_75t_L g1127 ( 
.A1(n_968),
.A2(n_1001),
.B1(n_989),
.B2(n_980),
.C(n_1009),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_937),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_1037),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1047),
.A2(n_1048),
.A3(n_1011),
.B(n_1002),
.Y(n_1130)
);

AOI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_989),
.A2(n_773),
.B1(n_674),
.B2(n_660),
.Y(n_1131)
);

INVx1_ASAP7_75t_SL g1132 ( 
.A(n_937),
.Y(n_1132)
);

AO31x2_ASAP7_75t_L g1133 ( 
.A1(n_1047),
.A2(n_1048),
.A3(n_1011),
.B(n_1002),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_934),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1020),
.B(n_773),
.Y(n_1135)
);

OR2x2_ASAP7_75t_L g1136 ( 
.A(n_962),
.B(n_506),
.Y(n_1136)
);

A2O1A1Ixp33_ASAP7_75t_L g1137 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.C(n_674),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.C(n_674),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1030),
.Y(n_1139)
);

A2O1A1Ixp33_ASAP7_75t_L g1140 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.C(n_674),
.Y(n_1140)
);

AOI22xp33_ASAP7_75t_L g1141 ( 
.A1(n_992),
.A2(n_674),
.B1(n_660),
.B2(n_989),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_1012),
.A2(n_972),
.B(n_1032),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1037),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1012),
.A2(n_972),
.B(n_1032),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_SL g1146 ( 
.A1(n_1009),
.A2(n_1006),
.B(n_978),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_969),
.B(n_617),
.Y(n_1147)
);

BUFx2_ASAP7_75t_SL g1148 ( 
.A(n_1021),
.Y(n_1148)
);

AO32x2_ASAP7_75t_L g1149 ( 
.A1(n_1002),
.A2(n_1004),
.A3(n_1000),
.B1(n_996),
.B2(n_874),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1030),
.Y(n_1150)
);

O2A1O1Ixp33_ASAP7_75t_SL g1151 ( 
.A1(n_1009),
.A2(n_1006),
.B(n_1035),
.C(n_968),
.Y(n_1151)
);

OA21x2_ASAP7_75t_L g1152 ( 
.A1(n_1019),
.A2(n_1011),
.B(n_1041),
.Y(n_1152)
);

INVx2_ASAP7_75t_SL g1153 ( 
.A(n_937),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1030),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1155)
);

INVxp67_ASAP7_75t_L g1156 ( 
.A(n_937),
.Y(n_1156)
);

INVx2_ASAP7_75t_SL g1157 ( 
.A(n_937),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1158)
);

BUFx10_ASAP7_75t_L g1159 ( 
.A(n_1016),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1012),
.A2(n_972),
.B(n_1032),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1012),
.A2(n_972),
.B(n_1032),
.Y(n_1161)
);

AO31x2_ASAP7_75t_L g1162 ( 
.A1(n_1047),
.A2(n_1048),
.A3(n_1011),
.B(n_1002),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1030),
.Y(n_1163)
);

AO21x1_ASAP7_75t_L g1164 ( 
.A1(n_1017),
.A2(n_773),
.B(n_978),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1047),
.A2(n_1048),
.A3(n_1011),
.B(n_1002),
.Y(n_1165)
);

OAI22xp5_ASAP7_75t_L g1166 ( 
.A1(n_1020),
.A2(n_773),
.B1(n_660),
.B2(n_799),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_962),
.B(n_506),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1168)
);

OAI21x1_ASAP7_75t_L g1169 ( 
.A1(n_1012),
.A2(n_972),
.B(n_1032),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_1030),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1030),
.Y(n_1171)
);

OA21x2_ASAP7_75t_L g1172 ( 
.A1(n_1019),
.A2(n_1011),
.B(n_1041),
.Y(n_1172)
);

O2A1O1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_989),
.A2(n_660),
.B(n_878),
.C(n_762),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1020),
.A2(n_773),
.B1(n_660),
.B2(n_799),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_937),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_989),
.A2(n_660),
.B(n_878),
.C(n_762),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_L g1180 ( 
.A(n_1020),
.B(n_773),
.Y(n_1180)
);

INVxp67_ASAP7_75t_L g1181 ( 
.A(n_937),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1037),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.C(n_674),
.Y(n_1183)
);

BUFx2_ASAP7_75t_L g1184 ( 
.A(n_962),
.Y(n_1184)
);

BUFx2_ASAP7_75t_R g1185 ( 
.A(n_952),
.Y(n_1185)
);

A2O1A1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.C(n_674),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_932),
.A2(n_972),
.B(n_1012),
.Y(n_1187)
);

AO22x2_ASAP7_75t_L g1188 ( 
.A1(n_996),
.A2(n_1000),
.B1(n_1004),
.B2(n_1002),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_989),
.A2(n_660),
.B(n_878),
.C(n_762),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_SL g1190 ( 
.A1(n_978),
.A2(n_797),
.B(n_1002),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1037),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_962),
.Y(n_1192)
);

OAI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1009),
.A2(n_773),
.B(n_660),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1020),
.B(n_773),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_962),
.Y(n_1195)
);

OA21x2_ASAP7_75t_L g1196 ( 
.A1(n_1019),
.A2(n_1011),
.B(n_1041),
.Y(n_1196)
);

CKINVDCx20_ASAP7_75t_R g1197 ( 
.A(n_1106),
.Y(n_1197)
);

OAI22xp5_ASAP7_75t_L g1198 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_1083),
.B2(n_1180),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_SL g1199 ( 
.A1(n_1188),
.A2(n_1135),
.B1(n_1194),
.B2(n_1193),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1075),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1188),
.A2(n_1166),
.B1(n_1174),
.B2(n_1087),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_1184),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1078),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1087),
.A2(n_1094),
.B1(n_1093),
.B2(n_1076),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1131),
.A2(n_1164),
.B1(n_1083),
.B2(n_1098),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1092),
.Y(n_1206)
);

BUFx4f_ASAP7_75t_L g1207 ( 
.A(n_1080),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1137),
.A2(n_1183),
.B1(n_1186),
.B2(n_1140),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1190),
.A2(n_1147),
.B1(n_1081),
.B2(n_1071),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_SL g1210 ( 
.A1(n_1094),
.A2(n_1062),
.B1(n_1067),
.B2(n_1074),
.Y(n_1210)
);

AOI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1077),
.A2(n_1096),
.B1(n_1068),
.B2(n_1085),
.Y(n_1211)
);

INVx1_ASAP7_75t_SL g1212 ( 
.A(n_1192),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_SL g1213 ( 
.A1(n_1070),
.A2(n_1086),
.B1(n_1189),
.B2(n_1173),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1088),
.Y(n_1214)
);

INVx6_ASAP7_75t_L g1215 ( 
.A(n_1088),
.Y(n_1215)
);

CKINVDCx11_ASAP7_75t_R g1216 ( 
.A(n_1104),
.Y(n_1216)
);

BUFx4_ASAP7_75t_SL g1217 ( 
.A(n_1124),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1063),
.A2(n_1125),
.B(n_1168),
.Y(n_1218)
);

BUFx8_ASAP7_75t_L g1219 ( 
.A(n_1195),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1071),
.A2(n_1114),
.B1(n_1123),
.B2(n_1182),
.Y(n_1220)
);

AOI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1123),
.A2(n_1102),
.B1(n_1191),
.B2(n_1129),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1143),
.B(n_1179),
.Y(n_1222)
);

AND2x4_ASAP7_75t_L g1223 ( 
.A(n_1111),
.B(n_1116),
.Y(n_1223)
);

CKINVDCx11_ASAP7_75t_R g1224 ( 
.A(n_1159),
.Y(n_1224)
);

BUFx10_ASAP7_75t_L g1225 ( 
.A(n_1153),
.Y(n_1225)
);

BUFx2_ASAP7_75t_SL g1226 ( 
.A(n_1157),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1175),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_SL g1228 ( 
.A1(n_1069),
.A2(n_1138),
.B1(n_1149),
.B2(n_1146),
.Y(n_1228)
);

OAI22xp33_ASAP7_75t_L g1229 ( 
.A1(n_1079),
.A2(n_1127),
.B1(n_1167),
.B2(n_1136),
.Y(n_1229)
);

AOI22xp33_ASAP7_75t_SL g1230 ( 
.A1(n_1069),
.A2(n_1149),
.B1(n_1095),
.B2(n_1100),
.Y(n_1230)
);

BUFx12f_ASAP7_75t_L g1231 ( 
.A(n_1159),
.Y(n_1231)
);

OAI22xp5_ASAP7_75t_L g1232 ( 
.A1(n_1132),
.A2(n_1113),
.B1(n_1156),
.B2(n_1082),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_SL g1233 ( 
.A1(n_1132),
.A2(n_1148),
.B1(n_1116),
.B2(n_1128),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1069),
.A2(n_1149),
.B1(n_1066),
.B2(n_1196),
.Y(n_1234)
);

AOI22xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1152),
.A2(n_1196),
.B1(n_1172),
.B2(n_1163),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1152),
.A2(n_1172),
.B1(n_1170),
.B2(n_1171),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1181),
.A2(n_1108),
.B1(n_1139),
.B2(n_1150),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1154),
.A2(n_1105),
.B1(n_1101),
.B2(n_1084),
.Y(n_1238)
);

AOI22xp5_ASAP7_75t_L g1239 ( 
.A1(n_1151),
.A2(n_1122),
.B1(n_1089),
.B2(n_1090),
.Y(n_1239)
);

BUFx12f_ASAP7_75t_L g1240 ( 
.A(n_1080),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1065),
.Y(n_1241)
);

INVx4_ASAP7_75t_L g1242 ( 
.A(n_1134),
.Y(n_1242)
);

CKINVDCx11_ASAP7_75t_R g1243 ( 
.A(n_1185),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1091),
.Y(n_1244)
);

NAND2x1p5_ASAP7_75t_L g1245 ( 
.A(n_1121),
.B(n_1107),
.Y(n_1245)
);

BUFx3_ASAP7_75t_L g1246 ( 
.A(n_1134),
.Y(n_1246)
);

INVx1_ASAP7_75t_SL g1247 ( 
.A(n_1117),
.Y(n_1247)
);

AOI22xp33_ASAP7_75t_L g1248 ( 
.A1(n_1103),
.A2(n_1115),
.B1(n_1073),
.B2(n_1097),
.Y(n_1248)
);

INVxp67_ASAP7_75t_L g1249 ( 
.A(n_1120),
.Y(n_1249)
);

BUFx4f_ASAP7_75t_SL g1250 ( 
.A(n_1118),
.Y(n_1250)
);

AOI21xp5_ASAP7_75t_L g1251 ( 
.A1(n_1144),
.A2(n_1187),
.B(n_1178),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1064),
.A2(n_1072),
.B1(n_1177),
.B2(n_1176),
.Y(n_1252)
);

CKINVDCx11_ASAP7_75t_R g1253 ( 
.A(n_1119),
.Y(n_1253)
);

INVxp67_ASAP7_75t_SL g1254 ( 
.A(n_1109),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1130),
.B(n_1165),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1061),
.A2(n_1155),
.B1(n_1158),
.B2(n_1099),
.Y(n_1256)
);

BUFx2_ASAP7_75t_SL g1257 ( 
.A(n_1112),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1133),
.B(n_1165),
.Y(n_1258)
);

INVx5_ASAP7_75t_L g1259 ( 
.A(n_1110),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_SL g1260 ( 
.A1(n_1112),
.A2(n_1161),
.B1(n_1169),
.B2(n_1142),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1162),
.B(n_1165),
.Y(n_1261)
);

OAI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1091),
.A2(n_1110),
.B1(n_1112),
.B2(n_1162),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1162),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1145),
.Y(n_1264)
);

OAI22xp5_ASAP7_75t_L g1265 ( 
.A1(n_1160),
.A2(n_1131),
.B1(n_773),
.B2(n_1141),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_1180),
.B2(n_1135),
.Y(n_1266)
);

BUFx2_ASAP7_75t_L g1267 ( 
.A(n_1184),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1147),
.B(n_1085),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_1180),
.B2(n_1135),
.Y(n_1269)
);

CKINVDCx11_ASAP7_75t_R g1270 ( 
.A(n_1104),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_SL g1271 ( 
.A1(n_1188),
.A2(n_325),
.B1(n_335),
.B2(n_327),
.Y(n_1271)
);

CKINVDCx20_ASAP7_75t_R g1272 ( 
.A(n_1106),
.Y(n_1272)
);

BUFx8_ASAP7_75t_SL g1273 ( 
.A(n_1106),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1135),
.B(n_1180),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1106),
.Y(n_1275)
);

CKINVDCx11_ASAP7_75t_R g1276 ( 
.A(n_1104),
.Y(n_1276)
);

INVx4_ASAP7_75t_L g1277 ( 
.A(n_1080),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1075),
.Y(n_1278)
);

BUFx2_ASAP7_75t_L g1279 ( 
.A(n_1184),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1147),
.B(n_1085),
.Y(n_1280)
);

INVx1_ASAP7_75t_SL g1281 ( 
.A(n_1184),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_1184),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_674),
.B2(n_989),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1184),
.Y(n_1284)
);

INVx6_ASAP7_75t_L g1285 ( 
.A(n_1088),
.Y(n_1285)
);

OAI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1131),
.A2(n_773),
.B1(n_1180),
.B2(n_1135),
.Y(n_1286)
);

CKINVDCx11_ASAP7_75t_R g1287 ( 
.A(n_1104),
.Y(n_1287)
);

CKINVDCx20_ASAP7_75t_R g1288 ( 
.A(n_1106),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1102),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1075),
.Y(n_1290)
);

INVx1_ASAP7_75t_SL g1291 ( 
.A(n_1184),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1075),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1135),
.B(n_1180),
.Y(n_1293)
);

CKINVDCx6p67_ASAP7_75t_R g1294 ( 
.A(n_1148),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1075),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1184),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1131),
.A2(n_773),
.B1(n_1141),
.B2(n_1083),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1184),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1131),
.A2(n_773),
.B1(n_1141),
.B2(n_1083),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_674),
.B2(n_989),
.Y(n_1300)
);

AOI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_674),
.B2(n_989),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1131),
.A2(n_1141),
.B1(n_674),
.B2(n_989),
.Y(n_1302)
);

BUFx2_ASAP7_75t_SL g1303 ( 
.A(n_1126),
.Y(n_1303)
);

BUFx10_ASAP7_75t_L g1304 ( 
.A(n_1067),
.Y(n_1304)
);

CKINVDCx11_ASAP7_75t_R g1305 ( 
.A(n_1104),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1228),
.B(n_1199),
.Y(n_1306)
);

OA21x2_ASAP7_75t_L g1307 ( 
.A1(n_1218),
.A2(n_1251),
.B(n_1255),
.Y(n_1307)
);

OA21x2_ASAP7_75t_L g1308 ( 
.A1(n_1218),
.A2(n_1251),
.B(n_1258),
.Y(n_1308)
);

OR2x2_ASAP7_75t_L g1309 ( 
.A(n_1261),
.B(n_1244),
.Y(n_1309)
);

INVx8_ASAP7_75t_L g1310 ( 
.A(n_1240),
.Y(n_1310)
);

CKINVDCx5p33_ASAP7_75t_R g1311 ( 
.A(n_1273),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1245),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1244),
.B(n_1257),
.Y(n_1313)
);

OAI221xp5_ASAP7_75t_L g1314 ( 
.A1(n_1283),
.A2(n_1301),
.B1(n_1300),
.B2(n_1302),
.C(n_1271),
.Y(n_1314)
);

BUFx6f_ASAP7_75t_L g1315 ( 
.A(n_1253),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1228),
.B(n_1199),
.Y(n_1316)
);

AND2x2_ASAP7_75t_L g1317 ( 
.A(n_1230),
.B(n_1201),
.Y(n_1317)
);

INVx2_ASAP7_75t_L g1318 ( 
.A(n_1200),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1203),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1206),
.Y(n_1320)
);

OR2x2_ASAP7_75t_L g1321 ( 
.A(n_1265),
.B(n_1208),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1212),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1263),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_1284),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1230),
.B(n_1201),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1262),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1274),
.B(n_1293),
.Y(n_1327)
);

CKINVDCx6p67_ASAP7_75t_R g1328 ( 
.A(n_1241),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1249),
.B(n_1239),
.Y(n_1329)
);

AND2x2_ASAP7_75t_L g1330 ( 
.A(n_1205),
.B(n_1234),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1205),
.B(n_1234),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1236),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1236),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1254),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1219),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_1243),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1297),
.A2(n_1299),
.B1(n_1198),
.B2(n_1271),
.Y(n_1337)
);

OAI21x1_ASAP7_75t_L g1338 ( 
.A1(n_1252),
.A2(n_1256),
.B(n_1248),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1249),
.B(n_1259),
.Y(n_1339)
);

CKINVDCx20_ASAP7_75t_R g1340 ( 
.A(n_1197),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1216),
.Y(n_1341)
);

OAI21x1_ASAP7_75t_L g1342 ( 
.A1(n_1254),
.A2(n_1238),
.B(n_1209),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1268),
.B(n_1280),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_L g1344 ( 
.A1(n_1209),
.A2(n_1237),
.B(n_1290),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1227),
.Y(n_1345)
);

BUFx2_ASAP7_75t_L g1346 ( 
.A(n_1259),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1278),
.Y(n_1347)
);

OR2x2_ASAP7_75t_L g1348 ( 
.A(n_1222),
.B(n_1229),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1292),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1250),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1270),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1219),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1295),
.Y(n_1353)
);

HB1xp67_ASAP7_75t_L g1354 ( 
.A(n_1247),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1229),
.B(n_1211),
.Y(n_1355)
);

INVx4_ASAP7_75t_SL g1356 ( 
.A(n_1250),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1235),
.Y(n_1357)
);

AOI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1286),
.A2(n_1269),
.B1(n_1266),
.B2(n_1210),
.Y(n_1358)
);

HB1xp67_ASAP7_75t_L g1359 ( 
.A(n_1232),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1235),
.Y(n_1360)
);

AND2x4_ASAP7_75t_L g1361 ( 
.A(n_1264),
.B(n_1223),
.Y(n_1361)
);

OR2x6_ASAP7_75t_L g1362 ( 
.A(n_1233),
.B(n_1285),
.Y(n_1362)
);

NOR2xp33_ASAP7_75t_L g1363 ( 
.A(n_1281),
.B(n_1291),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1260),
.Y(n_1364)
);

INVxp67_ASAP7_75t_L g1365 ( 
.A(n_1202),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1260),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1289),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1213),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1286),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1267),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1221),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1220),
.A2(n_1204),
.B(n_1285),
.Y(n_1372)
);

AND2x4_ASAP7_75t_SL g1373 ( 
.A(n_1294),
.B(n_1225),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1214),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1279),
.A2(n_1296),
.B(n_1298),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1282),
.B(n_1226),
.Y(n_1376)
);

NAND2x1p5_ASAP7_75t_L g1377 ( 
.A(n_1329),
.B(n_1207),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1343),
.B(n_1304),
.Y(n_1378)
);

NAND3xp33_ASAP7_75t_L g1379 ( 
.A(n_1337),
.B(n_1224),
.C(n_1277),
.Y(n_1379)
);

O2A1O1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1314),
.A2(n_1246),
.B(n_1217),
.C(n_1304),
.Y(n_1380)
);

INVx2_ASAP7_75t_L g1381 ( 
.A(n_1318),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1307),
.A2(n_1207),
.B(n_1242),
.Y(n_1382)
);

BUFx2_ASAP7_75t_L g1383 ( 
.A(n_1345),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1358),
.A2(n_1303),
.B(n_1215),
.C(n_1214),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1358),
.A2(n_1214),
.B(n_1215),
.C(n_1285),
.Y(n_1385)
);

OAI21xp5_ASAP7_75t_L g1386 ( 
.A1(n_1368),
.A2(n_1272),
.B(n_1275),
.Y(n_1386)
);

OA21x2_ASAP7_75t_L g1387 ( 
.A1(n_1338),
.A2(n_1215),
.B(n_1231),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1350),
.A2(n_1276),
.B1(n_1287),
.B2(n_1305),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1327),
.B(n_1288),
.Y(n_1389)
);

A2O1A1Ixp33_ASAP7_75t_L g1390 ( 
.A1(n_1355),
.A2(n_1321),
.B(n_1306),
.C(n_1316),
.Y(n_1390)
);

AO32x2_ASAP7_75t_L g1391 ( 
.A1(n_1326),
.A2(n_1348),
.A3(n_1309),
.B1(n_1313),
.B2(n_1350),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1355),
.A2(n_1321),
.B(n_1316),
.C(n_1306),
.Y(n_1392)
);

INVxp67_ASAP7_75t_L g1393 ( 
.A(n_1368),
.Y(n_1393)
);

CKINVDCx5p33_ASAP7_75t_R g1394 ( 
.A(n_1311),
.Y(n_1394)
);

BUFx4f_ASAP7_75t_SL g1395 ( 
.A(n_1340),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1370),
.B(n_1345),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1317),
.A2(n_1325),
.B1(n_1359),
.B2(n_1330),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1307),
.A2(n_1308),
.B(n_1338),
.Y(n_1398)
);

NAND2xp5_ASAP7_75t_L g1399 ( 
.A(n_1369),
.B(n_1354),
.Y(n_1399)
);

CKINVDCx20_ASAP7_75t_R g1400 ( 
.A(n_1336),
.Y(n_1400)
);

NOR2xp33_ASAP7_75t_L g1401 ( 
.A(n_1348),
.B(n_1329),
.Y(n_1401)
);

OR2x2_ASAP7_75t_L g1402 ( 
.A(n_1319),
.B(n_1320),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1344),
.B(n_1342),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1329),
.B(n_1375),
.Y(n_1404)
);

AO32x2_ASAP7_75t_L g1405 ( 
.A1(n_1326),
.A2(n_1313),
.A3(n_1350),
.B1(n_1366),
.B2(n_1364),
.Y(n_1405)
);

BUFx2_ASAP7_75t_L g1406 ( 
.A(n_1324),
.Y(n_1406)
);

AND4x1_ASAP7_75t_L g1407 ( 
.A(n_1363),
.B(n_1317),
.C(n_1325),
.D(n_1330),
.Y(n_1407)
);

INVx1_ASAP7_75t_SL g1408 ( 
.A(n_1322),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1362),
.A2(n_1356),
.B1(n_1371),
.B2(n_1372),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1307),
.A2(n_1308),
.B(n_1339),
.Y(n_1410)
);

AND2x4_ASAP7_75t_L g1411 ( 
.A(n_1361),
.B(n_1312),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1334),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1362),
.A2(n_1356),
.B1(n_1371),
.B2(n_1331),
.Y(n_1413)
);

INVxp67_ASAP7_75t_L g1414 ( 
.A(n_1347),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_L g1415 ( 
.A(n_1393),
.B(n_1365),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1412),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1391),
.B(n_1403),
.Y(n_1417)
);

OR2x2_ASAP7_75t_SL g1418 ( 
.A(n_1387),
.B(n_1315),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1393),
.B(n_1376),
.Y(n_1419)
);

BUFx2_ASAP7_75t_L g1420 ( 
.A(n_1391),
.Y(n_1420)
);

CKINVDCx20_ASAP7_75t_R g1421 ( 
.A(n_1400),
.Y(n_1421)
);

NOR2xp33_ASAP7_75t_SL g1422 ( 
.A(n_1384),
.B(n_1315),
.Y(n_1422)
);

AND2x2_ASAP7_75t_L g1423 ( 
.A(n_1391),
.B(n_1366),
.Y(n_1423)
);

OR2x2_ASAP7_75t_L g1424 ( 
.A(n_1403),
.B(n_1360),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1403),
.B(n_1357),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1381),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1381),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1405),
.B(n_1357),
.Y(n_1428)
);

HB1xp67_ASAP7_75t_L g1429 ( 
.A(n_1414),
.Y(n_1429)
);

NAND2xp5_ASAP7_75t_L g1430 ( 
.A(n_1404),
.B(n_1333),
.Y(n_1430)
);

AND2x2_ASAP7_75t_L g1431 ( 
.A(n_1405),
.B(n_1360),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1401),
.B(n_1376),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1404),
.B(n_1332),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1405),
.B(n_1332),
.Y(n_1434)
);

OAI22xp5_ASAP7_75t_L g1435 ( 
.A1(n_1390),
.A2(n_1392),
.B1(n_1397),
.B2(n_1379),
.Y(n_1435)
);

NAND2x1p5_ASAP7_75t_L g1436 ( 
.A(n_1387),
.B(n_1346),
.Y(n_1436)
);

AND2x2_ASAP7_75t_L g1437 ( 
.A(n_1410),
.B(n_1323),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1401),
.A2(n_1331),
.B1(n_1356),
.B2(n_1315),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1386),
.A2(n_1356),
.B1(n_1315),
.B2(n_1362),
.Y(n_1439)
);

BUFx3_ASAP7_75t_L g1440 ( 
.A(n_1418),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1417),
.A2(n_1398),
.B(n_1382),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1426),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1429),
.Y(n_1443)
);

HB1xp67_ASAP7_75t_L g1444 ( 
.A(n_1429),
.Y(n_1444)
);

AND3x1_ASAP7_75t_L g1445 ( 
.A(n_1422),
.B(n_1392),
.C(n_1390),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1420),
.B(n_1402),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1426),
.Y(n_1447)
);

OAI31xp33_ASAP7_75t_L g1448 ( 
.A1(n_1435),
.A2(n_1384),
.A3(n_1385),
.B(n_1380),
.Y(n_1448)
);

NOR3xp33_ASAP7_75t_L g1449 ( 
.A(n_1435),
.B(n_1385),
.C(n_1389),
.Y(n_1449)
);

INVx1_ASAP7_75t_SL g1450 ( 
.A(n_1424),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1436),
.B(n_1377),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1437),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1416),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1418),
.Y(n_1454)
);

INVx2_ASAP7_75t_SL g1455 ( 
.A(n_1427),
.Y(n_1455)
);

BUFx2_ASAP7_75t_L g1456 ( 
.A(n_1418),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1437),
.B(n_1411),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1437),
.Y(n_1458)
);

BUFx3_ASAP7_75t_L g1459 ( 
.A(n_1436),
.Y(n_1459)
);

NOR2xp33_ASAP7_75t_L g1460 ( 
.A(n_1430),
.B(n_1406),
.Y(n_1460)
);

OAI33xp33_ASAP7_75t_L g1461 ( 
.A1(n_1430),
.A2(n_1399),
.A3(n_1349),
.B1(n_1353),
.B2(n_1367),
.B3(n_1351),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1454),
.B(n_1423),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1454),
.B(n_1423),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1453),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1455),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1440),
.Y(n_1466)
);

AND2x4_ASAP7_75t_L g1467 ( 
.A(n_1440),
.B(n_1425),
.Y(n_1467)
);

INVx2_ASAP7_75t_SL g1468 ( 
.A(n_1440),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1453),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1440),
.Y(n_1470)
);

INVx2_ASAP7_75t_L g1471 ( 
.A(n_1455),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1454),
.B(n_1423),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_1443),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1474)
);

AND2x2_ASAP7_75t_L g1475 ( 
.A(n_1454),
.B(n_1428),
.Y(n_1475)
);

NOR2xp33_ASAP7_75t_L g1476 ( 
.A(n_1460),
.B(n_1461),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1440),
.B(n_1425),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1478)
);

AND2x2_ASAP7_75t_L g1479 ( 
.A(n_1456),
.B(n_1428),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1443),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1442),
.Y(n_1481)
);

AND2x2_ASAP7_75t_L g1482 ( 
.A(n_1456),
.B(n_1431),
.Y(n_1482)
);

CKINVDCx16_ASAP7_75t_R g1483 ( 
.A(n_1456),
.Y(n_1483)
);

INVx8_ASAP7_75t_L g1484 ( 
.A(n_1451),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1444),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1444),
.B(n_1433),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1445),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1455),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1442),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1442),
.Y(n_1490)
);

NAND2xp5_ASAP7_75t_L g1491 ( 
.A(n_1458),
.B(n_1434),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1447),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1458),
.B(n_1434),
.Y(n_1493)
);

INVx1_ASAP7_75t_SL g1494 ( 
.A(n_1466),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1465),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1464),
.Y(n_1497)
);

INVxp67_ASAP7_75t_L g1498 ( 
.A(n_1487),
.Y(n_1498)
);

HB1xp67_ASAP7_75t_L g1499 ( 
.A(n_1462),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1466),
.Y(n_1500)
);

INVxp67_ASAP7_75t_L g1501 ( 
.A(n_1487),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1464),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1469),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1483),
.B(n_1450),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1476),
.B(n_1460),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1474),
.B(n_1458),
.Y(n_1506)
);

INVx2_ASAP7_75t_SL g1507 ( 
.A(n_1466),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1474),
.B(n_1450),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1475),
.B(n_1478),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1469),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1473),
.Y(n_1511)
);

OR2x2_ASAP7_75t_L g1512 ( 
.A(n_1474),
.B(n_1446),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1473),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1480),
.Y(n_1514)
);

OR2x2_ASAP7_75t_L g1515 ( 
.A(n_1486),
.B(n_1446),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1475),
.B(n_1457),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1480),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1485),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1465),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1475),
.B(n_1478),
.Y(n_1520)
);

INVxp67_ASAP7_75t_L g1521 ( 
.A(n_1476),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1478),
.B(n_1479),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1486),
.B(n_1419),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1485),
.B(n_1419),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1465),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1491),
.B(n_1446),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1490),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1490),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1462),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1466),
.B(n_1459),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1468),
.B(n_1470),
.Y(n_1531)
);

A2O1A1Ixp33_ASAP7_75t_L g1532 ( 
.A1(n_1479),
.A2(n_1448),
.B(n_1449),
.C(n_1422),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1479),
.B(n_1432),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1492),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1491),
.B(n_1493),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1481),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1521),
.B(n_1449),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1499),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1503),
.Y(n_1539)
);

OAI21xp33_ASAP7_75t_L g1540 ( 
.A1(n_1505),
.A2(n_1445),
.B(n_1449),
.Y(n_1540)
);

INVxp67_ASAP7_75t_SL g1541 ( 
.A(n_1498),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1503),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1533),
.B(n_1493),
.Y(n_1543)
);

NOR2xp33_ASAP7_75t_L g1544 ( 
.A(n_1501),
.B(n_1341),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1523),
.B(n_1462),
.Y(n_1545)
);

OAI322xp33_ASAP7_75t_L g1546 ( 
.A1(n_1494),
.A2(n_1468),
.A3(n_1482),
.B1(n_1463),
.B2(n_1472),
.C1(n_1470),
.C2(n_1415),
.Y(n_1546)
);

AOI31xp33_ASAP7_75t_L g1547 ( 
.A1(n_1532),
.A2(n_1445),
.A3(n_1341),
.B(n_1351),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1510),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1510),
.Y(n_1549)
);

NOR3xp33_ASAP7_75t_SL g1550 ( 
.A(n_1511),
.B(n_1394),
.C(n_1311),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1500),
.B(n_1388),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1496),
.B(n_1448),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1496),
.B(n_1467),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1524),
.B(n_1432),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1511),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1504),
.B(n_1467),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1497),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1500),
.Y(n_1559)
);

OR2x2_ASAP7_75t_L g1560 ( 
.A(n_1529),
.B(n_1463),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1507),
.B(n_1415),
.Y(n_1561)
);

INVx3_ASAP7_75t_L g1562 ( 
.A(n_1531),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1502),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1507),
.B(n_1395),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1513),
.Y(n_1565)
);

INVxp67_ASAP7_75t_L g1566 ( 
.A(n_1514),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1515),
.B(n_1463),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1515),
.B(n_1472),
.Y(n_1568)
);

AOI21xp5_ASAP7_75t_L g1569 ( 
.A1(n_1531),
.A2(n_1448),
.B(n_1461),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1517),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1509),
.B(n_1520),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1518),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1541),
.B(n_1509),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1537),
.B(n_1310),
.Y(n_1574)
);

NAND4xp25_ASAP7_75t_L g1575 ( 
.A(n_1540),
.B(n_1439),
.C(n_1470),
.D(n_1438),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_SL g1576 ( 
.A(n_1547),
.B(n_1467),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1553),
.B(n_1520),
.Y(n_1577)
);

NAND2xp5_ASAP7_75t_SL g1578 ( 
.A(n_1550),
.B(n_1467),
.Y(n_1578)
);

OAI21xp33_ASAP7_75t_L g1579 ( 
.A1(n_1552),
.A2(n_1522),
.B(n_1468),
.Y(n_1579)
);

NOR4xp25_ASAP7_75t_SL g1580 ( 
.A(n_1541),
.B(n_1394),
.C(n_1528),
.D(n_1527),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1538),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1551),
.B(n_1522),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1559),
.B(n_1531),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1544),
.B(n_1400),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1538),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1556),
.B(n_1477),
.Y(n_1586)
);

O2A1O1Ixp33_ASAP7_75t_L g1587 ( 
.A1(n_1552),
.A2(n_1470),
.B(n_1482),
.C(n_1530),
.Y(n_1587)
);

HB1xp67_ASAP7_75t_L g1588 ( 
.A(n_1559),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1544),
.Y(n_1589)
);

OAI22xp5_ASAP7_75t_L g1590 ( 
.A1(n_1569),
.A2(n_1439),
.B1(n_1477),
.B2(n_1470),
.Y(n_1590)
);

AOI22xp5_ASAP7_75t_L g1591 ( 
.A1(n_1551),
.A2(n_1477),
.B1(n_1530),
.B2(n_1461),
.Y(n_1591)
);

NOR2x2_ASAP7_75t_L g1592 ( 
.A(n_1550),
.B(n_1451),
.Y(n_1592)
);

OAI21xp5_ASAP7_75t_L g1593 ( 
.A1(n_1564),
.A2(n_1530),
.B(n_1477),
.Y(n_1593)
);

XNOR2x1_ASAP7_75t_L g1594 ( 
.A(n_1557),
.B(n_1335),
.Y(n_1594)
);

OAI21xp33_ASAP7_75t_SL g1595 ( 
.A1(n_1571),
.A2(n_1516),
.B(n_1482),
.Y(n_1595)
);

OAI211xp5_ASAP7_75t_L g1596 ( 
.A1(n_1566),
.A2(n_1441),
.B(n_1472),
.C(n_1484),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1539),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1542),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1545),
.B(n_1535),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1582),
.B(n_1554),
.Y(n_1601)
);

INVx1_ASAP7_75t_SL g1602 ( 
.A(n_1584),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1588),
.Y(n_1603)
);

INVx1_ASAP7_75t_SL g1604 ( 
.A(n_1594),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1573),
.B(n_1561),
.Y(n_1605)
);

AOI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1580),
.A2(n_1546),
.B(n_1558),
.Y(n_1606)
);

NOR2xp33_ASAP7_75t_L g1607 ( 
.A(n_1575),
.B(n_1395),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1583),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1591),
.A2(n_1560),
.B1(n_1568),
.B2(n_1567),
.Y(n_1609)
);

AOI22xp5_ASAP7_75t_L g1610 ( 
.A1(n_1590),
.A2(n_1477),
.B1(n_1572),
.B2(n_1565),
.Y(n_1610)
);

NOR4xp25_ASAP7_75t_SL g1611 ( 
.A(n_1576),
.B(n_1555),
.C(n_1549),
.D(n_1548),
.Y(n_1611)
);

INVxp67_ASAP7_75t_SL g1612 ( 
.A(n_1581),
.Y(n_1612)
);

OAI21xp5_ASAP7_75t_L g1613 ( 
.A1(n_1587),
.A2(n_1570),
.B(n_1563),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1562),
.Y(n_1614)
);

OAI21xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1578),
.A2(n_1562),
.B(n_1516),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1577),
.B(n_1562),
.Y(n_1616)
);

OAI22xp5_ASAP7_75t_L g1617 ( 
.A1(n_1580),
.A2(n_1543),
.B1(n_1484),
.B2(n_1459),
.Y(n_1617)
);

NOR2xp67_ASAP7_75t_L g1618 ( 
.A(n_1615),
.B(n_1608),
.Y(n_1618)
);

AOI222xp33_ASAP7_75t_L g1619 ( 
.A1(n_1602),
.A2(n_1579),
.B1(n_1596),
.B2(n_1593),
.C1(n_1598),
.C2(n_1597),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1583),
.Y(n_1620)
);

AOI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1609),
.A2(n_1574),
.B1(n_1595),
.B2(n_1586),
.Y(n_1621)
);

NAND2xp33_ASAP7_75t_SL g1622 ( 
.A(n_1611),
.B(n_1315),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_L g1623 ( 
.A1(n_1612),
.A2(n_1574),
.B(n_1599),
.C(n_1352),
.Y(n_1623)
);

NOR3xp33_ASAP7_75t_L g1624 ( 
.A(n_1600),
.B(n_1352),
.C(n_1335),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1612),
.B(n_1574),
.Y(n_1625)
);

INVx1_ASAP7_75t_L g1626 ( 
.A(n_1614),
.Y(n_1626)
);

XOR2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1610),
.B(n_1592),
.Y(n_1627)
);

NAND3xp33_ASAP7_75t_L g1628 ( 
.A(n_1622),
.B(n_1606),
.C(n_1613),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_SL g1629 ( 
.A(n_1619),
.B(n_1604),
.Y(n_1629)
);

NOR2xp33_ASAP7_75t_L g1630 ( 
.A(n_1625),
.B(n_1607),
.Y(n_1630)
);

NAND4xp25_ASAP7_75t_L g1631 ( 
.A(n_1618),
.B(n_1606),
.C(n_1605),
.D(n_1601),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1623),
.A2(n_1617),
.B(n_1616),
.Y(n_1632)
);

NAND4xp25_ASAP7_75t_L g1633 ( 
.A(n_1624),
.B(n_1408),
.C(n_1438),
.D(n_1324),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1620),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1626),
.B(n_1421),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1621),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_L g1637 ( 
.A1(n_1628),
.A2(n_1627),
.B(n_1484),
.C(n_1310),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1634),
.Y(n_1638)
);

OAI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1629),
.A2(n_1508),
.B(n_1535),
.Y(n_1639)
);

AOI221xp5_ASAP7_75t_L g1640 ( 
.A1(n_1631),
.A2(n_1536),
.B1(n_1495),
.B2(n_1525),
.C(n_1519),
.Y(n_1640)
);

AOI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1636),
.A2(n_1484),
.B1(n_1328),
.B2(n_1441),
.Y(n_1641)
);

OAI21xp5_ASAP7_75t_L g1642 ( 
.A1(n_1637),
.A2(n_1635),
.B(n_1632),
.Y(n_1642)
);

OAI21xp5_ASAP7_75t_SL g1643 ( 
.A1(n_1639),
.A2(n_1630),
.B(n_1633),
.Y(n_1643)
);

OAI22xp5_ASAP7_75t_L g1644 ( 
.A1(n_1641),
.A2(n_1638),
.B1(n_1640),
.B2(n_1508),
.Y(n_1644)
);

NOR2xp67_ASAP7_75t_L g1645 ( 
.A(n_1637),
.B(n_1534),
.Y(n_1645)
);

OAI321xp33_ASAP7_75t_L g1646 ( 
.A1(n_1637),
.A2(n_1451),
.A3(n_1512),
.B1(n_1526),
.B2(n_1362),
.C(n_1506),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1638),
.Y(n_1647)
);

NOR3xp33_ASAP7_75t_L g1648 ( 
.A(n_1642),
.B(n_1328),
.C(n_1374),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1647),
.Y(n_1649)
);

AO211x2_ASAP7_75t_L g1650 ( 
.A1(n_1643),
.A2(n_1536),
.B(n_1373),
.C(n_1484),
.Y(n_1650)
);

NAND4xp75_ASAP7_75t_L g1651 ( 
.A(n_1645),
.B(n_1495),
.C(n_1525),
.D(n_1519),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1644),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1648),
.A2(n_1646),
.B(n_1373),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1652),
.A2(n_1310),
.B(n_1506),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1649),
.Y(n_1655)
);

OA22x2_ASAP7_75t_L g1656 ( 
.A1(n_1655),
.A2(n_1650),
.B1(n_1651),
.B2(n_1471),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1656),
.Y(n_1657)
);

A2O1A1Ixp33_ASAP7_75t_L g1658 ( 
.A1(n_1657),
.A2(n_1654),
.B(n_1653),
.C(n_1471),
.Y(n_1658)
);

XNOR2xp5_ASAP7_75t_SL g1659 ( 
.A(n_1657),
.B(n_1310),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1659),
.A2(n_1526),
.B(n_1512),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1658),
.B(n_1378),
.Y(n_1661)
);

HB1xp67_ASAP7_75t_L g1662 ( 
.A(n_1661),
.Y(n_1662)
);

OAI21xp5_ASAP7_75t_L g1663 ( 
.A1(n_1660),
.A2(n_1465),
.B(n_1471),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1662),
.B(n_1471),
.Y(n_1664)
);

OAI22xp5_ASAP7_75t_L g1665 ( 
.A1(n_1664),
.A2(n_1663),
.B1(n_1488),
.B2(n_1310),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1665),
.A2(n_1488),
.B1(n_1489),
.B2(n_1481),
.Y(n_1666)
);

OAI221xp5_ASAP7_75t_R g1667 ( 
.A1(n_1666),
.A2(n_1484),
.B1(n_1407),
.B2(n_1413),
.C(n_1409),
.Y(n_1667)
);

AOI211xp5_ASAP7_75t_L g1668 ( 
.A1(n_1667),
.A2(n_1374),
.B(n_1383),
.C(n_1396),
.Y(n_1668)
);


endmodule