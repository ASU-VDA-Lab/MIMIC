module real_jpeg_30265_n_32 (n_17, n_8, n_0, n_21, n_212, n_2, n_29, n_10, n_31, n_9, n_12, n_24, n_218, n_215, n_6, n_221, n_28, n_216, n_213, n_23, n_11, n_14, n_211, n_25, n_217, n_7, n_22, n_18, n_3, n_210, n_5, n_4, n_219, n_1, n_26, n_27, n_20, n_19, n_222, n_30, n_220, n_16, n_15, n_214, n_13, n_32);

input n_17;
input n_8;
input n_0;
input n_21;
input n_212;
input n_2;
input n_29;
input n_10;
input n_31;
input n_9;
input n_12;
input n_24;
input n_218;
input n_215;
input n_6;
input n_221;
input n_28;
input n_216;
input n_213;
input n_23;
input n_11;
input n_14;
input n_211;
input n_25;
input n_217;
input n_7;
input n_22;
input n_18;
input n_3;
input n_210;
input n_5;
input n_4;
input n_219;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_222;
input n_30;
input n_220;
input n_16;
input n_15;
input n_214;
input n_13;

output n_32;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_131;
wire n_47;
wire n_163;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_172;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_148;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_150;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_185;
wire n_125;
wire n_55;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_53;
wire n_127;
wire n_206;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_0),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g164 ( 
.A1(n_0),
.A2(n_100),
.A3(n_102),
.B1(n_105),
.B2(n_165),
.C1(n_167),
.C2(n_220),
.Y(n_164)
);

AOI221xp5_ASAP7_75t_L g125 ( 
.A1(n_1),
.A2(n_31),
.B1(n_126),
.B2(n_131),
.C(n_135),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_1),
.B(n_126),
.C(n_131),
.Y(n_138)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_2),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g34 ( 
.A(n_3),
.B(n_35),
.C(n_192),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_3),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_3),
.B(n_37),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_3),
.A2(n_43),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_4),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_6),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g44 ( 
.A(n_7),
.B(n_45),
.C(n_186),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_8),
.B(n_114),
.Y(n_113)
);

HAxp5_ASAP7_75t_SL g161 ( 
.A(n_8),
.B(n_162),
.CON(n_161),
.SN(n_161)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_9),
.B(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_10),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_10),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_11),
.B(n_68),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_12),
.B(n_78),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_13),
.Y(n_187)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_15),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_16),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_16),
.A2(n_47),
.B1(n_49),
.B2(n_171),
.Y(n_170)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_17),
.Y(n_148)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_18),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_19),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_20),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g181 ( 
.A(n_20),
.B(n_89),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_21),
.B(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_21),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_22),
.B(n_77),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_23),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_23),
.B(n_107),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_24),
.Y(n_42)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_25),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_156),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_26),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_27),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_27),
.B(n_83),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_29),
.B(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_30),
.B(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_30),
.Y(n_168)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_31),
.Y(n_137)
);

XOR2x2_ASAP7_75t_SL g32 ( 
.A(n_33),
.B(n_203),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_SL g33 ( 
.A(n_34),
.B(n_43),
.C(n_194),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_43),
.B(n_44),
.C(n_191),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_42),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_39),
.B(n_157),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_41),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_91),
.B(n_170),
.Y(n_45)
);

NAND4xp25_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_56),
.C(n_81),
.D(n_87),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_55),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_51),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_51),
.B(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_53),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR3xp33_ASAP7_75t_SL g56 ( 
.A(n_57),
.B(n_66),
.C(n_69),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_58),
.B(n_180),
.C(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_65),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_59),
.B(n_65),
.Y(n_174)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_66),
.Y(n_173)
);

OAI322xp33_ASAP7_75t_L g178 ( 
.A1(n_66),
.A2(n_71),
.A3(n_179),
.B1(n_182),
.B2(n_183),
.C1(n_184),
.C2(n_222),
.Y(n_178)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_68),
.B(n_211),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_70),
.A2(n_173),
.A3(n_174),
.B1(n_175),
.B2(n_178),
.C(n_221),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_72),
.Y(n_183)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_75),
.Y(n_130)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_76),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_80),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_82),
.A2(n_172),
.B(n_185),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_90),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AOI31xp67_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_119),
.A3(n_154),
.B(n_159),
.Y(n_91)
);

NOR3xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_104),
.C(n_113),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_93),
.A2(n_160),
.B(n_164),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NOR3xp33_ASAP7_75t_L g165 ( 
.A(n_95),
.B(n_113),
.C(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_96),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_103),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

OA21x2_ASAP7_75t_SL g160 ( 
.A1(n_104),
.A2(n_161),
.B(n_163),
.Y(n_160)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_112),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_109),
.Y(n_107)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_114),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_117),
.Y(n_201)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_148),
.C(n_149),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_121),
.A2(n_139),
.B(n_147),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_125),
.B1(n_137),
.B2(n_138),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_127),
.B(n_136),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_131),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_216),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_146),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_146),
.Y(n_147)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_161),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_188),
.B(n_193),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_202),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_199),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_207),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_210),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_212),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_213),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_214),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_215),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_217),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_218),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_219),
.Y(n_157)
);


endmodule