module fake_jpeg_894_n_349 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx6_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_13),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_12),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_51),
.Y(n_113)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_52),
.Y(n_138)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_54),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_55),
.B(n_56),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_17),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_17),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_64),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g141 ( 
.A(n_58),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_59),
.Y(n_133)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_60),
.Y(n_107)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_27),
.B(n_0),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_62),
.B(n_91),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_31),
.Y(n_63)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_66),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_67),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_40),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_83),
.Y(n_152)
);

OR2x2_ASAP7_75t_SL g69 ( 
.A(n_24),
.B(n_0),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_69),
.B(n_71),
.Y(n_144)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_22),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_72),
.Y(n_123)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_73),
.Y(n_134)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_48),
.Y(n_75)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_75),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_76),
.Y(n_120)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_77),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g78 ( 
.A(n_28),
.Y(n_78)
);

CKINVDCx6p67_ASAP7_75t_R g149 ( 
.A(n_78),
.Y(n_149)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_80),
.Y(n_156)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_24),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_85),
.B(n_95),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_86),
.Y(n_131)
);

INVx6_ASAP7_75t_SL g87 ( 
.A(n_32),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_87),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_88),
.Y(n_132)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_90),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_18),
.B(n_1),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_92),
.Y(n_127)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_34),
.Y(n_93)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_18),
.B(n_1),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_94),
.B(n_96),
.Y(n_142)
);

INVx5_ASAP7_75t_L g95 ( 
.A(n_37),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_20),
.B(n_3),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_33),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_97),
.B(n_98),
.Y(n_151)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_36),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_20),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_100),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_36),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_44),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_21),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_23),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

CKINVDCx6p67_ASAP7_75t_R g168 ( 
.A(n_105),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_49),
.B1(n_47),
.B2(n_46),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_108),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_78),
.A2(n_21),
.B1(n_45),
.B2(n_41),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_53),
.A2(n_26),
.B1(n_45),
.B2(n_41),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_51),
.A2(n_23),
.B1(n_29),
.B2(n_26),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_79),
.A2(n_29),
.B1(n_47),
.B2(n_46),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_118),
.A2(n_119),
.B1(n_125),
.B2(n_130),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_49),
.B1(n_43),
.B2(n_42),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_74),
.A2(n_43),
.B1(n_42),
.B2(n_7),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_4),
.B1(n_5),
.B2(n_9),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_54),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_136),
.A2(n_139),
.B1(n_143),
.B2(n_146),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_50),
.A2(n_67),
.B1(n_65),
.B2(n_63),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_103),
.A2(n_5),
.B1(n_9),
.B2(n_11),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_58),
.A2(n_14),
.B1(n_15),
.B2(n_52),
.Y(n_146)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_92),
.A2(n_100),
.B1(n_66),
.B2(n_77),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_125),
.B1(n_111),
.B2(n_105),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_58),
.A2(n_84),
.B1(n_86),
.B2(n_88),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_158),
.A2(n_119),
.B1(n_106),
.B2(n_146),
.Y(n_190)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_145),
.Y(n_161)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_151),
.B(n_89),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_170),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_142),
.B(n_155),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_163),
.B(n_179),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_121),
.B(n_160),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_164),
.B(n_176),
.Y(n_208)
);

OR2x4_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_149),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_165),
.A2(n_132),
.B(n_162),
.Y(n_230)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_152),
.Y(n_167)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_167),
.Y(n_202)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_113),
.Y(n_169)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_169),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_129),
.B(n_148),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_171),
.Y(n_231)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_138),
.Y(n_174)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_175),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_149),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_109),
.Y(n_178)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_178),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_140),
.B(n_144),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_149),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_187),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_114),
.B(n_156),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_181),
.B(n_185),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_107),
.B(n_134),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_182),
.B(n_195),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_123),
.B(n_130),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_192),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_120),
.B(n_159),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g215 ( 
.A(n_184),
.B(n_191),
.Y(n_215)
);

CKINVDCx12_ASAP7_75t_R g185 ( 
.A(n_141),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_186),
.A2(n_104),
.B1(n_135),
.B2(n_143),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_106),
.B(n_133),
.Y(n_187)
);

INVx6_ASAP7_75t_L g188 ( 
.A(n_109),
.Y(n_188)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_188),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_118),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_194),
.Y(n_212)
);

OA22x2_ASAP7_75t_L g223 ( 
.A1(n_190),
.A2(n_122),
.B1(n_128),
.B2(n_131),
.Y(n_223)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_112),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_153),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_112),
.B(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_193),
.B(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_110),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_147),
.Y(n_195)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_116),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_198),
.Y(n_227)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_117),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_199),
.B(n_200),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_126),
.B(n_131),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_124),
.B(n_132),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_168),
.B1(n_165),
.B2(n_186),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_192),
.A2(n_183),
.B1(n_177),
.B2(n_189),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_210),
.B(n_173),
.Y(n_233)
);

OA21x2_ASAP7_75t_L g217 ( 
.A1(n_168),
.A2(n_158),
.B(n_124),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_223),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_180),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_221),
.B(n_226),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

INVx5_ASAP7_75t_L g225 ( 
.A(n_174),
.Y(n_225)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_225),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_184),
.Y(n_226)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_169),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_229),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_219),
.B(n_227),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_233),
.A2(n_242),
.B(n_244),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_168),
.B1(n_166),
.B2(n_193),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_234),
.A2(n_235),
.B1(n_223),
.B2(n_207),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_206),
.A2(n_168),
.B1(n_164),
.B2(n_170),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_236),
.B(n_245),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_213),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_238),
.B(n_250),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_182),
.C(n_184),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_239),
.B(n_241),
.Y(n_274)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_215),
.Y(n_240)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_240),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_204),
.B(n_161),
.C(n_175),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_215),
.Y(n_243)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_243),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_206),
.A2(n_196),
.B(n_198),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_191),
.B1(n_188),
.B2(n_178),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_246),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_204),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_247),
.B(n_249),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_202),
.B(n_231),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_248),
.B(n_252),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_216),
.A2(n_230),
.B1(n_217),
.B2(n_223),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_203),
.C(n_215),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_L g251 ( 
.A1(n_217),
.A2(n_222),
.B(n_220),
.C(n_228),
.Y(n_251)
);

AOI21xp33_ASAP7_75t_L g271 ( 
.A1(n_251),
.A2(n_232),
.B(n_214),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_205),
.Y(n_252)
);

INVx3_ASAP7_75t_SL g256 ( 
.A(n_205),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_207),
.B(n_225),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_257),
.B(n_229),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_246),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_255),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_266),
.B(n_270),
.Y(n_294)
);

O2A1O1Ixp33_ASAP7_75t_L g267 ( 
.A1(n_251),
.A2(n_254),
.B(n_233),
.C(n_234),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_269),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_228),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_242),
.A2(n_232),
.B(n_214),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_272),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_273),
.B(n_277),
.Y(n_289)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_276),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_236),
.B(n_218),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_244),
.A2(n_246),
.B(n_254),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_278),
.B(n_256),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_273),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_279),
.B(n_280),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_250),
.Y(n_280)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_278),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_282),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_285),
.A2(n_260),
.B1(n_258),
.B2(n_284),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_265),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_288),
.C(n_290),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_274),
.B(n_239),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_265),
.B(n_241),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_268),
.A2(n_249),
.B1(n_238),
.B2(n_243),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_261),
.B1(n_258),
.B2(n_263),
.Y(n_305)
);

MAJx2_ASAP7_75t_L g292 ( 
.A(n_268),
.B(n_240),
.C(n_245),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g308 ( 
.A(n_292),
.B(n_262),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_270),
.B(n_237),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_272),
.C(n_263),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_275),
.Y(n_295)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_295),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_296),
.A2(n_284),
.B(n_271),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_277),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_308),
.C(n_309),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_299),
.B(n_304),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_285),
.B1(n_289),
.B2(n_286),
.Y(n_311)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_294),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_305),
.A2(n_310),
.B1(n_289),
.B2(n_261),
.Y(n_314)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_283),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_306),
.B(n_307),
.Y(n_320)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

AO22x1_ASAP7_75t_SL g310 ( 
.A1(n_285),
.A2(n_291),
.B1(n_267),
.B2(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g328 ( 
.A1(n_311),
.A2(n_316),
.B1(n_319),
.B2(n_310),
.Y(n_328)
);

OA21x2_ASAP7_75t_SL g312 ( 
.A1(n_298),
.A2(n_300),
.B(n_259),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_312),
.B(n_313),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_299),
.A2(n_267),
.B(n_286),
.Y(n_313)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_314),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_303),
.A2(n_262),
.B(n_276),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_287),
.C(n_290),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_297),
.C(n_308),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_303),
.A2(n_293),
.B1(n_292),
.B2(n_259),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_317),
.B(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_321),
.B(n_322),
.Y(n_329)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_320),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_316),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_323),
.B(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_326),
.B(n_328),
.Y(n_333)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_319),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_325),
.A2(n_313),
.B(n_315),
.Y(n_330)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_330),
.A2(n_331),
.B(n_309),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_325),
.A2(n_315),
.B(n_318),
.Y(n_331)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_310),
.Y(n_332)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_332),
.A2(n_311),
.B(n_324),
.Y(n_335)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_335),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_334),
.A2(n_324),
.B1(n_333),
.B2(n_328),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_336),
.B(n_339),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g340 ( 
.A(n_337),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_329),
.A2(n_266),
.B1(n_264),
.B2(n_269),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_338),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_255),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_336),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_344),
.Y(n_346)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_338),
.A3(n_264),
.B1(n_255),
.B2(n_211),
.C1(n_218),
.C2(n_256),
.Y(n_345)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_346),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_347),
.A2(n_340),
.B(n_341),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_345),
.Y(n_349)
);


endmodule