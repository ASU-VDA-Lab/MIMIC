module fake_jpeg_4354_n_300 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_300);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_300;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_288;
wire n_272;
wire n_284;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_294;
wire n_299;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_155;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx10_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_2),
.B(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_11),
.B(n_1),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_13),
.B(n_7),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_41),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_40),
.Y(n_52)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_25),
.B1(n_20),
.B2(n_32),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_39),
.Y(n_59)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_24),
.B(n_0),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp33_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g62 ( 
.A1(n_43),
.A2(n_21),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_46),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_45),
.A2(n_19),
.B(n_20),
.Y(n_92)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx5_ASAP7_75t_SL g48 ( 
.A(n_42),
.Y(n_48)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_50),
.B(n_51),
.Y(n_75)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_53),
.B(n_55),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_57),
.A2(n_65),
.B1(n_32),
.B2(n_26),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_62),
.A2(n_43),
.B(n_33),
.C(n_21),
.Y(n_68)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_40),
.A2(n_25),
.B1(n_27),
.B2(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_28),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_66),
.Y(n_77)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_68),
.A2(n_41),
.B(n_36),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_48),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_89),
.Y(n_97)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_59),
.B(n_35),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_17),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_62),
.B(n_60),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_73),
.B(n_1),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_38),
.B1(n_35),
.B2(n_40),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_74),
.A2(n_85),
.B1(n_39),
.B2(n_22),
.Y(n_120)
);

BUFx4f_ASAP7_75t_SL g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_76),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_79),
.A2(n_54),
.B1(n_16),
.B2(n_3),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_41),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_88),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_40),
.B1(n_35),
.B2(n_26),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_84),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_49),
.A2(n_41),
.B1(n_35),
.B2(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_44),
.B(n_41),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_41),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_36),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_92),
.A2(n_36),
.B(n_23),
.Y(n_113)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_55),
.Y(n_108)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_100),
.Y(n_126)
);

AND2x6_ASAP7_75t_L g98 ( 
.A(n_73),
.B(n_88),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g150 ( 
.A(n_98),
.B(n_105),
.C(n_58),
.Y(n_150)
);

OAI221xp5_ASAP7_75t_L g100 ( 
.A1(n_77),
.A2(n_36),
.B1(n_41),
.B2(n_50),
.C(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_102),
.Y(n_127)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_75),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_103),
.B(n_104),
.Y(n_135)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_71),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_109),
.Y(n_140)
);

INVx1_ASAP7_75t_SL g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_SL g142 ( 
.A(n_107),
.Y(n_142)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_82),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_82),
.Y(n_110)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_111),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_77),
.A2(n_64),
.B1(n_61),
.B2(n_51),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

OAI21xp33_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_118),
.B(n_94),
.Y(n_138)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_114),
.B(n_70),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_115),
.B(n_116),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_83),
.B(n_67),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_117),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_119),
.B(n_85),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_120),
.A2(n_76),
.B1(n_69),
.B2(n_91),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_90),
.C(n_74),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_123),
.B(n_99),
.C(n_105),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_124),
.B(n_39),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g125 ( 
.A(n_109),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_129),
.Y(n_162)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_130),
.A2(n_133),
.B1(n_149),
.B2(n_89),
.Y(n_152)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_132),
.Y(n_167)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_120),
.A2(n_121),
.B1(n_104),
.B2(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_136),
.B(n_137),
.Y(n_170)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_141),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_68),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_92),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_145),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_147),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_113),
.A2(n_93),
.B1(n_72),
.B2(n_91),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_148),
.A2(n_96),
.B1(n_101),
.B2(n_103),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_121),
.A2(n_72),
.B1(n_93),
.B2(n_69),
.Y(n_149)
);

XNOR2x1_ASAP7_75t_SL g176 ( 
.A(n_150),
.B(n_39),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_151),
.A2(n_155),
.B1(n_177),
.B2(n_125),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_152),
.A2(n_159),
.B1(n_168),
.B2(n_169),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_174),
.C(n_175),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_131),
.A2(n_114),
.B1(n_107),
.B2(n_95),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_124),
.A2(n_95),
.B(n_17),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_156),
.B(n_164),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_157),
.B(n_129),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_135),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_172),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_123),
.A2(n_87),
.B1(n_78),
.B2(n_86),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_132),
.A2(n_19),
.B(n_78),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_160),
.A2(n_161),
.B(n_171),
.Y(n_200)
);

AOI21xp33_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_106),
.B(n_17),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_L g164 ( 
.A1(n_136),
.A2(n_17),
.B(n_87),
.Y(n_164)
);

OAI32xp33_ASAP7_75t_L g165 ( 
.A1(n_137),
.A2(n_17),
.A3(n_22),
.B1(n_31),
.B2(n_23),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_173),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_47),
.Y(n_166)
);

XNOR2x1_ASAP7_75t_L g201 ( 
.A(n_166),
.B(n_34),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_144),
.A2(n_86),
.B1(n_31),
.B2(n_30),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_126),
.A2(n_19),
.B(n_39),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_127),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_133),
.A2(n_39),
.B(n_1),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_145),
.B(n_148),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_134),
.B(n_39),
.C(n_81),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_34),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_144),
.A2(n_39),
.B(n_22),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_140),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_179),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

OA21x2_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_143),
.B(n_130),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_181),
.A2(n_30),
.B(n_23),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_182),
.B(n_183),
.C(n_191),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_157),
.B(n_174),
.Y(n_183)
);

XOR2x2_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_176),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_SL g219 ( 
.A(n_184),
.B(n_190),
.Y(n_219)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_158),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_185),
.B(n_188),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_125),
.Y(n_186)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_186),
.Y(n_208)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_162),
.Y(n_188)
);

A2O1A1O1Ixp25_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_142),
.B(n_128),
.C(n_39),
.D(n_23),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_159),
.C(n_170),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_180),
.B(n_139),
.C(n_142),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_202),
.C(n_171),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_180),
.B(n_39),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_201),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_155),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_195),
.B(n_205),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_197),
.A2(n_204),
.B1(n_163),
.B2(n_169),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_165),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_153),
.B(n_81),
.C(n_122),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_122),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g204 ( 
.A1(n_151),
.A2(n_82),
.B1(n_34),
.B2(n_31),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_175),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_184),
.A2(n_160),
.B(n_177),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_209),
.A2(n_185),
.B(n_30),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_213),
.Y(n_232)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_212),
.B(n_214),
.Y(n_243)
);

MAJx2_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_164),
.C(n_169),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_206),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_192),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_218),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_216),
.B(n_223),
.C(n_224),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_195),
.A2(n_179),
.B1(n_163),
.B2(n_173),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_217),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_181),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_220),
.A2(n_194),
.B1(n_190),
.B2(n_181),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_201),
.A2(n_34),
.B1(n_31),
.B2(n_30),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_221),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_189),
.B(n_182),
.C(n_191),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_189),
.B(n_81),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_225),
.A2(n_56),
.B(n_2),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_193),
.A2(n_200),
.B1(n_198),
.B2(n_196),
.Y(n_226)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_226),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_187),
.B(n_202),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_229),
.B(n_2),
.C(n_3),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_239),
.Y(n_248)
);

BUFx12_ASAP7_75t_L g231 ( 
.A(n_213),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_246),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_240),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_237),
.A2(n_241),
.B1(n_219),
.B2(n_8),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_216),
.C(n_207),
.Y(n_249)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_219),
.B(n_3),
.CI(n_4),
.CON(n_239),
.SN(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_4),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_210),
.B1(n_227),
.B2(n_208),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_244),
.A2(n_221),
.B1(n_211),
.B2(n_225),
.Y(n_250)
);

NAND2x1_ASAP7_75t_L g245 ( 
.A(n_209),
.B(n_5),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_245),
.B(n_226),
.Y(n_251)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_228),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_247),
.B(n_222),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_249),
.B(n_238),
.C(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_250),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_234),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_223),
.C(n_224),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_253),
.C(n_257),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_235),
.B(n_229),
.C(n_222),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_254),
.B(n_256),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_5),
.C(n_9),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_16),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_240),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_236),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_259),
.B(n_260),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_245),
.A2(n_15),
.B1(n_10),
.B2(n_12),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_269),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_261),
.A2(n_243),
.B(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_263),
.Y(n_279)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_248),
.A2(n_245),
.B(n_237),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_251),
.B(n_239),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_267),
.B(n_272),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_232),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_231),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_257),
.B(n_246),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_255),
.Y(n_277)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_274),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_270),
.B(n_255),
.Y(n_276)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_277),
.B(n_278),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_271),
.B(n_239),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_266),
.B(n_249),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_231),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_275),
.B(n_268),
.C(n_269),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_286),
.B(n_290),
.C(n_280),
.Y(n_292)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_267),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_287),
.A2(n_283),
.B(n_280),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_279),
.A2(n_268),
.B1(n_272),
.B2(n_264),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_293),
.B1(n_287),
.B2(n_12),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_294),
.C(n_295),
.Y(n_296)
);

OR2x2_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_9),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_286),
.B(n_14),
.C(n_10),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_289),
.B(n_285),
.C(n_284),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_297),
.B(n_12),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_298),
.B(n_14),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_299),
.A2(n_296),
.B(n_14),
.Y(n_300)
);


endmodule