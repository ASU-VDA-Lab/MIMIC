module fake_jpeg_12809_n_565 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_565);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_565;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_7),
.B(n_4),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_5),
.B(n_0),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_16),
.Y(n_53)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_36),
.Y(n_54)
);

INVx1_ASAP7_75t_SL g168 ( 
.A(n_54),
.Y(n_168)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_56),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_57),
.Y(n_143)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_58),
.Y(n_125)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_59),
.Y(n_116)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_52),
.Y(n_60)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_61),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_48),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_62),
.B(n_53),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_63),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_64),
.Y(n_124)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g109 ( 
.A(n_65),
.Y(n_109)
);

BUFx12_ASAP7_75t_L g66 ( 
.A(n_20),
.Y(n_66)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_66),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_67),
.Y(n_130)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_68),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_69),
.B(n_77),
.Y(n_117)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g140 ( 
.A(n_70),
.Y(n_140)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_71),
.Y(n_134)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_25),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_75),
.Y(n_148)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_76),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_43),
.B(n_10),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_78),
.Y(n_136)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_52),
.Y(n_79)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_79),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_80),
.Y(n_151)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_20),
.Y(n_81)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_81),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_82),
.Y(n_158)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_83),
.Y(n_138)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_84),
.Y(n_162)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_85),
.Y(n_144)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_46),
.Y(n_86)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_86),
.Y(n_146)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_22),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_87),
.Y(n_172)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_88),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_89),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_90),
.Y(n_167)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_92),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_93),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_20),
.Y(n_95)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_96),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_97),
.Y(n_161)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_22),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_98),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_99),
.B(n_106),
.Y(n_170)
);

BUFx24_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_103),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_102),
.B(n_105),
.Y(n_113)
);

BUFx24_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_104),
.Y(n_166)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_44),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_44),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_44),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_40),
.B(n_10),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_48),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_114),
.B(n_132),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_127),
.B(n_33),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_63),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_76),
.A2(n_42),
.B1(n_51),
.B2(n_47),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_141),
.A2(n_149),
.B1(n_152),
.B2(n_155),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_84),
.B1(n_64),
.B2(n_73),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_76),
.A2(n_103),
.B1(n_100),
.B2(n_65),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_62),
.B(n_23),
.C(n_45),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_153),
.B(n_31),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_154),
.B(n_159),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_70),
.A2(n_42),
.B1(n_51),
.B2(n_47),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_92),
.B(n_53),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_156),
.B(n_165),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_80),
.A2(n_42),
.B1(n_106),
.B2(n_104),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_86),
.B(n_32),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_67),
.A2(n_51),
.B1(n_44),
.B2(n_47),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_L g163 ( 
.A1(n_74),
.A2(n_47),
.B1(n_38),
.B2(n_34),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_107),
.A2(n_30),
.B1(n_41),
.B2(n_32),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_72),
.B(n_30),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g173 ( 
.A1(n_149),
.A2(n_75),
.B1(n_94),
.B2(n_90),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_173),
.Y(n_270)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_123),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_174),
.Y(n_276)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_151),
.Y(n_175)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_175),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_113),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_176),
.B(n_195),
.Y(n_251)
);

INVx11_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g278 ( 
.A(n_177),
.Y(n_278)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_110),
.Y(n_178)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_178),
.Y(n_237)
);

AO22x1_ASAP7_75t_L g179 ( 
.A1(n_163),
.A2(n_19),
.B1(n_21),
.B2(n_29),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_179),
.A2(n_203),
.B(n_231),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_23),
.B1(n_39),
.B2(n_45),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g260 ( 
.A(n_180),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_181),
.B(n_190),
.Y(n_241)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_161),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g253 ( 
.A(n_182),
.Y(n_253)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_116),
.Y(n_183)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_183),
.Y(n_269)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_184),
.Y(n_283)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_134),
.Y(n_185)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g186 ( 
.A1(n_155),
.A2(n_101),
.B1(n_82),
.B2(n_88),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_186),
.A2(n_210),
.B1(n_227),
.B2(n_120),
.Y(n_240)
);

OA22x2_ASAP7_75t_L g188 ( 
.A1(n_160),
.A2(n_34),
.B1(n_26),
.B2(n_38),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_188),
.B(n_192),
.Y(n_245)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_117),
.B(n_41),
.Y(n_190)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_191),
.Y(n_261)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_193),
.Y(n_263)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_150),
.B(n_39),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g277 ( 
.A1(n_194),
.A2(n_229),
.B(n_12),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_113),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_150),
.A2(n_26),
.B1(n_29),
.B2(n_19),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_196),
.B(n_217),
.Y(n_254)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_197),
.Y(n_264)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_142),
.Y(n_198)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_198),
.Y(n_266)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_199),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_145),
.Y(n_200)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_201),
.Y(n_273)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_119),
.Y(n_202)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_202),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_170),
.A2(n_99),
.B1(n_86),
.B2(n_24),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_204),
.Y(n_282)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_119),
.Y(n_205)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_205),
.Y(n_285)
);

BUFx12f_ASAP7_75t_L g206 ( 
.A(n_143),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_206),
.B(n_207),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_152),
.Y(n_207)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_161),
.Y(n_209)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_209),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_141),
.A2(n_27),
.B1(n_31),
.B2(n_19),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_170),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_211),
.B(n_221),
.Y(n_247)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_171),
.Y(n_212)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_212),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_111),
.Y(n_213)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_213),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_111),
.Y(n_214)
);

NAND2xp33_ASAP7_75t_SL g281 ( 
.A(n_214),
.B(n_216),
.Y(n_281)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_115),
.Y(n_215)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_215),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_168),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_115),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_133),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_218),
.B(n_220),
.Y(n_275)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_133),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_138),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_224),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_125),
.A2(n_21),
.B1(n_169),
.B2(n_128),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_225),
.A2(n_139),
.B1(n_167),
.B2(n_158),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_144),
.B(n_27),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_226),
.B(n_232),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_120),
.A2(n_21),
.B1(n_33),
.B2(n_89),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_146),
.B(n_33),
.Y(n_228)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_228),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g229 ( 
.A(n_118),
.B(n_0),
.Y(n_229)
);

INVx5_ASAP7_75t_L g230 ( 
.A(n_118),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_230),
.Y(n_279)
);

OA22x2_ASAP7_75t_SL g231 ( 
.A1(n_140),
.A2(n_54),
.B1(n_81),
.B2(n_66),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_112),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_129),
.B(n_33),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_233),
.B(n_171),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_130),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_234),
.B(n_33),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g295 ( 
.A(n_236),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_121),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_238),
.B(n_274),
.C(n_8),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_207),
.A2(n_0),
.B(n_1),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_239),
.A2(n_0),
.B(n_1),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_240),
.B(n_257),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_208),
.A2(n_187),
.B1(n_186),
.B2(n_192),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g320 ( 
.A1(n_242),
.A2(n_248),
.B1(n_259),
.B2(n_265),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_179),
.A2(n_122),
.B1(n_135),
.B2(n_124),
.Y(n_243)
);

AO21x2_ASAP7_75t_L g326 ( 
.A1(n_243),
.A2(n_7),
.B(n_17),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_192),
.A2(n_173),
.B1(n_229),
.B2(n_188),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_188),
.A2(n_196),
.B1(n_231),
.B2(n_203),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_249),
.A2(n_250),
.B1(n_231),
.B2(n_182),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_173),
.A2(n_162),
.B1(n_112),
.B2(n_122),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_173),
.A2(n_162),
.B1(n_147),
.B2(n_124),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_229),
.A2(n_147),
.B1(n_135),
.B2(n_148),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_226),
.B(n_148),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_268),
.B(n_178),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_188),
.A2(n_167),
.B1(n_158),
.B2(n_151),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g335 ( 
.A1(n_271),
.A2(n_14),
.B1(n_17),
.B2(n_16),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_194),
.B(n_199),
.Y(n_274)
);

XNOR2x1_ASAP7_75t_L g290 ( 
.A(n_277),
.B(n_196),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_284),
.Y(n_298)
);

XNOR2x1_ASAP7_75t_L g353 ( 
.A(n_290),
.B(n_315),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_291),
.A2(n_300),
.B1(n_323),
.B2(n_326),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_241),
.B(n_222),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g366 ( 
.A(n_292),
.B(n_296),
.Y(n_366)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_293),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_242),
.A2(n_232),
.B1(n_223),
.B2(n_196),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_294),
.A2(n_299),
.B1(n_335),
.B2(n_250),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_238),
.B(n_213),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_247),
.B(n_234),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_297),
.B(n_303),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_248),
.A2(n_175),
.B1(n_193),
.B2(n_198),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_183),
.B1(n_184),
.B2(n_189),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_270),
.A2(n_191),
.B1(n_209),
.B2(n_206),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_301),
.Y(n_359)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_302),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_235),
.B(n_255),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_275),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_304),
.B(n_305),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_236),
.B(n_200),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_306),
.B(n_308),
.Y(n_350)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_273),
.Y(n_307)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_307),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_235),
.B(n_202),
.Y(n_308)
);

INVx3_ASAP7_75t_L g309 ( 
.A(n_256),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g369 ( 
.A(n_309),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_251),
.B(n_230),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_310),
.Y(n_358)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_273),
.Y(n_311)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_311),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_268),
.B(n_221),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_312),
.B(n_314),
.Y(n_360)
);

O2A1O1Ixp33_ASAP7_75t_L g313 ( 
.A1(n_254),
.A2(n_177),
.B(n_205),
.C(n_212),
.Y(n_313)
);

AO21x1_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_319),
.B(n_278),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_275),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_274),
.B(n_206),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_263),
.Y(n_316)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_316),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_282),
.B(n_96),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_317),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_254),
.B(n_0),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_318),
.B(n_324),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_96),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_321),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_256),
.Y(n_322)
);

INVx3_ASAP7_75t_L g348 ( 
.A(n_322),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_245),
.A2(n_89),
.B1(n_11),
.B2(n_12),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_254),
.B(n_1),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_327),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_245),
.B(n_284),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_245),
.B(n_1),
.C(n_2),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_331),
.C(n_281),
.Y(n_355)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_329),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_252),
.B(n_13),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_289),
.B(n_13),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_332),
.B(n_339),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_276),
.B(n_14),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_333),
.A2(n_295),
.B1(n_298),
.B2(n_332),
.Y(n_380)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_244),
.Y(n_334)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_337),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_6),
.Y(n_338)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_258),
.B(n_2),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_341),
.A2(n_342),
.B1(n_347),
.B2(n_373),
.Y(n_390)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_299),
.A2(n_286),
.B1(n_260),
.B2(n_253),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_295),
.A2(n_262),
.B(n_239),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g409 ( 
.A1(n_343),
.A2(n_362),
.B(n_319),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_320),
.A2(n_271),
.B1(n_240),
.B2(n_252),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g352 ( 
.A1(n_291),
.A2(n_259),
.B1(n_265),
.B2(n_286),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_352),
.A2(n_365),
.B1(n_371),
.B2(n_313),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_355),
.B(n_380),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_362),
.Y(n_385)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_322),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g365 ( 
.A1(n_320),
.A2(n_289),
.B1(n_244),
.B2(n_258),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_315),
.B(n_275),
.C(n_267),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_368),
.B(n_372),
.C(n_331),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_298),
.A2(n_279),
.B1(n_278),
.B2(n_267),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_325),
.B(n_246),
.C(n_287),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_330),
.A2(n_279),
.B1(n_287),
.B2(n_285),
.Y(n_373)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_293),
.Y(n_378)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_378),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g379 ( 
.A1(n_330),
.A2(n_285),
.B1(n_246),
.B2(n_272),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_379),
.A2(n_382),
.B1(n_300),
.B2(n_316),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_330),
.A2(n_272),
.B1(n_280),
.B2(n_283),
.Y(n_382)
);

XNOR2x1_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_368),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_374),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_388),
.C(n_393),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_387),
.A2(n_397),
.B1(n_399),
.B2(n_418),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_353),
.B(n_327),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g426 ( 
.A1(n_389),
.A2(n_412),
.B1(n_352),
.B2(n_341),
.Y(n_426)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_344),
.Y(n_392)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_392),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_370),
.B(n_360),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_350),
.B(n_306),
.Y(n_394)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_395),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_343),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_396),
.B(n_398),
.Y(n_427)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_365),
.A2(n_294),
.B1(n_335),
.B2(n_312),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_371),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g399 ( 
.A1(n_376),
.A2(n_324),
.B1(n_318),
.B2(n_314),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g400 ( 
.A(n_366),
.B(n_311),
.C(n_307),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_400),
.B(n_407),
.Y(n_435)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_344),
.Y(n_401)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_401),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_304),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_402),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_SL g403 ( 
.A(n_340),
.B(n_302),
.Y(n_403)
);

CKINVDCx14_ASAP7_75t_R g421 ( 
.A(n_403),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_290),
.C(n_334),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_414),
.C(n_415),
.Y(n_422)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_345),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_405),
.B(n_406),
.Y(n_442)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_345),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_360),
.Y(n_407)
);

INVxp33_ASAP7_75t_SL g408 ( 
.A(n_354),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_408),
.B(n_417),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_409),
.A2(n_283),
.B(n_269),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_358),
.B(n_339),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_410),
.B(n_411),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_350),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g412 ( 
.A1(n_347),
.A2(n_326),
.B1(n_323),
.B2(n_328),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_381),
.B(n_280),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_416),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_372),
.B(n_329),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_336),
.Y(n_415)
);

NAND3xp33_ASAP7_75t_L g416 ( 
.A(n_377),
.B(n_261),
.C(n_288),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_346),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_359),
.A2(n_309),
.B1(n_337),
.B2(n_326),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_356),
.B(n_326),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_419),
.B(n_349),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_355),
.C(n_374),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_448),
.C(n_422),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_425),
.B(n_404),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_426),
.A2(n_431),
.B1(n_432),
.B2(n_439),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_397),
.A2(n_398),
.B1(n_385),
.B2(n_387),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_430),
.A2(n_437),
.B1(n_447),
.B2(n_449),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_390),
.A2(n_359),
.B1(n_377),
.B2(n_378),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_385),
.A2(n_346),
.B1(n_349),
.B2(n_361),
.Y(n_432)
);

AOI22x1_ASAP7_75t_L g433 ( 
.A1(n_396),
.A2(n_382),
.B1(n_379),
.B2(n_361),
.Y(n_433)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_433),
.Y(n_455)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_434),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_399),
.A2(n_326),
.B1(n_357),
.B2(n_351),
.Y(n_437)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_412),
.A2(n_367),
.B1(n_357),
.B2(n_351),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_393),
.B(n_367),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_420),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g445 ( 
.A(n_402),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_445),
.B(n_391),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_419),
.A2(n_375),
.B1(n_363),
.B2(n_348),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_384),
.B(n_375),
.C(n_363),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_409),
.A2(n_348),
.B1(n_364),
.B2(n_369),
.Y(n_449)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_402),
.A2(n_369),
.B1(n_261),
.B2(n_288),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g477 ( 
.A1(n_450),
.A2(n_432),
.B1(n_440),
.B2(n_426),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g473 ( 
.A1(n_451),
.A2(n_418),
.B(n_269),
.Y(n_473)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_452),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_442),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_460),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_458),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_SL g486 ( 
.A(n_457),
.B(n_465),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_420),
.B(n_386),
.C(n_415),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_459),
.B(n_462),
.C(n_469),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_424),
.B(n_383),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_442),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_467),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_422),
.B(n_388),
.C(n_394),
.Y(n_462)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_444),
.Y(n_464)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_SL g465 ( 
.A(n_425),
.B(n_389),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_423),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_466),
.B(n_433),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_435),
.B(n_401),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_444),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_468),
.B(n_475),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_448),
.B(n_417),
.C(n_406),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_439),
.B(n_405),
.C(n_392),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_470),
.B(n_478),
.C(n_440),
.Y(n_487)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_429),
.Y(n_471)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_471),
.Y(n_485)
);

AOI21xp5_ASAP7_75t_L g500 ( 
.A1(n_473),
.A2(n_474),
.B(n_429),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g474 ( 
.A1(n_427),
.A2(n_237),
.B(n_15),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_424),
.B(n_237),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_428),
.B(n_6),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_476),
.B(n_421),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_477),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_447),
.B(n_2),
.C(n_3),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_430),
.B(n_6),
.Y(n_479)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_450),
.Y(n_491)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_463),
.A2(n_427),
.B(n_438),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_480),
.B(n_489),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_487),
.B(n_491),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_456),
.B(n_438),
.C(n_451),
.Y(n_489)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_463),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_466),
.B(n_446),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_493),
.B(n_495),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_462),
.B(n_436),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_496),
.B(n_497),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_459),
.B(n_433),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_498),
.B(n_481),
.Y(n_510)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_458),
.B(n_431),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_465),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g518 ( 
.A1(n_500),
.A2(n_471),
.B1(n_478),
.B2(n_474),
.Y(n_518)
);

O2A1O1Ixp33_ASAP7_75t_L g502 ( 
.A1(n_455),
.A2(n_434),
.B(n_443),
.C(n_437),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_502),
.A2(n_473),
.B1(n_449),
.B2(n_443),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_L g503 ( 
.A1(n_483),
.A2(n_453),
.B1(n_455),
.B2(n_454),
.Y(n_503)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_503),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_469),
.C(n_457),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_505),
.B(n_508),
.Y(n_524)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_507),
.B(n_520),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_484),
.B(n_470),
.C(n_472),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_494),
.B(n_472),
.C(n_477),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_509),
.B(n_511),
.C(n_512),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_SL g526 ( 
.A(n_510),
.B(n_516),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_494),
.B(n_453),
.C(n_464),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_499),
.B(n_461),
.C(n_468),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_513),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_497),
.C(n_489),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_515),
.B(n_487),
.C(n_501),
.Y(n_528)
);

CKINVDCx20_ASAP7_75t_R g516 ( 
.A(n_488),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g531 ( 
.A1(n_518),
.A2(n_502),
.B1(n_491),
.B2(n_482),
.Y(n_531)
);

AOI21x1_ASAP7_75t_L g520 ( 
.A1(n_480),
.A2(n_446),
.B(n_479),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_508),
.B(n_495),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_522),
.B(n_525),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_517),
.B(n_490),
.Y(n_523)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_523),
.Y(n_537)
);

OAI21xp5_ASAP7_75t_SL g525 ( 
.A1(n_514),
.A2(n_492),
.B(n_500),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_528),
.B(n_529),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_517),
.B(n_490),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_531),
.B(n_535),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_512),
.B(n_485),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_532),
.B(n_533),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_511),
.B(n_486),
.Y(n_533)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_509),
.A2(n_486),
.B1(n_16),
.B2(n_5),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_534),
.B(n_18),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_527),
.B(n_515),
.C(n_505),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_540),
.Y(n_548)
);

A2O1A1Ixp33_ASAP7_75t_L g538 ( 
.A1(n_525),
.A2(n_513),
.B(n_519),
.C(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_538),
.Y(n_551)
);

OAI21xp5_ASAP7_75t_SL g540 ( 
.A1(n_524),
.A2(n_504),
.B(n_506),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_535),
.Y(n_552)
);

MAJIxp5_ASAP7_75t_L g545 ( 
.A(n_527),
.B(n_504),
.C(n_506),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_545),
.B(n_546),
.Y(n_547)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_528),
.B(n_521),
.C(n_507),
.Y(n_546)
);

OAI21xp5_ASAP7_75t_L g549 ( 
.A1(n_541),
.A2(n_529),
.B(n_523),
.Y(n_549)
);

AOI21xp5_ASAP7_75t_L g555 ( 
.A1(n_549),
.A2(n_550),
.B(n_553),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g550 ( 
.A1(n_536),
.A2(n_534),
.B(n_531),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g556 ( 
.A(n_552),
.B(n_546),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_543),
.B(n_526),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_SL g554 ( 
.A1(n_548),
.A2(n_547),
.B(n_551),
.Y(n_554)
);

AOI21xp5_ASAP7_75t_L g559 ( 
.A1(n_554),
.A2(n_557),
.B(n_555),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g558 ( 
.A(n_556),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_SL g557 ( 
.A1(n_549),
.A2(n_542),
.B(n_545),
.Y(n_557)
);

NAND4xp25_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_537),
.C(n_539),
.D(n_538),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_560),
.B(n_561),
.C(n_530),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_530),
.Y(n_561)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_562),
.B(n_18),
.C(n_3),
.Y(n_563)
);

AOI21xp5_ASAP7_75t_L g564 ( 
.A1(n_563),
.A2(n_2),
.B(n_3),
.Y(n_564)
);

NOR3xp33_ASAP7_75t_SL g565 ( 
.A(n_564),
.B(n_3),
.C(n_4),
.Y(n_565)
);


endmodule