module real_jpeg_4111_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_516;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_470;
wire n_219;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_0),
.B(n_43),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_0),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_0),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_0),
.B(n_300),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_0),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_0),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_0),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_1),
.B(n_206),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_1),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_1),
.B(n_55),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_1),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_1),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_1),
.B(n_419),
.Y(n_418)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_2),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_2),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g321 ( 
.A(n_2),
.Y(n_321)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_2),
.Y(n_328)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_2),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_3),
.B(n_58),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_3),
.B(n_36),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_114),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_3),
.B(n_187),
.Y(n_186)
);

AND2x2_ASAP7_75t_SL g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_3),
.B(n_321),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_3),
.B(n_424),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_4),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_4),
.B(n_43),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_4),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_4),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_4),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_4),
.B(n_355),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_4),
.B(n_277),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_4),
.B(n_416),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_5),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_5),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_5),
.Y(n_208)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_5),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_6),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_6),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_6),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_6),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_6),
.B(n_124),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_6),
.B(n_201),
.Y(n_200)
);

AND2x2_ASAP7_75t_SL g221 ( 
.A(n_6),
.B(n_222),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_7),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_7),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_7),
.B(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_7),
.B(n_133),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_7),
.B(n_70),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_7),
.B(n_277),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_7),
.B(n_300),
.Y(n_299)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_7),
.B(n_266),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_8),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g102 ( 
.A(n_9),
.Y(n_102)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_9),
.Y(n_154)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_9),
.Y(n_185)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_10),
.Y(n_515)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_11),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g294 ( 
.A(n_11),
.Y(n_294)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_12),
.Y(n_73)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_13),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g220 ( 
.A(n_13),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_13),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_14),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_14),
.B(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_14),
.B(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_14),
.B(n_320),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g335 ( 
.A(n_14),
.B(n_336),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_14),
.B(n_65),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_14),
.B(n_386),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_14),
.B(n_413),
.Y(n_412)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_16),
.B(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_16),
.B(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_16),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_16),
.B(n_345),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_16),
.B(n_114),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_16),
.B(n_390),
.Y(n_389)
);

AND2x4_ASAP7_75t_SL g405 ( 
.A(n_16),
.B(n_406),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_17),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_17),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g82 ( 
.A(n_17),
.B(n_83),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_17),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_17),
.B(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_17),
.B(n_148),
.Y(n_147)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_19),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_19),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_19),
.B(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_19),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_19),
.B(n_264),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_513),
.B(n_516),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_167),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_166),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_105),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_25),
.B(n_105),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_85),
.B1(n_86),
.B2(n_104),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_26),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_56),
.C(n_74),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_27),
.A2(n_28),
.B1(n_163),
.B2(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_39),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_34),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_30),
.B(n_34),
.C(n_39),
.Y(n_103)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g133 ( 
.A(n_37),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_37),
.Y(n_227)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_38),
.Y(n_98)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_38),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_38),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_44),
.C(n_51),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_40),
.B(n_142),
.Y(n_141)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_44),
.A2(n_45),
.B1(n_51),
.B2(n_52),
.Y(n_142)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_48),
.Y(n_392)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g414 ( 
.A(n_50),
.Y(n_414)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_56),
.A2(n_74),
.B1(n_75),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_56),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_61),
.C(n_68),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_SL g158 ( 
.A(n_57),
.B(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_62),
.B1(n_135),
.B2(n_140),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_61),
.A2(n_62),
.B1(n_68),
.B2(n_69),
.Y(n_159)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_62),
.B(n_132),
.C(n_135),
.Y(n_160)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_66),
.Y(n_324)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_67),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_69),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_69),
.B(n_81),
.C(n_84),
.Y(n_92)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_72),
.Y(n_190)
);

INVx6_ASAP7_75t_L g361 ( 
.A(n_72),
.Y(n_361)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_73),
.Y(n_298)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_73),
.Y(n_387)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_79),
.B1(n_80),
.B2(n_84),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_81),
.A2(n_82),
.B1(n_95),
.B2(n_96),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_SL g86 ( 
.A(n_87),
.B(n_103),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_99),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_98),
.Y(n_390)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx3_ASAP7_75t_SL g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_102),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_157),
.C(n_162),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_106),
.A2(n_107),
.B1(n_498),
.B2(n_499),
.Y(n_497)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_141),
.C(n_143),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_108),
.B(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_118),
.C(n_131),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_109),
.A2(n_110),
.B1(n_118),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_111),
.B(n_113),
.C(n_115),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_114),
.Y(n_281)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_118),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_128),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_119),
.B(n_128),
.Y(n_240)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_123),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx8_ASAP7_75t_L g224 ( 
.A(n_126),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_127),
.Y(n_301)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_131),
.B(n_230),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_135),
.B(n_146),
.C(n_150),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_135),
.A2(n_140),
.B1(n_146),
.B2(n_147),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_139),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g502 ( 
.A(n_141),
.B(n_143),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_155),
.C(n_156),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_144),
.A2(n_145),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_147),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_146),
.B(n_200),
.C(n_238),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_149),
.Y(n_222)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_149),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_150),
.B(n_236),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_152),
.Y(n_150)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_154),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_155),
.A2(n_205),
.B1(n_209),
.B2(n_210),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_155),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_155),
.A2(n_156),
.B1(n_210),
.B2(n_246),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_155),
.B(n_209),
.C(n_248),
.Y(n_247)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_156),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g498 ( 
.A(n_157),
.B(n_162),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_161),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g503 ( 
.A(n_158),
.B(n_504),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_L g504 ( 
.A(n_160),
.B(n_161),
.Y(n_504)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_163),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_495),
.B(n_510),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_303),
.B(n_494),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_249),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_171),
.B(n_249),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_228),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g509 ( 
.A(n_172),
.B(n_229),
.C(n_232),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_203),
.C(n_212),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_173),
.B(n_252),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_181),
.C(n_193),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_174),
.B(n_480),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

INVx4_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_181),
.A2(n_182),
.B1(n_193),
.B2(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.C(n_191),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_183),
.B(n_191),
.Y(n_470)
);

INVx6_ASAP7_75t_L g407 ( 
.A(n_184),
.Y(n_407)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_186),
.B(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx5_ASAP7_75t_L g345 ( 
.A(n_190),
.Y(n_345)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_190),
.Y(n_419)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_193),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_194),
.Y(n_238)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_202),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_203),
.B(n_212),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_211),
.Y(n_203)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_205),
.Y(n_209)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_211),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_223),
.C(n_225),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_213),
.B(n_284),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.C(n_221),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_214),
.B(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_216),
.B(n_221),
.Y(n_261)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx5_ASAP7_75t_L g336 ( 
.A(n_220),
.Y(n_336)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_220),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_223),
.B(n_225),
.Y(n_284)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_232),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_241),
.B2(n_242),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_233),
.B(n_243),
.C(n_247),
.Y(n_505)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_235),
.B(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_239),
.Y(n_255)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_247),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.C(n_256),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_251),
.B(n_254),
.Y(n_490)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_256),
.B(n_490),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_282),
.C(n_285),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g482 ( 
.A(n_258),
.B(n_483),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_262),
.C(n_271),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_259),
.A2(n_260),
.B1(n_461),
.B2(n_462),
.Y(n_460)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g448 ( 
.A1(n_262),
.A2(n_263),
.B(n_267),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_262),
.B(n_271),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_267),
.Y(n_262)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx4_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

MAJx2_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.C(n_279),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g438 ( 
.A1(n_272),
.A2(n_273),
.B1(n_275),
.B2(n_276),
.Y(n_438)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_279),
.B(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_280),
.B(n_301),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_282),
.A2(n_283),
.B1(n_285),
.B2(n_484),
.Y(n_483)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_285),
.Y(n_484)
);

MAJx2_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_299),
.C(n_302),
.Y(n_285)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_287),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.C(n_295),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_288),
.B(n_450),
.Y(n_449)
);

INVx6_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g450 ( 
.A1(n_291),
.A2(n_295),
.B1(n_296),
.B2(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_SL g451 ( 
.A(n_291),
.Y(n_451)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx3_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_299),
.B(n_302),
.Y(n_472)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21x1_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_488),
.B(n_493),
.Y(n_303)
);

OAI21x1_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_475),
.B(n_487),
.Y(n_304)
);

AOI21x1_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_457),
.B(n_474),
.Y(n_305)
);

OAI21x1_ASAP7_75t_L g306 ( 
.A1(n_307),
.A2(n_431),
.B(n_456),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_396),
.B(n_430),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_367),
.B(n_395),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_347),
.B(n_366),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_311),
.A2(n_330),
.B(n_346),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_325),
.B(n_329),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_322),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_319),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_319),
.Y(n_331)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx5_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_318),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_331),
.B(n_332),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_333),
.A2(n_334),
.B1(n_339),
.B2(n_340),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_333),
.B(n_342),
.C(n_343),
.Y(n_365)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_337),
.Y(n_356)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_340),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_343),
.B2(n_344),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_344),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_348),
.B(n_365),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_348),
.B(n_365),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_357),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_356),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_350),
.B(n_356),
.C(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_354),
.Y(n_372)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_357),
.Y(n_369)
);

XOR2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_362),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_358),
.B(n_382),
.C(n_383),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx8_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVxp67_ASAP7_75t_L g382 ( 
.A(n_363),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_364),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_368),
.B(n_370),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_368),
.B(n_370),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_380),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_371),
.B(n_381),
.C(n_384),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_373),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_372),
.B(n_374),
.C(n_375),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_376),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.Y(n_375)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_376),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_377),
.B(n_379),
.Y(n_400)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_384),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

MAJx2_ASAP7_75t_L g428 ( 
.A(n_385),
.B(n_391),
.C(n_393),
.Y(n_428)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_389),
.A2(n_391),
.B1(n_393),
.B2(n_394),
.Y(n_388)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_389),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_391),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_397),
.B(n_429),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_397),
.B(n_429),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_409),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_408),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_399),
.B(n_408),
.C(n_455),
.Y(n_454)
);

XNOR2x1_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_401),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_400),
.B(n_445),
.C(n_446),
.Y(n_444)
);

XNOR2x1_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_402),
.Y(n_445)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_405),
.Y(n_446)
);

INVx3_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_409),
.Y(n_455)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_420),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_410),
.B(n_422),
.C(n_427),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_418),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_415),
.Y(n_411)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_412),
.B(n_415),
.C(n_418),
.Y(n_442)
);

INVx6_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx4_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_422),
.B1(n_427),
.B2(n_428),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_426),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_423),
.B(n_426),
.Y(n_441)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_428),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_454),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_432),
.B(n_454),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_443),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_434),
.B(n_435),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_434),
.B(n_435),
.C(n_443),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_436),
.A2(n_437),
.B1(n_439),
.B2(n_440),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_436),
.B(n_466),
.C(n_467),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_441),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g443 ( 
.A(n_444),
.B(n_447),
.Y(n_443)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_444),
.B(n_448),
.C(n_453),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_448),
.A2(n_449),
.B1(n_452),
.B2(n_453),
.Y(n_447)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_448),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_449),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_473),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_458),
.B(n_473),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_459),
.B(n_464),
.Y(n_458)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_460),
.B(n_463),
.C(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_461),
.Y(n_462)
);

INVxp67_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_SL g464 ( 
.A(n_465),
.B(n_468),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_465),
.B(n_469),
.C(n_471),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_471),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_476),
.B(n_485),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_476),
.B(n_485),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_478),
.Y(n_476)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_477),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_482),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_479),
.B(n_482),
.C(n_492),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g488 ( 
.A(n_489),
.B(n_491),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_489),
.B(n_491),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_506),
.Y(n_495)
);

OAI21xp33_ASAP7_75t_L g510 ( 
.A1(n_496),
.A2(n_511),
.B(n_512),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g496 ( 
.A(n_497),
.B(n_500),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_497),
.B(n_500),
.Y(n_512)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_498),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_503),
.C(n_505),
.Y(n_500)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_501),
.B(n_503),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g507 ( 
.A(n_505),
.B(n_508),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g506 ( 
.A(n_507),
.B(n_509),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_507),
.B(n_509),
.Y(n_511)
);

BUFx12f_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_514),
.Y(n_517)
);

INVx13_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_517),
.B(n_518),
.Y(n_516)
);


endmodule