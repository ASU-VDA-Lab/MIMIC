module fake_jpeg_19909_n_325 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_325);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_325;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx3_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_2),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx13_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_26),
.B(n_0),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_19),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_42),
.B(n_32),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_51),
.B(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_32),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_42),
.A2(n_33),
.B1(n_28),
.B2(n_17),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_58),
.Y(n_78)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_62),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_35),
.A2(n_17),
.B1(n_33),
.B2(n_22),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_64),
.A2(n_35),
.B1(n_41),
.B2(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_74),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_69),
.A2(n_88),
.B1(n_40),
.B2(n_63),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_35),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_71),
.B(n_83),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_49),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_76),
.B(n_91),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_77),
.B(n_27),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_SL g81 ( 
.A(n_58),
.B(n_64),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_90),
.C(n_92),
.Y(n_107)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_53),
.Y(n_82)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_57),
.A2(n_38),
.B(n_41),
.C(n_19),
.Y(n_83)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_65),
.A2(n_41),
.B1(n_44),
.B2(n_17),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_59),
.B1(n_53),
.B2(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_52),
.B(n_28),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_87),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_52),
.B(n_43),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_66),
.A2(n_17),
.B1(n_44),
.B2(n_33),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_45),
.B(n_43),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_61),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_45),
.B(n_43),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_78),
.A2(n_33),
.B1(n_19),
.B2(n_25),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_96),
.Y(n_124)
);

OAI22x1_ASAP7_75t_L g98 ( 
.A1(n_78),
.A2(n_20),
.B1(n_34),
.B2(n_31),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_99),
.B1(n_104),
.B2(n_115),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_73),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_100),
.B(n_101),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_102),
.B(n_103),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_70),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_81),
.A2(n_33),
.B1(n_40),
.B2(n_22),
.Y(n_104)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_105),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_92),
.B1(n_90),
.B2(n_67),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_108),
.B(n_111),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_109),
.Y(n_126)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_80),
.Y(n_111)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_114),
.B(n_119),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_69),
.B1(n_68),
.B2(n_87),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_116),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_117),
.Y(n_148)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_93),
.Y(n_118)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_118),
.Y(n_145)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

AOI32xp33_ASAP7_75t_L g120 ( 
.A1(n_79),
.A2(n_85),
.A3(n_77),
.B1(n_83),
.B2(n_91),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_31),
.Y(n_139)
);

MAJx2_ASAP7_75t_L g121 ( 
.A(n_85),
.B(n_34),
.C(n_20),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_121),
.A2(n_34),
.B(n_27),
.Y(n_136)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_122),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_131),
.B1(n_140),
.B2(n_144),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_56),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_110),
.A2(n_67),
.B1(n_72),
.B2(n_82),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_76),
.B1(n_74),
.B2(n_63),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_100),
.B1(n_108),
.B2(n_118),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_136),
.B(n_139),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_110),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_137),
.B(n_138),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_107),
.B(n_56),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_22),
.B1(n_40),
.B2(n_50),
.Y(n_140)
);

BUFx12_ASAP7_75t_L g141 ( 
.A(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_105),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_104),
.A2(n_75),
.B(n_27),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_34),
.B(n_20),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_22),
.B1(n_75),
.B2(n_25),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_96),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_116),
.Y(n_150)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

AND2x6_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_98),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_180),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_132),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_153),
.B(n_163),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_138),
.B(n_97),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_154),
.B(n_162),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_143),
.A2(n_121),
.B(n_94),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_157),
.A2(n_170),
.B(n_172),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_160),
.A2(n_144),
.B1(n_141),
.B2(n_147),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_99),
.B1(n_112),
.B2(n_113),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_161),
.A2(n_178),
.B1(n_134),
.B2(n_135),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_128),
.B(n_119),
.C(n_113),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

OAI22x1_ASAP7_75t_L g164 ( 
.A1(n_143),
.A2(n_20),
.B1(n_34),
.B2(n_39),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_164),
.A2(n_151),
.B1(n_163),
.B2(n_172),
.Y(n_195)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_124),
.Y(n_165)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_165),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_147),
.B(n_25),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_166),
.B(n_167),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_124),
.Y(n_167)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_168),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_30),
.Y(n_169)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_169),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_146),
.A2(n_136),
.B(n_142),
.Y(n_170)
);

INVxp67_ASAP7_75t_SL g173 ( 
.A(n_141),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_126),
.A2(n_34),
.B(n_114),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_175),
.A2(n_140),
.B(n_141),
.Y(n_199)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_129),
.Y(n_177)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_127),
.A2(n_61),
.B1(n_30),
.B2(n_29),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_149),
.Y(n_179)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_129),
.B(n_30),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_181),
.A2(n_184),
.B1(n_186),
.B2(n_192),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_158),
.A2(n_134),
.B1(n_152),
.B2(n_161),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_165),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_188),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_158),
.A2(n_148),
.B1(n_145),
.B2(n_126),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_176),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_178),
.A2(n_148),
.B1(n_145),
.B2(n_131),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_195),
.B(n_202),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_199),
.A2(n_208),
.B(n_157),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_174),
.A2(n_123),
.B1(n_1),
.B2(n_3),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_203),
.A2(n_204),
.B1(n_180),
.B2(n_4),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_174),
.A2(n_123),
.B1(n_3),
.B2(n_4),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_175),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_154),
.B(n_29),
.Y(n_206)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_206),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_177),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_207),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_170),
.A2(n_0),
.B(n_3),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_209),
.A2(n_203),
.B1(n_204),
.B2(n_205),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_156),
.C(n_162),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_213),
.C(n_217),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_200),
.B(n_156),
.C(n_155),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_214),
.Y(n_240)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_155),
.C(n_160),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_189),
.B(n_184),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_218),
.B(n_223),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_199),
.A2(n_179),
.B1(n_171),
.B2(n_159),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_219),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_169),
.Y(n_220)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_220),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_229),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_201),
.B1(n_182),
.B2(n_181),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_196),
.B(n_29),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_SL g224 ( 
.A(n_208),
.B(n_14),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_224),
.B(n_228),
.Y(n_248)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_194),
.Y(n_226)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_226),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_30),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_230),
.B(n_231),
.Y(n_239)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_191),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_232),
.B(n_29),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_190),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_233),
.B(n_221),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_211),
.B(n_186),
.C(n_193),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_238),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_235),
.B(n_252),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_198),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_236),
.A2(n_12),
.B(n_5),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_241),
.B1(n_250),
.B2(n_253),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_192),
.C(n_39),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_216),
.A2(n_212),
.B1(n_223),
.B2(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_244),
.B(n_39),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_212),
.A2(n_227),
.B1(n_215),
.B2(n_214),
.Y(n_250)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_251),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_217),
.B(n_24),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_13),
.B1(n_5),
.B2(n_7),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_236),
.B(n_224),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_257),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_249),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_240),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_258),
.B(n_267),
.Y(n_276)
);

A2O1A1O1Ixp25_ASAP7_75t_L g259 ( 
.A1(n_243),
.A2(n_209),
.B(n_218),
.C(n_219),
.D(n_228),
.Y(n_259)
);

OAI211xp5_ASAP7_75t_L g286 ( 
.A1(n_259),
.A2(n_15),
.B(n_8),
.C(n_9),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_243),
.A2(n_242),
.B1(n_245),
.B2(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_239),
.Y(n_263)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_246),
.Y(n_265)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_265),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g282 ( 
.A(n_266),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g267 ( 
.A1(n_248),
.A2(n_220),
.B1(n_24),
.B2(n_23),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_244),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_270),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_23),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_24),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_271),
.A2(n_14),
.B(n_7),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_254),
.C(n_247),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_280),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_254),
.C(n_247),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_274),
.B(n_277),
.C(n_265),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_262),
.B(n_248),
.C(n_39),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_269),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g279 ( 
.A1(n_264),
.A2(n_12),
.B(n_5),
.Y(n_279)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_279),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_259),
.A2(n_14),
.B(n_8),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_284),
.A2(n_286),
.B(n_271),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_287),
.B(n_292),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_282),
.B(n_260),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_288),
.B(n_290),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_255),
.Y(n_290)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_281),
.B(n_263),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_293),
.B(n_294),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_273),
.B(n_39),
.C(n_24),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_275),
.B(n_276),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_297),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_16),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_283),
.A2(n_16),
.B1(n_10),
.B2(n_11),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_298),
.A2(n_277),
.B1(n_285),
.B2(n_11),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_286),
.B(n_10),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_285),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_301),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g302 ( 
.A(n_292),
.B(n_18),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_306),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_289),
.C(n_287),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_10),
.B(n_11),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_307),
.A2(n_0),
.B(n_18),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_305),
.B(n_294),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_313),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_304),
.B(n_18),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_18),
.C(n_23),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_315),
.C(n_23),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_305),
.B(n_12),
.Y(n_315)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_316),
.B(n_309),
.C(n_39),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_308),
.B(n_302),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_317),
.Y(n_321)
);

OAI21xp33_ASAP7_75t_L g322 ( 
.A1(n_321),
.A2(n_311),
.B(n_319),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_310),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_320),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_324),
.B(n_318),
.Y(n_325)
);


endmodule