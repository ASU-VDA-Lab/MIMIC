module real_jpeg_27307_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_334, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_334;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

HB1xp67_ASAP7_75t_L g106 ( 
.A(n_0),
.Y(n_106)
);

INVx11_ASAP7_75t_L g111 ( 
.A(n_0),
.Y(n_111)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_0),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_1),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_1),
.A2(n_31),
.B1(n_33),
.B2(n_184),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_1),
.A2(n_45),
.B1(n_46),
.B2(n_184),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_1),
.A2(n_64),
.B1(n_66),
.B2(n_184),
.Y(n_268)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_3),
.A2(n_31),
.B1(n_33),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_3),
.A2(n_45),
.B1(n_46),
.B2(n_50),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_3),
.A2(n_50),
.B1(n_64),
.B2(n_66),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_4),
.A2(n_31),
.B1(n_33),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_4),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_4),
.A2(n_27),
.B1(n_28),
.B2(n_53),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_4),
.A2(n_53),
.B1(n_64),
.B2(n_66),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_4),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_6),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g178 ( 
.A1(n_6),
.A2(n_31),
.B1(n_33),
.B2(n_150),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_6),
.A2(n_45),
.B1(n_46),
.B2(n_150),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_6),
.A2(n_64),
.B1(n_66),
.B2(n_150),
.Y(n_260)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_45),
.B1(n_46),
.B2(n_48),
.Y(n_44)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_9),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_9),
.B(n_30),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_9),
.B(n_33),
.Y(n_220)
);

AOI21xp33_ASAP7_75t_L g224 ( 
.A1(n_9),
.A2(n_33),
.B(n_220),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_9),
.A2(n_45),
.B1(n_46),
.B2(n_182),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_9),
.A2(n_61),
.B(n_64),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_9),
.B(n_89),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_9),
.A2(n_129),
.B1(n_130),
.B2(n_268),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_10),
.A2(n_35),
.B1(n_45),
.B2(n_46),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_10),
.A2(n_31),
.B1(n_33),
.B2(n_35),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_35),
.B1(n_64),
.B2(n_66),
.Y(n_197)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_12),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_31),
.B1(n_33),
.B2(n_123),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_12),
.A2(n_45),
.B1(n_46),
.B2(n_123),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_12),
.A2(n_64),
.B1(n_66),
.B2(n_123),
.Y(n_255)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g36 ( 
.A1(n_14),
.A2(n_27),
.B1(n_28),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_14),
.A2(n_31),
.B1(n_33),
.B2(n_37),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_14),
.A2(n_37),
.B1(n_45),
.B2(n_46),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_14),
.A2(n_37),
.B1(n_64),
.B2(n_66),
.Y(n_140)
);

INVx11_ASAP7_75t_SL g65 ( 
.A(n_15),
.Y(n_65)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_96),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_94),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_81),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_19),
.B(n_81),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_71),
.C(n_75),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_20),
.A2(n_21),
.B1(n_71),
.B2(n_320),
.Y(n_324)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_40),
.B2(n_70),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_22),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_22)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_23),
.A2(n_122),
.B(n_124),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_23),
.A2(n_38),
.B1(n_122),
.B2(n_149),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_23),
.A2(n_38),
.B1(n_149),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_24),
.B(n_73),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_24),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_24),
.A2(n_86),
.B(n_125),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_24),
.A2(n_30),
.B1(n_181),
.B2(n_183),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_27),
.B(n_29),
.C(n_30),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B1(n_31),
.B2(n_33),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_25),
.B(n_33),
.Y(n_195)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

HAxp5_ASAP7_75t_SL g181 ( 
.A(n_27),
.B(n_182),
.CON(n_181),
.SN(n_181)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_29),
.A2(n_31),
.B1(n_181),
.B2(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_30),
.B(n_125),
.Y(n_124)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_31),
.A2(n_33),
.B1(n_48),
.B2(n_56),
.Y(n_55)
);

AOI32xp33_ASAP7_75t_L g218 ( 
.A1(n_31),
.A2(n_45),
.A3(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_218)
);

BUFx4f_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_34),
.A2(n_38),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_36),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_38),
.B(n_74),
.Y(n_86)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_58),
.B2(n_69),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_42),
.B(n_58),
.C(n_70),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_51),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_43),
.A2(n_77),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_49),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_44),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_44),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_44),
.A2(n_54),
.B1(n_79),
.B2(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_44),
.A2(n_54),
.B1(n_178),
.B2(n_179),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_44),
.A2(n_54),
.B1(n_178),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_44),
.A2(n_54),
.B1(n_206),
.B2(n_224),
.Y(n_223)
);

OAI22xp33_ASAP7_75t_L g60 ( 
.A1(n_45),
.A2(n_46),
.B1(n_61),
.B2(n_62),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp33_ASAP7_75t_SL g221 ( 
.A(n_46),
.B(n_56),
.Y(n_221)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_46),
.A2(n_62),
.B(n_182),
.C(n_247),
.Y(n_246)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_51),
.A2(n_89),
.B(n_119),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_54),
.Y(n_51)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_56),
.Y(n_219)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_58),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_58),
.A2(n_69),
.B1(n_76),
.B2(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_63),
.B(n_67),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_59),
.A2(n_63),
.B1(n_114),
.B2(n_115),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_59),
.A2(n_115),
.B(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_59),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_59),
.A2(n_67),
.B(n_133),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_59),
.A2(n_63),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_59),
.A2(n_156),
.B(n_228),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_59),
.A2(n_63),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_59),
.A2(n_63),
.B1(n_227),
.B2(n_245),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_63),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g63 ( 
.A1(n_61),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_63),
.A2(n_114),
.B(n_144),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_63),
.B(n_182),
.Y(n_266)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_66),
.B(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_66),
.B(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_68),
.B(n_135),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_71),
.C(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_71),
.A2(n_317),
.B1(n_319),
.B2(n_320),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_71),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_75),
.B(n_324),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_76),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B(n_80),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_77),
.A2(n_89),
.B(n_90),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_77),
.A2(n_80),
.B(n_90),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_83),
.A2(n_84),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_313),
.A3(n_325),
.B1(n_331),
.B2(n_332),
.C(n_334),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_167),
.B(n_312),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_151),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_99),
.B(n_151),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_126),
.C(n_137),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_100),
.A2(n_101),
.B1(n_126),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_116),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_102),
.B(n_118),
.C(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_113),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_103),
.B(n_113),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_109),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_104),
.A2(n_130),
.B(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_105),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_105),
.A2(n_112),
.B(n_142),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_105),
.A2(n_110),
.B1(n_259),
.B2(n_261),
.Y(n_258)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_106),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_130),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_109),
.A2(n_129),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_111),
.A2(n_129),
.B1(n_140),
.B2(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_112),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_119),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_126),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_132),
.B2(n_136),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_127),
.A2(n_128),
.B1(n_163),
.B2(n_164),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_132),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_128),
.A2(n_161),
.B(n_164),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B(n_131),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_129),
.A2(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_129),
.A2(n_130),
.B1(n_260),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_132),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_134),
.B(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_137),
.B(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_146),
.C(n_147),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_138),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_143),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_143),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_156),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_146),
.A2(n_147),
.B1(n_148),
.B2(n_302),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_146),
.Y(n_302)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_165),
.B2(n_166),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_154),
.B(n_160),
.C(n_166),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_157),
.B(n_159),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_157),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_159),
.B(n_315),
.C(n_321),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_159),
.A2(n_315),
.B1(n_316),
.B2(n_330),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_159),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_165),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_168),
.A2(n_306),
.B(n_311),
.Y(n_167)
);

O2A1O1Ixp33_ASAP7_75t_SL g168 ( 
.A1(n_169),
.A2(n_210),
.B(n_292),
.C(n_305),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_198),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_170),
.B(n_198),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_185),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_173),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_172),
.B(n_173),
.C(n_185),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_180),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_177),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_180),
.B(n_201),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_182),
.B(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_183),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_193),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_190),
.B2(n_191),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_187),
.B(n_191),
.C(n_193),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_202),
.C(n_204),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_199),
.A2(n_200),
.B1(n_287),
.B2(n_289),
.Y(n_286)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_202),
.A2(n_203),
.B1(n_204),
.B2(n_288),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_204),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_205),
.B(n_232),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_207),
.A2(n_208),
.B1(n_209),
.B2(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_211),
.B(n_291),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_284),
.B(n_290),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_238),
.B(n_283),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_229),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_214),
.B(n_229),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_222),
.C(n_225),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_215),
.A2(n_216),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_218),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_222),
.A2(n_223),
.B1(n_225),
.B2(n_226),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_285)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_277),
.B(n_282),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_240),
.A2(n_256),
.B(n_276),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_248),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_241),
.B(n_248),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_242),
.A2(n_243),
.B1(n_246),
.B2(n_263),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_246),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_253),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_253),
.C(n_254),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_255),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_264),
.B(n_275),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_262),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_258),
.B(n_262),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_265),
.A2(n_269),
.B(n_274),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_267),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_285),
.B(n_286),
.Y(n_290)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_287),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_293),
.B(n_294),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_303),
.B2(n_304),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_300),
.C(n_304),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_307),
.B(n_308),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_323),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_314),
.B(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_321),
.A2(n_322),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_326),
.B(n_327),
.Y(n_331)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);


endmodule