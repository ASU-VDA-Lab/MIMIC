module fake_ibex_103_n_1946 (n_151, n_85, n_395, n_84, n_64, n_171, n_103, n_389, n_204, n_274, n_387, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_193, n_108, n_350, n_165, n_86, n_70, n_255, n_175, n_398, n_59, n_28, n_125, n_304, n_191, n_5, n_62, n_71, n_153, n_194, n_249, n_334, n_312, n_239, n_94, n_134, n_371, n_403, n_357, n_88, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_176, n_58, n_43, n_216, n_33, n_166, n_163, n_114, n_236, n_34, n_376, n_377, n_15, n_24, n_189, n_280, n_317, n_340, n_375, n_105, n_187, n_1, n_154, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_117, n_265, n_158, n_259, n_276, n_339, n_210, n_348, n_220, n_91, n_287, n_54, n_243, n_19, n_228, n_147, n_251, n_384, n_373, n_244, n_73, n_343, n_310, n_323, n_143, n_106, n_386, n_8, n_224, n_183, n_67, n_333, n_110, n_306, n_400, n_47, n_169, n_10, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_7, n_109, n_127, n_121, n_48, n_325, n_57, n_301, n_296, n_120, n_168, n_155, n_315, n_13, n_122, n_116, n_370, n_0, n_289, n_12, n_150, n_286, n_321, n_133, n_51, n_215, n_279, n_49, n_374, n_235, n_22, n_136, n_261, n_30, n_367, n_221, n_355, n_407, n_102, n_52, n_99, n_269, n_156, n_126, n_356, n_25, n_104, n_45, n_141, n_222, n_186, n_349, n_295, n_331, n_230, n_96, n_185, n_388, n_352, n_290, n_174, n_157, n_219, n_246, n_31, n_146, n_207, n_167, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_139, n_275, n_98, n_129, n_267, n_245, n_229, n_209, n_347, n_335, n_82, n_263, n_27, n_353, n_359, n_299, n_87, n_262, n_75, n_137, n_338, n_173, n_363, n_402, n_180, n_369, n_201, n_14, n_351, n_368, n_257, n_77, n_44, n_401, n_66, n_305, n_307, n_192, n_140, n_365, n_4, n_6, n_100, n_179, n_354, n_206, n_392, n_329, n_26, n_188, n_200, n_199, n_410, n_308, n_135, n_283, n_366, n_397, n_111, n_36, n_18, n_322, n_53, n_227, n_115, n_11, n_248, n_92, n_101, n_190, n_138, n_409, n_214, n_238, n_332, n_211, n_218, n_314, n_132, n_277, n_337, n_225, n_360, n_272, n_23, n_223, n_381, n_382, n_95, n_405, n_285, n_288, n_247, n_320, n_379, n_55, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_148, n_2, n_342, n_233, n_385, n_118, n_378, n_164, n_38, n_198, n_264, n_217, n_324, n_391, n_78, n_20, n_69, n_390, n_39, n_178, n_303, n_362, n_93, n_162, n_240, n_282, n_61, n_266, n_42, n_294, n_112, n_46, n_284, n_80, n_172, n_250, n_313, n_345, n_408, n_119, n_361, n_72, n_319, n_195, n_212, n_311, n_406, n_97, n_197, n_181, n_131, n_123, n_260, n_302, n_344, n_393, n_297, n_41, n_252, n_396, n_83, n_32, n_107, n_149, n_399, n_254, n_213, n_271, n_241, n_68, n_292, n_394, n_79, n_81, n_35, n_364, n_159, n_202, n_231, n_298, n_160, n_184, n_56, n_232, n_380, n_281, n_1946);

input n_151;
input n_85;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_389;
input n_204;
input n_274;
input n_387;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_193;
input n_108;
input n_350;
input n_165;
input n_86;
input n_70;
input n_255;
input n_175;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_5;
input n_62;
input n_71;
input n_153;
input n_194;
input n_249;
input n_334;
input n_312;
input n_239;
input n_94;
input n_134;
input n_371;
input n_403;
input n_357;
input n_88;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_166;
input n_163;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_15;
input n_24;
input n_189;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_1;
input n_154;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_117;
input n_265;
input n_158;
input n_259;
input n_276;
input n_339;
input n_210;
input n_348;
input n_220;
input n_91;
input n_287;
input n_54;
input n_243;
input n_19;
input n_228;
input n_147;
input n_251;
input n_384;
input n_373;
input n_244;
input n_73;
input n_343;
input n_310;
input n_323;
input n_143;
input n_106;
input n_386;
input n_8;
input n_224;
input n_183;
input n_67;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_169;
input n_10;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_7;
input n_109;
input n_127;
input n_121;
input n_48;
input n_325;
input n_57;
input n_301;
input n_296;
input n_120;
input n_168;
input n_155;
input n_315;
input n_13;
input n_122;
input n_116;
input n_370;
input n_0;
input n_289;
input n_12;
input n_150;
input n_286;
input n_321;
input n_133;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_22;
input n_136;
input n_261;
input n_30;
input n_367;
input n_221;
input n_355;
input n_407;
input n_102;
input n_52;
input n_99;
input n_269;
input n_156;
input n_126;
input n_356;
input n_25;
input n_104;
input n_45;
input n_141;
input n_222;
input n_186;
input n_349;
input n_295;
input n_331;
input n_230;
input n_96;
input n_185;
input n_388;
input n_352;
input n_290;
input n_174;
input n_157;
input n_219;
input n_246;
input n_31;
input n_146;
input n_207;
input n_167;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_139;
input n_275;
input n_98;
input n_129;
input n_267;
input n_245;
input n_229;
input n_209;
input n_347;
input n_335;
input n_82;
input n_263;
input n_27;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_75;
input n_137;
input n_338;
input n_173;
input n_363;
input n_402;
input n_180;
input n_369;
input n_201;
input n_14;
input n_351;
input n_368;
input n_257;
input n_77;
input n_44;
input n_401;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_365;
input n_4;
input n_6;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_329;
input n_26;
input n_188;
input n_200;
input n_199;
input n_410;
input n_308;
input n_135;
input n_283;
input n_366;
input n_397;
input n_111;
input n_36;
input n_18;
input n_322;
input n_53;
input n_227;
input n_115;
input n_11;
input n_248;
input n_92;
input n_101;
input n_190;
input n_138;
input n_409;
input n_214;
input n_238;
input n_332;
input n_211;
input n_218;
input n_314;
input n_132;
input n_277;
input n_337;
input n_225;
input n_360;
input n_272;
input n_23;
input n_223;
input n_381;
input n_382;
input n_95;
input n_405;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_55;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_118;
input n_378;
input n_164;
input n_38;
input n_198;
input n_264;
input n_217;
input n_324;
input n_391;
input n_78;
input n_20;
input n_69;
input n_390;
input n_39;
input n_178;
input n_303;
input n_362;
input n_93;
input n_162;
input n_240;
input n_282;
input n_61;
input n_266;
input n_42;
input n_294;
input n_112;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_313;
input n_345;
input n_408;
input n_119;
input n_361;
input n_72;
input n_319;
input n_195;
input n_212;
input n_311;
input n_406;
input n_97;
input n_197;
input n_181;
input n_131;
input n_123;
input n_260;
input n_302;
input n_344;
input n_393;
input n_297;
input n_41;
input n_252;
input n_396;
input n_83;
input n_32;
input n_107;
input n_149;
input n_399;
input n_254;
input n_213;
input n_271;
input n_241;
input n_68;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_159;
input n_202;
input n_231;
input n_298;
input n_160;
input n_184;
input n_56;
input n_232;
input n_380;
input n_281;

output n_1946;

wire n_1084;
wire n_1474;
wire n_1295;
wire n_507;
wire n_992;
wire n_1582;
wire n_766;
wire n_1110;
wire n_1382;
wire n_1596;
wire n_926;
wire n_1079;
wire n_1100;
wire n_845;
wire n_446;
wire n_1930;
wire n_452;
wire n_1234;
wire n_1594;
wire n_1944;
wire n_1802;
wire n_773;
wire n_1469;
wire n_821;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_957;
wire n_1652;
wire n_969;
wire n_678;
wire n_1859;
wire n_1883;
wire n_1125;
wire n_733;
wire n_622;
wire n_1226;
wire n_1034;
wire n_1765;
wire n_872;
wire n_1873;
wire n_1619;
wire n_457;
wire n_1666;
wire n_494;
wire n_930;
wire n_1044;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_1722;
wire n_911;
wire n_652;
wire n_781;
wire n_475;
wire n_802;
wire n_1233;
wire n_1045;
wire n_1856;
wire n_500;
wire n_963;
wire n_1782;
wire n_531;
wire n_1308;
wire n_556;
wire n_1138;
wire n_498;
wire n_708;
wire n_1096;
wire n_1391;
wire n_884;
wire n_667;
wire n_850;
wire n_879;
wire n_723;
wire n_1144;
wire n_1392;
wire n_1268;
wire n_739;
wire n_853;
wire n_948;
wire n_504;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_481;
wire n_876;
wire n_497;
wire n_711;
wire n_1840;
wire n_671;
wire n_989;
wire n_1908;
wire n_1668;
wire n_1641;
wire n_829;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_1681;
wire n_939;
wire n_1636;
wire n_1687;
wire n_655;
wire n_1766;
wire n_550;
wire n_1922;
wire n_557;
wire n_641;
wire n_1937;
wire n_893;
wire n_527;
wire n_1654;
wire n_496;
wire n_434;
wire n_1258;
wire n_1344;
wire n_1929;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1195;
wire n_824;
wire n_1945;
wire n_441;
wire n_694;
wire n_787;
wire n_523;
wire n_614;
wire n_431;
wire n_1130;
wire n_1228;
wire n_1081;
wire n_538;
wire n_1155;
wire n_1292;
wire n_459;
wire n_1576;
wire n_1664;
wire n_518;
wire n_852;
wire n_1427;
wire n_1133;
wire n_1926;
wire n_904;
wire n_1778;
wire n_448;
wire n_646;
wire n_466;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_1496;
wire n_1910;
wire n_715;
wire n_530;
wire n_1663;
wire n_1214;
wire n_1274;
wire n_420;
wire n_1606;
wire n_769;
wire n_1595;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_1886;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_777;
wire n_917;
wire n_968;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_1493;
wire n_1313;
wire n_558;
wire n_666;
wire n_1638;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_793;
wire n_937;
wire n_1645;
wire n_973;
wire n_1038;
wire n_618;
wire n_1943;
wire n_1863;
wire n_1269;
wire n_662;
wire n_979;
wire n_1309;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_629;
wire n_1445;
wire n_573;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_433;
wire n_439;
wire n_1672;
wire n_1007;
wire n_643;
wire n_1276;
wire n_1637;
wire n_841;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_1588;
wire n_1301;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_554;
wire n_553;
wire n_1078;
wire n_1219;
wire n_713;
wire n_1865;
wire n_1252;
wire n_1170;
wire n_1927;
wire n_605;
wire n_539;
wire n_630;
wire n_1869;
wire n_567;
wire n_1853;
wire n_745;
wire n_447;
wire n_1753;
wire n_562;
wire n_564;
wire n_1322;
wire n_1305;
wire n_795;
wire n_592;
wire n_1248;
wire n_762;
wire n_1388;
wire n_800;
wire n_706;
wire n_784;
wire n_684;
wire n_1653;
wire n_1375;
wire n_1356;
wire n_894;
wire n_1118;
wire n_692;
wire n_1881;
wire n_709;
wire n_1296;
wire n_499;
wire n_702;
wire n_971;
wire n_1326;
wire n_1350;
wire n_451;
wire n_906;
wire n_1093;
wire n_1764;
wire n_978;
wire n_899;
wire n_579;
wire n_1799;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_1190;
wire n_1304;
wire n_744;
wire n_563;
wire n_1506;
wire n_881;
wire n_1702;
wire n_734;
wire n_1558;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_1370;
wire n_1209;
wire n_1708;
wire n_551;
wire n_1616;
wire n_729;
wire n_1569;
wire n_1434;
wire n_603;
wire n_1649;
wire n_422;
wire n_1936;
wire n_1717;
wire n_1609;
wire n_1613;
wire n_820;
wire n_805;
wire n_670;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_544;
wire n_1787;
wire n_1281;
wire n_1447;
wire n_695;
wire n_1549;
wire n_639;
wire n_1867;
wire n_1531;
wire n_1332;
wire n_482;
wire n_1424;
wire n_1742;
wire n_1818;
wire n_870;
wire n_1709;
wire n_1610;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_609;
wire n_1040;
wire n_476;
wire n_1159;
wire n_1368;
wire n_1154;
wire n_455;
wire n_1701;
wire n_1243;
wire n_1121;
wire n_693;
wire n_737;
wire n_606;
wire n_1571;
wire n_462;
wire n_1407;
wire n_1235;
wire n_1821;
wire n_1003;
wire n_889;
wire n_435;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_1543;
wire n_823;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_1441;
wire n_1924;
wire n_1921;
wire n_657;
wire n_1156;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_822;
wire n_1042;
wire n_1888;
wire n_743;
wire n_754;
wire n_1786;
wire n_1319;
wire n_1553;
wire n_1041;
wire n_1090;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_1731;
wire n_1905;
wire n_1031;
wire n_981;
wire n_1591;
wire n_583;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_663;
wire n_1377;
wire n_1583;
wire n_1521;
wire n_1152;
wire n_974;
wire n_1036;
wire n_1831;
wire n_608;
wire n_864;
wire n_412;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_449;
wire n_1733;
wire n_1634;
wire n_1932;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_1508;
wire n_421;
wire n_738;
wire n_1217;
wire n_1715;
wire n_1189;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_1255;
wire n_1700;
wire n_1218;
wire n_1181;
wire n_1140;
wire n_1772;
wire n_1056;
wire n_1283;
wire n_1446;
wire n_1487;
wire n_840;
wire n_1203;
wire n_1421;
wire n_561;
wire n_846;
wire n_471;
wire n_1793;
wire n_1237;
wire n_859;
wire n_965;
wire n_1109;
wire n_1633;
wire n_1711;
wire n_1051;
wire n_1008;
wire n_458;
wire n_1498;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_1032;
wire n_936;
wire n_469;
wire n_1884;
wire n_1825;
wire n_1589;
wire n_1210;
wire n_591;
wire n_1933;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_832;
wire n_1792;
wire n_1712;
wire n_590;
wire n_1568;
wire n_1877;
wire n_1184;
wire n_1477;
wire n_1724;
wire n_1364;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_929;
wire n_637;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_1918;
wire n_574;
wire n_515;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_907;
wire n_1179;
wire n_1153;
wire n_1751;
wire n_669;
wire n_1737;
wire n_521;
wire n_1117;
wire n_1273;
wire n_1748;
wire n_1083;
wire n_1014;
wire n_724;
wire n_437;
wire n_938;
wire n_1178;
wire n_474;
wire n_878;
wire n_594;
wire n_1464;
wire n_1566;
wire n_944;
wire n_1848;
wire n_623;
wire n_585;
wire n_1334;
wire n_483;
wire n_1695;
wire n_1418;
wire n_1137;
wire n_660;
wire n_524;
wire n_1200;
wire n_1120;
wire n_576;
wire n_1602;
wire n_1776;
wire n_1852;
wire n_1522;
wire n_1279;
wire n_931;
wire n_827;
wire n_607;
wire n_1064;
wire n_1408;
wire n_1028;
wire n_1264;
wire n_1935;
wire n_1146;
wire n_488;
wire n_705;
wire n_1548;
wire n_429;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_589;
wire n_1896;
wire n_472;
wire n_1704;
wire n_847;
wire n_1436;
wire n_413;
wire n_1069;
wire n_1485;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_679;
wire n_1345;
wire n_696;
wire n_837;
wire n_1590;
wire n_640;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_596;
wire n_1545;
wire n_456;
wire n_1471;
wire n_1738;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_801;
wire n_1479;
wire n_1046;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_651;
wire n_721;
wire n_814;
wire n_1864;
wire n_943;
wire n_1086;
wire n_1523;
wire n_1756;
wire n_1470;
wire n_444;
wire n_1761;
wire n_1836;
wire n_1593;
wire n_986;
wire n_495;
wire n_1420;
wire n_1750;
wire n_1775;
wire n_1699;
wire n_411;
wire n_927;
wire n_1563;
wire n_615;
wire n_803;
wire n_1875;
wire n_1615;
wire n_1087;
wire n_757;
wire n_1539;
wire n_712;
wire n_1400;
wire n_1599;
wire n_1806;
wire n_650;
wire n_1575;
wire n_1448;
wire n_517;
wire n_817;
wire n_555;
wire n_951;
wire n_468;
wire n_1580;
wire n_1574;
wire n_780;
wire n_502;
wire n_1705;
wire n_633;
wire n_1746;
wire n_726;
wire n_532;
wire n_1439;
wire n_863;
wire n_597;
wire n_1832;
wire n_1128;
wire n_1266;
wire n_1300;
wire n_807;
wire n_741;
wire n_430;
wire n_1785;
wire n_486;
wire n_1870;
wire n_1405;
wire n_997;
wire n_1428;
wire n_891;
wire n_1528;
wire n_1495;
wire n_717;
wire n_1357;
wire n_1512;
wire n_668;
wire n_871;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_485;
wire n_1315;
wire n_1413;
wire n_811;
wire n_808;
wire n_945;
wire n_460;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_1461;
wire n_461;
wire n_903;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_1378;
wire n_1048;
wire n_774;
wire n_1925;
wire n_588;
wire n_1430;
wire n_1251;
wire n_1247;
wire n_528;
wire n_836;
wire n_1475;
wire n_1263;
wire n_443;
wire n_1185;
wire n_1683;
wire n_436;
wire n_1122;
wire n_628;
wire n_890;
wire n_874;
wire n_1505;
wire n_1163;
wire n_677;
wire n_1514;
wire n_964;
wire n_916;
wire n_503;
wire n_895;
wire n_687;
wire n_1035;
wire n_1535;
wire n_751;
wire n_1127;
wire n_932;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_540;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_1437;
wire n_529;
wire n_626;
wire n_1707;
wire n_1941;
wire n_1679;
wire n_1497;
wire n_1578;
wire n_1143;
wire n_1783;
wire n_418;
wire n_510;
wire n_972;
wire n_1815;
wire n_601;
wire n_610;
wire n_1917;
wire n_1444;
wire n_920;
wire n_664;
wire n_1067;
wire n_994;
wire n_1857;
wire n_1920;
wire n_545;
wire n_887;
wire n_1162;
wire n_1894;
wire n_961;
wire n_634;
wire n_991;
wire n_1331;
wire n_1349;
wire n_1223;
wire n_1323;
wire n_578;
wire n_1739;
wire n_432;
wire n_1777;
wire n_1353;
wire n_423;
wire n_1429;
wire n_1546;
wire n_1432;
wire n_1320;
wire n_996;
wire n_915;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_1727;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_542;
wire n_1294;
wire n_1601;
wire n_900;
wire n_1351;
wire n_647;
wire n_1380;
wire n_1367;
wire n_1291;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_1830;
wire n_1629;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_1340;
wire n_1626;
wire n_674;
wire n_1850;
wire n_1660;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_552;
wire n_1112;
wire n_1267;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_1816;
wire n_1612;
wire n_703;
wire n_426;
wire n_1172;
wire n_1099;
wire n_598;
wire n_1422;
wire n_508;
wire n_453;
wire n_1527;
wire n_1055;
wire n_1524;
wire n_673;
wire n_798;
wire n_1754;
wire n_1177;
wire n_1025;
wire n_1517;
wire n_690;
wire n_1225;
wire n_982;
wire n_1624;
wire n_785;
wire n_604;
wire n_1598;
wire n_977;
wire n_1895;
wire n_719;
wire n_1491;
wire n_1860;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_642;
wire n_1607;
wire n_1625;
wire n_933;
wire n_1774;
wire n_1797;
wire n_1037;
wire n_1899;
wire n_464;
wire n_1348;
wire n_838;
wire n_1289;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_742;
wire n_1191;
wire n_1503;
wire n_1052;
wire n_789;
wire n_1942;
wire n_656;
wire n_602;
wire n_842;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_636;
wire n_1259;
wire n_490;
wire n_595;
wire n_1001;
wire n_570;
wire n_1396;
wire n_1224;
wire n_1923;
wire n_1538;
wire n_487;
wire n_454;
wire n_1017;
wire n_730;
wire n_1456;
wire n_1889;
wire n_625;
wire n_619;
wire n_1124;
wire n_611;
wire n_1690;
wire n_1673;
wire n_922;
wire n_1790;
wire n_851;
wire n_993;
wire n_1725;
wire n_1135;
wire n_1820;
wire n_1800;
wire n_541;
wire n_613;
wire n_659;
wire n_1494;
wire n_1550;
wire n_1066;
wire n_1169;
wire n_571;
wire n_648;
wire n_1726;
wire n_1938;
wire n_830;
wire n_473;
wire n_1241;
wire n_445;
wire n_1072;
wire n_1231;
wire n_1173;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_826;
wire n_1337;
wire n_1906;
wire n_1647;
wire n_1901;
wire n_768;
wire n_839;
wire n_1278;
wire n_796;
wire n_797;
wire n_1006;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_1063;
wire n_1270;
wire n_834;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_1054;
wire n_722;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_804;
wire n_484;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_480;
wire n_1057;
wire n_1473;
wire n_516;
wire n_1403;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_506;
wire n_868;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_1457;
wire n_905;
wire n_975;
wire n_675;
wire n_463;
wire n_624;
wire n_520;
wire n_934;
wire n_775;
wire n_512;
wire n_950;
wire n_685;
wire n_1222;
wire n_1630;
wire n_1879;
wire n_1198;
wire n_1311;
wire n_1261;
wire n_776;
wire n_1114;
wire n_818;
wire n_1167;
wire n_1282;
wire n_1321;
wire n_700;
wire n_1779;
wire n_1770;
wire n_1107;
wire n_1846;
wire n_1573;
wire n_525;
wire n_815;
wire n_919;
wire n_535;
wire n_681;
wire n_415;
wire n_1718;
wire n_1411;
wire n_1139;
wire n_1018;
wire n_858;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_782;
wire n_616;
wire n_1885;
wire n_1740;
wire n_1838;
wire n_833;
wire n_1343;
wire n_1801;
wire n_1371;
wire n_1513;
wire n_728;
wire n_1788;
wire n_786;
wire n_505;
wire n_1621;
wire n_1919;
wire n_1342;
wire n_501;
wire n_752;
wire n_958;
wire n_1175;
wire n_1416;
wire n_1659;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_1435;
wire n_1688;
wire n_792;
wire n_1314;
wire n_1433;
wire n_575;
wire n_1242;
wire n_1119;
wire n_1085;
wire n_419;
wire n_1907;
wire n_885;
wire n_1530;
wire n_513;
wire n_877;
wire n_1088;
wire n_896;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_631;
wire n_794;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_428;
wire n_697;
wire n_1105;
wire n_1459;
wire n_912;
wire n_1893;
wire n_1570;
wire n_424;
wire n_701;
wire n_995;
wire n_1000;
wire n_1931;
wire n_1256;
wire n_587;
wire n_1303;
wire n_1771;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_812;
wire n_1050;
wire n_599;
wire n_1769;
wire n_1060;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_1632;
wire n_688;
wire n_1542;
wire n_946;
wire n_1586;
wire n_707;
wire n_1362;
wire n_1547;
wire n_1097;
wire n_1909;
wire n_621;
wire n_956;
wire n_790;
wire n_1541;
wire n_1812;
wire n_586;
wire n_1330;
wire n_638;
wire n_1697;
wire n_1872;
wire n_1940;
wire n_593;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_1767;
wire n_1939;
wire n_1768;
wire n_1443;
wire n_478;
wire n_1585;
wire n_1861;
wire n_1564;
wire n_1631;
wire n_1623;
wire n_861;
wire n_1828;
wire n_1389;
wire n_1131;
wire n_547;
wire n_1798;
wire n_727;
wire n_1077;
wire n_1554;
wire n_1481;
wire n_1584;
wire n_1928;
wire n_828;
wire n_1438;
wire n_753;
wire n_747;
wire n_645;
wire n_1147;
wire n_1363;
wire n_1691;
wire n_1098;
wire n_584;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_1693;
wire n_698;
wire n_1892;
wire n_1061;
wire n_682;
wire n_1373;
wire n_1686;
wire n_1302;
wire n_886;
wire n_1010;
wire n_883;
wire n_417;
wire n_755;
wire n_1029;
wire n_470;
wire n_770;
wire n_1635;
wire n_1572;
wire n_941;
wire n_1245;
wire n_1317;
wire n_632;
wire n_1329;
wire n_854;
wire n_714;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_1734;
wire n_1876;
wire n_740;
wire n_549;
wire n_533;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_967;
wire n_736;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_465;
wire n_1486;
wire n_1068;
wire n_617;
wire n_1833;
wire n_914;
wire n_526;
wire n_1024;
wire n_1141;
wire n_1197;
wire n_1168;
wire n_865;
wire n_569;
wire n_600;
wire n_1556;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_1759;
wire n_987;
wire n_750;
wire n_1299;
wire n_665;
wire n_1101;
wire n_1720;
wire n_880;
wire n_654;
wire n_1911;
wire n_731;
wire n_1336;
wire n_758;
wire n_1166;
wire n_710;
wire n_720;
wire n_1390;
wire n_1023;
wire n_568;
wire n_1358;
wire n_813;
wire n_1211;
wire n_1397;
wire n_1284;
wire n_1359;
wire n_1116;
wire n_1758;
wire n_791;
wire n_1532;
wire n_1419;
wire n_543;
wire n_580;
wire n_1784;
wire n_1685;
wire n_1082;
wire n_1213;
wire n_1193;
wire n_980;
wire n_849;
wire n_1488;
wire n_1074;
wire n_759;
wire n_1379;
wire n_1721;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_536;
wire n_1866;
wire n_1220;
wire n_467;
wire n_1398;
wire n_427;
wire n_1262;
wire n_1904;
wire n_442;
wire n_1692;
wire n_438;
wire n_1012;
wire n_1805;
wire n_689;
wire n_960;
wire n_1022;
wire n_1760;
wire n_676;
wire n_1240;
wire n_1183;
wire n_1204;
wire n_1151;
wire n_1814;
wire n_771;
wire n_999;
wire n_514;
wire n_1092;
wire n_1808;
wire n_560;
wire n_1658;
wire n_1386;
wire n_910;
wire n_635;
wire n_844;
wire n_1728;
wire n_1020;
wire n_783;
wire n_1385;
wire n_1142;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_1499;
wire n_1500;
wire n_1868;
wire n_966;
wire n_949;
wire n_704;
wire n_924;
wire n_1600;
wire n_477;
wire n_1661;
wire n_1757;
wire n_699;
wire n_918;
wire n_1913;
wire n_672;
wire n_1039;
wire n_1043;
wire n_1402;
wire n_735;
wire n_1450;
wire n_566;
wire n_416;
wire n_581;
wire n_1365;
wire n_1472;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_548;
wire n_1158;
wire n_763;
wire n_1882;
wire n_1915;
wire n_940;
wire n_1762;
wire n_1404;
wire n_546;
wire n_788;
wire n_1736;
wire n_1160;
wire n_1442;
wire n_658;
wire n_1216;
wire n_1891;
wire n_1026;
wire n_1454;
wire n_1033;
wire n_627;
wire n_990;
wire n_1383;
wire n_888;
wire n_1325;
wire n_582;
wire n_1483;
wire n_1703;
wire n_653;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1059;
wire n_799;
wire n_691;
wire n_1804;
wire n_1581;
wire n_522;
wire n_479;
wire n_534;
wire n_1837;
wire n_511;
wire n_1744;
wire n_1414;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_1111;
wire n_1819;
wire n_1341;
wire n_1807;
wire n_1310;
wire n_1745;
wire n_1714;
wire n_612;
wire n_1611;
wire n_955;
wire n_440;
wire n_1333;
wire n_1916;
wire n_414;
wire n_952;
wire n_1675;
wire n_1640;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_1511;
wire n_1791;
wire n_537;
wire n_1113;
wire n_1651;
wire n_1468;
wire n_913;
wire n_509;
wire n_1164;
wire n_1732;
wire n_1354;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_680;
wire n_1355;
wire n_809;
wire n_856;
wire n_779;
wire n_1559;
wire n_1579;
wire n_1280;
wire n_493;
wire n_1335;
wire n_1934;
wire n_1900;
wire n_519;
wire n_1843;
wire n_1665;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_1287;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_661;
wire n_1902;
wire n_683;
wire n_1194;
wire n_1150;
wire n_620;
wire n_1399;
wire n_450;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_686;
wire n_572;
wire n_867;
wire n_983;
wire n_1417;
wire n_644;
wire n_577;
wire n_970;
wire n_491;
wire n_921;
wire n_489;
wire n_1534;
wire n_908;
wire n_1346;
wire n_565;
wire n_1123;
wire n_1272;
wire n_1393;
wire n_984;
wire n_1655;
wire n_1410;
wire n_988;
wire n_760;
wire n_1157;
wire n_806;
wire n_1186;
wire n_1743;
wire n_492;
wire n_649;
wire n_1854;
wire n_866;
wire n_559;
wire n_425;

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_29),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_43),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_260),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_331),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_15),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_318),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_201),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_333),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_263),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_71),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_353),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_314),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_248),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_305),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_206),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_292),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_357),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_388),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_35),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_407),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_54),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_241),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_268),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_112),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_370),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_209),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_313),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_258),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_233),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_327),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_14),
.Y(n_441)
);

INVx1_ASAP7_75t_SL g442 ( 
.A(n_141),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_378),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_185),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_315),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_51),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_328),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_59),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_7),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_157),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_42),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g452 ( 
.A(n_65),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_214),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_15),
.Y(n_454)
);

INVx2_ASAP7_75t_SL g455 ( 
.A(n_223),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_301),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_170),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_335),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_403),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_251),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_227),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_81),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_128),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_0),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_347),
.Y(n_465)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_289),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_332),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_280),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_138),
.Y(n_469)
);

INVxp67_ASAP7_75t_SL g470 ( 
.A(n_190),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_218),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_358),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_9),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_143),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_146),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_380),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_7),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_57),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_44),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_341),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_202),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_229),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_192),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_25),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_277),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_212),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_25),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_283),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_180),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_343),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_326),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_176),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_298),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_46),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_5),
.Y(n_495)
);

BUFx2_ASAP7_75t_L g496 ( 
.A(n_33),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_220),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_340),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_322),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_193),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_155),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_196),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_171),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_266),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_320),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_390),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_97),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_352),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_96),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_372),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_395),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_400),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_257),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_130),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_312),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_371),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_150),
.Y(n_519)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_177),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_368),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_293),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_344),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_396),
.Y(n_524)
);

BUFx10_ASAP7_75t_L g525 ( 
.A(n_237),
.Y(n_525)
);

BUFx10_ASAP7_75t_L g526 ( 
.A(n_195),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_244),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_104),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_383),
.Y(n_529)
);

BUFx8_ASAP7_75t_SL g530 ( 
.A(n_200),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_21),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_389),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_279),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_342),
.Y(n_534)
);

BUFx3_ASAP7_75t_L g535 ( 
.A(n_178),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_6),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_31),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_99),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_363),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_19),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_88),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_348),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_294),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_346),
.Y(n_544)
);

BUFx10_ASAP7_75t_L g545 ( 
.A(n_338),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_198),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_26),
.Y(n_547)
);

CKINVDCx5p33_ASAP7_75t_R g548 ( 
.A(n_304),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_336),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_167),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_325),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_361),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_21),
.Y(n_553)
);

BUFx5_ASAP7_75t_L g554 ( 
.A(n_95),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_19),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_53),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_107),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_356),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_387),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_273),
.Y(n_560)
);

INVx2_ASAP7_75t_SL g561 ( 
.A(n_360),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_120),
.Y(n_562)
);

BUFx5_ASAP7_75t_L g563 ( 
.A(n_225),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_30),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g565 ( 
.A(n_115),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_13),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_375),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_73),
.Y(n_568)
);

CKINVDCx5p33_ASAP7_75t_R g569 ( 
.A(n_310),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_119),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_345),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_27),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_84),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_228),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_291),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_392),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_307),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_165),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_286),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_391),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_169),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_369),
.Y(n_582)
);

INVxp33_ASAP7_75t_L g583 ( 
.A(n_37),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_409),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_9),
.Y(n_585)
);

CKINVDCx5p33_ASAP7_75t_R g586 ( 
.A(n_393),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_152),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_408),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_238),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_324),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_88),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_309),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_367),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_284),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_36),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_50),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_239),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_203),
.Y(n_598)
);

BUFx3_ASAP7_75t_L g599 ( 
.A(n_104),
.Y(n_599)
);

CKINVDCx5p33_ASAP7_75t_R g600 ( 
.A(n_379),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_97),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_337),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_354),
.Y(n_603)
);

INVxp67_ASAP7_75t_L g604 ( 
.A(n_174),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_40),
.Y(n_605)
);

CKINVDCx5p33_ASAP7_75t_R g606 ( 
.A(n_191),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_316),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_17),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_394),
.Y(n_609)
);

CKINVDCx5p33_ASAP7_75t_R g610 ( 
.A(n_319),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_153),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_134),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_339),
.Y(n_613)
);

CKINVDCx5p33_ASAP7_75t_R g614 ( 
.A(n_137),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_99),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_131),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_82),
.Y(n_617)
);

INVx1_ASAP7_75t_SL g618 ( 
.A(n_311),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_133),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_351),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_208),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_69),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_140),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_269),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_87),
.Y(n_625)
);

CKINVDCx5p33_ASAP7_75t_R g626 ( 
.A(n_401),
.Y(n_626)
);

INVx1_ASAP7_75t_SL g627 ( 
.A(n_221),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_105),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_382),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_84),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_53),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_359),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_355),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_302),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_82),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_317),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_102),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_329),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_232),
.Y(n_639)
);

CKINVDCx5p33_ASAP7_75t_R g640 ( 
.A(n_385),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_386),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_235),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_303),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_321),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_323),
.Y(n_645)
);

CKINVDCx20_ASAP7_75t_R g646 ( 
.A(n_362),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_373),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_300),
.Y(n_648)
);

BUFx6f_ASAP7_75t_L g649 ( 
.A(n_350),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g650 ( 
.A(n_120),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_274),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_374),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_14),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_166),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_308),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_265),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_183),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_384),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_366),
.Y(n_659)
);

BUFx6f_ASAP7_75t_L g660 ( 
.A(n_290),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_399),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_164),
.Y(n_662)
);

BUFx2_ASAP7_75t_L g663 ( 
.A(n_365),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_80),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_127),
.Y(n_665)
);

CKINVDCx5p33_ASAP7_75t_R g666 ( 
.A(n_48),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_114),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_299),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_349),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_282),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_5),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_376),
.Y(n_672)
);

BUFx2_ASAP7_75t_L g673 ( 
.A(n_330),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_398),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_404),
.Y(n_675)
);

CKINVDCx20_ASAP7_75t_R g676 ( 
.A(n_240),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_364),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_199),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_297),
.Y(n_679)
);

CKINVDCx5p33_ASAP7_75t_R g680 ( 
.A(n_295),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_377),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_158),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_4),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_90),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_207),
.Y(n_685)
);

CKINVDCx14_ASAP7_75t_R g686 ( 
.A(n_23),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_55),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_296),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_59),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_45),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_249),
.Y(n_691)
);

CKINVDCx5p33_ASAP7_75t_R g692 ( 
.A(n_306),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_41),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_397),
.Y(n_694)
);

CKINVDCx20_ASAP7_75t_R g695 ( 
.A(n_83),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_406),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_162),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_334),
.Y(n_698)
);

BUFx3_ASAP7_75t_L g699 ( 
.A(n_121),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_402),
.Y(n_700)
);

CKINVDCx20_ASAP7_75t_R g701 ( 
.A(n_46),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_231),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_103),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_245),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_410),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_278),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_530),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_496),
.B(n_0),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_432),
.Y(n_709)
);

BUFx2_ASAP7_75t_SL g710 ( 
.A(n_423),
.Y(n_710)
);

CKINVDCx16_ASAP7_75t_R g711 ( 
.A(n_686),
.Y(n_711)
);

HB1xp67_ASAP7_75t_L g712 ( 
.A(n_540),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_458),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_439),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_520),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_529),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_499),
.Y(n_717)
);

CKINVDCx20_ASAP7_75t_R g718 ( 
.A(n_434),
.Y(n_718)
);

XOR2xp5_ASAP7_75t_L g719 ( 
.A(n_479),
.B(n_1),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_683),
.B(n_1),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_673),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_452),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_452),
.Y(n_724)
);

CKINVDCx20_ASAP7_75t_R g725 ( 
.A(n_565),
.Y(n_725)
);

CKINVDCx20_ASAP7_75t_R g726 ( 
.A(n_695),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_599),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_599),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_699),
.Y(n_729)
);

CKINVDCx5p33_ASAP7_75t_R g730 ( 
.A(n_467),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_701),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_472),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_567),
.Y(n_733)
);

HB1xp67_ASAP7_75t_L g734 ( 
.A(n_699),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_587),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_525),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_633),
.Y(n_737)
);

INVxp67_ASAP7_75t_SL g738 ( 
.A(n_583),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_646),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_554),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_554),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_658),
.Y(n_742)
);

CKINVDCx20_ASAP7_75t_R g743 ( 
.A(n_676),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_466),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_554),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_427),
.B(n_2),
.Y(n_746)
);

CKINVDCx16_ASAP7_75t_R g747 ( 
.A(n_525),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_411),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_554),
.Y(n_749)
);

INVxp67_ASAP7_75t_L g750 ( 
.A(n_412),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_554),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_554),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_415),
.Y(n_753)
);

CKINVDCx16_ASAP7_75t_R g754 ( 
.A(n_526),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_526),
.Y(n_755)
);

INVxp67_ASAP7_75t_SL g756 ( 
.A(n_650),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_420),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_429),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_446),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_431),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_448),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_464),
.Y(n_762)
);

CKINVDCx20_ASAP7_75t_R g763 ( 
.A(n_441),
.Y(n_763)
);

INVxp67_ASAP7_75t_SL g764 ( 
.A(n_473),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_494),
.Y(n_765)
);

INVxp67_ASAP7_75t_SL g766 ( 
.A(n_538),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_449),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_553),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_451),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_454),
.Y(n_770)
);

INVxp67_ASAP7_75t_SL g771 ( 
.A(n_555),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_L g772 ( 
.A(n_455),
.B(n_2),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_557),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_545),
.B(n_3),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_561),
.B(n_3),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_604),
.B(n_4),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_566),
.B(n_6),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_591),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_462),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_601),
.Y(n_780)
);

CKINVDCx20_ASAP7_75t_R g781 ( 
.A(n_477),
.Y(n_781)
);

CKINVDCx16_ASAP7_75t_R g782 ( 
.A(n_545),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_478),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_608),
.Y(n_784)
);

CKINVDCx16_ASAP7_75t_R g785 ( 
.A(n_491),
.Y(n_785)
);

BUFx10_ASAP7_75t_L g786 ( 
.A(n_418),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_491),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_622),
.B(n_8),
.Y(n_788)
);

NOR2xp67_ASAP7_75t_L g789 ( 
.A(n_625),
.B(n_8),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_563),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_498),
.B(n_10),
.Y(n_791)
);

CKINVDCx20_ASAP7_75t_R g792 ( 
.A(n_484),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_563),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_630),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_487),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_495),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_671),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_511),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_684),
.B(n_687),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_690),
.Y(n_800)
);

CKINVDCx20_ASAP7_75t_R g801 ( 
.A(n_528),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_537),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_541),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_417),
.B(n_10),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_547),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_693),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_417),
.B(n_11),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_584),
.B(n_11),
.Y(n_808)
);

CKINVDCx20_ASAP7_75t_R g809 ( 
.A(n_718),
.Y(n_809)
);

CKINVDCx20_ASAP7_75t_R g810 ( 
.A(n_718),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_713),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_734),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_723),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_741),
.Y(n_814)
);

INVx4_ASAP7_75t_L g815 ( 
.A(n_736),
.Y(n_815)
);

AND2x4_ASAP7_75t_L g816 ( 
.A(n_709),
.B(n_509),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_741),
.Y(n_817)
);

AND2x4_ASAP7_75t_L g818 ( 
.A(n_714),
.B(n_509),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_724),
.Y(n_819)
);

AND2x4_ASAP7_75t_L g820 ( 
.A(n_715),
.B(n_509),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_740),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_727),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_730),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_712),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_733),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_737),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_739),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_736),
.B(n_419),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_728),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_738),
.B(n_556),
.Y(n_830)
);

INVxp67_ASAP7_75t_L g831 ( 
.A(n_710),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_786),
.Y(n_832)
);

XNOR2xp5_ASAP7_75t_L g833 ( 
.A(n_725),
.B(n_562),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_729),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_745),
.Y(n_835)
);

HB1xp67_ASAP7_75t_L g836 ( 
.A(n_757),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_760),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_749),
.Y(n_838)
);

BUFx6f_ASAP7_75t_L g839 ( 
.A(n_790),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_751),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_752),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_790),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_756),
.A2(n_564),
.B1(n_570),
.B2(n_568),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_767),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_793),
.Y(n_845)
);

OA21x2_ASAP7_75t_L g846 ( 
.A1(n_793),
.A2(n_657),
.B(n_584),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_R g847 ( 
.A(n_707),
.B(n_413),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_753),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_758),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_716),
.B(n_572),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_742),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_732),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_735),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_759),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_743),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_807),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_786),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_748),
.Y(n_858)
);

NOR2xp67_ASAP7_75t_L g859 ( 
.A(n_761),
.B(n_414),
.Y(n_859)
);

AND2x6_ASAP7_75t_L g860 ( 
.A(n_774),
.B(n_508),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_762),
.Y(n_861)
);

CKINVDCx5p33_ASAP7_75t_R g862 ( 
.A(n_748),
.Y(n_862)
);

CKINVDCx20_ASAP7_75t_R g863 ( 
.A(n_726),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_765),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_768),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_785),
.B(n_416),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_781),
.Y(n_867)
);

BUFx6f_ASAP7_75t_L g868 ( 
.A(n_791),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_746),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_711),
.B(n_573),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_773),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_781),
.Y(n_872)
);

BUFx8_ASAP7_75t_L g873 ( 
.A(n_788),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_778),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_792),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_780),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_784),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_797),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_731),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_787),
.B(n_421),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_800),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_792),
.Y(n_882)
);

CKINVDCx16_ASAP7_75t_R g883 ( 
.A(n_747),
.Y(n_883)
);

BUFx6f_ASAP7_75t_L g884 ( 
.A(n_806),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_717),
.B(n_585),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_764),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_766),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_754),
.B(n_595),
.Y(n_888)
);

CKINVDCx5p33_ASAP7_75t_R g889 ( 
.A(n_763),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_799),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_795),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_769),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_721),
.B(n_596),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_R g894 ( 
.A(n_744),
.B(n_605),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_771),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_798),
.Y(n_896)
);

CKINVDCx5p33_ASAP7_75t_R g897 ( 
.A(n_801),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_722),
.B(n_424),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_720),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_803),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_770),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_772),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_779),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_783),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_750),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_796),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_802),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_772),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_775),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_805),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_775),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_755),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_794),
.Y(n_913)
);

AND2x4_ASAP7_75t_L g914 ( 
.A(n_777),
.B(n_789),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_782),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_804),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_804),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_719),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_808),
.Y(n_919)
);

OAI22xp5_ASAP7_75t_L g920 ( 
.A1(n_708),
.A2(n_615),
.B1(n_628),
.B2(n_617),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_776),
.B(n_631),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_776),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_808),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_734),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_734),
.Y(n_925)
);

AND2x4_ASAP7_75t_L g926 ( 
.A(n_709),
.B(n_509),
.Y(n_926)
);

AND3x1_ASAP7_75t_L g927 ( 
.A(n_774),
.B(n_435),
.C(n_426),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_741),
.Y(n_928)
);

INVx3_ASAP7_75t_L g929 ( 
.A(n_736),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_738),
.B(n_635),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_734),
.Y(n_931)
);

INVx6_ASAP7_75t_L g932 ( 
.A(n_786),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_713),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_741),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_741),
.Y(n_935)
);

INVx3_ASAP7_75t_L g936 ( 
.A(n_736),
.Y(n_936)
);

BUFx8_ASAP7_75t_L g937 ( 
.A(n_774),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_734),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_738),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_741),
.Y(n_940)
);

CKINVDCx20_ASAP7_75t_R g941 ( 
.A(n_718),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_734),
.Y(n_942)
);

OA21x2_ASAP7_75t_L g943 ( 
.A1(n_790),
.A2(n_675),
.B(n_657),
.Y(n_943)
);

OAI21x1_ASAP7_75t_L g944 ( 
.A1(n_790),
.A2(n_675),
.B(n_438),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_713),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_741),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_734),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_713),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_709),
.B(n_536),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_713),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_734),
.Y(n_951)
);

CKINVDCx20_ASAP7_75t_R g952 ( 
.A(n_718),
.Y(n_952)
);

BUFx10_ASAP7_75t_L g953 ( 
.A(n_744),
.Y(n_953)
);

AND2x4_ASAP7_75t_L g954 ( 
.A(n_709),
.B(n_536),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_734),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_741),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_741),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_741),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_734),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_734),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_R g961 ( 
.A(n_707),
.B(n_422),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_R g962 ( 
.A(n_707),
.B(n_425),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_718),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_712),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_734),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_734),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_785),
.B(n_428),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_741),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_816),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_932),
.Y(n_970)
);

BUFx6f_ASAP7_75t_L g971 ( 
.A(n_932),
.Y(n_971)
);

INVx5_ASAP7_75t_L g972 ( 
.A(n_884),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_890),
.B(n_430),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_884),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_889),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_L g976 ( 
.A(n_860),
.B(n_857),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_884),
.Y(n_977)
);

OR2x6_ASAP7_75t_L g978 ( 
.A(n_912),
.B(n_536),
.Y(n_978)
);

INVx4_ASAP7_75t_SL g979 ( 
.A(n_860),
.Y(n_979)
);

INVxp67_ASAP7_75t_SL g980 ( 
.A(n_824),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_891),
.Y(n_981)
);

INVx2_ASAP7_75t_L g982 ( 
.A(n_839),
.Y(n_982)
);

AND2x6_ASAP7_75t_L g983 ( 
.A(n_832),
.B(n_508),
.Y(n_983)
);

NOR2xp33_ASAP7_75t_L g984 ( 
.A(n_815),
.B(n_442),
.Y(n_984)
);

AND2x6_ASAP7_75t_L g985 ( 
.A(n_832),
.B(n_916),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_846),
.Y(n_986)
);

INVx3_ASAP7_75t_L g987 ( 
.A(n_816),
.Y(n_987)
);

OAI22xp33_ASAP7_75t_L g988 ( 
.A1(n_964),
.A2(n_637),
.B1(n_666),
.B2(n_664),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_846),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_943),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_815),
.B(n_500),
.Y(n_991)
);

INVx4_ASAP7_75t_L g992 ( 
.A(n_881),
.Y(n_992)
);

AND2x2_ASAP7_75t_L g993 ( 
.A(n_905),
.B(n_667),
.Y(n_993)
);

AOI22xp33_ASAP7_75t_L g994 ( 
.A1(n_902),
.A2(n_536),
.B1(n_436),
.B2(n_460),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_913),
.B(n_437),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_818),
.Y(n_996)
);

OR2x6_ASAP7_75t_L g997 ( 
.A(n_836),
.B(n_450),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_818),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_839),
.Y(n_999)
);

INVx2_ASAP7_75t_L g1000 ( 
.A(n_839),
.Y(n_1000)
);

AND2x6_ASAP7_75t_L g1001 ( 
.A(n_917),
.B(n_535),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_820),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_845),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_820),
.Y(n_1004)
);

INVx6_ASAP7_75t_L g1005 ( 
.A(n_953),
.Y(n_1005)
);

NAND2xp5_ASAP7_75t_L g1006 ( 
.A(n_881),
.B(n_440),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_926),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_926),
.Y(n_1008)
);

NOR2xp33_ASAP7_75t_L g1009 ( 
.A(n_939),
.B(n_543),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_869),
.Y(n_1010)
);

INVxp67_ASAP7_75t_SL g1011 ( 
.A(n_856),
.Y(n_1011)
);

INVx5_ASAP7_75t_L g1012 ( 
.A(n_860),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_845),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_929),
.B(n_618),
.Y(n_1014)
);

CKINVDCx5p33_ASAP7_75t_R g1015 ( 
.A(n_896),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_868),
.B(n_443),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_929),
.B(n_620),
.Y(n_1017)
);

INVx4_ASAP7_75t_SL g1018 ( 
.A(n_860),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_949),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_L g1020 ( 
.A(n_812),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_868),
.B(n_444),
.Y(n_1021)
);

INVx1_ASAP7_75t_L g1022 ( 
.A(n_949),
.Y(n_1022)
);

INVx5_ASAP7_75t_L g1023 ( 
.A(n_845),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_888),
.B(n_689),
.Y(n_1024)
);

BUFx6f_ASAP7_75t_L g1025 ( 
.A(n_856),
.Y(n_1025)
);

AND2x6_ASAP7_75t_L g1026 ( 
.A(n_919),
.B(n_535),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_868),
.B(n_445),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_954),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_856),
.B(n_447),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_936),
.B(n_531),
.Y(n_1030)
);

AND2x2_ASAP7_75t_L g1031 ( 
.A(n_843),
.B(n_703),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_869),
.B(n_453),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_944),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_935),
.Y(n_1034)
);

OR2x2_ASAP7_75t_L g1035 ( 
.A(n_883),
.B(n_653),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_935),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_869),
.B(n_456),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_922),
.B(n_457),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_943),
.Y(n_1039)
);

AND2x6_ASAP7_75t_L g1040 ( 
.A(n_908),
.B(n_463),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_954),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_901),
.Y(n_1042)
);

BUFx6f_ASAP7_75t_L g1043 ( 
.A(n_953),
.Y(n_1043)
);

INVx3_ASAP7_75t_L g1044 ( 
.A(n_936),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_897),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_899),
.B(n_470),
.Y(n_1046)
);

AO22x2_ASAP7_75t_L g1047 ( 
.A1(n_924),
.A2(n_476),
.B1(n_481),
.B2(n_468),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_813),
.Y(n_1048)
);

AO21x2_ASAP7_75t_L g1049 ( 
.A1(n_909),
.A2(n_483),
.B(n_482),
.Y(n_1049)
);

INVx2_ASAP7_75t_L g1050 ( 
.A(n_935),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_819),
.Y(n_1051)
);

OR2x2_ASAP7_75t_L g1052 ( 
.A(n_925),
.B(n_12),
.Y(n_1052)
);

HB1xp67_ASAP7_75t_L g1053 ( 
.A(n_837),
.Y(n_1053)
);

NOR2xp33_ASAP7_75t_L g1054 ( 
.A(n_911),
.B(n_627),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_923),
.B(n_459),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_822),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_829),
.Y(n_1057)
);

NOR2xp33_ASAP7_75t_L g1058 ( 
.A(n_886),
.B(n_632),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_834),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_914),
.B(n_486),
.Y(n_1060)
);

BUFx2_ASAP7_75t_L g1061 ( 
.A(n_903),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_830),
.B(n_461),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_914),
.Y(n_1063)
);

OR2x6_ASAP7_75t_L g1064 ( 
.A(n_844),
.B(n_488),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_864),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_871),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_843),
.B(n_706),
.Y(n_1067)
);

INVx4_ASAP7_75t_L g1068 ( 
.A(n_904),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_874),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_906),
.Y(n_1070)
);

INVx5_ASAP7_75t_L g1071 ( 
.A(n_842),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_907),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_848),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_910),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_870),
.Y(n_1075)
);

NOR2xp33_ASAP7_75t_L g1076 ( 
.A(n_887),
.B(n_465),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_849),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_931),
.B(n_938),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_854),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_942),
.B(n_469),
.Y(n_1080)
);

INVx1_ASAP7_75t_SL g1081 ( 
.A(n_892),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_915),
.Y(n_1082)
);

NAND3x1_ASAP7_75t_L g1083 ( 
.A(n_863),
.B(n_501),
.C(n_497),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_921),
.B(n_471),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_937),
.Y(n_1085)
);

INVxp67_ASAP7_75t_SL g1086 ( 
.A(n_831),
.Y(n_1086)
);

AOI22xp33_ASAP7_75t_L g1087 ( 
.A1(n_895),
.A2(n_506),
.B1(n_512),
.B2(n_503),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_861),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_930),
.B(n_474),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_865),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_SL g1091 ( 
.A(n_927),
.B(n_475),
.Y(n_1091)
);

BUFx6f_ASAP7_75t_L g1092 ( 
.A(n_876),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_877),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_885),
.B(n_480),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_947),
.B(n_517),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_878),
.B(n_485),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_828),
.Y(n_1097)
);

AND2x4_ASAP7_75t_L g1098 ( 
.A(n_951),
.B(n_955),
.Y(n_1098)
);

INVx2_ASAP7_75t_L g1099 ( 
.A(n_814),
.Y(n_1099)
);

AND2x4_ASAP7_75t_L g1100 ( 
.A(n_959),
.B(n_518),
.Y(n_1100)
);

BUFx4f_ASAP7_75t_L g1101 ( 
.A(n_960),
.Y(n_1101)
);

HB1xp67_ASAP7_75t_L g1102 ( 
.A(n_900),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_965),
.B(n_966),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_817),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_850),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_859),
.B(n_489),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_928),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_893),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_L g1109 ( 
.A(n_866),
.B(n_880),
.Y(n_1109)
);

INVx2_ASAP7_75t_L g1110 ( 
.A(n_934),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_967),
.B(n_490),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_859),
.B(n_492),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_898),
.Y(n_1113)
);

NOR2x1_ASAP7_75t_L g1114 ( 
.A(n_920),
.B(n_521),
.Y(n_1114)
);

INVx4_ASAP7_75t_L g1115 ( 
.A(n_821),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_SL g1116 ( 
.A(n_927),
.B(n_493),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_968),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_847),
.B(n_505),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_838),
.B(n_524),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_858),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_840),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_841),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_940),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_835),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_937),
.B(n_507),
.Y(n_1125)
);

INVx2_ASAP7_75t_SL g1126 ( 
.A(n_873),
.Y(n_1126)
);

INVx2_ASAP7_75t_SL g1127 ( 
.A(n_873),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_946),
.Y(n_1128)
);

NOR2xp67_ASAP7_75t_L g1129 ( 
.A(n_811),
.B(n_12),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_L g1130 ( 
.A(n_823),
.B(n_510),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_825),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_956),
.Y(n_1132)
);

NAND3xp33_ASAP7_75t_SL g1133 ( 
.A(n_826),
.B(n_514),
.C(n_513),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_957),
.B(n_516),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_958),
.Y(n_1135)
);

CKINVDCx20_ASAP7_75t_R g1136 ( 
.A(n_809),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_961),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_962),
.Y(n_1138)
);

INVx2_ASAP7_75t_L g1139 ( 
.A(n_827),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_879),
.Y(n_1140)
);

BUFx3_ASAP7_75t_L g1141 ( 
.A(n_851),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_933),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_862),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_945),
.Y(n_1144)
);

INVx1_ASAP7_75t_SL g1145 ( 
.A(n_867),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_948),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_950),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_872),
.B(n_519),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_875),
.Y(n_1149)
);

INVx4_ASAP7_75t_L g1150 ( 
.A(n_882),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_833),
.B(n_852),
.Y(n_1151)
);

AND2x6_ASAP7_75t_L g1152 ( 
.A(n_894),
.B(n_539),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_853),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_855),
.B(n_522),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_810),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_918),
.B(n_523),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_941),
.Y(n_1157)
);

BUFx4f_ASAP7_75t_L g1158 ( 
.A(n_952),
.Y(n_1158)
);

INVx5_ASAP7_75t_L g1159 ( 
.A(n_963),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_927),
.A2(n_558),
.B1(n_571),
.B2(n_546),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_884),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_832),
.B(n_527),
.Y(n_1162)
);

INVx4_ASAP7_75t_L g1163 ( 
.A(n_932),
.Y(n_1163)
);

INVx8_ASAP7_75t_L g1164 ( 
.A(n_860),
.Y(n_1164)
);

INVx3_ASAP7_75t_L g1165 ( 
.A(n_932),
.Y(n_1165)
);

AND2x2_ASAP7_75t_SL g1166 ( 
.A(n_883),
.B(n_575),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_932),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_832),
.B(n_532),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_815),
.B(n_533),
.Y(n_1169)
);

NOR2xp33_ASAP7_75t_L g1170 ( 
.A(n_815),
.B(n_534),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_890),
.B(n_542),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_932),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_932),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_824),
.B(n_544),
.Y(n_1174)
);

OR2x6_ASAP7_75t_L g1175 ( 
.A(n_912),
.B(n_577),
.Y(n_1175)
);

BUFx6f_ASAP7_75t_L g1176 ( 
.A(n_932),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_890),
.B(n_548),
.Y(n_1177)
);

OAI221xp5_ASAP7_75t_L g1178 ( 
.A1(n_843),
.A2(n_582),
.B1(n_588),
.B2(n_579),
.C(n_578),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_932),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_884),
.Y(n_1180)
);

CKINVDCx6p67_ASAP7_75t_R g1181 ( 
.A(n_883),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_890),
.B(n_549),
.Y(n_1182)
);

AND2x2_ASAP7_75t_SL g1183 ( 
.A(n_883),
.B(n_592),
.Y(n_1183)
);

INVx3_ASAP7_75t_L g1184 ( 
.A(n_932),
.Y(n_1184)
);

INVx2_ASAP7_75t_L g1185 ( 
.A(n_884),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_R g1186 ( 
.A(n_915),
.B(n_550),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_846),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_832),
.B(n_551),
.Y(n_1188)
);

NOR2xp33_ASAP7_75t_SL g1189 ( 
.A(n_901),
.B(n_552),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_846),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_884),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_846),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_832),
.B(n_559),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_890),
.B(n_560),
.Y(n_1194)
);

AND2x6_ASAP7_75t_L g1195 ( 
.A(n_832),
.B(n_602),
.Y(n_1195)
);

INVx4_ASAP7_75t_L g1196 ( 
.A(n_932),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_815),
.B(n_569),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_884),
.Y(n_1198)
);

AND2x4_ASAP7_75t_L g1199 ( 
.A(n_832),
.B(n_616),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_L g1200 ( 
.A1(n_1105),
.A2(n_623),
.B1(n_639),
.B2(n_624),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1090),
.B(n_574),
.Y(n_1201)
);

NOR2xp33_ASAP7_75t_L g1202 ( 
.A(n_980),
.B(n_576),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1025),
.Y(n_1203)
);

INVx2_ASAP7_75t_L g1204 ( 
.A(n_1025),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1081),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_L g1206 ( 
.A(n_1108),
.B(n_580),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1113),
.B(n_581),
.Y(n_1207)
);

NAND2x1_ASAP7_75t_L g1208 ( 
.A(n_992),
.B(n_433),
.Y(n_1208)
);

OAI22xp33_ASAP7_75t_L g1209 ( 
.A1(n_1061),
.A2(n_589),
.B1(n_590),
.B2(n_586),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1119),
.B(n_593),
.Y(n_1210)
);

NOR2xp67_ASAP7_75t_SL g1211 ( 
.A(n_1043),
.B(n_594),
.Y(n_1211)
);

CKINVDCx20_ASAP7_75t_R g1212 ( 
.A(n_1181),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1093),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1119),
.B(n_597),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_992),
.B(n_1189),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_L g1216 ( 
.A1(n_1098),
.A2(n_648),
.B1(n_655),
.B2(n_652),
.Y(n_1216)
);

INVx2_ASAP7_75t_SL g1217 ( 
.A(n_978),
.Y(n_1217)
);

NAND2xp5_ASAP7_75t_L g1218 ( 
.A(n_1097),
.B(n_598),
.Y(n_1218)
);

NOR2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1068),
.B(n_1085),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1093),
.B(n_600),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1078),
.B(n_603),
.Y(n_1221)
);

BUFx3_ASAP7_75t_L g1222 ( 
.A(n_1005),
.Y(n_1222)
);

NOR2xp67_ASAP7_75t_L g1223 ( 
.A(n_1012),
.B(n_122),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1088),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_SL g1225 ( 
.A1(n_1054),
.A2(n_705),
.B(n_662),
.C(n_669),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1088),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1115),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1047),
.A2(n_659),
.B1(n_679),
.B2(n_670),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1040),
.B(n_1092),
.Y(n_1229)
);

OR2x6_ASAP7_75t_L g1230 ( 
.A(n_1005),
.B(n_681),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1040),
.B(n_606),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1040),
.B(n_607),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1073),
.Y(n_1233)
);

NAND2x1p5_ASAP7_75t_L g1234 ( 
.A(n_1043),
.B(n_682),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1077),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_978),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1053),
.B(n_13),
.Y(n_1237)
);

OAI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1115),
.A2(n_691),
.B1(n_704),
.B2(n_688),
.Y(n_1238)
);

AOI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_986),
.A2(n_610),
.B(n_609),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1098),
.A2(n_563),
.B1(n_612),
.B2(n_611),
.Y(n_1240)
);

NOR2xp67_ASAP7_75t_L g1241 ( 
.A(n_1012),
.B(n_123),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1095),
.A2(n_563),
.B1(n_614),
.B2(n_613),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_SL g1243 ( 
.A(n_1092),
.B(n_619),
.Y(n_1243)
);

NAND2xp5_ASAP7_75t_L g1244 ( 
.A(n_1095),
.B(n_621),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1100),
.B(n_626),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1121),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_1061),
.Y(n_1247)
);

AOI22xp5_ASAP7_75t_L g1248 ( 
.A1(n_1047),
.A2(n_1122),
.B1(n_1049),
.B2(n_1056),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_SL g1249 ( 
.A(n_1012),
.B(n_702),
.Y(n_1249)
);

A2O1A1Ixp33_ASAP7_75t_SL g1250 ( 
.A1(n_1094),
.A2(n_1089),
.B(n_1017),
.C(n_1014),
.Y(n_1250)
);

INVx2_ASAP7_75t_L g1251 ( 
.A(n_1069),
.Y(n_1251)
);

NOR2xp33_ASAP7_75t_SL g1252 ( 
.A(n_1068),
.B(n_629),
.Y(n_1252)
);

NAND2x1_ASAP7_75t_L g1253 ( 
.A(n_985),
.B(n_433),
.Y(n_1253)
);

AOI22xp5_ASAP7_75t_L g1254 ( 
.A1(n_1048),
.A2(n_1059),
.B1(n_1079),
.B2(n_1100),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_993),
.B(n_634),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1069),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1163),
.B(n_16),
.Y(n_1257)
);

INVx2_ASAP7_75t_SL g1258 ( 
.A(n_971),
.Y(n_1258)
);

AOI22xp5_ASAP7_75t_L g1259 ( 
.A1(n_1103),
.A2(n_563),
.B1(n_638),
.B2(n_636),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1063),
.B(n_640),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1199),
.B(n_641),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1199),
.B(n_642),
.Y(n_1262)
);

INVxp67_ASAP7_75t_L g1263 ( 
.A(n_1175),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1145),
.B(n_1035),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1195),
.B(n_1114),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1195),
.B(n_643),
.Y(n_1266)
);

AND2x2_ASAP7_75t_L g1267 ( 
.A(n_1031),
.B(n_16),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1195),
.B(n_1065),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_987),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_996),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1007),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_SL g1272 ( 
.A(n_1020),
.B(n_700),
.Y(n_1272)
);

NOR2xp33_ASAP7_75t_SL g1273 ( 
.A(n_1042),
.B(n_644),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1066),
.B(n_645),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1051),
.B(n_647),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1057),
.B(n_651),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1117),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_969),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1178),
.A2(n_563),
.B1(n_656),
.B2(n_654),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1101),
.B(n_698),
.Y(n_1280)
);

AOI22xp5_ASAP7_75t_L g1281 ( 
.A1(n_1160),
.A2(n_665),
.B1(n_668),
.B2(n_661),
.Y(n_1281)
);

INVx2_ASAP7_75t_SL g1282 ( 
.A(n_971),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1063),
.B(n_672),
.Y(n_1283)
);

AOI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1067),
.A2(n_677),
.B1(n_680),
.B2(n_674),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1174),
.B(n_685),
.Y(n_1285)
);

INVx3_ASAP7_75t_L g1286 ( 
.A(n_1071),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_997),
.B(n_17),
.Y(n_1287)
);

NOR2x2_ASAP7_75t_L g1288 ( 
.A(n_1175),
.B(n_18),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1046),
.A2(n_694),
.B1(n_696),
.B2(n_692),
.Y(n_1289)
);

NOR2x2_ASAP7_75t_L g1290 ( 
.A(n_997),
.B(n_18),
.Y(n_1290)
);

INVx2_ASAP7_75t_SL g1291 ( 
.A(n_1176),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1024),
.B(n_697),
.Y(n_1292)
);

INVx1_ASAP7_75t_SL g1293 ( 
.A(n_970),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1117),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1080),
.B(n_20),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_998),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_SL g1297 ( 
.A(n_1176),
.B(n_433),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1058),
.B(n_20),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1009),
.B(n_22),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1010),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_L g1301 ( 
.A(n_1109),
.B(n_22),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1124),
.Y(n_1302)
);

OAI221xp5_ASAP7_75t_L g1303 ( 
.A1(n_1087),
.A2(n_504),
.B1(n_515),
.B2(n_502),
.C(n_433),
.Y(n_1303)
);

NOR2xp33_ASAP7_75t_L g1304 ( 
.A(n_1086),
.B(n_1148),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_973),
.B(n_23),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1002),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1171),
.B(n_24),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_986),
.A2(n_504),
.B(n_502),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_989),
.A2(n_504),
.B(n_502),
.Y(n_1309)
);

NAND2x1_ASAP7_75t_L g1310 ( 
.A(n_985),
.B(n_502),
.Y(n_1310)
);

AND2x2_ASAP7_75t_SL g1311 ( 
.A(n_1158),
.B(n_504),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_989),
.A2(n_649),
.B(n_515),
.Y(n_1312)
);

AND2x4_ASAP7_75t_L g1313 ( 
.A(n_1163),
.B(n_24),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_990),
.A2(n_1187),
.B(n_1039),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_SL g1315 ( 
.A(n_1070),
.B(n_515),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1177),
.B(n_26),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_L g1317 ( 
.A(n_1182),
.B(n_27),
.Y(n_1317)
);

NAND2x1_ASAP7_75t_L g1318 ( 
.A(n_985),
.B(n_515),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1011),
.A2(n_660),
.B1(n_678),
.B2(n_649),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1099),
.Y(n_1320)
);

INVx2_ASAP7_75t_SL g1321 ( 
.A(n_1173),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1194),
.B(n_28),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1104),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1196),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1004),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1046),
.A2(n_1116),
.B1(n_1091),
.B2(n_1060),
.Y(n_1326)
);

NOR2xp33_ASAP7_75t_L g1327 ( 
.A(n_1196),
.B(n_28),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1030),
.B(n_29),
.Y(n_1328)
);

BUFx8_ASAP7_75t_L g1329 ( 
.A(n_1126),
.Y(n_1329)
);

NAND2xp5_ASAP7_75t_L g1330 ( 
.A(n_1030),
.B(n_30),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1082),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_990),
.A2(n_1187),
.B(n_1039),
.Y(n_1332)
);

BUFx3_ASAP7_75t_L g1333 ( 
.A(n_1072),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1107),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1075),
.B(n_31),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1060),
.B(n_32),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1008),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1110),
.Y(n_1338)
);

NAND2xp5_ASAP7_75t_L g1339 ( 
.A(n_1076),
.B(n_32),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1019),
.Y(n_1340)
);

OR2x2_ASAP7_75t_L g1341 ( 
.A(n_1157),
.B(n_33),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_SL g1342 ( 
.A1(n_1166),
.A2(n_660),
.B1(n_678),
.B2(n_649),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1064),
.B(n_1141),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_SL g1344 ( 
.A(n_1071),
.B(n_1169),
.Y(n_1344)
);

BUFx6f_ASAP7_75t_L g1345 ( 
.A(n_1164),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1022),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_SL g1347 ( 
.A(n_1071),
.B(n_649),
.Y(n_1347)
);

A2O1A1Ixp33_ASAP7_75t_L g1348 ( 
.A1(n_1190),
.A2(n_678),
.B(n_660),
.C(n_36),
.Y(n_1348)
);

AND2x6_ASAP7_75t_L g1349 ( 
.A(n_1190),
.B(n_1192),
.Y(n_1349)
);

OAI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1064),
.A2(n_678),
.B1(n_660),
.B2(n_37),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_L g1351 ( 
.A(n_984),
.B(n_34),
.Y(n_1351)
);

NOR2xp33_ASAP7_75t_L g1352 ( 
.A(n_1075),
.B(n_34),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1123),
.Y(n_1353)
);

NOR2xp33_ASAP7_75t_L g1354 ( 
.A(n_1154),
.B(n_35),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_SL g1355 ( 
.A(n_1170),
.B(n_38),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1052),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1356)
);

NAND2xp33_ASAP7_75t_L g1357 ( 
.A(n_1164),
.B(n_124),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1028),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1137),
.B(n_39),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1072),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_991),
.B(n_41),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1062),
.B(n_42),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1128),
.A2(n_45),
.B1(n_43),
.B2(n_44),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1001),
.B(n_1026),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_SL g1365 ( 
.A(n_1197),
.B(n_47),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_988),
.B(n_979),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1192),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1132),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1001),
.B(n_49),
.Y(n_1369)
);

O2A1O1Ixp5_ASAP7_75t_L g1370 ( 
.A1(n_1106),
.A2(n_126),
.B(n_129),
.C(n_125),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1041),
.A2(n_52),
.B1(n_50),
.B2(n_51),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1135),
.Y(n_1372)
);

AOI22xp5_ASAP7_75t_L g1373 ( 
.A1(n_1152),
.A2(n_55),
.B1(n_52),
.B2(n_54),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1152),
.A2(n_1001),
.B1(n_1026),
.B2(n_983),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1044),
.Y(n_1375)
);

A2O1A1Ixp33_ASAP7_75t_SL g1376 ( 
.A1(n_1111),
.A2(n_135),
.B(n_136),
.C(n_132),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1029),
.Y(n_1377)
);

CKINVDCx11_ASAP7_75t_R g1378 ( 
.A(n_1136),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1026),
.B(n_983),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_974),
.Y(n_1380)
);

AND2x2_ASAP7_75t_L g1381 ( 
.A(n_1137),
.B(n_56),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1033),
.A2(n_142),
.B(n_139),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_979),
.B(n_56),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_983),
.B(n_57),
.Y(n_1384)
);

INVx3_ASAP7_75t_L g1385 ( 
.A(n_972),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_977),
.Y(n_1386)
);

INVx4_ASAP7_75t_L g1387 ( 
.A(n_1018),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1096),
.B(n_58),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1161),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1016),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_994),
.A2(n_61),
.B1(n_58),
.B2(n_60),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1006),
.B(n_60),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1021),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1254),
.B(n_1233),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1213),
.Y(n_1395)
);

INVx5_ASAP7_75t_L g1396 ( 
.A(n_1230),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1205),
.Y(n_1397)
);

NOR3xp33_ASAP7_75t_SL g1398 ( 
.A(n_1209),
.B(n_981),
.C(n_975),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1235),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1378),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1254),
.B(n_1152),
.Y(n_1401)
);

INVxp67_ASAP7_75t_SL g1402 ( 
.A(n_1329),
.Y(n_1402)
);

OR2x6_ASAP7_75t_L g1403 ( 
.A(n_1230),
.B(n_1127),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1264),
.B(n_1155),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1219),
.B(n_1018),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_SL g1406 ( 
.A(n_1252),
.B(n_1074),
.Y(n_1406)
);

BUFx8_ASAP7_75t_SL g1407 ( 
.A(n_1212),
.Y(n_1407)
);

INVx3_ASAP7_75t_L g1408 ( 
.A(n_1387),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1246),
.B(n_1074),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1302),
.Y(n_1410)
);

HB1xp67_ASAP7_75t_L g1411 ( 
.A(n_1247),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1368),
.Y(n_1412)
);

AND2x4_ASAP7_75t_L g1413 ( 
.A(n_1230),
.B(n_1167),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1329),
.Y(n_1414)
);

INVx2_ASAP7_75t_L g1415 ( 
.A(n_1372),
.Y(n_1415)
);

INVx3_ASAP7_75t_L g1416 ( 
.A(n_1387),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1278),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1296),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1222),
.Y(n_1419)
);

AND2x2_ASAP7_75t_L g1420 ( 
.A(n_1287),
.B(n_1183),
.Y(n_1420)
);

AND2x4_ASAP7_75t_L g1421 ( 
.A(n_1377),
.B(n_1172),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1267),
.B(n_1131),
.Y(n_1422)
);

INVxp33_ASAP7_75t_L g1423 ( 
.A(n_1343),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_1306),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1304),
.B(n_1139),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1221),
.B(n_1156),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1331),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1320),
.Y(n_1428)
);

CKINVDCx20_ASAP7_75t_R g1429 ( 
.A(n_1333),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1227),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1248),
.B(n_1142),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_1360),
.Y(n_1432)
);

HB1xp67_ASAP7_75t_L g1433 ( 
.A(n_1263),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_SL g1434 ( 
.A(n_1273),
.B(n_1150),
.Y(n_1434)
);

BUFx3_ASAP7_75t_L g1435 ( 
.A(n_1321),
.Y(n_1435)
);

HB1xp67_ASAP7_75t_L g1436 ( 
.A(n_1257),
.Y(n_1436)
);

INVx5_ASAP7_75t_L g1437 ( 
.A(n_1345),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1325),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_1311),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1257),
.Y(n_1440)
);

CKINVDCx5p33_ASAP7_75t_R g1441 ( 
.A(n_1293),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1337),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_R g1443 ( 
.A(n_1315),
.B(n_1140),
.Y(n_1443)
);

INVx3_ASAP7_75t_L g1444 ( 
.A(n_1227),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1340),
.Y(n_1445)
);

NOR3xp33_ASAP7_75t_SL g1446 ( 
.A(n_1335),
.B(n_1045),
.C(n_1015),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1323),
.Y(n_1447)
);

INVx3_ASAP7_75t_L g1448 ( 
.A(n_1345),
.Y(n_1448)
);

AND2x4_ASAP7_75t_SL g1449 ( 
.A(n_1313),
.B(n_1150),
.Y(n_1449)
);

O2A1O1Ixp33_ASAP7_75t_L g1450 ( 
.A1(n_1225),
.A2(n_1120),
.B(n_1102),
.C(n_1144),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1345),
.Y(n_1451)
);

INVx3_ASAP7_75t_L g1452 ( 
.A(n_1385),
.Y(n_1452)
);

BUFx12f_ASAP7_75t_L g1453 ( 
.A(n_1341),
.Y(n_1453)
);

NAND2xp5_ASAP7_75t_L g1454 ( 
.A(n_1248),
.B(n_1146),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1390),
.B(n_1165),
.Y(n_1455)
);

BUFx4f_ASAP7_75t_L g1456 ( 
.A(n_1217),
.Y(n_1456)
);

INVx2_ASAP7_75t_L g1457 ( 
.A(n_1334),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1237),
.B(n_1130),
.Y(n_1458)
);

INVx3_ASAP7_75t_L g1459 ( 
.A(n_1385),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_1313),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1346),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1338),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1284),
.B(n_1153),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1228),
.B(n_1147),
.Y(n_1464)
);

A2O1A1Ixp33_ASAP7_75t_L g1465 ( 
.A1(n_1301),
.A2(n_976),
.B(n_1129),
.C(n_1112),
.Y(n_1465)
);

INVx5_ASAP7_75t_L g1466 ( 
.A(n_1349),
.Y(n_1466)
);

AND2x6_ASAP7_75t_L g1467 ( 
.A(n_1229),
.B(n_1138),
.Y(n_1467)
);

AND2x4_ASAP7_75t_L g1468 ( 
.A(n_1393),
.B(n_1179),
.Y(n_1468)
);

AOI21xp5_ASAP7_75t_L g1469 ( 
.A1(n_1314),
.A2(n_1033),
.B(n_1134),
.Y(n_1469)
);

INVx1_ASAP7_75t_SL g1470 ( 
.A(n_1359),
.Y(n_1470)
);

BUFx2_ASAP7_75t_L g1471 ( 
.A(n_1236),
.Y(n_1471)
);

AND2x2_ASAP7_75t_L g1472 ( 
.A(n_1228),
.B(n_1184),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1200),
.B(n_995),
.Y(n_1473)
);

CKINVDCx20_ASAP7_75t_R g1474 ( 
.A(n_1258),
.Y(n_1474)
);

OAI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1363),
.A2(n_1159),
.B1(n_1143),
.B2(n_1149),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1326),
.B(n_1084),
.Y(n_1476)
);

AND2x4_ASAP7_75t_L g1477 ( 
.A(n_1375),
.B(n_1032),
.Y(n_1477)
);

BUFx6f_ASAP7_75t_L g1478 ( 
.A(n_1349),
.Y(n_1478)
);

INVx3_ASAP7_75t_L g1479 ( 
.A(n_1286),
.Y(n_1479)
);

INVx2_ASAP7_75t_L g1480 ( 
.A(n_1353),
.Y(n_1480)
);

INVx3_ASAP7_75t_L g1481 ( 
.A(n_1286),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1358),
.Y(n_1482)
);

NOR3xp33_ASAP7_75t_SL g1483 ( 
.A(n_1352),
.B(n_1186),
.C(n_1133),
.Y(n_1483)
);

AND2x4_ASAP7_75t_SL g1484 ( 
.A(n_1374),
.B(n_1324),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_SL g1485 ( 
.A(n_1202),
.B(n_1159),
.Y(n_1485)
);

AO22x1_ASAP7_75t_L g1486 ( 
.A1(n_1290),
.A2(n_1159),
.B1(n_1151),
.B2(n_1125),
.Y(n_1486)
);

BUFx10_ASAP7_75t_L g1487 ( 
.A(n_1327),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1366),
.B(n_1162),
.Y(n_1488)
);

BUFx3_ASAP7_75t_L g1489 ( 
.A(n_1282),
.Y(n_1489)
);

INVx1_ASAP7_75t_SL g1490 ( 
.A(n_1381),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1332),
.Y(n_1491)
);

INVx2_ASAP7_75t_SL g1492 ( 
.A(n_1234),
.Y(n_1492)
);

BUFx10_ASAP7_75t_L g1493 ( 
.A(n_1291),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1300),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1328),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1292),
.B(n_1055),
.Y(n_1496)
);

BUFx2_ASAP7_75t_L g1497 ( 
.A(n_1288),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1330),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1336),
.B(n_1083),
.Y(n_1499)
);

NOR3xp33_ASAP7_75t_SL g1500 ( 
.A(n_1238),
.B(n_1118),
.C(n_1272),
.Y(n_1500)
);

HB1xp67_ASAP7_75t_L g1501 ( 
.A(n_1268),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1269),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1215),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1384),
.Y(n_1504)
);

BUFx3_ASAP7_75t_L g1505 ( 
.A(n_1251),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1342),
.B(n_1037),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1349),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1270),
.Y(n_1508)
);

INVx3_ASAP7_75t_L g1509 ( 
.A(n_1224),
.Y(n_1509)
);

NAND2xp5_ASAP7_75t_L g1510 ( 
.A(n_1206),
.B(n_1038),
.Y(n_1510)
);

BUFx2_ASAP7_75t_L g1511 ( 
.A(n_1349),
.Y(n_1511)
);

BUFx12f_ASAP7_75t_L g1512 ( 
.A(n_1211),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1281),
.B(n_1027),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1271),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1216),
.B(n_1168),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1363),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1392),
.Y(n_1517)
);

INVx4_ASAP7_75t_L g1518 ( 
.A(n_1226),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1203),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1204),
.Y(n_1520)
);

BUFx2_ASAP7_75t_L g1521 ( 
.A(n_1369),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1305),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_R g1523 ( 
.A(n_1364),
.B(n_61),
.Y(n_1523)
);

INVx4_ASAP7_75t_L g1524 ( 
.A(n_1256),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1295),
.B(n_1188),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1265),
.B(n_1193),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1307),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1316),
.Y(n_1528)
);

BUFx6f_ASAP7_75t_L g1529 ( 
.A(n_1253),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1380),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1386),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1281),
.A2(n_1180),
.B1(n_1191),
.B2(n_1185),
.Y(n_1532)
);

BUFx12f_ASAP7_75t_L g1533 ( 
.A(n_1350),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1389),
.Y(n_1534)
);

INVx3_ASAP7_75t_L g1535 ( 
.A(n_1277),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1201),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1294),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1208),
.Y(n_1538)
);

BUFx2_ASAP7_75t_L g1539 ( 
.A(n_1261),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1279),
.B(n_972),
.Y(n_1540)
);

INVxp67_ASAP7_75t_L g1541 ( 
.A(n_1244),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1207),
.B(n_972),
.Y(n_1542)
);

OAI21x1_ASAP7_75t_L g1543 ( 
.A1(n_1469),
.A2(n_1309),
.B(n_1308),
.Y(n_1543)
);

AOI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1465),
.A2(n_1250),
.B(n_1312),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_1410),
.Y(n_1545)
);

OA21x2_ASAP7_75t_L g1546 ( 
.A1(n_1491),
.A2(n_1348),
.B(n_1370),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1491),
.A2(n_1319),
.B(n_1382),
.Y(n_1547)
);

OAI21x1_ASAP7_75t_L g1548 ( 
.A1(n_1538),
.A2(n_1318),
.B(n_1310),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1516),
.B(n_1255),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1399),
.Y(n_1550)
);

INVx8_ASAP7_75t_L g1551 ( 
.A(n_1407),
.Y(n_1551)
);

A2O1A1Ixp33_ASAP7_75t_L g1552 ( 
.A1(n_1522),
.A2(n_1354),
.B(n_1362),
.C(n_1317),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1429),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1210),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1399),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1464),
.B(n_1214),
.Y(n_1556)
);

O2A1O1Ixp5_ASAP7_75t_L g1557 ( 
.A1(n_1506),
.A2(n_1355),
.B(n_1365),
.C(n_1344),
.Y(n_1557)
);

AOI21xp5_ASAP7_75t_L g1558 ( 
.A1(n_1522),
.A2(n_1357),
.B(n_1322),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1527),
.A2(n_1376),
.B(n_1388),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1397),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_SL g1561 ( 
.A(n_1396),
.B(n_1439),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1527),
.A2(n_1361),
.B(n_1351),
.Y(n_1562)
);

OAI21x1_ASAP7_75t_L g1563 ( 
.A1(n_1535),
.A2(n_1241),
.B(n_1223),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1394),
.B(n_1426),
.Y(n_1564)
);

AO31x2_ASAP7_75t_L g1565 ( 
.A1(n_1431),
.A2(n_1367),
.A3(n_1391),
.B(n_1371),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1395),
.B(n_1245),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1528),
.A2(n_1339),
.B(n_1299),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1414),
.Y(n_1568)
);

NAND2xp5_ASAP7_75t_L g1569 ( 
.A(n_1395),
.B(n_1259),
.Y(n_1569)
);

NAND2x1p5_ASAP7_75t_L g1570 ( 
.A(n_1396),
.B(n_1023),
.Y(n_1570)
);

NOR2xp67_ASAP7_75t_SL g1571 ( 
.A(n_1396),
.B(n_1379),
.Y(n_1571)
);

AO31x2_ASAP7_75t_L g1572 ( 
.A1(n_1454),
.A2(n_1298),
.A3(n_1239),
.B(n_1198),
.Y(n_1572)
);

OAI22xp5_ASAP7_75t_L g1573 ( 
.A1(n_1440),
.A2(n_1470),
.B1(n_1490),
.B2(n_1436),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1528),
.A2(n_1517),
.B(n_1473),
.Y(n_1574)
);

NOR2xp33_ASAP7_75t_L g1575 ( 
.A(n_1475),
.B(n_1285),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1460),
.A2(n_1356),
.B1(n_1259),
.B2(n_1373),
.Y(n_1576)
);

OA21x2_ASAP7_75t_L g1577 ( 
.A1(n_1517),
.A2(n_1319),
.B(n_1303),
.Y(n_1577)
);

OAI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1425),
.A2(n_1218),
.B(n_1220),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1472),
.B(n_1262),
.Y(n_1579)
);

OAI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1535),
.A2(n_1241),
.B(n_1223),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1525),
.A2(n_1383),
.B(n_1274),
.Y(n_1581)
);

NAND2x1_ASAP7_75t_L g1582 ( 
.A(n_1507),
.B(n_982),
.Y(n_1582)
);

BUFx2_ASAP7_75t_L g1583 ( 
.A(n_1403),
.Y(n_1583)
);

INVx2_ASAP7_75t_L g1584 ( 
.A(n_1415),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1513),
.B(n_1242),
.Y(n_1585)
);

AO21x1_ASAP7_75t_L g1586 ( 
.A1(n_1401),
.A2(n_1347),
.B(n_1297),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1509),
.A2(n_1000),
.B(n_999),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1412),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1420),
.B(n_1289),
.Y(n_1589)
);

AO31x2_ASAP7_75t_L g1590 ( 
.A1(n_1495),
.A2(n_1013),
.A3(n_1034),
.B(n_1003),
.Y(n_1590)
);

AOI21x1_ASAP7_75t_SL g1591 ( 
.A1(n_1540),
.A2(n_1476),
.B(n_1488),
.Y(n_1591)
);

INVxp67_ASAP7_75t_SL g1592 ( 
.A(n_1411),
.Y(n_1592)
);

AND2x4_ASAP7_75t_L g1593 ( 
.A(n_1405),
.B(n_1243),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1510),
.A2(n_1542),
.B(n_1515),
.Y(n_1594)
);

AOI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1511),
.A2(n_1249),
.B(n_1275),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1536),
.B(n_1260),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_L g1597 ( 
.A1(n_1498),
.A2(n_1276),
.B(n_1232),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1417),
.Y(n_1598)
);

INVx3_ASAP7_75t_L g1599 ( 
.A(n_1451),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1409),
.B(n_1283),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1509),
.A2(n_1050),
.B(n_1036),
.Y(n_1601)
);

NAND2xp5_ASAP7_75t_SL g1602 ( 
.A(n_1443),
.B(n_1231),
.Y(n_1602)
);

OAI21x1_ASAP7_75t_L g1603 ( 
.A1(n_1479),
.A2(n_1266),
.B(n_1240),
.Y(n_1603)
);

OAI21x1_ASAP7_75t_L g1604 ( 
.A1(n_1479),
.A2(n_1280),
.B(n_1023),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1418),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1424),
.B(n_1023),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1450),
.A2(n_145),
.B(n_144),
.Y(n_1607)
);

AOI21xp33_ASAP7_75t_L g1608 ( 
.A1(n_1463),
.A2(n_62),
.B(n_63),
.Y(n_1608)
);

INVx3_ASAP7_75t_L g1609 ( 
.A(n_1451),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1438),
.B(n_62),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1405),
.B(n_63),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1451),
.Y(n_1612)
);

AOI22xp5_ASAP7_75t_L g1613 ( 
.A1(n_1404),
.A2(n_66),
.B1(n_64),
.B2(n_65),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1481),
.A2(n_148),
.B(n_147),
.Y(n_1614)
);

OAI21x1_ASAP7_75t_L g1615 ( 
.A1(n_1481),
.A2(n_151),
.B(n_149),
.Y(n_1615)
);

AOI21xp5_ASAP7_75t_L g1616 ( 
.A1(n_1488),
.A2(n_156),
.B(n_154),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1519),
.A2(n_160),
.B(n_159),
.Y(n_1617)
);

AOI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1530),
.A2(n_163),
.B(n_161),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1403),
.B(n_1441),
.Y(n_1619)
);

OAI21x1_ASAP7_75t_L g1620 ( 
.A1(n_1520),
.A2(n_172),
.B(n_168),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1442),
.B(n_64),
.Y(n_1621)
);

OAI21x1_ASAP7_75t_L g1622 ( 
.A1(n_1452),
.A2(n_175),
.B(n_173),
.Y(n_1622)
);

OAI21x1_ASAP7_75t_L g1623 ( 
.A1(n_1452),
.A2(n_181),
.B(n_179),
.Y(n_1623)
);

INVx4_ASAP7_75t_L g1624 ( 
.A(n_1437),
.Y(n_1624)
);

AO31x2_ASAP7_75t_L g1625 ( 
.A1(n_1507),
.A2(n_68),
.A3(n_66),
.B(n_67),
.Y(n_1625)
);

AOI211x1_ASAP7_75t_L g1626 ( 
.A1(n_1486),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1626)
);

O2A1O1Ixp5_ASAP7_75t_L g1627 ( 
.A1(n_1485),
.A2(n_184),
.B(n_186),
.C(n_182),
.Y(n_1627)
);

OAI21x1_ASAP7_75t_L g1628 ( 
.A1(n_1459),
.A2(n_188),
.B(n_187),
.Y(n_1628)
);

INVx2_ASAP7_75t_SL g1629 ( 
.A(n_1437),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1402),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_SL g1631 ( 
.A(n_1413),
.B(n_70),
.Y(n_1631)
);

OAI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1541),
.A2(n_70),
.B(n_71),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1445),
.B(n_72),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_L g1634 ( 
.A(n_1461),
.B(n_72),
.Y(n_1634)
);

AOI22xp5_ASAP7_75t_L g1635 ( 
.A1(n_1575),
.A2(n_1533),
.B1(n_1458),
.B2(n_1422),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1598),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1598),
.Y(n_1637)
);

NAND2x1p5_ASAP7_75t_L g1638 ( 
.A(n_1624),
.B(n_1437),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1545),
.Y(n_1639)
);

AO31x2_ASAP7_75t_L g1640 ( 
.A1(n_1544),
.A2(n_1534),
.A3(n_1531),
.B(n_1447),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1605),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1559),
.A2(n_1543),
.B(n_1563),
.Y(n_1642)
);

OAI21x1_ASAP7_75t_L g1643 ( 
.A1(n_1591),
.A2(n_1459),
.B(n_1444),
.Y(n_1643)
);

INVx3_ASAP7_75t_SL g1644 ( 
.A(n_1551),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1580),
.A2(n_1601),
.B(n_1587),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1605),
.Y(n_1646)
);

OAI21x1_ASAP7_75t_L g1647 ( 
.A1(n_1617),
.A2(n_1444),
.B(n_1430),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1624),
.B(n_1466),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1584),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1589),
.B(n_1409),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1560),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_L g1652 ( 
.A1(n_1576),
.A2(n_1497),
.B1(n_1499),
.B2(n_1539),
.Y(n_1652)
);

AOI21xp5_ASAP7_75t_L g1653 ( 
.A1(n_1558),
.A2(n_1466),
.B(n_1478),
.Y(n_1653)
);

OA21x2_ASAP7_75t_L g1654 ( 
.A1(n_1562),
.A2(n_1532),
.B(n_1537),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1550),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1656)
);

OAI21x1_ASAP7_75t_SL g1657 ( 
.A1(n_1632),
.A2(n_1492),
.B(n_1466),
.Y(n_1657)
);

BUFx3_ASAP7_75t_L g1658 ( 
.A(n_1568),
.Y(n_1658)
);

AOI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1564),
.A2(n_1482),
.B1(n_1496),
.B2(n_1423),
.C(n_1421),
.Y(n_1659)
);

OAI21x1_ASAP7_75t_L g1660 ( 
.A1(n_1620),
.A2(n_1430),
.B(n_1416),
.Y(n_1660)
);

HB1xp67_ASAP7_75t_L g1661 ( 
.A(n_1592),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1551),
.Y(n_1662)
);

OAI21x1_ASAP7_75t_L g1663 ( 
.A1(n_1614),
.A2(n_1416),
.B(n_1408),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1588),
.Y(n_1664)
);

OAI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1594),
.A2(n_1500),
.B(n_1504),
.Y(n_1665)
);

NOR2xp33_ASAP7_75t_L g1666 ( 
.A(n_1630),
.B(n_1453),
.Y(n_1666)
);

OAI22xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1583),
.A2(n_1400),
.B1(n_1499),
.B2(n_1474),
.Y(n_1667)
);

O2A1O1Ixp33_ASAP7_75t_SL g1668 ( 
.A1(n_1608),
.A2(n_1434),
.B(n_1406),
.C(n_1503),
.Y(n_1668)
);

OAI22xp33_ASAP7_75t_L g1669 ( 
.A1(n_1613),
.A2(n_1523),
.B1(n_1478),
.B2(n_1521),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1615),
.A2(n_1408),
.B(n_1428),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1610),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1622),
.A2(n_1462),
.B(n_1457),
.Y(n_1672)
);

OAI21x1_ASAP7_75t_SL g1673 ( 
.A1(n_1569),
.A2(n_1518),
.B(n_1524),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1570),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1552),
.A2(n_1526),
.B(n_1483),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1629),
.B(n_1456),
.Y(n_1676)
);

OAI21x1_ASAP7_75t_L g1677 ( 
.A1(n_1623),
.A2(n_1480),
.B(n_1448),
.Y(n_1677)
);

CKINVDCx20_ASAP7_75t_R g1678 ( 
.A(n_1553),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1619),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1621),
.Y(n_1680)
);

OAI21xp5_ASAP7_75t_L g1681 ( 
.A1(n_1556),
.A2(n_1526),
.B(n_1508),
.Y(n_1681)
);

BUFx10_ASAP7_75t_L g1682 ( 
.A(n_1611),
.Y(n_1682)
);

OAI21x1_ASAP7_75t_L g1683 ( 
.A1(n_1628),
.A2(n_1448),
.B(n_1494),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1554),
.B(n_1501),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1664),
.Y(n_1685)
);

CKINVDCx8_ASAP7_75t_R g1686 ( 
.A(n_1674),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1636),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1639),
.Y(n_1688)
);

AOI22xp33_ASAP7_75t_L g1689 ( 
.A1(n_1659),
.A2(n_1585),
.B1(n_1579),
.B2(n_1549),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1650),
.B(n_1611),
.Y(n_1690)
);

OAI22xp33_ASAP7_75t_L g1691 ( 
.A1(n_1635),
.A2(n_1661),
.B1(n_1684),
.B2(n_1659),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1637),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1641),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1661),
.B(n_1573),
.Y(n_1694)
);

AOI22xp33_ASAP7_75t_SL g1695 ( 
.A1(n_1682),
.A2(n_1449),
.B1(n_1596),
.B2(n_1413),
.Y(n_1695)
);

AOI21xp5_ASAP7_75t_L g1696 ( 
.A1(n_1653),
.A2(n_1607),
.B(n_1567),
.Y(n_1696)
);

INVx2_ASAP7_75t_L g1697 ( 
.A(n_1649),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1646),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1655),
.Y(n_1699)
);

CKINVDCx11_ASAP7_75t_R g1700 ( 
.A(n_1644),
.Y(n_1700)
);

NAND2xp33_ASAP7_75t_R g1701 ( 
.A(n_1679),
.B(n_1398),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1651),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1651),
.B(n_1600),
.Y(n_1703)
);

AND2x2_ASAP7_75t_SL g1704 ( 
.A(n_1648),
.B(n_1478),
.Y(n_1704)
);

AO31x2_ASAP7_75t_L g1705 ( 
.A1(n_1656),
.A2(n_1586),
.A3(n_1581),
.B(n_1616),
.Y(n_1705)
);

OAI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1684),
.A2(n_1631),
.B1(n_1634),
.B2(n_1633),
.Y(n_1706)
);

OAI211xp5_ASAP7_75t_L g1707 ( 
.A1(n_1652),
.A2(n_1626),
.B(n_1446),
.C(n_1602),
.Y(n_1707)
);

AOI22xp33_ASAP7_75t_L g1708 ( 
.A1(n_1675),
.A2(n_1578),
.B1(n_1566),
.B2(n_1577),
.Y(n_1708)
);

AOI22xp33_ASAP7_75t_L g1709 ( 
.A1(n_1675),
.A2(n_1577),
.B1(n_1487),
.B2(n_1597),
.Y(n_1709)
);

AOI22xp33_ASAP7_75t_L g1710 ( 
.A1(n_1671),
.A2(n_1487),
.B1(n_1467),
.B2(n_1561),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1656),
.Y(n_1711)
);

AND2x4_ASAP7_75t_L g1712 ( 
.A(n_1648),
.B(n_1599),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1640),
.Y(n_1713)
);

OAI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1669),
.A2(n_1606),
.B1(n_1512),
.B2(n_1456),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1682),
.B(n_73),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1680),
.Y(n_1716)
);

AOI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1665),
.A2(n_1557),
.B(n_1571),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1638),
.B(n_74),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1681),
.Y(n_1719)
);

AO31x2_ASAP7_75t_L g1720 ( 
.A1(n_1696),
.A2(n_1713),
.A3(n_1719),
.B(n_1711),
.Y(n_1720)
);

OAI22xp5_ASAP7_75t_L g1721 ( 
.A1(n_1691),
.A2(n_1665),
.B1(n_1681),
.B2(n_1638),
.Y(n_1721)
);

OAI211xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1707),
.A2(n_1666),
.B(n_1427),
.C(n_1433),
.Y(n_1722)
);

OAI211xp5_ASAP7_75t_L g1723 ( 
.A1(n_1695),
.A2(n_1668),
.B(n_1658),
.C(n_1662),
.Y(n_1723)
);

AO21x2_ASAP7_75t_L g1724 ( 
.A1(n_1717),
.A2(n_1706),
.B(n_1691),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1703),
.B(n_1625),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1685),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1706),
.A2(n_1421),
.B1(n_1468),
.B2(n_1455),
.C(n_1502),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_L g1728 ( 
.A1(n_1714),
.A2(n_1467),
.B1(n_1657),
.B2(n_1667),
.Y(n_1728)
);

AOI222xp33_ASAP7_75t_L g1729 ( 
.A1(n_1689),
.A2(n_1593),
.B1(n_1678),
.B2(n_1471),
.C1(n_1477),
.C2(n_1468),
.Y(n_1729)
);

BUFx6f_ASAP7_75t_L g1730 ( 
.A(n_1686),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1689),
.A2(n_1676),
.B1(n_1674),
.B2(n_1653),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1714),
.A2(n_1690),
.B1(n_1694),
.B2(n_1718),
.Y(n_1732)
);

AOI21xp33_ASAP7_75t_SL g1733 ( 
.A1(n_1701),
.A2(n_1676),
.B(n_1432),
.Y(n_1733)
);

AO21x2_ASAP7_75t_L g1734 ( 
.A1(n_1702),
.A2(n_1673),
.B(n_1670),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1716),
.B(n_1625),
.Y(n_1735)
);

BUFx2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1699),
.Y(n_1737)
);

AOI222xp33_ASAP7_75t_L g1738 ( 
.A1(n_1700),
.A2(n_1593),
.B1(n_1477),
.B2(n_1455),
.C1(n_1514),
.C2(n_1484),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1688),
.B(n_1697),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1687),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1692),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1693),
.B(n_1625),
.Y(n_1742)
);

OR2x2_ASAP7_75t_L g1743 ( 
.A(n_1698),
.B(n_1674),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1708),
.B(n_1565),
.Y(n_1744)
);

AOI21xp33_ASAP7_75t_L g1745 ( 
.A1(n_1708),
.A2(n_1642),
.B(n_1654),
.Y(n_1745)
);

AND2x4_ASAP7_75t_L g1746 ( 
.A(n_1712),
.B(n_1643),
.Y(n_1746)
);

INVxp67_ASAP7_75t_SL g1747 ( 
.A(n_1709),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1715),
.Y(n_1748)
);

AOI22xp33_ASAP7_75t_L g1749 ( 
.A1(n_1709),
.A2(n_1467),
.B1(n_1654),
.B2(n_1603),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1739),
.B(n_1710),
.Y(n_1750)
);

INVx3_ASAP7_75t_L g1751 ( 
.A(n_1746),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1725),
.B(n_1710),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1726),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1746),
.B(n_1705),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1720),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1737),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1741),
.B(n_1705),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1720),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1736),
.B(n_1704),
.Y(n_1759)
);

INVxp67_ASAP7_75t_SL g1760 ( 
.A(n_1743),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1740),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1742),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1730),
.Y(n_1763)
);

AOI22xp33_ASAP7_75t_L g1764 ( 
.A1(n_1729),
.A2(n_1695),
.B1(n_1704),
.B2(n_1467),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1735),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1748),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1730),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1744),
.B(n_1705),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1720),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1734),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1724),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1724),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1721),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1753),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1760),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1763),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1756),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1764),
.A2(n_1732),
.B1(n_1728),
.B2(n_1730),
.Y(n_1778)
);

AOI22xp5_ASAP7_75t_L g1779 ( 
.A1(n_1773),
.A2(n_1721),
.B1(n_1722),
.B2(n_1729),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1764),
.A2(n_1723),
.B1(n_1747),
.B2(n_1738),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1760),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1757),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1769),
.Y(n_1783)
);

INVx3_ASAP7_75t_L g1784 ( 
.A(n_1751),
.Y(n_1784)
);

AOI22xp33_ASAP7_75t_L g1785 ( 
.A1(n_1766),
.A2(n_1727),
.B1(n_1738),
.B2(n_1731),
.Y(n_1785)
);

NAND4xp25_ASAP7_75t_SL g1786 ( 
.A(n_1759),
.B(n_1733),
.C(n_1749),
.D(n_1745),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1751),
.B(n_1734),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1762),
.B(n_1731),
.Y(n_1788)
);

INVxp67_ASAP7_75t_SL g1789 ( 
.A(n_1755),
.Y(n_1789)
);

OAI31xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1771),
.A2(n_1745),
.A3(n_1663),
.B(n_1683),
.Y(n_1790)
);

OR2x2_ASAP7_75t_L g1791 ( 
.A(n_1781),
.B(n_1768),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1774),
.Y(n_1792)
);

CKINVDCx16_ASAP7_75t_R g1793 ( 
.A(n_1776),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1775),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1781),
.B(n_1765),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1784),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1782),
.Y(n_1797)
);

INVx2_ASAP7_75t_SL g1798 ( 
.A(n_1784),
.Y(n_1798)
);

HB1xp67_ASAP7_75t_L g1799 ( 
.A(n_1782),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1788),
.B(n_1754),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1787),
.B(n_1754),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1777),
.B(n_1761),
.Y(n_1802)
);

INVx1_ASAP7_75t_SL g1803 ( 
.A(n_1778),
.Y(n_1803)
);

AND2x4_ASAP7_75t_SL g1804 ( 
.A(n_1785),
.B(n_1763),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1779),
.B(n_1772),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1783),
.B(n_1752),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1783),
.B(n_1750),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1789),
.B(n_1754),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1789),
.B(n_1755),
.Y(n_1809)
);

NOR2x1_ASAP7_75t_L g1810 ( 
.A(n_1786),
.B(n_1770),
.Y(n_1810)
);

INVx2_ASAP7_75t_L g1811 ( 
.A(n_1780),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1801),
.B(n_1790),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1795),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1801),
.B(n_1767),
.Y(n_1814)
);

OAI21xp5_ASAP7_75t_L g1815 ( 
.A1(n_1803),
.A2(n_1785),
.B(n_1767),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1802),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1800),
.B(n_1770),
.Y(n_1817)
);

NAND2xp33_ASAP7_75t_L g1818 ( 
.A(n_1794),
.B(n_1419),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_L g1819 ( 
.A(n_1813),
.B(n_1811),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1818),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1815),
.A2(n_1811),
.B1(n_1804),
.B2(n_1805),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1818),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1819),
.B(n_1816),
.Y(n_1823)
);

NAND4xp75_ASAP7_75t_L g1824 ( 
.A(n_1820),
.B(n_1810),
.C(n_1812),
.D(n_1808),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1823),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1824),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1824),
.A2(n_1821),
.B1(n_1822),
.B2(n_1812),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1824),
.B(n_1793),
.Y(n_1828)
);

INVx1_ASAP7_75t_L g1829 ( 
.A(n_1825),
.Y(n_1829)
);

INVxp67_ASAP7_75t_L g1830 ( 
.A(n_1826),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1827),
.Y(n_1831)
);

O2A1O1Ixp33_ASAP7_75t_L g1832 ( 
.A1(n_1828),
.A2(n_1794),
.B(n_1435),
.C(n_1798),
.Y(n_1832)
);

NAND3xp33_ASAP7_75t_SL g1833 ( 
.A(n_1826),
.B(n_1791),
.C(n_1808),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1828),
.B(n_1794),
.Y(n_1834)
);

INVx1_ASAP7_75t_L g1835 ( 
.A(n_1825),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1829),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1835),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_L g1838 ( 
.A1(n_1831),
.A2(n_1798),
.B1(n_1796),
.B2(n_1791),
.C(n_1809),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_L g1839 ( 
.A(n_1830),
.B(n_1489),
.C(n_1809),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_SL g1840 ( 
.A(n_1832),
.B(n_1804),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1833),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1834),
.B(n_1814),
.C(n_1796),
.D(n_1800),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1831),
.B(n_1817),
.Y(n_1843)
);

NOR2x1_ASAP7_75t_L g1844 ( 
.A(n_1831),
.B(n_1796),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1831),
.B(n_1814),
.Y(n_1845)
);

NAND3xp33_ASAP7_75t_SL g1846 ( 
.A(n_1830),
.B(n_1806),
.C(n_1807),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1829),
.Y(n_1847)
);

BUFx2_ASAP7_75t_L g1848 ( 
.A(n_1844),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1836),
.Y(n_1849)
);

INVxp67_ASAP7_75t_L g1850 ( 
.A(n_1837),
.Y(n_1850)
);

O2A1O1Ixp33_ASAP7_75t_L g1851 ( 
.A1(n_1847),
.A2(n_1799),
.B(n_1627),
.C(n_1792),
.Y(n_1851)
);

O2A1O1Ixp33_ASAP7_75t_L g1852 ( 
.A1(n_1841),
.A2(n_1797),
.B(n_1599),
.C(n_1612),
.Y(n_1852)
);

AOI22xp5_ASAP7_75t_L g1853 ( 
.A1(n_1845),
.A2(n_1797),
.B1(n_1758),
.B2(n_1493),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_SL g1854 ( 
.A1(n_1838),
.A2(n_76),
.B(n_74),
.C(n_75),
.Y(n_1854)
);

OAI21xp5_ASAP7_75t_SL g1855 ( 
.A1(n_1843),
.A2(n_1612),
.B(n_1609),
.Y(n_1855)
);

AOI211x1_ASAP7_75t_SL g1856 ( 
.A1(n_1839),
.A2(n_1758),
.B(n_77),
.C(n_75),
.Y(n_1856)
);

AOI211x1_ASAP7_75t_L g1857 ( 
.A1(n_1840),
.A2(n_1595),
.B(n_1618),
.C(n_78),
.Y(n_1857)
);

OAI21xp5_ASAP7_75t_SL g1858 ( 
.A1(n_1846),
.A2(n_1609),
.B(n_76),
.Y(n_1858)
);

OAI221xp5_ASAP7_75t_L g1859 ( 
.A1(n_1842),
.A2(n_1582),
.B1(n_78),
.B2(n_79),
.C(n_80),
.Y(n_1859)
);

AOI21xp33_ASAP7_75t_L g1860 ( 
.A1(n_1847),
.A2(n_77),
.B(n_79),
.Y(n_1860)
);

NAND4xp75_ASAP7_75t_L g1861 ( 
.A(n_1844),
.B(n_85),
.C(n_81),
.D(n_83),
.Y(n_1861)
);

NAND4xp25_ASAP7_75t_L g1862 ( 
.A(n_1845),
.B(n_87),
.C(n_85),
.D(n_86),
.Y(n_1862)
);

AOI221xp5_ASAP7_75t_L g1863 ( 
.A1(n_1841),
.A2(n_1505),
.B1(n_1518),
.B2(n_1524),
.C(n_91),
.Y(n_1863)
);

AOI221xp5_ASAP7_75t_L g1864 ( 
.A1(n_1841),
.A2(n_86),
.B1(n_89),
.B2(n_90),
.C(n_91),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1861),
.Y(n_1865)
);

INVxp67_ASAP7_75t_L g1866 ( 
.A(n_1848),
.Y(n_1866)
);

HB1xp67_ASAP7_75t_L g1867 ( 
.A(n_1850),
.Y(n_1867)
);

AOI32xp33_ASAP7_75t_L g1868 ( 
.A1(n_1854),
.A2(n_1604),
.A3(n_1493),
.B1(n_1660),
.B2(n_1677),
.Y(n_1868)
);

AOI221xp5_ASAP7_75t_L g1869 ( 
.A1(n_1857),
.A2(n_89),
.B1(n_92),
.B2(n_93),
.C(n_94),
.Y(n_1869)
);

OAI21xp5_ASAP7_75t_L g1870 ( 
.A1(n_1858),
.A2(n_1672),
.B(n_1548),
.Y(n_1870)
);

AOI221xp5_ASAP7_75t_L g1871 ( 
.A1(n_1863),
.A2(n_92),
.B1(n_93),
.B2(n_94),
.C(n_95),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1856),
.B(n_96),
.Y(n_1872)
);

XOR2xp5_ASAP7_75t_L g1873 ( 
.A(n_1862),
.B(n_98),
.Y(n_1873)
);

XNOR2x1_ASAP7_75t_L g1874 ( 
.A(n_1849),
.B(n_98),
.Y(n_1874)
);

INVx2_ASAP7_75t_SL g1875 ( 
.A(n_1853),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1860),
.B(n_100),
.Y(n_1876)
);

AOI222xp33_ASAP7_75t_L g1877 ( 
.A1(n_1859),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.C1(n_103),
.C2(n_105),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1852),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1864),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1855),
.B(n_101),
.Y(n_1880)
);

AOI221xp5_ASAP7_75t_L g1881 ( 
.A1(n_1851),
.A2(n_106),
.B1(n_107),
.B2(n_108),
.C(n_109),
.Y(n_1881)
);

NAND4xp75_ASAP7_75t_L g1882 ( 
.A(n_1865),
.B(n_106),
.C(n_108),
.D(n_109),
.Y(n_1882)
);

HB1xp67_ASAP7_75t_L g1883 ( 
.A(n_1866),
.Y(n_1883)
);

AND3x1_ASAP7_75t_L g1884 ( 
.A(n_1880),
.B(n_110),
.C(n_111),
.Y(n_1884)
);

NAND3xp33_ASAP7_75t_SL g1885 ( 
.A(n_1877),
.B(n_110),
.C(n_111),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1875),
.Y(n_1886)
);

AOI221xp5_ASAP7_75t_L g1887 ( 
.A1(n_1869),
.A2(n_112),
.B1(n_113),
.B2(n_114),
.C(n_115),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1874),
.B(n_113),
.Y(n_1888)
);

NOR3xp33_ASAP7_75t_L g1889 ( 
.A(n_1867),
.B(n_116),
.C(n_117),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1873),
.A2(n_1642),
.B1(n_1546),
.B2(n_1547),
.Y(n_1890)
);

OR2x2_ASAP7_75t_L g1891 ( 
.A(n_1872),
.B(n_116),
.Y(n_1891)
);

NAND2xp33_ASAP7_75t_SL g1892 ( 
.A(n_1879),
.B(n_117),
.Y(n_1892)
);

AND2x4_ASAP7_75t_SL g1893 ( 
.A(n_1876),
.B(n_1529),
.Y(n_1893)
);

OAI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1881),
.A2(n_118),
.B(n_119),
.Y(n_1894)
);

AND2x2_ASAP7_75t_SL g1895 ( 
.A(n_1871),
.B(n_1529),
.Y(n_1895)
);

NOR3xp33_ASAP7_75t_L g1896 ( 
.A(n_1878),
.B(n_118),
.C(n_121),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1870),
.B(n_1529),
.Y(n_1897)
);

INVxp67_ASAP7_75t_L g1898 ( 
.A(n_1868),
.Y(n_1898)
);

NAND3xp33_ASAP7_75t_L g1899 ( 
.A(n_1866),
.B(n_1547),
.C(n_1546),
.Y(n_1899)
);

NAND3xp33_ASAP7_75t_SL g1900 ( 
.A(n_1889),
.B(n_189),
.C(n_194),
.Y(n_1900)
);

AOI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1885),
.A2(n_197),
.B(n_204),
.C(n_205),
.Y(n_1901)
);

OAI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1886),
.A2(n_1705),
.B1(n_1565),
.B2(n_1572),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1883),
.B(n_1882),
.Y(n_1903)
);

AOI22xp33_ASAP7_75t_L g1904 ( 
.A1(n_1892),
.A2(n_1647),
.B1(n_1645),
.B2(n_1565),
.Y(n_1904)
);

AND4x2_ASAP7_75t_L g1905 ( 
.A(n_1888),
.B(n_1887),
.C(n_1884),
.D(n_1897),
.Y(n_1905)
);

OR3x1_ASAP7_75t_L g1906 ( 
.A(n_1894),
.B(n_210),
.C(n_211),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1891),
.Y(n_1907)
);

OAI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1898),
.A2(n_1572),
.B1(n_1640),
.B2(n_1590),
.Y(n_1908)
);

OR3x2_ASAP7_75t_L g1909 ( 
.A(n_1896),
.B(n_213),
.C(n_215),
.Y(n_1909)
);

OAI211xp5_ASAP7_75t_SL g1910 ( 
.A1(n_1895),
.A2(n_216),
.B(n_217),
.C(n_219),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1893),
.B(n_1640),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1899),
.A2(n_222),
.B(n_224),
.Y(n_1912)
);

NOR2x1_ASAP7_75t_L g1913 ( 
.A(n_1903),
.B(n_1906),
.Y(n_1913)
);

CKINVDCx20_ASAP7_75t_R g1914 ( 
.A(n_1907),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1905),
.Y(n_1915)
);

BUFx2_ASAP7_75t_SL g1916 ( 
.A(n_1901),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1911),
.Y(n_1917)
);

CKINVDCx20_ASAP7_75t_R g1918 ( 
.A(n_1900),
.Y(n_1918)
);

NAND4xp25_ASAP7_75t_L g1919 ( 
.A(n_1910),
.B(n_1890),
.C(n_230),
.D(n_234),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1912),
.B(n_226),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1908),
.B(n_236),
.Y(n_1921)
);

AOI221xp5_ASAP7_75t_SL g1922 ( 
.A1(n_1909),
.A2(n_1572),
.B1(n_1590),
.B2(n_246),
.C(n_247),
.Y(n_1922)
);

XNOR2xp5_ASAP7_75t_L g1923 ( 
.A(n_1913),
.B(n_1902),
.Y(n_1923)
);

BUFx2_ASAP7_75t_L g1924 ( 
.A(n_1914),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1919),
.A2(n_1904),
.B1(n_243),
.B2(n_250),
.C(n_252),
.Y(n_1925)
);

HB1xp67_ASAP7_75t_L g1926 ( 
.A(n_1915),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1917),
.Y(n_1927)
);

AND2x2_ASAP7_75t_L g1928 ( 
.A(n_1916),
.B(n_242),
.Y(n_1928)
);

NAND3xp33_ASAP7_75t_L g1929 ( 
.A(n_1920),
.B(n_253),
.C(n_254),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1918),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1927),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1930),
.A2(n_1922),
.B1(n_1921),
.B2(n_1590),
.Y(n_1932)
);

OAI22xp5_ASAP7_75t_L g1933 ( 
.A1(n_1926),
.A2(n_255),
.B1(n_256),
.B2(n_259),
.Y(n_1933)
);

INVx1_ASAP7_75t_L g1934 ( 
.A(n_1924),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1931),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1934),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1932),
.Y(n_1937)
);

XNOR2xp5_ASAP7_75t_L g1938 ( 
.A(n_1936),
.B(n_1925),
.Y(n_1938)
);

NAND2xp5_ASAP7_75t_SL g1939 ( 
.A(n_1935),
.B(n_1923),
.Y(n_1939)
);

OAI21xp5_ASAP7_75t_SL g1940 ( 
.A1(n_1938),
.A2(n_1928),
.B(n_1937),
.Y(n_1940)
);

AOI22xp5_ASAP7_75t_L g1941 ( 
.A1(n_1939),
.A2(n_1929),
.B1(n_1933),
.B2(n_264),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1938),
.Y(n_1942)
);

AOI222xp33_ASAP7_75t_L g1943 ( 
.A1(n_1942),
.A2(n_1940),
.B1(n_1941),
.B2(n_267),
.C1(n_270),
.C2(n_271),
.Y(n_1943)
);

AOI22xp33_ASAP7_75t_L g1944 ( 
.A1(n_1942),
.A2(n_261),
.B1(n_262),
.B2(n_272),
.Y(n_1944)
);

OAI221xp5_ASAP7_75t_L g1945 ( 
.A1(n_1943),
.A2(n_275),
.B1(n_276),
.B2(n_281),
.C(n_285),
.Y(n_1945)
);

AOI211xp5_ASAP7_75t_L g1946 ( 
.A1(n_1945),
.A2(n_1944),
.B(n_287),
.C(n_288),
.Y(n_1946)
);


endmodule