module fake_netlist_6_1582_n_2012 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2012);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2012;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1413;
wire n_1330;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_683;
wire n_474;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_934;
wire n_482;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_814;
wire n_389;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g206 ( 
.A(n_114),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_25),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_139),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_47),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_107),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_88),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_22),
.Y(n_213)
);

INVxp33_ASAP7_75t_R g214 ( 
.A(n_74),
.Y(n_214)
);

BUFx10_ASAP7_75t_L g215 ( 
.A(n_172),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_57),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_119),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_168),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_33),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_58),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_30),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_176),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_26),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_74),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_71),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_11),
.Y(n_226)
);

BUFx10_ASAP7_75t_L g227 ( 
.A(n_48),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_1),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_154),
.Y(n_229)
);

INVxp33_ASAP7_75t_R g230 ( 
.A(n_83),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_164),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_178),
.Y(n_233)
);

BUFx8_ASAP7_75t_SL g234 ( 
.A(n_42),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_57),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_46),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_138),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

INVx2_ASAP7_75t_SL g239 ( 
.A(n_79),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_82),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_15),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_121),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_21),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_60),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_4),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_200),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_81),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_113),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_64),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_150),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_89),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_105),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_28),
.Y(n_254)
);

BUFx5_ASAP7_75t_L g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_122),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_33),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_108),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_163),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_158),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_111),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_64),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_148),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_36),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_81),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_153),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_190),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_100),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_40),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_143),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_79),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_71),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_80),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_87),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_136),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_102),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_125),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_191),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_28),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_117),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_59),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_118),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_126),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_26),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_155),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_94),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_38),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g289 ( 
.A(n_62),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_132),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_51),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_35),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g293 ( 
.A(n_53),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_110),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_175),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_43),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_39),
.Y(n_297)
);

BUFx10_ASAP7_75t_L g298 ( 
.A(n_202),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_2),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_120),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_47),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_203),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_174),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_128),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_6),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_11),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_101),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_15),
.Y(n_309)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_165),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_189),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_43),
.Y(n_312)
);

CKINVDCx16_ASAP7_75t_R g313 ( 
.A(n_72),
.Y(n_313)
);

BUFx2_ASAP7_75t_SL g314 ( 
.A(n_131),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_35),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_124),
.Y(n_316)
);

BUFx2_ASAP7_75t_L g317 ( 
.A(n_184),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_40),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_116),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_56),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_58),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_44),
.Y(n_322)
);

BUFx3_ASAP7_75t_L g323 ( 
.A(n_72),
.Y(n_323)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_134),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_18),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_48),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_56),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_78),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_5),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_50),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_80),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_106),
.Y(n_332)
);

BUFx10_ASAP7_75t_L g333 ( 
.A(n_6),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_73),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_16),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g336 ( 
.A(n_192),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_115),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_109),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_144),
.Y(n_339)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_23),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_179),
.Y(n_341)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_181),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_129),
.Y(n_343)
);

BUFx5_ASAP7_75t_L g344 ( 
.A(n_61),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_17),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_103),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_18),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_180),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_137),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_193),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_70),
.Y(n_351)
);

BUFx10_ASAP7_75t_L g352 ( 
.A(n_135),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_183),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_41),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_50),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_159),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_196),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_142),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_66),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_36),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_166),
.Y(n_361)
);

BUFx10_ASAP7_75t_L g362 ( 
.A(n_97),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_68),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_133),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_140),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_187),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_62),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_156),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_146),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_95),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_27),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_73),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_32),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_52),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g375 ( 
.A(n_0),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_162),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_38),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_186),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_173),
.Y(n_379)
);

CKINVDCx16_ASAP7_75t_R g380 ( 
.A(n_171),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_54),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_22),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g383 ( 
.A(n_23),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_7),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_78),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_39),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_86),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_75),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_60),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_63),
.Y(n_390)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_61),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_16),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_198),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_104),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_194),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_68),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_31),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_177),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_65),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_182),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_76),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_157),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_7),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_149),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_14),
.Y(n_405)
);

BUFx3_ASAP7_75t_L g406 ( 
.A(n_96),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_59),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_161),
.Y(n_408)
);

BUFx6f_ASAP7_75t_SL g409 ( 
.A(n_215),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_211),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_234),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

NOR2xp67_ASAP7_75t_L g413 ( 
.A(n_324),
.B(n_0),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_231),
.Y(n_414)
);

BUFx2_ASAP7_75t_L g415 ( 
.A(n_323),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_344),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_233),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_344),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_344),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_344),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_344),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_223),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_223),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_335),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_255),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_335),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_255),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_209),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_209),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_213),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_317),
.B(n_1),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_320),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_324),
.B(n_2),
.Y(n_436)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_213),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_251),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_302),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_237),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_308),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_216),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_238),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_216),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_219),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_242),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_219),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_252),
.Y(n_448)
);

CKINVDCx16_ASAP7_75t_R g449 ( 
.A(n_375),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_235),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_253),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_257),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_317),
.B(n_3),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_235),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_259),
.Y(n_455)
);

CKINVDCx16_ASAP7_75t_R g456 ( 
.A(n_320),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_260),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_240),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_262),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_267),
.B(n_3),
.Y(n_460)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_240),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_269),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_267),
.B(n_5),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_248),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_248),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_250),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_311),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_369),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_255),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_275),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_313),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_250),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_254),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_254),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_270),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_255),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_283),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_284),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_398),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_249),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_270),
.Y(n_481)
);

INVxp67_ASAP7_75t_SL g482 ( 
.A(n_342),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_282),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_255),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_282),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_287),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_301),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_301),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_307),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_290),
.Y(n_490)
);

BUFx3_ASAP7_75t_L g491 ( 
.A(n_342),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_380),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_307),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_325),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_325),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_327),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_294),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_295),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_327),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_351),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_351),
.B(n_8),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_393),
.Y(n_502)
);

BUFx2_ASAP7_75t_L g503 ( 
.A(n_323),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_355),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_303),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_207),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_355),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_206),
.B(n_9),
.Y(n_508)
);

INVxp67_ASAP7_75t_SL g509 ( 
.A(n_376),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_206),
.B(n_9),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_359),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_304),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_431),
.Y(n_513)
);

AND2x4_ASAP7_75t_L g514 ( 
.A(n_413),
.B(n_376),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_435),
.Y(n_515)
);

AND2x6_ASAP7_75t_L g516 ( 
.A(n_412),
.B(n_324),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_482),
.B(n_310),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_509),
.B(n_336),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_431),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_456),
.A2(n_210),
.B1(n_312),
.B2(n_226),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_432),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_428),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_471),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_491),
.B(n_406),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_491),
.B(n_406),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_414),
.Y(n_526)
);

AND3x2_ASAP7_75t_L g527 ( 
.A(n_434),
.B(n_334),
.C(n_263),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_412),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_SL g529 ( 
.A(n_449),
.B(n_215),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_413),
.B(n_222),
.Y(n_530)
);

BUFx6f_ASAP7_75t_L g531 ( 
.A(n_428),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_432),
.Y(n_532)
);

NAND2x1p5_ASAP7_75t_L g533 ( 
.A(n_436),
.B(n_247),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_415),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g535 ( 
.A(n_415),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_463),
.B(n_416),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_501),
.A2(n_322),
.B1(n_326),
.B2(n_318),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_433),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_410),
.B(n_439),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_416),
.B(n_222),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_417),
.B(n_286),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_417),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_503),
.B(n_340),
.Y(n_543)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_503),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_433),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_430),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_444),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_449),
.B(n_215),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_430),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_506),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_419),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_419),
.B(n_340),
.Y(n_552)
);

AND2x4_ASAP7_75t_L g553 ( 
.A(n_420),
.B(n_286),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_469),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_456),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_420),
.B(n_338),
.Y(n_556)
);

AND2x4_ASAP7_75t_L g557 ( 
.A(n_421),
.B(n_319),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_421),
.B(n_319),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_422),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_422),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_423),
.B(n_339),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_469),
.Y(n_563)
);

OA21x2_ASAP7_75t_L g564 ( 
.A1(n_423),
.A2(n_371),
.B(n_359),
.Y(n_564)
);

BUFx6f_ASAP7_75t_L g565 ( 
.A(n_476),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_453),
.B(n_215),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_445),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_418),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_445),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_424),
.B(n_343),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_424),
.B(n_367),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_508),
.B(n_348),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g573 ( 
.A1(n_476),
.A2(n_361),
.B(n_332),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_447),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_484),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_447),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_484),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_450),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_450),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_454),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_425),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_425),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_426),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_426),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_454),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_427),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_427),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_429),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_501),
.B(n_239),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_429),
.B(n_367),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_458),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_510),
.B(n_349),
.Y(n_592)
);

INVx3_ASAP7_75t_L g593 ( 
.A(n_458),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_464),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

BUFx10_ASAP7_75t_L g596 ( 
.A(n_526),
.Y(n_596)
);

BUFx4f_ASAP7_75t_L g597 ( 
.A(n_564),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_522),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_556),
.B(n_440),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_539),
.Y(n_600)
);

BUFx10_ASAP7_75t_L g601 ( 
.A(n_568),
.Y(n_601)
);

NOR2x1p5_ASAP7_75t_L g602 ( 
.A(n_589),
.B(n_411),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_564),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_556),
.B(n_562),
.Y(n_604)
);

AND2x2_ASAP7_75t_SL g605 ( 
.A(n_530),
.B(n_332),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_552),
.B(n_571),
.Y(n_606)
);

AND2x2_ASAP7_75t_SL g607 ( 
.A(n_530),
.B(n_361),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_566),
.A2(n_438),
.B1(n_460),
.B2(n_293),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_566),
.B(n_443),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_522),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_575),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_575),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_517),
.B(n_446),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_575),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_564),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_522),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_577),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_543),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_577),
.Y(n_619)
);

AND2x2_ASAP7_75t_L g620 ( 
.A(n_552),
.B(n_466),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_564),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_564),
.Y(n_622)
);

OR2x2_ASAP7_75t_L g623 ( 
.A(n_534),
.B(n_448),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_577),
.Y(n_624)
);

AOI21x1_ASAP7_75t_L g625 ( 
.A1(n_536),
.A2(n_541),
.B(n_540),
.Y(n_625)
);

BUFx10_ASAP7_75t_L g626 ( 
.A(n_514),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_528),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_522),
.Y(n_628)
);

AND2x2_ASAP7_75t_L g629 ( 
.A(n_552),
.B(n_571),
.Y(n_629)
);

BUFx6f_ASAP7_75t_SL g630 ( 
.A(n_530),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_572),
.B(n_451),
.Y(n_631)
);

AO22x2_ASAP7_75t_L g632 ( 
.A1(n_537),
.A2(n_548),
.B1(n_529),
.B2(n_589),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g633 ( 
.A1(n_537),
.A2(n_360),
.B1(n_397),
.B2(n_390),
.Y(n_633)
);

NOR2xp33_ASAP7_75t_L g634 ( 
.A(n_572),
.B(n_452),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_528),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_562),
.B(n_455),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_570),
.B(n_457),
.Y(n_637)
);

INVx5_ASAP7_75t_L g638 ( 
.A(n_516),
.Y(n_638)
);

NOR2xp33_ASAP7_75t_L g639 ( 
.A(n_592),
.B(n_459),
.Y(n_639)
);

AND2x6_ASAP7_75t_L g640 ( 
.A(n_530),
.B(n_366),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_529),
.B(n_314),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_570),
.B(n_517),
.Y(n_642)
);

INVx8_ASAP7_75t_L g643 ( 
.A(n_516),
.Y(n_643)
);

AND2x2_ASAP7_75t_L g644 ( 
.A(n_571),
.B(n_466),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_528),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_564),
.Y(n_646)
);

INVx2_ASAP7_75t_SL g647 ( 
.A(n_543),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_516),
.Y(n_648)
);

AND2x4_ASAP7_75t_L g649 ( 
.A(n_514),
.B(n_208),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_542),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_542),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_561),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_518),
.B(n_462),
.Y(n_653)
);

AOI22xp33_ASAP7_75t_L g654 ( 
.A1(n_530),
.A2(n_293),
.B1(n_309),
.B2(n_239),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_542),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_561),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_555),
.Y(n_657)
);

AOI22xp5_ASAP7_75t_L g658 ( 
.A1(n_548),
.A2(n_401),
.B1(n_391),
.B2(n_289),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_536),
.A2(n_212),
.B1(n_218),
.B2(n_208),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_518),
.B(n_470),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_561),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_477),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_524),
.B(n_472),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_561),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_514),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_592),
.B(n_478),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_555),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_522),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_514),
.B(n_486),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_551),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_551),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_551),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_543),
.B(n_490),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_524),
.B(n_497),
.Y(n_674)
);

BUFx6f_ASAP7_75t_L g675 ( 
.A(n_522),
.Y(n_675)
);

BUFx10_ASAP7_75t_L g676 ( 
.A(n_550),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_589),
.B(n_498),
.Y(n_677)
);

INVxp33_ASAP7_75t_L g678 ( 
.A(n_515),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_560),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_560),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_560),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_549),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_550),
.B(n_505),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_540),
.B(n_366),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_539),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_540),
.B(n_212),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_525),
.B(n_512),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_549),
.Y(n_688)
);

NAND2xp33_ASAP7_75t_L g689 ( 
.A(n_516),
.B(n_247),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_522),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_549),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_549),
.Y(n_692)
);

NAND3xp33_ASAP7_75t_L g693 ( 
.A(n_534),
.B(n_442),
.C(n_437),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_540),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_525),
.B(n_480),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_549),
.Y(n_696)
);

BUFx6f_ASAP7_75t_L g697 ( 
.A(n_522),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_540),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_525),
.B(n_341),
.Y(n_699)
);

OAI22xp5_ASAP7_75t_L g700 ( 
.A1(n_535),
.A2(n_492),
.B1(n_502),
.B2(n_383),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_531),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_541),
.B(n_353),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_541),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_541),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_541),
.B(n_465),
.C(n_461),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_581),
.Y(n_706)
);

OAI22xp33_ASAP7_75t_L g707 ( 
.A1(n_535),
.A2(n_329),
.B1(n_272),
.B2(n_407),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_531),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_531),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_581),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_553),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_581),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_409),
.Y(n_713)
);

BUFx3_ASAP7_75t_L g714 ( 
.A(n_553),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_553),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_553),
.B(n_557),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_520),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_553),
.B(n_356),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_581),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_557),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_544),
.B(n_217),
.Y(n_721)
);

INVx2_ASAP7_75t_SL g722 ( 
.A(n_515),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_531),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_531),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_523),
.B(n_409),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_SL g726 ( 
.A1(n_520),
.A2(n_409),
.B1(n_479),
.B2(n_468),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_557),
.Y(n_727)
);

AND2x2_ASAP7_75t_SL g728 ( 
.A(n_557),
.B(n_387),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_557),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_558),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_558),
.B(n_357),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_581),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_581),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_523),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_531),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_590),
.B(n_472),
.Y(n_736)
);

INVx4_ASAP7_75t_L g737 ( 
.A(n_531),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_SL g738 ( 
.A(n_523),
.B(n_309),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_558),
.A2(n_374),
.B1(n_371),
.B2(n_405),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_581),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_558),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_590),
.B(n_314),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_558),
.A2(n_374),
.B1(n_381),
.B2(n_405),
.Y(n_743)
);

OR2x6_ASAP7_75t_L g744 ( 
.A(n_590),
.B(n_218),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_593),
.B(n_217),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_631),
.B(n_441),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_606),
.B(n_593),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_604),
.B(n_642),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_634),
.B(n_467),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_605),
.B(n_247),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_714),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_639),
.B(n_593),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_605),
.B(n_247),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_606),
.B(n_593),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_629),
.B(n_531),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_629),
.B(n_546),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_599),
.B(n_230),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_603),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_605),
.B(n_247),
.Y(n_760)
);

INVxp33_ASAP7_75t_SL g761 ( 
.A(n_700),
.Y(n_761)
);

AO22x2_ASAP7_75t_L g762 ( 
.A1(n_632),
.A2(n_229),
.B1(n_261),
.B2(n_244),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_618),
.B(n_527),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_714),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_694),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_636),
.B(n_527),
.Y(n_766)
);

BUFx6f_ASAP7_75t_SL g767 ( 
.A(n_596),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_694),
.Y(n_768)
);

OAI22xp33_ASAP7_75t_L g769 ( 
.A1(n_641),
.A2(n_658),
.B1(n_744),
.B2(n_647),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_637),
.B(n_214),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_603),
.Y(n_771)
);

NOR2xp33_ASAP7_75t_SL g772 ( 
.A(n_596),
.B(n_217),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_615),
.Y(n_773)
);

INVx2_ASAP7_75t_L g774 ( 
.A(n_615),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_607),
.B(n_546),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_607),
.B(n_546),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_698),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_626),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_607),
.B(n_546),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_728),
.B(n_546),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_698),
.Y(n_781)
);

BUFx6f_ASAP7_75t_L g782 ( 
.A(n_626),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_728),
.B(n_546),
.Y(n_783)
);

NOR2xp67_ASAP7_75t_SL g784 ( 
.A(n_638),
.B(n_229),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_693),
.B(n_513),
.Y(n_785)
);

OAI21xp5_ASAP7_75t_L g786 ( 
.A1(n_597),
.A2(n_622),
.B(n_621),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_728),
.B(n_546),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_703),
.Y(n_788)
);

AOI21xp5_ASAP7_75t_L g789 ( 
.A1(n_716),
.A2(n_554),
.B(n_546),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_621),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_653),
.B(n_554),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_L g792 ( 
.A(n_660),
.B(n_264),
.Y(n_792)
);

NAND2x1p5_ASAP7_75t_L g793 ( 
.A(n_638),
.B(n_573),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_638),
.B(n_554),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_652),
.B(n_554),
.Y(n_795)
);

NOR2xp67_ASAP7_75t_L g796 ( 
.A(n_623),
.B(n_513),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_638),
.B(n_554),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_703),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_638),
.B(n_554),
.Y(n_799)
);

AND2x4_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_519),
.Y(n_800)
);

AND2x2_ASAP7_75t_SL g801 ( 
.A(n_597),
.B(n_387),
.Y(n_801)
);

OAI22xp33_ASAP7_75t_L g802 ( 
.A1(n_641),
.A2(n_261),
.B1(n_268),
.B2(n_244),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_652),
.B(n_554),
.Y(n_803)
);

INVxp67_ASAP7_75t_L g804 ( 
.A(n_677),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_656),
.B(n_554),
.Y(n_805)
);

O2A1O1Ixp33_ASAP7_75t_L g806 ( 
.A1(n_659),
.A2(n_622),
.B(n_646),
.C(n_618),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_638),
.B(n_563),
.Y(n_807)
);

OAI221xp5_ASAP7_75t_L g808 ( 
.A1(n_608),
.A2(n_654),
.B1(n_739),
.B2(n_743),
.C(n_658),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_646),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_704),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_704),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_647),
.A2(n_271),
.B1(n_276),
.B2(n_268),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_656),
.B(n_563),
.Y(n_813)
);

INVxp33_ASAP7_75t_L g814 ( 
.A(n_678),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_711),
.Y(n_815)
);

OAI22xp33_ASAP7_75t_L g816 ( 
.A1(n_641),
.A2(n_276),
.B1(n_277),
.B2(n_271),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_661),
.B(n_563),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_648),
.B(n_563),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_667),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_643),
.B(n_516),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_648),
.B(n_563),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_663),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_715),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_641),
.A2(n_516),
.B1(n_370),
.B2(n_364),
.Y(n_824)
);

BUFx6f_ASAP7_75t_L g825 ( 
.A(n_626),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_661),
.B(n_563),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_611),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_611),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_563),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_648),
.B(n_597),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_648),
.B(n_563),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_664),
.B(n_565),
.Y(n_832)
);

OR2x2_ASAP7_75t_SL g833 ( 
.A(n_623),
.B(n_381),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_620),
.B(n_565),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_620),
.B(n_519),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_612),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_644),
.B(n_521),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_648),
.B(n_565),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_644),
.B(n_521),
.Y(n_839)
);

NOR2xp33_ASAP7_75t_L g840 ( 
.A(n_666),
.B(n_220),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_736),
.B(n_532),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_649),
.B(n_565),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_649),
.B(n_565),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_649),
.B(n_565),
.Y(n_844)
);

AND2x4_ASAP7_75t_SL g845 ( 
.A(n_596),
.B(n_217),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_649),
.B(n_565),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_715),
.B(n_565),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_612),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_722),
.B(n_532),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_648),
.B(n_255),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_625),
.A2(n_573),
.B(n_516),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_720),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_L g853 ( 
.A(n_674),
.B(n_221),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_720),
.B(n_516),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_736),
.B(n_538),
.Y(n_855)
);

AO21x1_ASAP7_75t_L g856 ( 
.A1(n_659),
.A2(n_533),
.B(n_278),
.Y(n_856)
);

BUFx3_ASAP7_75t_L g857 ( 
.A(n_727),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_614),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_727),
.B(n_729),
.Y(n_859)
);

OAI22xp5_ASAP7_75t_L g860 ( 
.A1(n_641),
.A2(n_408),
.B1(n_316),
.B2(n_402),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_626),
.B(n_255),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_730),
.B(n_741),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_730),
.B(n_516),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_741),
.Y(n_864)
);

BUFx6f_ASAP7_75t_L g865 ( 
.A(n_665),
.Y(n_865)
);

BUFx6f_ASAP7_75t_L g866 ( 
.A(n_665),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_734),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_614),
.Y(n_868)
);

INVx2_ASAP7_75t_SL g869 ( 
.A(n_742),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_722),
.B(n_538),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_665),
.B(n_625),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_746),
.Y(n_872)
);

INVx2_ASAP7_75t_SL g873 ( 
.A(n_742),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_662),
.B(n_533),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_687),
.B(n_224),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_744),
.B(n_545),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_665),
.B(n_255),
.Y(n_877)
);

AND2x6_ASAP7_75t_SL g878 ( 
.A(n_725),
.B(n_382),
.Y(n_878)
);

OAI22xp5_ASAP7_75t_L g879 ( 
.A1(n_742),
.A2(n_400),
.B1(n_278),
.B2(n_279),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_669),
.B(n_533),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_L g881 ( 
.A1(n_699),
.A2(n_579),
.B(n_594),
.C(n_591),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_746),
.B(n_533),
.Y(n_882)
);

OAI221xp5_ASAP7_75t_L g883 ( 
.A1(n_705),
.A2(n_388),
.B1(n_384),
.B2(n_382),
.C(n_585),
.Y(n_883)
);

NOR2x1p5_ASAP7_75t_L g884 ( 
.A(n_657),
.B(n_225),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_686),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_686),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_686),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_686),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_L g889 ( 
.A(n_613),
.B(n_228),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_617),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_617),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_609),
.B(n_232),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_619),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_619),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_724),
.B(n_584),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_670),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_744),
.B(n_545),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_670),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_702),
.B(n_584),
.Y(n_899)
);

AOI22xp5_ASAP7_75t_L g900 ( 
.A1(n_632),
.A2(n_395),
.B1(n_358),
.B2(n_365),
.Y(n_900)
);

AOI22xp33_ASAP7_75t_L g901 ( 
.A1(n_640),
.A2(n_337),
.B1(n_402),
.B2(n_277),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_624),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_734),
.B(n_547),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_671),
.Y(n_904)
);

OAI22xp5_ASAP7_75t_L g905 ( 
.A1(n_742),
.A2(n_279),
.B1(n_281),
.B2(n_300),
.Y(n_905)
);

AO22x1_ASAP7_75t_L g906 ( 
.A1(n_713),
.A2(n_717),
.B1(n_388),
.B2(n_384),
.Y(n_906)
);

BUFx5_ASAP7_75t_L g907 ( 
.A(n_640),
.Y(n_907)
);

NOR2xp33_ASAP7_75t_L g908 ( 
.A(n_673),
.B(n_236),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_SL g909 ( 
.A(n_643),
.B(n_255),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_632),
.A2(n_378),
.B1(n_404),
.B2(n_394),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_718),
.B(n_584),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_744),
.B(n_547),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_624),
.Y(n_913)
);

CKINVDCx20_ASAP7_75t_R g914 ( 
.A(n_600),
.Y(n_914)
);

AOI22xp33_ASAP7_75t_L g915 ( 
.A1(n_640),
.A2(n_408),
.B1(n_281),
.B2(n_350),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_731),
.B(n_598),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_749),
.B(n_792),
.Y(n_917)
);

NOR2x1_ASAP7_75t_L g918 ( 
.A(n_766),
.B(n_602),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_775),
.A2(n_643),
.B(n_628),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_748),
.B(n_744),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_827),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_819),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_857),
.Y(n_923)
);

AOI21xp5_ASAP7_75t_L g924 ( 
.A1(n_776),
.A2(n_643),
.B(n_628),
.Y(n_924)
);

NOR2xp33_ASAP7_75t_L g925 ( 
.A(n_804),
.B(n_695),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_857),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_748),
.B(n_632),
.Y(n_927)
);

O2A1O1Ixp33_ASAP7_75t_L g928 ( 
.A1(n_806),
.A2(n_745),
.B(n_742),
.C(n_721),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_755),
.B(n_640),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_864),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_SL g931 ( 
.A(n_801),
.B(n_643),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_755),
.B(n_640),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_822),
.B(n_640),
.Y(n_933)
);

A2O1A1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_808),
.A2(n_705),
.B(n_633),
.C(n_717),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_867),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_864),
.Y(n_936)
);

NOR2xp33_ASAP7_75t_L g937 ( 
.A(n_758),
.B(n_683),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_801),
.B(n_596),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_779),
.A2(n_737),
.B(n_628),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_822),
.B(n_640),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_835),
.B(n_679),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_778),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_L g943 ( 
.A(n_770),
.B(n_667),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_835),
.B(n_681),
.Y(n_944)
);

BUFx2_ASAP7_75t_L g945 ( 
.A(n_914),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_786),
.A2(n_681),
.B(n_573),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_907),
.B(n_601),
.Y(n_947)
);

NAND3xp33_ASAP7_75t_L g948 ( 
.A(n_840),
.B(n_633),
.C(n_738),
.Y(n_948)
);

OAI21xp5_ASAP7_75t_L g949 ( 
.A1(n_756),
.A2(n_635),
.B(n_627),
.Y(n_949)
);

HB1xp67_ASAP7_75t_L g950 ( 
.A(n_903),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_837),
.B(n_598),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_765),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_778),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_778),
.B(n_598),
.Y(n_954)
);

AND2x2_ASAP7_75t_L g955 ( 
.A(n_849),
.B(n_676),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_827),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_837),
.B(n_839),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_780),
.A2(n_871),
.B(n_820),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_839),
.B(n_610),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_768),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_871),
.A2(n_820),
.B(n_787),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_841),
.B(n_610),
.Y(n_962)
);

O2A1O1Ixp5_ASAP7_75t_L g963 ( 
.A1(n_751),
.A2(n_616),
.B(n_668),
.C(n_610),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_841),
.B(n_616),
.Y(n_964)
);

AOI21xp5_ASAP7_75t_L g965 ( 
.A1(n_783),
.A2(n_737),
.B(n_689),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_783),
.A2(n_737),
.B(n_697),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_787),
.A2(n_697),
.B(n_675),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_747),
.B(n_601),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_750),
.B(n_601),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_757),
.A2(n_697),
.B(n_675),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_753),
.B(n_616),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_777),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_853),
.B(n_668),
.Y(n_973)
);

O2A1O1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_860),
.A2(n_707),
.B(n_635),
.C(n_645),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_791),
.A2(n_697),
.B(n_675),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_834),
.A2(n_645),
.B(n_627),
.Y(n_976)
);

NAND2x1p5_ASAP7_75t_L g977 ( 
.A(n_778),
.B(n_668),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_907),
.B(n_601),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_855),
.Y(n_979)
);

INVx2_ASAP7_75t_SL g980 ( 
.A(n_870),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_830),
.A2(n_697),
.B(n_675),
.Y(n_981)
);

HB1xp67_ASAP7_75t_L g982 ( 
.A(n_876),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_875),
.B(n_690),
.Y(n_983)
);

AO21x1_ASAP7_75t_L g984 ( 
.A1(n_751),
.A2(n_316),
.B(n_300),
.Y(n_984)
);

AO21x1_ASAP7_75t_L g985 ( 
.A1(n_754),
.A2(n_760),
.B(n_769),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_830),
.A2(n_916),
.B(n_843),
.Y(n_986)
);

AO21x1_ASAP7_75t_L g987 ( 
.A1(n_754),
.A2(n_346),
.B(n_337),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_842),
.A2(n_675),
.B(n_690),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_855),
.B(n_701),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_763),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_855),
.B(n_701),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_844),
.A2(n_708),
.B(n_701),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_846),
.A2(n_709),
.B(n_708),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_861),
.A2(n_651),
.B(n_650),
.Y(n_994)
);

CKINVDCx5p33_ASAP7_75t_R g995 ( 
.A(n_767),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_899),
.A2(n_709),
.B(n_708),
.Y(n_996)
);

INVx2_ASAP7_75t_SL g997 ( 
.A(n_884),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_800),
.B(n_709),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_800),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_907),
.B(n_676),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_911),
.A2(n_735),
.B(n_723),
.Y(n_1001)
);

AND2x2_ASAP7_75t_L g1002 ( 
.A(n_796),
.B(n_676),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_800),
.B(n_723),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_874),
.A2(n_735),
.B(n_723),
.Y(n_1004)
);

AND2x4_ASAP7_75t_L g1005 ( 
.A(n_876),
.B(n_897),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_SL g1006 ( 
.A1(n_760),
.A2(n_400),
.B(n_346),
.C(n_379),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_828),
.Y(n_1007)
);

OAI21xp33_ASAP7_75t_SL g1008 ( 
.A1(n_759),
.A2(n_602),
.B(n_379),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_781),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_880),
.A2(n_710),
.B(n_706),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_788),
.Y(n_1011)
);

OAI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_851),
.A2(n_651),
.B(n_650),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_895),
.A2(n_710),
.B(n_706),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_828),
.Y(n_1014)
);

AOI33xp33_ASAP7_75t_L g1015 ( 
.A1(n_802),
.A2(n_473),
.A3(n_511),
.B1(n_474),
.B2(n_475),
.B3(n_481),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_771),
.B(n_655),
.Y(n_1016)
);

BUFx8_ASAP7_75t_L g1017 ( 
.A(n_767),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_771),
.B(n_655),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_773),
.A2(n_630),
.B1(n_657),
.B2(n_726),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_SL g1020 ( 
.A(n_907),
.B(n_676),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_854),
.A2(n_719),
.B(n_712),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_773),
.B(n_672),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_863),
.A2(n_733),
.B(n_732),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_774),
.B(n_672),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_847),
.A2(n_733),
.B(n_732),
.Y(n_1025)
);

CKINVDCx10_ASAP7_75t_R g1026 ( 
.A(n_767),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_882),
.A2(n_740),
.B(n_680),
.Y(n_1027)
);

BUFx12f_ASAP7_75t_L g1028 ( 
.A(n_833),
.Y(n_1028)
);

A2O1A1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_900),
.A2(n_350),
.B(n_569),
.C(n_567),
.Y(n_1029)
);

INVx1_ASAP7_75t_SL g1030 ( 
.A(n_814),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_789),
.A2(n_740),
.B(n_680),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_774),
.B(n_684),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_859),
.A2(n_862),
.B(n_803),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_782),
.Y(n_1034)
);

AND2x2_ASAP7_75t_SL g1035 ( 
.A(n_772),
.B(n_473),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_795),
.A2(n_688),
.B(n_682),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_907),
.B(n_682),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_805),
.A2(n_691),
.B(n_688),
.Y(n_1038)
);

HB1xp67_ASAP7_75t_L g1039 ( 
.A(n_897),
.Y(n_1039)
);

NAND2xp5_ASAP7_75t_L g1040 ( 
.A(n_790),
.B(n_684),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_798),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_813),
.A2(n_692),
.B(n_691),
.Y(n_1042)
);

INVxp33_ASAP7_75t_SL g1043 ( 
.A(n_889),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_817),
.A2(n_696),
.B(n_692),
.Y(n_1044)
);

OAI22xp5_ASAP7_75t_L g1045 ( 
.A1(n_809),
.A2(n_630),
.B1(n_368),
.B2(n_696),
.Y(n_1045)
);

A2O1A1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_910),
.A2(n_567),
.B(n_559),
.C(n_594),
.Y(n_1046)
);

O2A1O1Ixp33_ASAP7_75t_L g1047 ( 
.A1(n_816),
.A2(n_559),
.B(n_569),
.C(n_579),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_892),
.B(n_685),
.C(n_243),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_826),
.A2(n_595),
.B(n_684),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_829),
.A2(n_832),
.B(n_825),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_810),
.Y(n_1051)
);

AOI21xp5_ASAP7_75t_L g1052 ( 
.A1(n_782),
.A2(n_595),
.B(n_684),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_782),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_836),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_809),
.B(n_684),
.Y(n_1055)
);

NAND2xp33_ASAP7_75t_L g1056 ( 
.A(n_782),
.B(n_684),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_SL g1057 ( 
.A(n_907),
.B(n_581),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_825),
.A2(n_595),
.B(n_684),
.Y(n_1058)
);

O2A1O1Ixp33_ASAP7_75t_SL g1059 ( 
.A1(n_879),
.A2(n_905),
.B(n_877),
.C(n_812),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_811),
.B(n_584),
.Y(n_1060)
);

AND2x2_ASAP7_75t_L g1061 ( 
.A(n_845),
.B(n_685),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_883),
.A2(n_578),
.B(n_591),
.C(n_574),
.Y(n_1062)
);

AND2x2_ASAP7_75t_L g1063 ( 
.A(n_845),
.B(n_574),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_825),
.A2(n_595),
.B(n_578),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_761),
.B(n_241),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_836),
.Y(n_1066)
);

AO21x1_ASAP7_75t_L g1067 ( 
.A1(n_877),
.A2(n_580),
.B(n_576),
.Y(n_1067)
);

AO21x1_ASAP7_75t_L g1068 ( 
.A1(n_872),
.A2(n_580),
.B(n_576),
.Y(n_1068)
);

HB1xp67_ASAP7_75t_L g1069 ( 
.A(n_912),
.Y(n_1069)
);

AOI21xp5_ASAP7_75t_L g1070 ( 
.A1(n_825),
.A2(n_866),
.B(n_865),
.Y(n_1070)
);

NAND2xp5_ASAP7_75t_L g1071 ( 
.A(n_815),
.B(n_585),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_823),
.B(n_586),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_852),
.B(n_586),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_912),
.B(n_586),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_865),
.A2(n_588),
.B(n_587),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_909),
.A2(n_587),
.B(n_588),
.Y(n_1076)
);

AOI22xp33_ASAP7_75t_L g1077 ( 
.A1(n_762),
.A2(n_227),
.B1(n_333),
.B2(n_362),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_752),
.B(n_588),
.Y(n_1078)
);

NOR2xp33_ASAP7_75t_R g1079 ( 
.A(n_914),
.B(n_245),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_865),
.A2(n_587),
.B(n_583),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_764),
.B(n_885),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_907),
.B(n_582),
.Y(n_1082)
);

INVxp67_ASAP7_75t_SL g1083 ( 
.A(n_865),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_886),
.B(n_582),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_887),
.B(n_474),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_L g1086 ( 
.A1(n_909),
.A2(n_475),
.B(n_481),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_888),
.B(n_582),
.Y(n_1087)
);

BUFx2_ASAP7_75t_L g1088 ( 
.A(n_762),
.Y(n_1088)
);

AOI21xp5_ASAP7_75t_L g1089 ( 
.A1(n_866),
.A2(n_583),
.B(n_582),
.Y(n_1089)
);

INVx2_ASAP7_75t_SL g1090 ( 
.A(n_906),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_848),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_896),
.B(n_582),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_848),
.Y(n_1093)
);

NAND2x1p5_ASAP7_75t_L g1094 ( 
.A(n_866),
.B(n_582),
.Y(n_1094)
);

AND2x4_ASAP7_75t_L g1095 ( 
.A(n_785),
.B(n_483),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_898),
.Y(n_1096)
);

OAI22xp5_ASAP7_75t_L g1097 ( 
.A1(n_869),
.A2(n_246),
.B1(n_256),
.B2(n_258),
.Y(n_1097)
);

OR2x2_ASAP7_75t_L g1098 ( 
.A(n_908),
.B(n_483),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_866),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_869),
.B(n_582),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_793),
.A2(n_583),
.B(n_582),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_793),
.A2(n_583),
.B(n_511),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_917),
.B(n_762),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_957),
.B(n_873),
.Y(n_1104)
);

OAI22xp33_ASAP7_75t_L g1105 ( 
.A1(n_1043),
.A2(n_948),
.B1(n_761),
.B2(n_1065),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_1033),
.A2(n_873),
.B(n_797),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_922),
.Y(n_1107)
);

AOI22x1_ASAP7_75t_L g1108 ( 
.A1(n_1010),
.A2(n_1004),
.B1(n_961),
.B2(n_1049),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_SL g1109 ( 
.A(n_968),
.B(n_298),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_942),
.Y(n_1110)
);

BUFx2_ASAP7_75t_L g1111 ( 
.A(n_1030),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_952),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_L g1113 ( 
.A1(n_937),
.A2(n_856),
.B1(n_915),
.B2(n_901),
.Y(n_1113)
);

NOR2xp33_ASAP7_75t_L g1114 ( 
.A(n_1065),
.B(n_878),
.Y(n_1114)
);

AOI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_919),
.A2(n_797),
.B(n_794),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_927),
.B(n_941),
.Y(n_1116)
);

AOI221x1_ASAP7_75t_L g1117 ( 
.A1(n_1029),
.A2(n_904),
.B1(n_913),
.B2(n_902),
.C(n_894),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_944),
.B(n_858),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_924),
.A2(n_799),
.B(n_794),
.Y(n_1119)
);

NOR2xp33_ASAP7_75t_L g1120 ( 
.A(n_968),
.B(n_824),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1098),
.B(n_881),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1091),
.Y(n_1122)
);

O2A1O1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_934),
.A2(n_913),
.B(n_902),
.C(n_894),
.Y(n_1123)
);

INVx3_ASAP7_75t_SL g1124 ( 
.A(n_995),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_1056),
.A2(n_831),
.B(n_799),
.Y(n_1125)
);

NAND3xp33_ASAP7_75t_SL g1126 ( 
.A(n_937),
.B(n_372),
.C(n_266),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_960),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_950),
.B(n_227),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_972),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_958),
.A2(n_931),
.B(n_973),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_955),
.B(n_868),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_951),
.B(n_959),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_R g1133 ( 
.A(n_969),
.B(n_868),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_950),
.B(n_890),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_943),
.A2(n_784),
.B(n_891),
.C(n_890),
.Y(n_1135)
);

NOR3xp33_ASAP7_75t_SL g1136 ( 
.A(n_934),
.B(n_1019),
.C(n_943),
.Y(n_1136)
);

INVxp67_ASAP7_75t_L g1137 ( 
.A(n_935),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1009),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1002),
.B(n_891),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_1035),
.A2(n_893),
.B1(n_385),
.B2(n_377),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_931),
.A2(n_821),
.B(n_838),
.Y(n_1141)
);

BUFx6f_ASAP7_75t_L g1142 ( 
.A(n_942),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_921),
.Y(n_1143)
);

INVxp67_ASAP7_75t_L g1144 ( 
.A(n_945),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_942),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_969),
.B(n_893),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1011),
.Y(n_1147)
);

AND2x4_ASAP7_75t_L g1148 ( 
.A(n_979),
.B(n_807),
.Y(n_1148)
);

A2O1A1Ixp33_ASAP7_75t_L g1149 ( 
.A1(n_925),
.A2(n_850),
.B(n_831),
.C(n_818),
.Y(n_1149)
);

OAI21xp5_ASAP7_75t_L g1150 ( 
.A1(n_986),
.A2(n_850),
.B(n_818),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_1035),
.B(n_298),
.Y(n_1151)
);

AOI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_983),
.A2(n_807),
.B(n_583),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_SL g1153 ( 
.A1(n_1028),
.A2(n_331),
.B1(n_330),
.B2(n_328),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_939),
.A2(n_583),
.B(n_507),
.Y(n_1154)
);

NAND2xp33_ASAP7_75t_R g1155 ( 
.A(n_1079),
.B(n_84),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_942),
.Y(n_1156)
);

NAND2xp5_ASAP7_75t_SL g1157 ( 
.A(n_925),
.B(n_298),
.Y(n_1157)
);

OAI22xp5_ASAP7_75t_L g1158 ( 
.A1(n_1077),
.A2(n_363),
.B1(n_274),
.B2(n_280),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_SL g1159 ( 
.A(n_979),
.B(n_298),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1041),
.B(n_583),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_953),
.B(n_583),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_999),
.B(n_352),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_1026),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1051),
.B(n_265),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1029),
.A2(n_507),
.B(n_504),
.C(n_500),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_921),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1050),
.A2(n_504),
.B(n_500),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_929),
.A2(n_499),
.B(n_496),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_932),
.A2(n_499),
.B(n_496),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_965),
.A2(n_495),
.B(n_494),
.Y(n_1170)
);

O2A1O1Ixp33_ASAP7_75t_L g1171 ( 
.A1(n_1046),
.A2(n_495),
.B(n_494),
.C(n_493),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_1096),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_980),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1085),
.Y(n_1174)
);

O2A1O1Ixp5_ASAP7_75t_L g1175 ( 
.A1(n_1068),
.A2(n_493),
.B(n_489),
.C(n_488),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_SL g1176 ( 
.A(n_999),
.B(n_352),
.Y(n_1176)
);

BUFx4f_ASAP7_75t_SL g1177 ( 
.A(n_1017),
.Y(n_1177)
);

AND2x4_ASAP7_75t_L g1178 ( 
.A(n_1005),
.B(n_982),
.Y(n_1178)
);

NOR2xp33_ASAP7_75t_L g1179 ( 
.A(n_1090),
.B(n_982),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_1085),
.Y(n_1180)
);

A2O1A1Ixp33_ASAP7_75t_L g1181 ( 
.A1(n_928),
.A2(n_345),
.B(n_273),
.C(n_285),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1032),
.A2(n_489),
.B(n_488),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_923),
.B(n_288),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1079),
.Y(n_1184)
);

AND2x6_ASAP7_75t_L g1185 ( 
.A(n_1034),
.B(n_487),
.Y(n_1185)
);

OR2x6_ASAP7_75t_SL g1186 ( 
.A(n_1048),
.B(n_291),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1005),
.B(n_485),
.Y(n_1187)
);

A2O1A1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1046),
.A2(n_292),
.B(n_305),
.C(n_403),
.Y(n_1188)
);

O2A1O1Ixp33_ASAP7_75t_L g1189 ( 
.A1(n_938),
.A2(n_487),
.B(n_485),
.C(n_352),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1039),
.B(n_296),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1040),
.A2(n_93),
.B(n_205),
.Y(n_1191)
);

O2A1O1Ixp33_ASAP7_75t_L g1192 ( 
.A1(n_938),
.A2(n_352),
.B(n_362),
.C(n_227),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1077),
.A2(n_399),
.B1(n_396),
.B2(n_392),
.Y(n_1193)
);

AOI22xp33_ASAP7_75t_L g1194 ( 
.A1(n_985),
.A2(n_362),
.B1(n_227),
.B2(n_333),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1088),
.A2(n_389),
.B1(n_386),
.B2(n_373),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_956),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_1017),
.Y(n_1197)
);

A2O1A1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_920),
.A2(n_321),
.B(n_354),
.C(n_347),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1007),
.Y(n_1199)
);

A2O1A1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1008),
.A2(n_315),
.B(n_306),
.C(n_299),
.Y(n_1200)
);

BUFx6f_ASAP7_75t_L g1201 ( 
.A(n_1034),
.Y(n_1201)
);

O2A1O1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1059),
.A2(n_362),
.B(n_333),
.C(n_297),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_962),
.B(n_204),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_946),
.A2(n_152),
.B(n_201),
.Y(n_1204)
);

AOI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1055),
.A2(n_199),
.B(n_197),
.Y(n_1205)
);

AOI21xp5_ASAP7_75t_L g1206 ( 
.A1(n_975),
.A2(n_195),
.B(n_188),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_964),
.B(n_185),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_971),
.A2(n_170),
.B(n_169),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1034),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1074),
.B(n_1039),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1007),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1014),
.Y(n_1212)
);

NOR2xp33_ASAP7_75t_SL g1213 ( 
.A(n_1061),
.B(n_333),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1069),
.B(n_167),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_970),
.A2(n_160),
.B(n_151),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1071),
.B(n_145),
.Y(n_1216)
);

A2O1A1Ixp33_ASAP7_75t_L g1217 ( 
.A1(n_974),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_1217)
);

INVx1_ASAP7_75t_L g1218 ( 
.A(n_1014),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_1054),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_SL g1220 ( 
.A(n_926),
.B(n_130),
.Y(n_1220)
);

AND2x4_ASAP7_75t_L g1221 ( 
.A(n_990),
.B(n_127),
.Y(n_1221)
);

AOI21xp5_ASAP7_75t_L g1222 ( 
.A1(n_1070),
.A2(n_123),
.B(n_112),
.Y(n_1222)
);

NAND2xp5_ASAP7_75t_L g1223 ( 
.A(n_1054),
.B(n_99),
.Y(n_1223)
);

O2A1O1Ixp33_ASAP7_75t_L g1224 ( 
.A1(n_1059),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_1224)
);

INVx2_ASAP7_75t_L g1225 ( 
.A(n_1093),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_966),
.A2(n_98),
.B(n_92),
.Y(n_1226)
);

AND2x6_ASAP7_75t_L g1227 ( 
.A(n_1034),
.B(n_90),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_930),
.B(n_85),
.Y(n_1228)
);

AOI22x1_ASAP7_75t_L g1229 ( 
.A1(n_1027),
.A2(n_14),
.B1(n_17),
.B2(n_19),
.Y(n_1229)
);

NOR2xp33_ASAP7_75t_L g1230 ( 
.A(n_1063),
.B(n_19),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1093),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1012),
.A2(n_20),
.B(n_21),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_997),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1099),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_989),
.B(n_20),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1095),
.B(n_24),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1097),
.A2(n_24),
.B(n_25),
.C(n_29),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1095),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_991),
.B(n_29),
.Y(n_1239)
);

INVx2_ASAP7_75t_L g1240 ( 
.A(n_1066),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1099),
.Y(n_1241)
);

O2A1O1Ixp33_ASAP7_75t_L g1242 ( 
.A1(n_1047),
.A2(n_34),
.B(n_37),
.C(n_41),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_998),
.B(n_34),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_918),
.B(n_37),
.Y(n_1244)
);

AND2x2_ASAP7_75t_L g1245 ( 
.A(n_936),
.B(n_42),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1003),
.B(n_45),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1083),
.A2(n_45),
.B1(n_46),
.B2(n_49),
.Y(n_1247)
);

O2A1O1Ixp33_ASAP7_75t_L g1248 ( 
.A1(n_1081),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_933),
.A2(n_82),
.B1(n_54),
.B2(n_55),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1016),
.B(n_53),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_SL g1251 ( 
.A(n_1099),
.B(n_55),
.Y(n_1251)
);

INVx4_ASAP7_75t_L g1252 ( 
.A(n_1099),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1037),
.A2(n_1082),
.B(n_1057),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1037),
.A2(n_77),
.B(n_65),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1086),
.B(n_63),
.Y(n_1255)
);

INVxp67_ASAP7_75t_L g1256 ( 
.A(n_1078),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_953),
.B(n_66),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_1057),
.A2(n_76),
.B(n_69),
.Y(n_1258)
);

INVx2_ASAP7_75t_SL g1259 ( 
.A(n_1100),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1082),
.A2(n_67),
.B(n_69),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1120),
.A2(n_1105),
.B1(n_1114),
.B2(n_1136),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1187),
.B(n_1015),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1108),
.A2(n_994),
.B(n_1101),
.Y(n_1263)
);

AO21x1_ASAP7_75t_L g1264 ( 
.A1(n_1232),
.A2(n_1020),
.B(n_1000),
.Y(n_1264)
);

AO22x2_ASAP7_75t_L g1265 ( 
.A1(n_1151),
.A2(n_1020),
.B1(n_1000),
.B2(n_978),
.Y(n_1265)
);

NOR2xp33_ASAP7_75t_SL g1266 ( 
.A(n_1109),
.B(n_1053),
.Y(n_1266)
);

AO31x2_ASAP7_75t_L g1267 ( 
.A1(n_1117),
.A2(n_1067),
.A3(n_984),
.B(n_987),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1106),
.A2(n_1013),
.B(n_1025),
.Y(n_1268)
);

NAND3x1_ASAP7_75t_L g1269 ( 
.A(n_1230),
.B(n_1015),
.C(n_940),
.Y(n_1269)
);

AOI21xp5_ASAP7_75t_L g1270 ( 
.A1(n_1130),
.A2(n_978),
.B(n_947),
.Y(n_1270)
);

INVx2_ASAP7_75t_L g1271 ( 
.A(n_1143),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1187),
.B(n_1062),
.Y(n_1272)
);

AOI22xp33_ASAP7_75t_L g1273 ( 
.A1(n_1126),
.A2(n_1238),
.B1(n_1180),
.B2(n_1174),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1115),
.A2(n_1031),
.B(n_1001),
.Y(n_1274)
);

AOI221x1_ASAP7_75t_L g1275 ( 
.A1(n_1217),
.A2(n_1045),
.B1(n_996),
.B2(n_967),
.C(n_1064),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1116),
.B(n_1024),
.Y(n_1276)
);

AOI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1132),
.A2(n_947),
.B(n_1053),
.Y(n_1277)
);

AO31x2_ASAP7_75t_L g1278 ( 
.A1(n_1181),
.A2(n_1102),
.A3(n_1075),
.B(n_981),
.Y(n_1278)
);

OAI21x1_ASAP7_75t_L g1279 ( 
.A1(n_1119),
.A2(n_992),
.B(n_993),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_1166),
.Y(n_1280)
);

BUFx8_ASAP7_75t_L g1281 ( 
.A(n_1107),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1132),
.A2(n_1052),
.B(n_1058),
.Y(n_1282)
);

BUFx4_ASAP7_75t_SL g1283 ( 
.A(n_1197),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1146),
.A2(n_949),
.B(n_976),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1121),
.A2(n_988),
.B(n_963),
.Y(n_1285)
);

NOR2xp33_ASAP7_75t_L g1286 ( 
.A(n_1111),
.B(n_1072),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1178),
.B(n_1100),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1150),
.A2(n_1152),
.B(n_1141),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1210),
.B(n_1073),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1253),
.A2(n_1021),
.B(n_1023),
.Y(n_1290)
);

OR2x6_ASAP7_75t_L g1291 ( 
.A(n_1178),
.B(n_954),
.Y(n_1291)
);

OAI21x1_ASAP7_75t_L g1292 ( 
.A1(n_1154),
.A2(n_1038),
.B(n_1044),
.Y(n_1292)
);

AOI221xp5_ASAP7_75t_SL g1293 ( 
.A1(n_1224),
.A2(n_1060),
.B1(n_1022),
.B2(n_1018),
.C(n_1076),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1203),
.A2(n_1094),
.B(n_954),
.Y(n_1294)
);

CKINVDCx5p33_ASAP7_75t_R g1295 ( 
.A(n_1163),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_SL g1296 ( 
.A1(n_1204),
.A2(n_1087),
.B(n_1084),
.C(n_1092),
.Y(n_1296)
);

A2O1A1Ixp33_ASAP7_75t_L g1297 ( 
.A1(n_1202),
.A2(n_1042),
.B(n_1036),
.C(n_1080),
.Y(n_1297)
);

AO31x2_ASAP7_75t_L g1298 ( 
.A1(n_1188),
.A2(n_1149),
.A3(n_1170),
.B(n_1167),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1175),
.A2(n_1089),
.B(n_1006),
.Y(n_1299)
);

A2O1A1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1204),
.A2(n_1006),
.B(n_977),
.C(n_75),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1203),
.A2(n_67),
.B(n_70),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1116),
.B(n_1210),
.Y(n_1302)
);

BUFx3_ASAP7_75t_L g1303 ( 
.A(n_1233),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1207),
.A2(n_1125),
.B(n_1118),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1207),
.A2(n_1118),
.B(n_1216),
.Y(n_1305)
);

INVx3_ASAP7_75t_L g1306 ( 
.A(n_1252),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1216),
.A2(n_1139),
.B(n_1104),
.Y(n_1307)
);

NAND3x1_ASAP7_75t_L g1308 ( 
.A(n_1236),
.B(n_1179),
.C(n_1249),
.Y(n_1308)
);

AOI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1250),
.A2(n_1235),
.B(n_1239),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_L g1310 ( 
.A1(n_1123),
.A2(n_1135),
.B(n_1131),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1127),
.Y(n_1311)
);

NAND3x1_ASAP7_75t_L g1312 ( 
.A(n_1245),
.B(n_1190),
.C(n_1128),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1223),
.A2(n_1226),
.B(n_1160),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1244),
.B(n_1184),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1144),
.B(n_1252),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1223),
.A2(n_1206),
.B(n_1215),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_SL g1317 ( 
.A1(n_1220),
.A2(n_1228),
.B(n_1255),
.C(n_1103),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1256),
.B(n_1134),
.Y(n_1318)
);

AOI221x1_ASAP7_75t_L g1319 ( 
.A1(n_1254),
.A2(n_1260),
.B1(n_1258),
.B2(n_1247),
.C(n_1198),
.Y(n_1319)
);

NOR2xp33_ASAP7_75t_L g1320 ( 
.A(n_1137),
.B(n_1213),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1113),
.A2(n_1192),
.B(n_1189),
.C(n_1157),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_L g1322 ( 
.A1(n_1214),
.A2(n_1208),
.B(n_1205),
.Y(n_1322)
);

BUFx4f_ASAP7_75t_SL g1323 ( 
.A(n_1124),
.Y(n_1323)
);

BUFx6f_ASAP7_75t_L g1324 ( 
.A(n_1110),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1214),
.A2(n_1191),
.B(n_1222),
.Y(n_1325)
);

NOR2xp33_ASAP7_75t_L g1326 ( 
.A(n_1173),
.B(n_1164),
.Y(n_1326)
);

OR2x2_ASAP7_75t_L g1327 ( 
.A(n_1183),
.B(n_1147),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1129),
.B(n_1172),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1168),
.A2(n_1169),
.B(n_1182),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_1177),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1186),
.B(n_1138),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_SL g1332 ( 
.A(n_1133),
.B(n_1221),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1196),
.B(n_1219),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1199),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1211),
.B(n_1218),
.Y(n_1335)
);

O2A1O1Ixp33_ASAP7_75t_SL g1336 ( 
.A1(n_1235),
.A2(n_1246),
.B(n_1243),
.C(n_1239),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1225),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1195),
.B(n_1159),
.Y(n_1338)
);

AOI21xp5_ASAP7_75t_L g1339 ( 
.A1(n_1162),
.A2(n_1176),
.B(n_1250),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1231),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1110),
.Y(n_1341)
);

AOI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1243),
.A2(n_1246),
.B(n_1259),
.Y(n_1342)
);

INVx3_ASAP7_75t_L g1343 ( 
.A(n_1110),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1212),
.A2(n_1148),
.B(n_1257),
.Y(n_1344)
);

NAND2x1_ASAP7_75t_L g1345 ( 
.A(n_1185),
.B(n_1145),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_SL g1346 ( 
.A(n_1227),
.B(n_1242),
.Y(n_1346)
);

AO21x1_ASAP7_75t_L g1347 ( 
.A1(n_1237),
.A2(n_1248),
.B(n_1251),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1161),
.A2(n_1240),
.B(n_1122),
.Y(n_1348)
);

AOI221xp5_ASAP7_75t_SL g1349 ( 
.A1(n_1194),
.A2(n_1193),
.B1(n_1158),
.B2(n_1140),
.C(n_1200),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1148),
.A2(n_1161),
.B(n_1142),
.Y(n_1350)
);

OAI21xp5_ASAP7_75t_L g1351 ( 
.A1(n_1140),
.A2(n_1171),
.B(n_1229),
.Y(n_1351)
);

BUFx6f_ASAP7_75t_L g1352 ( 
.A(n_1142),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1165),
.A2(n_1185),
.B(n_1195),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1145),
.Y(n_1354)
);

AO31x2_ASAP7_75t_L g1355 ( 
.A1(n_1158),
.A2(n_1193),
.A3(n_1185),
.B(n_1227),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1142),
.Y(n_1356)
);

NAND3xp33_ASAP7_75t_L g1357 ( 
.A(n_1155),
.B(n_1241),
.C(n_1156),
.Y(n_1357)
);

OAI21x1_ASAP7_75t_L g1358 ( 
.A1(n_1209),
.A2(n_1185),
.B(n_1227),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1156),
.Y(n_1359)
);

AO31x2_ASAP7_75t_L g1360 ( 
.A1(n_1227),
.A2(n_1209),
.A3(n_1156),
.B(n_1201),
.Y(n_1360)
);

A2O1A1Ixp33_ASAP7_75t_L g1361 ( 
.A1(n_1201),
.A2(n_1234),
.B(n_1241),
.C(n_1153),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1201),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1234),
.B(n_1241),
.Y(n_1363)
);

BUFx6f_ASAP7_75t_L g1364 ( 
.A(n_1234),
.Y(n_1364)
);

AO31x2_ASAP7_75t_L g1365 ( 
.A1(n_1117),
.A2(n_985),
.A3(n_1068),
.B(n_1181),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1366)
);

OAI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1120),
.A2(n_917),
.B1(n_749),
.B2(n_1043),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1117),
.A2(n_1130),
.B(n_1175),
.Y(n_1368)
);

AOI21xp5_ASAP7_75t_L g1369 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1107),
.Y(n_1370)
);

A2O1A1Ixp33_ASAP7_75t_L g1371 ( 
.A1(n_1120),
.A2(n_917),
.B(n_937),
.C(n_948),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1373)
);

BUFx10_ASAP7_75t_L g1374 ( 
.A(n_1163),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1130),
.A2(n_1117),
.B(n_1106),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_SL g1376 ( 
.A(n_1105),
.B(n_1043),
.Y(n_1376)
);

OAI21x1_ASAP7_75t_L g1377 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1377)
);

INVx5_ASAP7_75t_L g1378 ( 
.A(n_1110),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1143),
.Y(n_1380)
);

NAND3x1_ASAP7_75t_L g1381 ( 
.A(n_1114),
.B(n_633),
.C(n_658),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1382)
);

NOR2x1_ASAP7_75t_L g1383 ( 
.A(n_1252),
.B(n_1111),
.Y(n_1383)
);

AO21x2_ASAP7_75t_L g1384 ( 
.A1(n_1130),
.A2(n_1181),
.B(n_1135),
.Y(n_1384)
);

A2O1A1Ixp33_ASAP7_75t_L g1385 ( 
.A1(n_1120),
.A2(n_917),
.B(n_937),
.C(n_948),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1116),
.B(n_749),
.Y(n_1386)
);

AO31x2_ASAP7_75t_L g1387 ( 
.A1(n_1117),
.A2(n_985),
.A3(n_1068),
.B(n_1181),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1116),
.B(n_749),
.Y(n_1388)
);

AOI21xp5_ASAP7_75t_L g1389 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1389)
);

CKINVDCx5p33_ASAP7_75t_R g1390 ( 
.A(n_1163),
.Y(n_1390)
);

O2A1O1Ixp5_ASAP7_75t_SL g1391 ( 
.A1(n_1157),
.A2(n_566),
.B(n_1151),
.C(n_1162),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1116),
.B(n_749),
.Y(n_1392)
);

AOI21xp5_ASAP7_75t_L g1393 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1393)
);

O2A1O1Ixp33_ASAP7_75t_SL g1394 ( 
.A1(n_1217),
.A2(n_1029),
.B(n_1204),
.C(n_1188),
.Y(n_1394)
);

INVx1_ASAP7_75t_SL g1395 ( 
.A(n_1111),
.Y(n_1395)
);

AO32x2_ASAP7_75t_L g1396 ( 
.A1(n_1247),
.A2(n_860),
.A3(n_1140),
.B1(n_812),
.B2(n_905),
.Y(n_1396)
);

AOI21xp5_ASAP7_75t_L g1397 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1397)
);

INVx3_ASAP7_75t_SL g1398 ( 
.A(n_1197),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1105),
.B(n_1043),
.Y(n_1399)
);

AOI21xp5_ASAP7_75t_L g1400 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1400)
);

AOI21xp5_ASAP7_75t_L g1401 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1112),
.Y(n_1402)
);

OAI21x1_ASAP7_75t_L g1403 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1403)
);

O2A1O1Ixp33_ASAP7_75t_L g1404 ( 
.A1(n_1105),
.A2(n_1043),
.B(n_917),
.C(n_804),
.Y(n_1404)
);

AOI21xp5_ASAP7_75t_L g1405 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1112),
.Y(n_1406)
);

AOI21xp5_ASAP7_75t_L g1407 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1120),
.A2(n_1043),
.B1(n_761),
.B2(n_1065),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1130),
.A2(n_749),
.B(n_917),
.Y(n_1409)
);

A2O1A1Ixp33_ASAP7_75t_L g1410 ( 
.A1(n_1120),
.A2(n_917),
.B(n_937),
.C(n_948),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1112),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1120),
.A2(n_917),
.B(n_937),
.C(n_948),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1210),
.B(n_917),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1112),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1415)
);

NOR2x1_ASAP7_75t_R g1416 ( 
.A(n_1163),
.B(n_685),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1120),
.A2(n_1105),
.B1(n_1114),
.B2(n_1065),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1105),
.B(n_1043),
.Y(n_1418)
);

O2A1O1Ixp33_ASAP7_75t_L g1419 ( 
.A1(n_1105),
.A2(n_1043),
.B(n_917),
.C(n_804),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1112),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1108),
.A2(n_1106),
.B(n_1010),
.Y(n_1421)
);

CKINVDCx16_ASAP7_75t_R g1422 ( 
.A(n_1374),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1261),
.B2(n_1367),
.Y(n_1423)
);

CKINVDCx11_ASAP7_75t_R g1424 ( 
.A(n_1374),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_1367),
.B2(n_1399),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1413),
.B(n_1371),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1418),
.A2(n_1346),
.B1(n_1338),
.B2(n_1266),
.Y(n_1427)
);

AOI22xp33_ASAP7_75t_L g1428 ( 
.A1(n_1376),
.A2(n_1346),
.B1(n_1347),
.B2(n_1331),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1385),
.A2(n_1410),
.B1(n_1412),
.B2(n_1388),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1323),
.Y(n_1430)
);

AOI22xp5_ASAP7_75t_L g1431 ( 
.A1(n_1381),
.A2(n_1312),
.B1(n_1320),
.B2(n_1326),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1311),
.Y(n_1432)
);

INVx6_ASAP7_75t_L g1433 ( 
.A(n_1281),
.Y(n_1433)
);

OAI21xp5_ASAP7_75t_SL g1434 ( 
.A1(n_1404),
.A2(n_1419),
.B(n_1319),
.Y(n_1434)
);

INVxp67_ASAP7_75t_SL g1435 ( 
.A(n_1302),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1280),
.Y(n_1436)
);

BUFx4f_ASAP7_75t_SL g1437 ( 
.A(n_1281),
.Y(n_1437)
);

OAI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1386),
.A2(n_1392),
.B1(n_1388),
.B2(n_1266),
.Y(n_1438)
);

OAI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1386),
.A2(n_1392),
.B1(n_1302),
.B2(n_1327),
.Y(n_1439)
);

BUFx10_ASAP7_75t_L g1440 ( 
.A(n_1295),
.Y(n_1440)
);

OAI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1318),
.A2(n_1357),
.B1(n_1289),
.B2(n_1276),
.Y(n_1441)
);

OAI21xp5_ASAP7_75t_SL g1442 ( 
.A1(n_1321),
.A2(n_1353),
.B(n_1301),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1308),
.A2(n_1332),
.B1(n_1272),
.B2(n_1314),
.Y(n_1443)
);

OAI21xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1353),
.A2(n_1273),
.B(n_1351),
.Y(n_1444)
);

BUFx2_ASAP7_75t_SL g1445 ( 
.A(n_1303),
.Y(n_1445)
);

CKINVDCx11_ASAP7_75t_R g1446 ( 
.A(n_1398),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1380),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_L g1448 ( 
.A1(n_1351),
.A2(n_1262),
.B1(n_1318),
.B2(n_1379),
.Y(n_1448)
);

INVx4_ASAP7_75t_L g1449 ( 
.A(n_1378),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1357),
.A2(n_1284),
.B1(n_1396),
.B2(n_1286),
.Y(n_1450)
);

INVx6_ASAP7_75t_L g1451 ( 
.A(n_1378),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_L g1452 ( 
.A1(n_1395),
.A2(n_1315),
.B1(n_1269),
.B2(n_1370),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1276),
.A2(n_1402),
.B1(n_1411),
.B2(n_1414),
.Y(n_1453)
);

BUFx3_ASAP7_75t_L g1454 ( 
.A(n_1330),
.Y(n_1454)
);

CKINVDCx11_ASAP7_75t_R g1455 ( 
.A(n_1283),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1366),
.A2(n_1382),
.B1(n_1393),
.B2(n_1397),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1390),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1369),
.A2(n_1407),
.B1(n_1389),
.B2(n_1401),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1406),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1315),
.A2(n_1420),
.B1(n_1291),
.B2(n_1383),
.Y(n_1460)
);

CKINVDCx11_ASAP7_75t_R g1461 ( 
.A(n_1416),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1400),
.A2(n_1409),
.B1(n_1405),
.B2(n_1344),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1324),
.Y(n_1463)
);

CKINVDCx20_ASAP7_75t_R g1464 ( 
.A(n_1363),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1349),
.A2(n_1291),
.B1(n_1361),
.B2(n_1339),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1334),
.A2(n_1337),
.B1(n_1340),
.B2(n_1305),
.Y(n_1466)
);

AOI22xp33_ASAP7_75t_SL g1467 ( 
.A1(n_1396),
.A2(n_1265),
.B1(n_1349),
.B2(n_1394),
.Y(n_1467)
);

INVx4_ASAP7_75t_L g1468 ( 
.A(n_1324),
.Y(n_1468)
);

OAI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1333),
.A2(n_1335),
.B1(n_1291),
.B2(n_1396),
.Y(n_1469)
);

OAI22xp5_ASAP7_75t_L g1470 ( 
.A1(n_1265),
.A2(n_1300),
.B1(n_1333),
.B2(n_1335),
.Y(n_1470)
);

INVx3_ASAP7_75t_L g1471 ( 
.A(n_1360),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1354),
.Y(n_1472)
);

INVx6_ASAP7_75t_L g1473 ( 
.A(n_1341),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_SL g1474 ( 
.A1(n_1384),
.A2(n_1355),
.B1(n_1329),
.B2(n_1358),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1362),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1348),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1343),
.Y(n_1477)
);

BUFx12f_ASAP7_75t_L g1478 ( 
.A(n_1341),
.Y(n_1478)
);

INVx6_ASAP7_75t_L g1479 ( 
.A(n_1341),
.Y(n_1479)
);

OAI21xp33_ASAP7_75t_SL g1480 ( 
.A1(n_1391),
.A2(n_1316),
.B(n_1313),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1307),
.A2(n_1342),
.B1(n_1309),
.B2(n_1310),
.Y(n_1481)
);

OAI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1350),
.A2(n_1277),
.B1(n_1306),
.B2(n_1322),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1306),
.A2(n_1304),
.B1(n_1345),
.B2(n_1294),
.Y(n_1483)
);

OAI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1275),
.A2(n_1285),
.B1(n_1325),
.B2(n_1329),
.Y(n_1484)
);

OAI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1356),
.A2(n_1359),
.B1(n_1282),
.B2(n_1368),
.Y(n_1485)
);

AOI22x1_ASAP7_75t_SL g1486 ( 
.A1(n_1359),
.A2(n_1355),
.B1(n_1317),
.B2(n_1336),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1264),
.A2(n_1384),
.B1(n_1299),
.B2(n_1270),
.Y(n_1487)
);

BUFx2_ASAP7_75t_SL g1488 ( 
.A(n_1352),
.Y(n_1488)
);

CKINVDCx6p67_ASAP7_75t_R g1489 ( 
.A(n_1364),
.Y(n_1489)
);

BUFx2_ASAP7_75t_R g1490 ( 
.A(n_1293),
.Y(n_1490)
);

INVx2_ASAP7_75t_L g1491 ( 
.A(n_1364),
.Y(n_1491)
);

AOI22xp33_ASAP7_75t_SL g1492 ( 
.A1(n_1368),
.A2(n_1288),
.B1(n_1299),
.B2(n_1293),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1365),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1365),
.Y(n_1494)
);

OAI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1375),
.A2(n_1387),
.B1(n_1296),
.B2(n_1298),
.Y(n_1495)
);

BUFx3_ASAP7_75t_L g1496 ( 
.A(n_1278),
.Y(n_1496)
);

OAI21xp5_ASAP7_75t_SL g1497 ( 
.A1(n_1297),
.A2(n_1298),
.B(n_1387),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1290),
.A2(n_1421),
.B1(n_1415),
.B2(n_1372),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_SL g1499 ( 
.A1(n_1373),
.A2(n_1377),
.B1(n_1403),
.B2(n_1263),
.Y(n_1499)
);

BUFx3_ASAP7_75t_L g1500 ( 
.A(n_1279),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1292),
.A2(n_1274),
.B1(n_1268),
.B2(n_1267),
.Y(n_1501)
);

BUFx3_ASAP7_75t_L g1502 ( 
.A(n_1267),
.Y(n_1502)
);

INVx6_ASAP7_75t_L g1503 ( 
.A(n_1281),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_SL g1505 ( 
.A1(n_1399),
.A2(n_1109),
.B1(n_761),
.B2(n_632),
.Y(n_1505)
);

CKINVDCx11_ASAP7_75t_R g1506 ( 
.A(n_1374),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1507)
);

CKINVDCx6p67_ASAP7_75t_R g1508 ( 
.A(n_1398),
.Y(n_1508)
);

BUFx4f_ASAP7_75t_SL g1509 ( 
.A(n_1281),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1417),
.A2(n_750),
.B1(n_747),
.B2(n_1043),
.Y(n_1510)
);

CKINVDCx20_ASAP7_75t_R g1511 ( 
.A(n_1323),
.Y(n_1511)
);

INVx3_ASAP7_75t_L g1512 ( 
.A(n_1360),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1328),
.Y(n_1513)
);

OAI22xp5_ASAP7_75t_L g1514 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1514)
);

AND2x4_ASAP7_75t_L g1515 ( 
.A(n_1287),
.B(n_1178),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1367),
.B(n_917),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1271),
.Y(n_1517)
);

INVx2_ASAP7_75t_L g1518 ( 
.A(n_1271),
.Y(n_1518)
);

CKINVDCx11_ASAP7_75t_R g1519 ( 
.A(n_1374),
.Y(n_1519)
);

CKINVDCx11_ASAP7_75t_R g1520 ( 
.A(n_1374),
.Y(n_1520)
);

AOI22xp33_ASAP7_75t_L g1521 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1399),
.A2(n_1109),
.B1(n_761),
.B2(n_632),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1523)
);

AOI21xp33_ASAP7_75t_L g1524 ( 
.A1(n_1417),
.A2(n_969),
.B(n_968),
.Y(n_1524)
);

INVx2_ASAP7_75t_SL g1525 ( 
.A(n_1303),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1328),
.Y(n_1526)
);

OAI22xp5_ASAP7_75t_L g1527 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1528)
);

INVx6_ASAP7_75t_L g1529 ( 
.A(n_1281),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1367),
.B(n_917),
.Y(n_1530)
);

BUFx2_ASAP7_75t_L g1531 ( 
.A(n_1370),
.Y(n_1531)
);

AOI22xp33_ASAP7_75t_L g1532 ( 
.A1(n_1417),
.A2(n_1114),
.B1(n_1043),
.B2(n_1408),
.Y(n_1532)
);

INVx6_ASAP7_75t_L g1533 ( 
.A(n_1281),
.Y(n_1533)
);

INVx1_ASAP7_75t_SL g1534 ( 
.A(n_1395),
.Y(n_1534)
);

OAI22xp5_ASAP7_75t_L g1535 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1535)
);

CKINVDCx11_ASAP7_75t_R g1536 ( 
.A(n_1374),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1537)
);

OAI21xp5_ASAP7_75t_SL g1538 ( 
.A1(n_1417),
.A2(n_750),
.B(n_747),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1328),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1271),
.Y(n_1540)
);

INVx2_ASAP7_75t_SL g1541 ( 
.A(n_1303),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1367),
.B(n_917),
.Y(n_1542)
);

INVx6_ASAP7_75t_L g1543 ( 
.A(n_1281),
.Y(n_1543)
);

CKINVDCx11_ASAP7_75t_R g1544 ( 
.A(n_1374),
.Y(n_1544)
);

OAI22xp33_ASAP7_75t_L g1545 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_1109),
.B2(n_1367),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1328),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1417),
.A2(n_1261),
.B1(n_632),
.B2(n_1367),
.Y(n_1549)
);

BUFx8_ASAP7_75t_L g1550 ( 
.A(n_1314),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_SL g1551 ( 
.A1(n_1399),
.A2(n_1109),
.B1(n_761),
.B2(n_632),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1408),
.A2(n_1417),
.B1(n_1043),
.B2(n_1261),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1328),
.Y(n_1553)
);

AOI22xp33_ASAP7_75t_SL g1554 ( 
.A1(n_1399),
.A2(n_1109),
.B1(n_761),
.B2(n_632),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1328),
.Y(n_1555)
);

NAND2x1_ASAP7_75t_L g1556 ( 
.A(n_1306),
.B(n_953),
.Y(n_1556)
);

CKINVDCx11_ASAP7_75t_R g1557 ( 
.A(n_1374),
.Y(n_1557)
);

BUFx2_ASAP7_75t_L g1558 ( 
.A(n_1370),
.Y(n_1558)
);

BUFx4f_ASAP7_75t_SL g1559 ( 
.A(n_1281),
.Y(n_1559)
);

CKINVDCx20_ASAP7_75t_R g1560 ( 
.A(n_1323),
.Y(n_1560)
);

INVx2_ASAP7_75t_SL g1561 ( 
.A(n_1303),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1516),
.B(n_1530),
.Y(n_1562)
);

BUFx3_ASAP7_75t_L g1563 ( 
.A(n_1478),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1432),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1493),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1494),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1502),
.Y(n_1567)
);

OR2x6_ASAP7_75t_L g1568 ( 
.A(n_1497),
.B(n_1442),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1471),
.Y(n_1569)
);

INVx2_ASAP7_75t_SL g1570 ( 
.A(n_1451),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1450),
.B(n_1467),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1459),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1531),
.Y(n_1573)
);

AOI21x1_ASAP7_75t_L g1574 ( 
.A1(n_1482),
.A2(n_1483),
.B(n_1429),
.Y(n_1574)
);

OAI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1498),
.A2(n_1501),
.B(n_1458),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1512),
.Y(n_1576)
);

OR2x6_ASAP7_75t_L g1577 ( 
.A(n_1444),
.B(n_1496),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1450),
.B(n_1467),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1453),
.Y(n_1579)
);

AOI21x1_ASAP7_75t_L g1580 ( 
.A1(n_1542),
.A2(n_1470),
.B(n_1426),
.Y(n_1580)
);

INVx3_ASAP7_75t_L g1581 ( 
.A(n_1500),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1453),
.Y(n_1582)
);

OA21x2_ASAP7_75t_L g1583 ( 
.A1(n_1456),
.A2(n_1458),
.B(n_1487),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1476),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1469),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1534),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1435),
.B(n_1448),
.Y(n_1587)
);

OAI21x1_ASAP7_75t_L g1588 ( 
.A1(n_1498),
.A2(n_1501),
.B(n_1456),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1469),
.Y(n_1589)
);

OAI21x1_ASAP7_75t_L g1590 ( 
.A1(n_1462),
.A2(n_1466),
.B(n_1448),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1455),
.Y(n_1591)
);

AND2x4_ASAP7_75t_L g1592 ( 
.A(n_1465),
.B(n_1435),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1439),
.B(n_1423),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1495),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1495),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1439),
.B(n_1441),
.Y(n_1596)
);

A2O1A1Ixp33_ASAP7_75t_L g1597 ( 
.A1(n_1538),
.A2(n_1510),
.B(n_1524),
.C(n_1425),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1464),
.B(n_1443),
.Y(n_1598)
);

INVx1_ASAP7_75t_SL g1599 ( 
.A(n_1558),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1486),
.Y(n_1600)
);

OAI21x1_ASAP7_75t_L g1601 ( 
.A1(n_1462),
.A2(n_1466),
.B(n_1460),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1545),
.A2(n_1535),
.B(n_1537),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1485),
.Y(n_1603)
);

NAND2xp33_ASAP7_75t_R g1604 ( 
.A(n_1515),
.B(n_1477),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1513),
.Y(n_1605)
);

INVx1_ASAP7_75t_SL g1606 ( 
.A(n_1445),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1485),
.Y(n_1607)
);

OAI21xp33_ASAP7_75t_SL g1608 ( 
.A1(n_1504),
.A2(n_1507),
.B(n_1549),
.Y(n_1608)
);

OAI21x1_ASAP7_75t_L g1609 ( 
.A1(n_1434),
.A2(n_1452),
.B(n_1428),
.Y(n_1609)
);

BUFx3_ASAP7_75t_L g1610 ( 
.A(n_1463),
.Y(n_1610)
);

INVx3_ASAP7_75t_L g1611 ( 
.A(n_1526),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1481),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1481),
.Y(n_1613)
);

OAI21x1_ASAP7_75t_L g1614 ( 
.A1(n_1539),
.A2(n_1555),
.B(n_1553),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1548),
.Y(n_1615)
);

INVxp67_ASAP7_75t_L g1616 ( 
.A(n_1525),
.Y(n_1616)
);

A2O1A1Ixp33_ASAP7_75t_L g1617 ( 
.A1(n_1425),
.A2(n_1427),
.B(n_1514),
.C(n_1552),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1492),
.Y(n_1618)
);

OAI21x1_ASAP7_75t_L g1619 ( 
.A1(n_1499),
.A2(n_1475),
.B(n_1528),
.Y(n_1619)
);

AND2x4_ASAP7_75t_L g1620 ( 
.A(n_1436),
.B(n_1447),
.Y(n_1620)
);

OAI21x1_ASAP7_75t_L g1621 ( 
.A1(n_1499),
.A2(n_1549),
.B(n_1504),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1492),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1507),
.B(n_1521),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1474),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1523),
.B(n_1527),
.Y(n_1625)
);

INVx2_ASAP7_75t_L g1626 ( 
.A(n_1517),
.Y(n_1626)
);

AO21x2_ASAP7_75t_L g1627 ( 
.A1(n_1484),
.A2(n_1438),
.B(n_1545),
.Y(n_1627)
);

INVx1_ASAP7_75t_L g1628 ( 
.A(n_1474),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1546),
.B(n_1433),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1521),
.B(n_1528),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1433),
.B(n_1503),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1480),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1484),
.Y(n_1633)
);

HB1xp67_ASAP7_75t_L g1634 ( 
.A(n_1472),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1441),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1518),
.Y(n_1636)
);

INVxp67_ASAP7_75t_L g1637 ( 
.A(n_1541),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1540),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1438),
.Y(n_1639)
);

BUFx3_ASAP7_75t_L g1640 ( 
.A(n_1550),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1532),
.B(n_1427),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1515),
.B(n_1431),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1547),
.B(n_1505),
.Y(n_1644)
);

AO31x2_ASAP7_75t_L g1645 ( 
.A1(n_1490),
.A2(n_1554),
.A3(n_1522),
.B(n_1551),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1491),
.Y(n_1646)
);

AND2x2_ASAP7_75t_L g1647 ( 
.A(n_1522),
.B(n_1554),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1550),
.Y(n_1648)
);

OA21x2_ASAP7_75t_L g1649 ( 
.A1(n_1561),
.A2(n_1556),
.B(n_1449),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1433),
.B(n_1503),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1422),
.B(n_1468),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1488),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1473),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1489),
.A2(n_1479),
.B(n_1533),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1503),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1529),
.Y(n_1656)
);

INVx4_ASAP7_75t_L g1657 ( 
.A(n_1529),
.Y(n_1657)
);

BUFx2_ASAP7_75t_L g1658 ( 
.A(n_1529),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1533),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1533),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_L g1661 ( 
.A(n_1543),
.B(n_1508),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1454),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1543),
.Y(n_1663)
);

AOI21x1_ASAP7_75t_L g1664 ( 
.A1(n_1543),
.A2(n_1509),
.B(n_1559),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1440),
.B(n_1424),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1437),
.A2(n_1559),
.B1(n_1509),
.B2(n_1511),
.Y(n_1666)
);

INVx1_ASAP7_75t_SL g1667 ( 
.A(n_1457),
.Y(n_1667)
);

AO21x2_ASAP7_75t_L g1668 ( 
.A1(n_1632),
.A2(n_1437),
.B(n_1519),
.Y(n_1668)
);

INVx2_ASAP7_75t_SL g1669 ( 
.A(n_1573),
.Y(n_1669)
);

INVx5_ASAP7_75t_L g1670 ( 
.A(n_1631),
.Y(n_1670)
);

A2O1A1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1597),
.A2(n_1430),
.B(n_1560),
.C(n_1536),
.Y(n_1671)
);

A2O1A1Ixp33_ASAP7_75t_L g1672 ( 
.A1(n_1617),
.A2(n_1557),
.B(n_1506),
.C(n_1520),
.Y(n_1672)
);

AO32x2_ASAP7_75t_L g1673 ( 
.A1(n_1570),
.A2(n_1544),
.A3(n_1446),
.B1(n_1440),
.B2(n_1461),
.Y(n_1673)
);

AOI22xp5_ASAP7_75t_L g1674 ( 
.A1(n_1602),
.A2(n_1625),
.B1(n_1641),
.B2(n_1629),
.Y(n_1674)
);

OAI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1580),
.A2(n_1590),
.B(n_1609),
.Y(n_1675)
);

OA21x2_ASAP7_75t_L g1676 ( 
.A1(n_1575),
.A2(n_1588),
.B(n_1609),
.Y(n_1676)
);

A2O1A1Ixp33_ASAP7_75t_L g1677 ( 
.A1(n_1608),
.A2(n_1596),
.B(n_1593),
.C(n_1598),
.Y(n_1677)
);

NAND4xp25_ASAP7_75t_L g1678 ( 
.A(n_1562),
.B(n_1635),
.C(n_1596),
.D(n_1633),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_SL g1679 ( 
.A(n_1568),
.B(n_1577),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1573),
.Y(n_1680)
);

AOI221x1_ASAP7_75t_SL g1681 ( 
.A1(n_1635),
.A2(n_1643),
.B1(n_1589),
.B2(n_1585),
.C(n_1639),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1565),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1644),
.A2(n_1647),
.B1(n_1593),
.B2(n_1623),
.Y(n_1683)
);

A2O1A1Ixp33_ASAP7_75t_L g1684 ( 
.A1(n_1590),
.A2(n_1601),
.B(n_1621),
.C(n_1644),
.Y(n_1684)
);

AOI221xp5_ASAP7_75t_L g1685 ( 
.A1(n_1647),
.A2(n_1630),
.B1(n_1623),
.B2(n_1633),
.C(n_1639),
.Y(n_1685)
);

OR2x2_ASAP7_75t_L g1686 ( 
.A(n_1589),
.B(n_1564),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1583),
.A2(n_1627),
.B(n_1601),
.Y(n_1687)
);

OAI21xp5_ASAP7_75t_L g1688 ( 
.A1(n_1580),
.A2(n_1574),
.B(n_1621),
.Y(n_1688)
);

AOI22xp5_ASAP7_75t_L g1689 ( 
.A1(n_1629),
.A2(n_1600),
.B1(n_1592),
.B2(n_1642),
.Y(n_1689)
);

A2O1A1Ixp33_ASAP7_75t_L g1690 ( 
.A1(n_1630),
.A2(n_1571),
.B(n_1578),
.C(n_1600),
.Y(n_1690)
);

AOI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1583),
.A2(n_1627),
.B(n_1612),
.Y(n_1691)
);

OAI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1571),
.A2(n_1578),
.B1(n_1592),
.B2(n_1629),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1574),
.A2(n_1575),
.B(n_1588),
.Y(n_1693)
);

AND2x2_ASAP7_75t_SL g1694 ( 
.A(n_1583),
.B(n_1592),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1632),
.A2(n_1595),
.B(n_1594),
.Y(n_1695)
);

OAI22xp5_ASAP7_75t_L g1696 ( 
.A1(n_1629),
.A2(n_1582),
.B1(n_1579),
.B2(n_1586),
.Y(n_1696)
);

OAI21xp5_ASAP7_75t_L g1697 ( 
.A1(n_1612),
.A2(n_1613),
.B(n_1582),
.Y(n_1697)
);

O2A1O1Ixp33_ASAP7_75t_SL g1698 ( 
.A1(n_1606),
.A2(n_1591),
.B(n_1661),
.C(n_1651),
.Y(n_1698)
);

AO21x1_ASAP7_75t_L g1699 ( 
.A1(n_1604),
.A2(n_1567),
.B(n_1579),
.Y(n_1699)
);

A2O1A1Ixp33_ASAP7_75t_L g1700 ( 
.A1(n_1613),
.A2(n_1587),
.B(n_1628),
.C(n_1624),
.Y(n_1700)
);

NOR2x1_ASAP7_75t_SL g1701 ( 
.A(n_1650),
.B(n_1627),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_L g1702 ( 
.A(n_1599),
.B(n_1618),
.C(n_1622),
.D(n_1603),
.Y(n_1702)
);

OAI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1583),
.A2(n_1619),
.B(n_1614),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1572),
.B(n_1634),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1611),
.B(n_1638),
.Y(n_1705)
);

CKINVDCx5p33_ASAP7_75t_R g1706 ( 
.A(n_1666),
.Y(n_1706)
);

AOI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1614),
.A2(n_1615),
.B(n_1605),
.Y(n_1707)
);

NAND2xp33_ASAP7_75t_L g1708 ( 
.A(n_1665),
.B(n_1656),
.Y(n_1708)
);

OR2x6_ASAP7_75t_L g1709 ( 
.A(n_1650),
.B(n_1619),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1607),
.A2(n_1628),
.B(n_1624),
.Y(n_1710)
);

A2O1A1Ixp33_ASAP7_75t_L g1711 ( 
.A1(n_1607),
.A2(n_1618),
.B(n_1622),
.C(n_1648),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1615),
.B(n_1611),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1565),
.Y(n_1713)
);

A2O1A1Ixp33_ASAP7_75t_L g1714 ( 
.A1(n_1640),
.A2(n_1648),
.B(n_1655),
.C(n_1663),
.Y(n_1714)
);

A2O1A1Ixp33_ASAP7_75t_L g1715 ( 
.A1(n_1640),
.A2(n_1655),
.B(n_1663),
.C(n_1660),
.Y(n_1715)
);

OAI21xp5_ASAP7_75t_L g1716 ( 
.A1(n_1620),
.A2(n_1654),
.B(n_1616),
.Y(n_1716)
);

AOI22xp5_ASAP7_75t_L g1717 ( 
.A1(n_1660),
.A2(n_1656),
.B1(n_1662),
.B2(n_1659),
.Y(n_1717)
);

CKINVDCx20_ASAP7_75t_R g1718 ( 
.A(n_1667),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1566),
.Y(n_1719)
);

A2O1A1Ixp33_ASAP7_75t_L g1720 ( 
.A1(n_1658),
.A2(n_1637),
.B(n_1563),
.C(n_1652),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1581),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1698),
.B(n_1706),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1716),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1682),
.Y(n_1724)
);

HB1xp67_ASAP7_75t_L g1725 ( 
.A(n_1682),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1713),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1719),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1716),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1707),
.Y(n_1729)
);

AOI22xp33_ASAP7_75t_L g1730 ( 
.A1(n_1674),
.A2(n_1658),
.B1(n_1659),
.B2(n_1657),
.Y(n_1730)
);

CKINVDCx5p33_ASAP7_75t_R g1731 ( 
.A(n_1718),
.Y(n_1731)
);

OR2x2_ASAP7_75t_SL g1732 ( 
.A(n_1676),
.B(n_1649),
.Y(n_1732)
);

INVx2_ASAP7_75t_SL g1733 ( 
.A(n_1670),
.Y(n_1733)
);

AND2x4_ASAP7_75t_L g1734 ( 
.A(n_1709),
.B(n_1581),
.Y(n_1734)
);

HB1xp67_ASAP7_75t_L g1735 ( 
.A(n_1695),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1694),
.B(n_1569),
.Y(n_1736)
);

AOI22xp33_ASAP7_75t_L g1737 ( 
.A1(n_1678),
.A2(n_1659),
.B1(n_1657),
.B2(n_1665),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1697),
.B(n_1704),
.Y(n_1738)
);

NOR2x1_ASAP7_75t_L g1739 ( 
.A(n_1668),
.B(n_1720),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1680),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1694),
.B(n_1576),
.Y(n_1741)
);

BUFx3_ASAP7_75t_L g1742 ( 
.A(n_1668),
.Y(n_1742)
);

HB1xp67_ASAP7_75t_L g1743 ( 
.A(n_1695),
.Y(n_1743)
);

OAI222xp33_ASAP7_75t_L g1744 ( 
.A1(n_1683),
.A2(n_1664),
.B1(n_1645),
.B2(n_1646),
.C1(n_1636),
.C2(n_1626),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1676),
.B(n_1569),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1703),
.B(n_1576),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1703),
.B(n_1584),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1712),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1684),
.B(n_1584),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1712),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1693),
.B(n_1687),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1707),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1726),
.Y(n_1753)
);

OR2x2_ASAP7_75t_L g1754 ( 
.A(n_1723),
.B(n_1691),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1725),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1739),
.A2(n_1672),
.B1(n_1671),
.B2(n_1677),
.C(n_1690),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_1701),
.Y(n_1757)
);

OAI22xp5_ASAP7_75t_L g1758 ( 
.A1(n_1722),
.A2(n_1685),
.B1(n_1683),
.B2(n_1700),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1726),
.Y(n_1759)
);

NOR2xp33_ASAP7_75t_L g1760 ( 
.A(n_1738),
.B(n_1669),
.Y(n_1760)
);

AND2x2_ASAP7_75t_L g1761 ( 
.A(n_1736),
.B(n_1675),
.Y(n_1761)
);

NAND4xp25_ASAP7_75t_L g1762 ( 
.A(n_1739),
.B(n_1681),
.C(n_1685),
.D(n_1691),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

OAI33xp33_ASAP7_75t_L g1764 ( 
.A1(n_1724),
.A2(n_1696),
.A3(n_1702),
.B1(n_1692),
.B2(n_1686),
.B3(n_1681),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1735),
.Y(n_1765)
);

INVx2_ASAP7_75t_L g1766 ( 
.A(n_1745),
.Y(n_1766)
);

OR2x6_ASAP7_75t_L g1767 ( 
.A(n_1733),
.B(n_1734),
.Y(n_1767)
);

OAI31xp33_ASAP7_75t_L g1768 ( 
.A1(n_1744),
.A2(n_1711),
.A3(n_1692),
.B(n_1696),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1732),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1736),
.B(n_1688),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1741),
.B(n_1688),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1741),
.B(n_1723),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_SL g1773 ( 
.A(n_1742),
.B(n_1699),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1731),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1728),
.B(n_1705),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1748),
.B(n_1710),
.Y(n_1776)
);

NAND4xp25_ASAP7_75t_L g1777 ( 
.A(n_1737),
.B(n_1717),
.C(n_1714),
.D(n_1689),
.Y(n_1777)
);

INVx1_ASAP7_75t_L g1778 ( 
.A(n_1724),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1732),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1734),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1746),
.Y(n_1781)
);

AOI21xp5_ASAP7_75t_L g1782 ( 
.A1(n_1729),
.A2(n_1670),
.B(n_1679),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1746),
.Y(n_1783)
);

BUFx6f_ASAP7_75t_L g1784 ( 
.A(n_1751),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1746),
.Y(n_1785)
);

NOR3xp33_ASAP7_75t_SL g1786 ( 
.A(n_1744),
.B(n_1715),
.C(n_1653),
.Y(n_1786)
);

HB1xp67_ASAP7_75t_L g1787 ( 
.A(n_1725),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1781),
.B(n_1735),
.Y(n_1788)
);

BUFx3_ASAP7_75t_L g1789 ( 
.A(n_1769),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1781),
.B(n_1743),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1766),
.Y(n_1791)
);

BUFx3_ASAP7_75t_L g1792 ( 
.A(n_1769),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1776),
.B(n_1748),
.Y(n_1794)
);

INVxp67_ASAP7_75t_L g1795 ( 
.A(n_1773),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1776),
.B(n_1750),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1783),
.B(n_1743),
.Y(n_1797)
);

NAND3x1_ASAP7_75t_L g1798 ( 
.A(n_1768),
.B(n_1664),
.C(n_1673),
.Y(n_1798)
);

AND2x2_ASAP7_75t_L g1799 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1766),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1766),
.Y(n_1801)
);

NAND2x1p5_ASAP7_75t_L g1802 ( 
.A(n_1773),
.B(n_1670),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1753),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1753),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1755),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1767),
.B(n_1734),
.Y(n_1807)
);

AND2x4_ASAP7_75t_L g1808 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1783),
.B(n_1749),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1759),
.Y(n_1810)
);

INVxp67_ASAP7_75t_SL g1811 ( 
.A(n_1765),
.Y(n_1811)
);

AND2x4_ASAP7_75t_L g1812 ( 
.A(n_1767),
.B(n_1721),
.Y(n_1812)
);

OR2x2_ASAP7_75t_L g1813 ( 
.A(n_1785),
.B(n_1729),
.Y(n_1813)
);

HB1xp67_ASAP7_75t_L g1814 ( 
.A(n_1755),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1759),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1759),
.Y(n_1816)
);

AND2x2_ASAP7_75t_L g1817 ( 
.A(n_1780),
.B(n_1769),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1763),
.Y(n_1818)
);

HB1xp67_ASAP7_75t_L g1819 ( 
.A(n_1787),
.Y(n_1819)
);

AND2x2_ASAP7_75t_SL g1820 ( 
.A(n_1754),
.B(n_1772),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1747),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1793),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1793),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1795),
.Y(n_1824)
);

INVxp67_ASAP7_75t_SL g1825 ( 
.A(n_1795),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1803),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1803),
.Y(n_1827)
);

NOR2x1_ASAP7_75t_L g1828 ( 
.A(n_1789),
.B(n_1762),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1820),
.B(n_1780),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1804),
.Y(n_1830)
);

NOR2xp33_ASAP7_75t_L g1831 ( 
.A(n_1794),
.B(n_1774),
.Y(n_1831)
);

AOI21xp5_ASAP7_75t_L g1832 ( 
.A1(n_1802),
.A2(n_1756),
.B(n_1768),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1791),
.Y(n_1833)
);

INVxp67_ASAP7_75t_L g1834 ( 
.A(n_1789),
.Y(n_1834)
);

INVx5_ASAP7_75t_L g1835 ( 
.A(n_1789),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1791),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

INVx2_ASAP7_75t_L g1838 ( 
.A(n_1791),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1810),
.Y(n_1839)
);

OR2x2_ASAP7_75t_L g1840 ( 
.A(n_1794),
.B(n_1754),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1820),
.B(n_1772),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1820),
.B(n_1817),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1791),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1800),
.Y(n_1844)
);

OR2x2_ASAP7_75t_L g1845 ( 
.A(n_1796),
.B(n_1754),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1800),
.Y(n_1846)
);

NAND2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1789),
.B(n_1742),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_SL g1848 ( 
.A(n_1820),
.B(n_1768),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1810),
.Y(n_1849)
);

INVx2_ASAP7_75t_SL g1850 ( 
.A(n_1792),
.Y(n_1850)
);

AND2x2_ASAP7_75t_L g1851 ( 
.A(n_1817),
.B(n_1772),
.Y(n_1851)
);

OR2x2_ASAP7_75t_L g1852 ( 
.A(n_1796),
.B(n_1775),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1817),
.B(n_1808),
.Y(n_1853)
);

INVx2_ASAP7_75t_SL g1854 ( 
.A(n_1792),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1800),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1808),
.B(n_1757),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1815),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1815),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1800),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1801),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1805),
.B(n_1778),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1816),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1798),
.A2(n_1756),
.B1(n_1758),
.B2(n_1786),
.Y(n_1863)
);

INVxp67_ASAP7_75t_SL g1864 ( 
.A(n_1802),
.Y(n_1864)
);

NOR2xp33_ASAP7_75t_L g1865 ( 
.A(n_1808),
.B(n_1774),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1816),
.Y(n_1866)
);

INVxp67_ASAP7_75t_L g1867 ( 
.A(n_1792),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1818),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1828),
.B(n_1825),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1850),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1824),
.B(n_1813),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1828),
.Y(n_1872)
);

NAND2xp5_ASAP7_75t_L g1873 ( 
.A(n_1824),
.B(n_1770),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1842),
.B(n_1792),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1842),
.B(n_1821),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1850),
.Y(n_1876)
);

INVx2_ASAP7_75t_SL g1877 ( 
.A(n_1835),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1863),
.B(n_1770),
.Y(n_1878)
);

NOR2xp33_ASAP7_75t_L g1879 ( 
.A(n_1831),
.B(n_1764),
.Y(n_1879)
);

INVx3_ASAP7_75t_L g1880 ( 
.A(n_1835),
.Y(n_1880)
);

OR2x2_ASAP7_75t_L g1881 ( 
.A(n_1852),
.B(n_1813),
.Y(n_1881)
);

HB1xp67_ASAP7_75t_L g1882 ( 
.A(n_1834),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1863),
.B(n_1770),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1822),
.Y(n_1884)
);

AOI221xp5_ASAP7_75t_L g1885 ( 
.A1(n_1848),
.A2(n_1764),
.B1(n_1758),
.B2(n_1762),
.C(n_1779),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1822),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1823),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1832),
.B(n_1771),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1852),
.B(n_1813),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1832),
.B(n_1834),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1867),
.B(n_1771),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_SL g1892 ( 
.A1(n_1867),
.A2(n_1798),
.B(n_1708),
.C(n_1811),
.Y(n_1892)
);

AND2x2_ASAP7_75t_L g1893 ( 
.A(n_1841),
.B(n_1821),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1835),
.B(n_1807),
.Y(n_1894)
);

NAND2xp5_ASAP7_75t_L g1895 ( 
.A(n_1851),
.B(n_1771),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1841),
.B(n_1821),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1829),
.B(n_1808),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1823),
.Y(n_1898)
);

INVx1_ASAP7_75t_SL g1899 ( 
.A(n_1835),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1829),
.B(n_1808),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1840),
.B(n_1805),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1840),
.B(n_1814),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1851),
.B(n_1760),
.Y(n_1903)
);

OAI32xp33_ASAP7_75t_L g1904 ( 
.A1(n_1847),
.A2(n_1802),
.A3(n_1798),
.B1(n_1779),
.B2(n_1814),
.Y(n_1904)
);

NAND2x1p5_ASAP7_75t_L g1905 ( 
.A(n_1835),
.B(n_1742),
.Y(n_1905)
);

OAI221xp5_ASAP7_75t_L g1906 ( 
.A1(n_1872),
.A2(n_1802),
.B1(n_1786),
.B2(n_1847),
.C(n_1864),
.Y(n_1906)
);

AOI321xp33_ASAP7_75t_L g1907 ( 
.A1(n_1885),
.A2(n_1865),
.A3(n_1853),
.B1(n_1811),
.B2(n_1752),
.C(n_1779),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1880),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1879),
.B(n_1854),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1890),
.B(n_1854),
.Y(n_1910)
);

OA22x2_ASAP7_75t_L g1911 ( 
.A1(n_1869),
.A2(n_1779),
.B1(n_1853),
.B2(n_1819),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1884),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1880),
.Y(n_1913)
);

AOI322xp5_ASAP7_75t_L g1914 ( 
.A1(n_1888),
.A2(n_1761),
.A3(n_1806),
.B1(n_1809),
.B2(n_1799),
.C1(n_1819),
.C2(n_1856),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1884),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1882),
.B(n_1835),
.Y(n_1916)
);

OAI322xp33_ASAP7_75t_L g1917 ( 
.A1(n_1878),
.A2(n_1847),
.A3(n_1845),
.B1(n_1861),
.B2(n_1788),
.C1(n_1790),
.C2(n_1797),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1874),
.B(n_1835),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1903),
.B(n_1845),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1874),
.B(n_1799),
.Y(n_1920)
);

AOI22xp5_ASAP7_75t_L g1921 ( 
.A1(n_1883),
.A2(n_1777),
.B1(n_1812),
.B2(n_1808),
.Y(n_1921)
);

OAI222xp33_ASAP7_75t_L g1922 ( 
.A1(n_1873),
.A2(n_1740),
.B1(n_1861),
.B2(n_1761),
.C1(n_1765),
.C2(n_1782),
.Y(n_1922)
);

OAI21xp33_ASAP7_75t_L g1923 ( 
.A1(n_1892),
.A2(n_1777),
.B(n_1760),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1886),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1871),
.B(n_1775),
.Y(n_1925)
);

OR2x2_ASAP7_75t_L g1926 ( 
.A(n_1871),
.B(n_1775),
.Y(n_1926)
);

A2O1A1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1892),
.A2(n_1782),
.B(n_1752),
.C(n_1761),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1880),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1886),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1887),
.Y(n_1930)
);

INVxp67_ASAP7_75t_L g1931 ( 
.A(n_1870),
.Y(n_1931)
);

NAND3xp33_ASAP7_75t_L g1932 ( 
.A(n_1870),
.B(n_1827),
.C(n_1826),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1907),
.B(n_1877),
.Y(n_1933)
);

AOI21xp33_ASAP7_75t_SL g1934 ( 
.A1(n_1923),
.A2(n_1904),
.B(n_1905),
.Y(n_1934)
);

CKINVDCx14_ASAP7_75t_R g1935 ( 
.A(n_1909),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1910),
.B(n_1875),
.Y(n_1936)
);

OAI21xp5_ASAP7_75t_L g1937 ( 
.A1(n_1927),
.A2(n_1904),
.B(n_1905),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1912),
.Y(n_1938)
);

AOI221xp5_ASAP7_75t_L g1939 ( 
.A1(n_1917),
.A2(n_1875),
.B1(n_1876),
.B2(n_1893),
.C(n_1896),
.Y(n_1939)
);

AOI21xp5_ASAP7_75t_L g1940 ( 
.A1(n_1927),
.A2(n_1899),
.B(n_1877),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1915),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1924),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1918),
.B(n_1893),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1931),
.B(n_1876),
.Y(n_1944)
);

OAI22xp33_ASAP7_75t_L g1945 ( 
.A1(n_1906),
.A2(n_1905),
.B1(n_1899),
.B2(n_1891),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1929),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1930),
.Y(n_1947)
);

AOI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1906),
.A2(n_1896),
.B1(n_1894),
.B2(n_1900),
.Y(n_1948)
);

INVx1_ASAP7_75t_L g1949 ( 
.A(n_1931),
.Y(n_1949)
);

AND2x2_ASAP7_75t_L g1950 ( 
.A(n_1920),
.B(n_1897),
.Y(n_1950)
);

OAI211xp5_ASAP7_75t_SL g1951 ( 
.A1(n_1921),
.A2(n_1902),
.B(n_1901),
.C(n_1898),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1919),
.B(n_1895),
.Y(n_1952)
);

AOI222xp33_ASAP7_75t_L g1953 ( 
.A1(n_1922),
.A2(n_1932),
.B1(n_1916),
.B2(n_1913),
.C1(n_1908),
.C2(n_1894),
.Y(n_1953)
);

INVx2_ASAP7_75t_L g1954 ( 
.A(n_1943),
.Y(n_1954)
);

BUFx6f_ASAP7_75t_L g1955 ( 
.A(n_1949),
.Y(n_1955)
);

O2A1O1Ixp33_ASAP7_75t_L g1956 ( 
.A1(n_1934),
.A2(n_1922),
.B(n_1928),
.C(n_1902),
.Y(n_1956)
);

NOR2xp33_ASAP7_75t_L g1957 ( 
.A(n_1935),
.B(n_1925),
.Y(n_1957)
);

AOI22xp33_ASAP7_75t_L g1958 ( 
.A1(n_1953),
.A2(n_1911),
.B1(n_1894),
.B2(n_1897),
.Y(n_1958)
);

OAI221xp5_ASAP7_75t_L g1959 ( 
.A1(n_1937),
.A2(n_1911),
.B1(n_1914),
.B2(n_1928),
.C(n_1901),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1944),
.Y(n_1960)
);

INVxp67_ASAP7_75t_L g1961 ( 
.A(n_1936),
.Y(n_1961)
);

OAI321xp33_ASAP7_75t_L g1962 ( 
.A1(n_1945),
.A2(n_1926),
.A3(n_1900),
.B1(n_1881),
.B2(n_1889),
.C(n_1898),
.Y(n_1962)
);

INVxp67_ASAP7_75t_SL g1963 ( 
.A(n_1945),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1948),
.B(n_1894),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_SL g1965 ( 
.A1(n_1939),
.A2(n_1889),
.B1(n_1881),
.B2(n_1887),
.C(n_1856),
.Y(n_1965)
);

NOR2x1_ASAP7_75t_L g1966 ( 
.A(n_1955),
.B(n_1933),
.Y(n_1966)
);

AND3x1_ASAP7_75t_L g1967 ( 
.A(n_1957),
.B(n_1940),
.C(n_1938),
.Y(n_1967)
);

NAND3xp33_ASAP7_75t_SL g1968 ( 
.A(n_1956),
.B(n_1933),
.C(n_1952),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1955),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1955),
.Y(n_1970)
);

AOI22xp5_ASAP7_75t_L g1971 ( 
.A1(n_1963),
.A2(n_1951),
.B1(n_1942),
.B2(n_1947),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1954),
.B(n_1950),
.Y(n_1972)
);

AO21x1_ASAP7_75t_L g1973 ( 
.A1(n_1964),
.A2(n_1946),
.B(n_1941),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1961),
.B(n_1960),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1958),
.B(n_1799),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1959),
.Y(n_1976)
);

AOI221x1_ASAP7_75t_L g1977 ( 
.A1(n_1976),
.A2(n_1951),
.B1(n_1962),
.B2(n_1959),
.C(n_1965),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1969),
.B(n_1806),
.Y(n_1978)
);

AO221x1_ASAP7_75t_L g1979 ( 
.A1(n_1970),
.A2(n_1784),
.B1(n_1826),
.B2(n_1866),
.C(n_1862),
.Y(n_1979)
);

AOI221xp5_ASAP7_75t_L g1980 ( 
.A1(n_1968),
.A2(n_1838),
.B1(n_1833),
.B2(n_1836),
.C(n_1860),
.Y(n_1980)
);

A2O1A1Ixp33_ASAP7_75t_L g1981 ( 
.A1(n_1966),
.A2(n_1868),
.B(n_1866),
.C(n_1862),
.Y(n_1981)
);

AOI221xp5_ASAP7_75t_L g1982 ( 
.A1(n_1967),
.A2(n_1838),
.B1(n_1860),
.B2(n_1859),
.C(n_1833),
.Y(n_1982)
);

AOI211xp5_ASAP7_75t_L g1983 ( 
.A1(n_1978),
.A2(n_1973),
.B(n_1971),
.C(n_1972),
.Y(n_1983)
);

OAI211xp5_ASAP7_75t_SL g1984 ( 
.A1(n_1981),
.A2(n_1971),
.B(n_1975),
.C(n_1974),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1979),
.Y(n_1985)
);

AOI211xp5_ASAP7_75t_L g1986 ( 
.A1(n_1977),
.A2(n_1980),
.B(n_1982),
.C(n_1563),
.Y(n_1986)
);

INVx1_ASAP7_75t_SL g1987 ( 
.A(n_1978),
.Y(n_1987)
);

AOI22xp5_ASAP7_75t_L g1988 ( 
.A1(n_1978),
.A2(n_1868),
.B1(n_1849),
.B2(n_1827),
.Y(n_1988)
);

OAI321xp33_ASAP7_75t_L g1989 ( 
.A1(n_1978),
.A2(n_1860),
.A3(n_1859),
.B1(n_1833),
.B2(n_1836),
.C(n_1838),
.Y(n_1989)
);

XNOR2xp5_ASAP7_75t_L g1990 ( 
.A(n_1983),
.B(n_1673),
.Y(n_1990)
);

OAI22xp5_ASAP7_75t_SL g1991 ( 
.A1(n_1987),
.A2(n_1673),
.B1(n_1740),
.B2(n_1837),
.Y(n_1991)
);

NOR2x1_ASAP7_75t_L g1992 ( 
.A(n_1984),
.B(n_1830),
.Y(n_1992)
);

INVx2_ASAP7_75t_L g1993 ( 
.A(n_1985),
.Y(n_1993)
);

OR2x2_ASAP7_75t_L g1994 ( 
.A(n_1988),
.B(n_1830),
.Y(n_1994)
);

NAND4xp75_ASAP7_75t_L g1995 ( 
.A(n_1986),
.B(n_1673),
.C(n_1858),
.D(n_1839),
.Y(n_1995)
);

AOI21xp5_ASAP7_75t_L g1996 ( 
.A1(n_1990),
.A2(n_1989),
.B(n_1843),
.Y(n_1996)
);

NAND4xp75_ASAP7_75t_L g1997 ( 
.A(n_1993),
.B(n_1849),
.C(n_1858),
.D(n_1837),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1991),
.B(n_1836),
.Y(n_1998)
);

AOI21xp5_ASAP7_75t_SL g1999 ( 
.A1(n_1998),
.A2(n_1994),
.B(n_1995),
.Y(n_1999)
);

OAI22xp5_ASAP7_75t_L g2000 ( 
.A1(n_1999),
.A2(n_1992),
.B1(n_1996),
.B2(n_1997),
.Y(n_2000)
);

AOI221xp5_ASAP7_75t_L g2001 ( 
.A1(n_2000),
.A2(n_1859),
.B1(n_1843),
.B2(n_1855),
.C(n_1846),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_2000),
.B(n_1843),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_2002),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_2001),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_2003),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_2004),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_2005),
.A2(n_1846),
.B(n_1844),
.Y(n_2007)
);

OAI21xp5_ASAP7_75t_SL g2008 ( 
.A1(n_2006),
.A2(n_1846),
.B(n_1844),
.Y(n_2008)
);

AO21x2_ASAP7_75t_L g2009 ( 
.A1(n_2007),
.A2(n_1855),
.B(n_1844),
.Y(n_2009)
);

HB1xp67_ASAP7_75t_L g2010 ( 
.A(n_2009),
.Y(n_2010)
);

OAI221xp5_ASAP7_75t_R g2011 ( 
.A1(n_2010),
.A2(n_2008),
.B1(n_1730),
.B2(n_1855),
.C(n_1857),
.Y(n_2011)
);

AOI211xp5_ASAP7_75t_L g2012 ( 
.A1(n_2011),
.A2(n_1857),
.B(n_1839),
.C(n_1610),
.Y(n_2012)
);


endmodule