module fake_jpeg_30037_n_60 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_60);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_60;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_37;
wire n_29;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_7),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_SL g10 ( 
.A(n_4),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_6),
.B(n_2),
.Y(n_12)
);

AOI22xp5_ASAP7_75t_L g13 ( 
.A1(n_0),
.A2(n_2),
.B1(n_6),
.B2(n_3),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_4),
.B(n_5),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_23),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_15),
.A2(n_0),
.B(n_1),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_21),
.B(n_13),
.Y(n_27)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_0),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_9),
.B(n_2),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_10),
.B(n_3),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_26),
.B(n_10),
.Y(n_28)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_28),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_20),
.B(n_10),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_35),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_8),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

OAI21xp33_ASAP7_75t_SL g37 ( 
.A1(n_19),
.A2(n_13),
.B(n_11),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_37),
.A2(n_11),
.B1(n_16),
.B2(n_17),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_27),
.A2(n_22),
.B1(n_11),
.B2(n_16),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_45),
.B1(n_16),
.B2(n_17),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_36),
.C(n_27),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.C(n_34),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.C(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_51),
.C(n_44),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.C(n_42),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_50),
.A2(n_42),
.B1(n_40),
.B2(n_46),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_38),
.Y(n_51)
);

AOI21xp5_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_54),
.B(n_51),
.Y(n_56)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_53),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_56),
.B(n_49),
.C(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_55),
.B(n_39),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_57),
.A2(n_58),
.B(n_17),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g60 ( 
.A1(n_59),
.A2(n_8),
.B(n_15),
.Y(n_60)
);


endmodule