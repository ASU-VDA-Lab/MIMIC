module fake_jpeg_7663_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx12_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_5),
.B(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_9),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_25),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_36),
.B(n_46),
.Y(n_58)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_37),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_29),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_41),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_0),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_48),
.B(n_50),
.Y(n_70)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_54),
.B(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_56),
.B(n_59),
.Y(n_89)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_61),
.B(n_74),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g62 ( 
.A1(n_47),
.A2(n_25),
.B1(n_32),
.B2(n_17),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_62),
.A2(n_63),
.B1(n_73),
.B2(n_76),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_32),
.B1(n_25),
.B2(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_26),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_71),
.Y(n_116)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_44),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_72),
.B(n_78),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_43),
.A2(n_32),
.B1(n_19),
.B2(n_33),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_48),
.B(n_35),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_35),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_19),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_17),
.B1(n_23),
.B2(n_34),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_39),
.B(n_34),
.Y(n_80)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_80),
.Y(n_87)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_81),
.Y(n_130)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_83),
.B(n_84),
.Y(n_119)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_88),
.B(n_98),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_19),
.B(n_33),
.C(n_30),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_90),
.A2(n_93),
.B1(n_95),
.B2(n_114),
.Y(n_132)
);

OAI21xp33_ASAP7_75t_L g91 ( 
.A1(n_54),
.A2(n_0),
.B(n_1),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_91),
.A2(n_22),
.B(n_18),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g93 ( 
.A1(n_64),
.A2(n_21),
.B1(n_18),
.B2(n_30),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_52),
.Y(n_94)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_94),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_53),
.A2(n_17),
.B1(n_23),
.B2(n_27),
.Y(n_95)
);

BUFx2_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_60),
.Y(n_98)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_99),
.B(n_100),
.Y(n_134)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_79),
.Y(n_101)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_101),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_102),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_69),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

OR2x2_ASAP7_75t_SL g145 ( 
.A(n_104),
.B(n_105),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_33),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_109),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_55),
.B(n_27),
.Y(n_107)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_56),
.B(n_30),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_58),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_110),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_22),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_66),
.Y(n_125)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_113),
.Y(n_138)
);

AO22x1_ASAP7_75t_SL g114 ( 
.A1(n_64),
.A2(n_21),
.B1(n_26),
.B2(n_42),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_117),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_22),
.C(n_18),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_118),
.B(n_14),
.Y(n_126)
);

AND2x4_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_21),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_122),
.A2(n_124),
.B(n_141),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_125),
.B(n_87),
.Y(n_163)
);

OAI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_126),
.A2(n_136),
.B(n_24),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_82),
.B(n_57),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_89),
.B(n_57),
.Y(n_128)
);

AOI32xp33_ASAP7_75t_L g136 ( 
.A1(n_114),
.A2(n_69),
.A3(n_51),
.B1(n_79),
.B2(n_26),
.Y(n_136)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_149),
.Y(n_158)
);

NOR2x1_ASAP7_75t_SL g141 ( 
.A(n_91),
.B(n_51),
.Y(n_141)
);

AND2x4_ASAP7_75t_SL g142 ( 
.A(n_105),
.B(n_85),
.Y(n_142)
);

MAJx2_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_28),
.C(n_24),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_92),
.B(n_26),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_86),
.Y(n_162)
);

OA22x2_ASAP7_75t_L g148 ( 
.A1(n_83),
.A2(n_71),
.B1(n_28),
.B2(n_24),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_148),
.A2(n_93),
.B1(n_116),
.B2(n_108),
.Y(n_175)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_90),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_128),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_151),
.B(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_141),
.A2(n_99),
.B1(n_122),
.B2(n_108),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_153),
.A2(n_183),
.B1(n_132),
.B2(n_148),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_125),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_157),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_149),
.A2(n_94),
.B(n_28),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_156),
.A2(n_159),
.B(n_173),
.Y(n_197)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_121),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_122),
.A2(n_142),
.B(n_147),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_160),
.B(n_167),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_161),
.A2(n_175),
.B1(n_142),
.B2(n_137),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_163),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_117),
.Y(n_164)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_117),
.Y(n_165)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_165),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_138),
.B(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_166),
.Y(n_208)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_131),
.B(n_88),
.Y(n_169)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_169),
.Y(n_210)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVx2_ASAP7_75t_SL g196 ( 
.A(n_170),
.Y(n_196)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_119),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_171),
.B(n_174),
.Y(n_216)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_120),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_172),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_133),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_148),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_176),
.A2(n_28),
.B(n_98),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_145),
.Y(n_177)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_177),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_1),
.Y(n_178)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_178),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_24),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_179),
.B(n_139),
.C(n_130),
.Y(n_198)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_135),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_145),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g186 ( 
.A(n_181),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_131),
.B(n_98),
.Y(n_182)
);

NAND2xp33_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_124),
.Y(n_193)
);

OAI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_122),
.A2(n_116),
.B1(n_115),
.B2(n_102),
.Y(n_183)
);

INVx6_ASAP7_75t_L g184 ( 
.A(n_144),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_184),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_189),
.B(n_193),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_123),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_198),
.C(n_199),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_168),
.A2(n_138),
.B(n_130),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_194),
.A2(n_213),
.B(n_181),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_159),
.B(n_132),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_158),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_156),
.A2(n_143),
.B1(n_135),
.B2(n_146),
.Y(n_201)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_201),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_177),
.B(n_173),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_175),
.A2(n_146),
.B1(n_126),
.B2(n_115),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_205),
.A2(n_217),
.B1(n_178),
.B2(n_170),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_155),
.C(n_150),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_207),
.B(n_209),
.C(n_215),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_126),
.C(n_86),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_24),
.B1(n_28),
.B2(n_97),
.Y(n_212)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_212),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_9),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_180),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_218),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_249)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_199),
.A2(n_151),
.B1(n_176),
.B2(n_162),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_221),
.A2(n_189),
.B1(n_213),
.B2(n_198),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_222),
.B(n_6),
.Y(n_266)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_223),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_211),
.B1(n_186),
.B2(n_202),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_190),
.B(n_171),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_234),
.C(n_240),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_227),
.B(n_230),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_195),
.B(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_229),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_231),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_2),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_184),
.C(n_157),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_191),
.B(n_172),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_187),
.Y(n_236)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_236),
.Y(n_262)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_196),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_237),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_191),
.B(n_160),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_242),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_197),
.A2(n_3),
.B(n_6),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_194),
.B(n_10),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_202),
.B(n_3),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_216),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_203),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_196),
.B1(n_3),
.B2(n_7),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_246),
.A2(n_253),
.B1(n_260),
.B2(n_238),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_255),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_224),
.A2(n_192),
.B1(n_204),
.B2(n_203),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_219),
.B(n_209),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_219),
.B(n_215),
.C(n_205),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_263),
.C(n_267),
.Y(n_269)
);

NOR2xp67_ASAP7_75t_SL g257 ( 
.A(n_221),
.B(n_208),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_240),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_218),
.A2(n_217),
.B1(n_210),
.B2(n_214),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_228),
.B1(n_245),
.B2(n_223),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_241),
.A2(n_220),
.B1(n_221),
.B2(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_185),
.C(n_196),
.Y(n_263)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_264),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_239),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_233),
.B(n_6),
.C(n_8),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_252),
.B(n_229),
.Y(n_270)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_270),
.Y(n_288)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_251),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_274),
.Y(n_295)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_235),
.Y(n_275)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_275),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_285),
.Y(n_291)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_246),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_277),
.A2(n_278),
.B(n_281),
.Y(n_290)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_279),
.A2(n_282),
.B1(n_284),
.B2(n_281),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_280),
.A2(n_286),
.B1(n_261),
.B2(n_242),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_259),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_258),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_256),
.Y(n_296)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_255),
.B(n_234),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_254),
.A2(n_248),
.B(n_232),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_268),
.B(n_243),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_237),
.Y(n_297)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_285),
.B(n_263),
.C(n_247),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_300),
.C(n_269),
.Y(n_306)
);

AO22x1_ASAP7_75t_L g293 ( 
.A1(n_280),
.A2(n_232),
.B1(n_260),
.B2(n_222),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_293),
.A2(n_302),
.B(n_297),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_296),
.B(n_271),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_297),
.B(n_8),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_298),
.Y(n_308)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_9),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_247),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_272),
.A2(n_250),
.B1(n_266),
.B2(n_265),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_301),
.A2(n_302),
.B1(n_290),
.B2(n_293),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_286),
.A2(n_262),
.B1(n_236),
.B2(n_233),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_303),
.B(n_304),
.C(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_300),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_267),
.Y(n_305)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_283),
.B1(n_276),
.B2(n_269),
.Y(n_309)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_309),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_310),
.B(n_311),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_288),
.B(n_8),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_312),
.B(n_315),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_313),
.B(n_314),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_294),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_291),
.Y(n_322)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_292),
.C(n_291),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_323),
.B(n_15),
.C(n_318),
.Y(n_330)
);

NOR2x1_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_15),
.Y(n_324)
);

NOR2xp67_ASAP7_75t_SL g327 ( 
.A(n_324),
.B(n_10),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_318),
.B(n_304),
.C(n_303),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_326),
.B(n_330),
.C(n_323),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_327),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_308),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_321),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_319),
.A2(n_309),
.B(n_14),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_329),
.B(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_332),
.B(n_334),
.Y(n_335)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_335),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_316),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_336),
.B(n_333),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_317),
.B(n_325),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_15),
.Y(n_341)
);


endmodule