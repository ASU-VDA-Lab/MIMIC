module fake_ariane_1150_n_1541 (n_295, n_356, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_332, n_294, n_197, n_176, n_34, n_172, n_347, n_183, n_299, n_12, n_133, n_66, n_205, n_341, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_345, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_349, n_346, n_214, n_348, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_327, n_77, n_15, n_23, n_87, n_279, n_207, n_354, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_338, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_336, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_339, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_331, n_267, n_335, n_350, n_291, n_344, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_326, n_227, n_48, n_188, n_323, n_330, n_11, n_129, n_126, n_282, n_328, n_277, n_248, n_301, n_293, n_228, n_325, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_352, n_238, n_136, n_334, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_333, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_343, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_355, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_324, n_337, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_342, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_353, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_351, n_39, n_155, n_127, n_1541);

input n_295;
input n_356;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_332;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_347;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_345;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_349;
input n_346;
input n_214;
input n_348;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_327;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_354;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_338;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_336;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_339;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_331;
input n_267;
input n_335;
input n_350;
input n_291;
input n_344;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_326;
input n_227;
input n_48;
input n_188;
input n_323;
input n_330;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_325;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_238;
input n_136;
input n_334;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_333;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_343;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_324;
input n_337;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_342;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_353;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_351;
input n_39;
input n_155;
input n_127;

output n_1541;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_559;
wire n_495;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_1495;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_436;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_604;
wire n_439;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_1035;
wire n_1143;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_914;
wire n_689;
wire n_400;
wire n_1116;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_718;
wire n_1434;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_71),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_199),
.Y(n_358)
);

BUFx2_ASAP7_75t_L g359 ( 
.A(n_266),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_243),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_218),
.Y(n_361)
);

INVx1_ASAP7_75t_SL g362 ( 
.A(n_281),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_326),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_107),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_193),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_178),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_146),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_347),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_310),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_231),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_320),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_53),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_329),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_260),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_187),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_235),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_90),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_162),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_160),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_48),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_295),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_276),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_81),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_51),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_195),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_134),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_215),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_204),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_52),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_142),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_318),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_344),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_263),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_76),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_130),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_214),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_212),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_153),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_105),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_203),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_17),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_124),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_346),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_336),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_70),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_13),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_249),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_280),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_229),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_300),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_340),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_39),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_48),
.Y(n_414)
);

BUFx3_ASAP7_75t_L g415 ( 
.A(n_256),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_298),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_251),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_190),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_8),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_108),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_8),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_13),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_135),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g424 ( 
.A(n_328),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_339),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_296),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_301),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_337),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_99),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g430 ( 
.A(n_221),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_308),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_29),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_19),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_4),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_27),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_335),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_61),
.Y(n_437)
);

BUFx10_ASAP7_75t_L g438 ( 
.A(n_314),
.Y(n_438)
);

INVx2_ASAP7_75t_L g439 ( 
.A(n_89),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_41),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_10),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_253),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_282),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_68),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_197),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_36),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_23),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_332),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_145),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_45),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_262),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_72),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_74),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_288),
.Y(n_454)
);

BUFx10_ASAP7_75t_L g455 ( 
.A(n_59),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_118),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_311),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_7),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_224),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_246),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_324),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_25),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_159),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_16),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_45),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_91),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_104),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_312),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_258),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_127),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g471 ( 
.A(n_10),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_11),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_88),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_66),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_194),
.Y(n_475)
);

BUFx10_ASAP7_75t_L g476 ( 
.A(n_27),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_32),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_333),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_175),
.Y(n_479)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_87),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_49),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_163),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_43),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_352),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_309),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_131),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_278),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_226),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_35),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_100),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_2),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_22),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_18),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_355),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_28),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_176),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_242),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_22),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_141),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_101),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_171),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_112),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_327),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_341),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_351),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_275),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_16),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_150),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_168),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_14),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_232),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_56),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_181),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_230),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_225),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_237),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_38),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_183),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_267),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_121),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_299),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_338),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_319),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_247),
.Y(n_524)
);

BUFx2_ASAP7_75t_L g525 ( 
.A(n_140),
.Y(n_525)
);

CKINVDCx14_ASAP7_75t_R g526 ( 
.A(n_303),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_169),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_184),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_177),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_35),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_3),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_349),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_9),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_44),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_58),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_7),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_5),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_0),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_265),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_321),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_55),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_334),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g543 ( 
.A(n_192),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_79),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_302),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_73),
.Y(n_546)
);

CKINVDCx16_ASAP7_75t_R g547 ( 
.A(n_206),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_129),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_19),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_24),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_493),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_493),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_373),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_371),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_373),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_485),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_380),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_377),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_540),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_386),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_540),
.Y(n_562)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_413),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_419),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_406),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_419),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_419),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_419),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_419),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g570 ( 
.A(n_430),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_442),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_480),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_497),
.Y(n_573)
);

CKINVDCx20_ASAP7_75t_R g574 ( 
.A(n_502),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_419),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_532),
.Y(n_576)
);

INVxp67_ASAP7_75t_SL g577 ( 
.A(n_507),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_414),
.Y(n_578)
);

CKINVDCx16_ASAP7_75t_R g579 ( 
.A(n_390),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_440),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_359),
.B(n_0),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_458),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_384),
.Y(n_583)
);

INVxp33_ASAP7_75t_SL g584 ( 
.A(n_402),
.Y(n_584)
);

BUFx3_ASAP7_75t_L g585 ( 
.A(n_415),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_477),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_389),
.Y(n_587)
);

INVx1_ASAP7_75t_SL g588 ( 
.A(n_495),
.Y(n_588)
);

CKINVDCx20_ASAP7_75t_R g589 ( 
.A(n_538),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_421),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_507),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_489),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_422),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_432),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_434),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_435),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_491),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_498),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_530),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_476),
.Y(n_600)
);

BUFx8_ASAP7_75t_SL g601 ( 
.A(n_399),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_476),
.Y(n_602)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_441),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_533),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_446),
.Y(n_605)
);

CKINVDCx20_ASAP7_75t_R g606 ( 
.A(n_447),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_450),
.Y(n_607)
);

INVxp67_ASAP7_75t_SL g608 ( 
.A(n_507),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_507),
.Y(n_609)
);

INVxp33_ASAP7_75t_SL g610 ( 
.A(n_462),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_526),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_526),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_534),
.Y(n_613)
);

CKINVDCx20_ASAP7_75t_R g614 ( 
.A(n_547),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_464),
.Y(n_615)
);

INVxp67_ASAP7_75t_SL g616 ( 
.A(n_550),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_438),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g618 ( 
.A(n_407),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_465),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_472),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_481),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_516),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_525),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_438),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_483),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_455),
.Y(n_626)
);

INVxp67_ASAP7_75t_SL g627 ( 
.A(n_415),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_455),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_514),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_514),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_370),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_374),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_R g633 ( 
.A(n_357),
.B(n_54),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_535),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_378),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_492),
.Y(n_636)
);

CKINVDCx20_ASAP7_75t_R g637 ( 
.A(n_510),
.Y(n_637)
);

CKINVDCx5p33_ASAP7_75t_R g638 ( 
.A(n_517),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_531),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_392),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_395),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_433),
.B(n_1),
.Y(n_642)
);

CKINVDCx5p33_ASAP7_75t_R g643 ( 
.A(n_536),
.Y(n_643)
);

INVxp67_ASAP7_75t_SL g644 ( 
.A(n_396),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_537),
.Y(n_645)
);

INVxp67_ASAP7_75t_SL g646 ( 
.A(n_404),
.Y(n_646)
);

NOR2xp67_ASAP7_75t_L g647 ( 
.A(n_549),
.B(n_1),
.Y(n_647)
);

CKINVDCx20_ASAP7_75t_R g648 ( 
.A(n_471),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_360),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_411),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_412),
.B(n_2),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_361),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_363),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_416),
.B(n_3),
.Y(n_654)
);

CKINVDCx16_ASAP7_75t_R g655 ( 
.A(n_358),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_417),
.Y(n_656)
);

NOR2xp33_ASAP7_75t_R g657 ( 
.A(n_364),
.B(n_57),
.Y(n_657)
);

CKINVDCx20_ASAP7_75t_R g658 ( 
.A(n_365),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_418),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_420),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_426),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_427),
.Y(n_662)
);

INVxp67_ASAP7_75t_SL g663 ( 
.A(n_431),
.Y(n_663)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_366),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_655),
.B(n_383),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_577),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_585),
.B(n_358),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_648),
.A2(n_456),
.B1(n_461),
.B2(n_444),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_608),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_585),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_564),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_554),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_566),
.B(n_463),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_624),
.B(n_379),
.Y(n_674)
);

HB1xp67_ASAP7_75t_L g675 ( 
.A(n_583),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_567),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_568),
.B(n_469),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_591),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_575),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_569),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_569),
.Y(n_681)
);

BUFx6f_ASAP7_75t_L g682 ( 
.A(n_591),
.Y(n_682)
);

INVxp67_ASAP7_75t_L g683 ( 
.A(n_557),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_578),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_581),
.B(n_437),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_580),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_582),
.Y(n_687)
);

BUFx2_ASAP7_75t_L g688 ( 
.A(n_637),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_626),
.B(n_473),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_590),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_627),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_609),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_586),
.Y(n_693)
);

BUFx6f_ASAP7_75t_L g694 ( 
.A(n_609),
.Y(n_694)
);

INVx3_ASAP7_75t_L g695 ( 
.A(n_551),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_628),
.B(n_475),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_592),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_597),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_552),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_598),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_629),
.B(n_478),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_588),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_649),
.B(n_652),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_599),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_604),
.Y(n_705)
);

OA21x2_ASAP7_75t_L g706 ( 
.A1(n_654),
.A2(n_503),
.B(n_484),
.Y(n_706)
);

OAI21x1_ASAP7_75t_L g707 ( 
.A1(n_631),
.A2(n_509),
.B(n_504),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_613),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_632),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_616),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_640),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_639),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_650),
.B(n_513),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_656),
.B(n_515),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_659),
.Y(n_717)
);

INVx1_ASAP7_75t_SL g718 ( 
.A(n_648),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_660),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_630),
.B(n_518),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_593),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_622),
.B(n_519),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_661),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_644),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_646),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_579),
.B(n_548),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_553),
.Y(n_727)
);

INVx3_ASAP7_75t_L g728 ( 
.A(n_555),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_663),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_623),
.B(n_556),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_651),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_618),
.Y(n_732)
);

OA21x2_ASAP7_75t_L g733 ( 
.A1(n_662),
.A2(n_528),
.B(n_527),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_563),
.Y(n_734)
);

BUFx6f_ASAP7_75t_L g735 ( 
.A(n_642),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_634),
.B(n_529),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_L g737 ( 
.A(n_653),
.B(n_539),
.Y(n_737)
);

INVx1_ASAP7_75t_SL g738 ( 
.A(n_603),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_559),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_560),
.B(n_362),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_562),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_594),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_595),
.B(n_424),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_596),
.B(n_439),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_605),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_607),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_615),
.Y(n_747)
);

OA21x2_ASAP7_75t_L g748 ( 
.A1(n_647),
.A2(n_544),
.B(n_541),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_619),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_633),
.B(n_358),
.Y(n_750)
);

BUFx6f_ASAP7_75t_L g751 ( 
.A(n_621),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_625),
.B(n_545),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_636),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_638),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_643),
.Y(n_755)
);

BUFx6f_ASAP7_75t_L g756 ( 
.A(n_645),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_584),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_678),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_678),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_699),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_678),
.Y(n_761)
);

BUFx4f_ASAP7_75t_L g762 ( 
.A(n_751),
.Y(n_762)
);

INVx4_ASAP7_75t_L g763 ( 
.A(n_670),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_691),
.B(n_610),
.Y(n_764)
);

AND2x6_ASAP7_75t_L g765 ( 
.A(n_751),
.B(n_358),
.Y(n_765)
);

INVx4_ASAP7_75t_L g766 ( 
.A(n_670),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_705),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

AND2x2_ASAP7_75t_SL g769 ( 
.A(n_751),
.B(n_601),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_682),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_682),
.Y(n_771)
);

AND2x4_ASAP7_75t_L g772 ( 
.A(n_735),
.B(n_658),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_717),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_702),
.B(n_558),
.Y(n_774)
);

BUFx6f_ASAP7_75t_L g775 ( 
.A(n_682),
.Y(n_775)
);

BUFx4f_ASAP7_75t_L g776 ( 
.A(n_756),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_684),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_686),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_694),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_687),
.Y(n_781)
);

INVxp67_ASAP7_75t_L g782 ( 
.A(n_702),
.Y(n_782)
);

AND2x4_ASAP7_75t_L g783 ( 
.A(n_735),
.B(n_658),
.Y(n_783)
);

BUFx6f_ASAP7_75t_L g784 ( 
.A(n_694),
.Y(n_784)
);

AOI22xp33_ASAP7_75t_L g785 ( 
.A1(n_750),
.A2(n_612),
.B1(n_611),
.B2(n_606),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_743),
.B(n_664),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_694),
.Y(n_787)
);

AND2x4_ASAP7_75t_L g788 ( 
.A(n_735),
.B(n_727),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_738),
.Y(n_789)
);

BUFx6f_ASAP7_75t_L g790 ( 
.A(n_700),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_680),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_L g792 ( 
.A(n_736),
.B(n_606),
.C(n_603),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_731),
.B(n_543),
.Y(n_793)
);

INVxp67_ASAP7_75t_SL g794 ( 
.A(n_680),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_672),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_672),
.Y(n_796)
);

INVx4_ASAP7_75t_L g797 ( 
.A(n_756),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_693),
.Y(n_798)
);

AND2x2_ASAP7_75t_SL g799 ( 
.A(n_756),
.B(n_601),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_731),
.B(n_657),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_681),
.Y(n_801)
);

NAND2xp33_ASAP7_75t_L g802 ( 
.A(n_750),
.B(n_746),
.Y(n_802)
);

AND2x4_ASAP7_75t_L g803 ( 
.A(n_727),
.B(n_614),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_692),
.Y(n_804)
);

NAND3xp33_ASAP7_75t_L g805 ( 
.A(n_736),
.B(n_620),
.C(n_368),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_737),
.B(n_671),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_683),
.B(n_617),
.Y(n_807)
);

INVx4_ASAP7_75t_SL g808 ( 
.A(n_667),
.Y(n_808)
);

INVx4_ASAP7_75t_L g809 ( 
.A(n_739),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_737),
.B(n_676),
.Y(n_810)
);

INVx4_ASAP7_75t_L g811 ( 
.A(n_739),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_697),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_683),
.B(n_561),
.Y(n_813)
);

AND2x2_ASAP7_75t_SL g814 ( 
.A(n_726),
.B(n_445),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_752),
.B(n_746),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_688),
.Y(n_816)
);

INVxp67_ASAP7_75t_L g817 ( 
.A(n_713),
.Y(n_817)
);

INVx4_ASAP7_75t_L g818 ( 
.A(n_739),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_698),
.Y(n_819)
);

AND2x6_ASAP7_75t_L g820 ( 
.A(n_747),
.B(n_742),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_679),
.B(n_657),
.Y(n_821)
);

AO22x2_ASAP7_75t_L g822 ( 
.A1(n_718),
.A2(n_738),
.B1(n_722),
.B2(n_740),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_724),
.B(n_367),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_700),
.Y(n_824)
);

AND2x6_ASAP7_75t_L g825 ( 
.A(n_747),
.B(n_449),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_734),
.B(n_565),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_700),
.Y(n_827)
);

BUFx6f_ASAP7_75t_L g828 ( 
.A(n_707),
.Y(n_828)
);

NOR2xp33_ASAP7_75t_L g829 ( 
.A(n_755),
.B(n_571),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_724),
.B(n_369),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_675),
.B(n_572),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_752),
.B(n_745),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_750),
.B(n_372),
.Y(n_833)
);

BUFx3_ASAP7_75t_L g834 ( 
.A(n_666),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_704),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_675),
.Y(n_836)
);

BUFx6f_ASAP7_75t_L g837 ( 
.A(n_723),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_695),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_708),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_723),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_695),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_709),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_750),
.B(n_375),
.Y(n_843)
);

AND3x2_ASAP7_75t_L g844 ( 
.A(n_690),
.B(n_470),
.C(n_466),
.Y(n_844)
);

BUFx8_ASAP7_75t_SL g845 ( 
.A(n_757),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_690),
.Y(n_846)
);

AND2x4_ASAP7_75t_L g847 ( 
.A(n_797),
.B(n_710),
.Y(n_847)
);

OAI221xp5_ASAP7_75t_L g848 ( 
.A1(n_764),
.A2(n_685),
.B1(n_744),
.B2(n_729),
.C(n_725),
.Y(n_848)
);

HB1xp67_ASAP7_75t_L g849 ( 
.A(n_782),
.Y(n_849)
);

BUFx6f_ASAP7_75t_SL g850 ( 
.A(n_769),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_778),
.Y(n_851)
);

OAI221xp5_ASAP7_75t_L g852 ( 
.A1(n_806),
.A2(n_685),
.B1(n_744),
.B2(n_716),
.C(n_715),
.Y(n_852)
);

AO22x2_ASAP7_75t_L g853 ( 
.A1(n_792),
.A2(n_718),
.B1(n_668),
.B2(n_665),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_779),
.Y(n_854)
);

NOR3xp33_ASAP7_75t_L g855 ( 
.A(n_836),
.B(n_703),
.C(n_721),
.Y(n_855)
);

BUFx8_ASAP7_75t_L g856 ( 
.A(n_831),
.Y(n_856)
);

NAND2x1p5_ASAP7_75t_L g857 ( 
.A(n_762),
.B(n_776),
.Y(n_857)
);

NAND2x1p5_ASAP7_75t_L g858 ( 
.A(n_797),
.B(n_703),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_809),
.B(n_749),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_837),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_781),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_798),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_813),
.B(n_774),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_812),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_837),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_819),
.Y(n_866)
);

BUFx8_ASAP7_75t_L g867 ( 
.A(n_807),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_810),
.B(n_750),
.Y(n_868)
);

BUFx3_ASAP7_75t_L g869 ( 
.A(n_795),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_837),
.Y(n_870)
);

CKINVDCx5p33_ASAP7_75t_R g871 ( 
.A(n_796),
.Y(n_871)
);

AO22x2_ASAP7_75t_L g872 ( 
.A1(n_805),
.A2(n_665),
.B1(n_722),
.B2(n_674),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_800),
.B(n_793),
.Y(n_873)
);

AO22x2_ASAP7_75t_L g874 ( 
.A1(n_772),
.A2(n_674),
.B1(n_741),
.B2(n_696),
.Y(n_874)
);

AND2x4_ASAP7_75t_L g875 ( 
.A(n_789),
.B(n_570),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_835),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_839),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_760),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_763),
.B(n_766),
.Y(n_879)
);

AO22x2_ASAP7_75t_L g880 ( 
.A1(n_772),
.A2(n_696),
.B1(n_701),
.B2(n_689),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_767),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_845),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_788),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_846),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_788),
.Y(n_885)
);

AO22x2_ASAP7_75t_L g886 ( 
.A1(n_783),
.A2(n_701),
.B1(n_720),
.B2(n_689),
.Y(n_886)
);

AO22x2_ASAP7_75t_L g887 ( 
.A1(n_783),
.A2(n_786),
.B1(n_803),
.B2(n_822),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_814),
.A2(n_733),
.B1(n_748),
.B2(n_706),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_816),
.Y(n_889)
);

NAND2x1p5_ASAP7_75t_L g890 ( 
.A(n_809),
.B(n_811),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_801),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_826),
.B(n_721),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_803),
.A2(n_720),
.B1(n_576),
.B2(n_574),
.Y(n_893)
);

NOR2xp33_ASAP7_75t_L g894 ( 
.A(n_815),
.B(n_753),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_834),
.Y(n_895)
);

AND2x2_ASAP7_75t_SL g896 ( 
.A(n_799),
.B(n_754),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_842),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_842),
.Y(n_898)
);

AO22x2_ASAP7_75t_L g899 ( 
.A1(n_822),
.A2(n_832),
.B1(n_817),
.B2(n_785),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_829),
.B(n_573),
.Y(n_900)
);

NAND2x1p5_ASAP7_75t_L g901 ( 
.A(n_811),
.B(n_728),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_763),
.B(n_669),
.Y(n_902)
);

NAND2x1p5_ASAP7_75t_L g903 ( 
.A(n_818),
.B(n_728),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_818),
.B(n_620),
.Y(n_904)
);

AO22x2_ASAP7_75t_L g905 ( 
.A1(n_768),
.A2(n_587),
.B1(n_589),
.B2(n_730),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_804),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_790),
.B(n_712),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_790),
.B(n_714),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_766),
.B(n_733),
.Y(n_909)
);

NAND2x1p5_ASAP7_75t_L g910 ( 
.A(n_790),
.B(n_719),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_820),
.B(n_711),
.Y(n_911)
);

HAxp5_ASAP7_75t_SL g912 ( 
.A(n_773),
.B(n_600),
.CON(n_912),
.SN(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_841),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_840),
.Y(n_914)
);

AO22x2_ASAP7_75t_L g915 ( 
.A1(n_777),
.A2(n_600),
.B1(n_602),
.B2(n_732),
.Y(n_915)
);

AO22x2_ASAP7_75t_L g916 ( 
.A1(n_827),
.A2(n_602),
.B1(n_716),
.B2(n_715),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_840),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_840),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_791),
.Y(n_919)
);

INVx3_ASAP7_75t_L g920 ( 
.A(n_824),
.Y(n_920)
);

BUFx3_ASAP7_75t_L g921 ( 
.A(n_765),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_823),
.A2(n_673),
.B1(n_677),
.B2(n_706),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_838),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_765),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_794),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_824),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_824),
.Y(n_927)
);

BUFx8_ASAP7_75t_L g928 ( 
.A(n_765),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_761),
.Y(n_929)
);

AO22x2_ASAP7_75t_L g930 ( 
.A1(n_830),
.A2(n_844),
.B1(n_833),
.B2(n_843),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_820),
.B(n_673),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_820),
.B(n_677),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_761),
.Y(n_933)
);

AO22x2_ASAP7_75t_L g934 ( 
.A1(n_808),
.A2(n_821),
.B1(n_759),
.B2(n_771),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_761),
.Y(n_935)
);

AND2x4_ASAP7_75t_L g936 ( 
.A(n_808),
.B(n_667),
.Y(n_936)
);

INVxp67_ASAP7_75t_L g937 ( 
.A(n_758),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_802),
.B(n_748),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_780),
.Y(n_939)
);

NOR2xp67_ASAP7_75t_L g940 ( 
.A(n_787),
.B(n_376),
.Y(n_940)
);

AO22x2_ASAP7_75t_L g941 ( 
.A1(n_825),
.A2(n_542),
.B1(n_6),
.B2(n_4),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_770),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_770),
.Y(n_943)
);

AO22x2_ASAP7_75t_L g944 ( 
.A1(n_825),
.A2(n_9),
.B1(n_5),
.B2(n_6),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_770),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_892),
.B(n_775),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_863),
.B(n_828),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_847),
.B(n_775),
.Y(n_948)
);

NAND2xp33_ASAP7_75t_SL g949 ( 
.A(n_871),
.B(n_828),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_900),
.B(n_775),
.Y(n_950)
);

NAND2xp33_ASAP7_75t_SL g951 ( 
.A(n_884),
.B(n_889),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_SL g952 ( 
.A(n_894),
.B(n_784),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_855),
.B(n_784),
.Y(n_953)
);

NAND2xp33_ASAP7_75t_SL g954 ( 
.A(n_851),
.B(n_854),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_847),
.B(n_784),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_873),
.B(n_825),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_SL g957 ( 
.A(n_904),
.B(n_381),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_858),
.B(n_382),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_869),
.B(n_385),
.Y(n_959)
);

NAND2xp33_ASAP7_75t_SL g960 ( 
.A(n_861),
.B(n_387),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_883),
.B(n_885),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_931),
.B(n_388),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_SL g963 ( 
.A(n_931),
.B(n_932),
.Y(n_963)
);

NAND2xp33_ASAP7_75t_SL g964 ( 
.A(n_862),
.B(n_864),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_866),
.B(n_667),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_SL g966 ( 
.A(n_932),
.B(n_391),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_895),
.B(n_667),
.Y(n_967)
);

NAND2xp33_ASAP7_75t_SL g968 ( 
.A(n_876),
.B(n_393),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_857),
.B(n_394),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_896),
.B(n_849),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_868),
.B(n_397),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_SL g972 ( 
.A(n_859),
.B(n_398),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_SL g973 ( 
.A(n_901),
.B(n_400),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_903),
.B(n_401),
.Y(n_974)
);

NAND2xp33_ASAP7_75t_SL g975 ( 
.A(n_877),
.B(n_403),
.Y(n_975)
);

NAND2xp33_ASAP7_75t_SL g976 ( 
.A(n_879),
.B(n_405),
.Y(n_976)
);

NAND2xp33_ASAP7_75t_SL g977 ( 
.A(n_923),
.B(n_408),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_SL g978 ( 
.A(n_902),
.B(n_409),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_911),
.B(n_410),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_SL g980 ( 
.A(n_856),
.B(n_423),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_890),
.B(n_425),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_852),
.B(n_667),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_936),
.B(n_11),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_SL g984 ( 
.A(n_913),
.B(n_428),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_920),
.B(n_429),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_848),
.B(n_436),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_878),
.B(n_443),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_SL g988 ( 
.A(n_935),
.B(n_448),
.Y(n_988)
);

NAND2xp33_ASAP7_75t_SL g989 ( 
.A(n_850),
.B(n_546),
.Y(n_989)
);

NAND2xp33_ASAP7_75t_SL g990 ( 
.A(n_882),
.B(n_451),
.Y(n_990)
);

NAND2xp33_ASAP7_75t_SL g991 ( 
.A(n_897),
.B(n_524),
.Y(n_991)
);

NAND2xp33_ASAP7_75t_SL g992 ( 
.A(n_898),
.B(n_452),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_909),
.B(n_453),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_SL g994 ( 
.A(n_867),
.B(n_454),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_875),
.B(n_12),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_881),
.B(n_457),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_SL g997 ( 
.A(n_940),
.B(n_459),
.Y(n_997)
);

NAND2xp33_ASAP7_75t_SL g998 ( 
.A(n_926),
.B(n_523),
.Y(n_998)
);

NAND2xp33_ASAP7_75t_SL g999 ( 
.A(n_927),
.B(n_460),
.Y(n_999)
);

NAND2xp33_ASAP7_75t_SL g1000 ( 
.A(n_942),
.B(n_467),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_SL g1001 ( 
.A(n_914),
.B(n_468),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_860),
.B(n_474),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_925),
.B(n_479),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_865),
.B(n_482),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_870),
.B(n_917),
.Y(n_1005)
);

NAND2xp33_ASAP7_75t_SL g1006 ( 
.A(n_943),
.B(n_486),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_918),
.B(n_945),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_SL g1008 ( 
.A(n_936),
.B(n_487),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_872),
.B(n_488),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_907),
.B(n_490),
.Y(n_1010)
);

NAND2xp33_ASAP7_75t_SL g1011 ( 
.A(n_929),
.B(n_494),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_SL g1012 ( 
.A(n_908),
.B(n_496),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_SL g1013 ( 
.A(n_910),
.B(n_499),
.Y(n_1013)
);

OR2x2_ASAP7_75t_L g1014 ( 
.A(n_891),
.B(n_12),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_933),
.B(n_500),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_SL g1016 ( 
.A(n_921),
.B(n_924),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_937),
.B(n_501),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_SL g1018 ( 
.A(n_939),
.B(n_505),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_888),
.B(n_506),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_906),
.B(n_508),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_928),
.B(n_511),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_872),
.B(n_853),
.Y(n_1022)
);

NAND2xp33_ASAP7_75t_SL g1023 ( 
.A(n_938),
.B(n_919),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_SL g1024 ( 
.A(n_880),
.B(n_512),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_880),
.B(n_520),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_886),
.B(n_521),
.Y(n_1026)
);

OR2x2_ASAP7_75t_L g1027 ( 
.A(n_970),
.B(n_912),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_946),
.B(n_886),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_948),
.B(n_853),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_961),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_948),
.B(n_887),
.Y(n_1031)
);

INVx1_ASAP7_75t_SL g1032 ( 
.A(n_951),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_1019),
.A2(n_934),
.B(n_922),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_963),
.Y(n_1034)
);

NAND2xp5_ASAP7_75t_L g1035 ( 
.A(n_961),
.B(n_899),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_995),
.B(n_874),
.Y(n_1036)
);

OAI21x1_ASAP7_75t_L g1037 ( 
.A1(n_947),
.A2(n_930),
.B(n_941),
.Y(n_1037)
);

AOI21xp33_ASAP7_75t_L g1038 ( 
.A1(n_986),
.A2(n_899),
.B(n_874),
.Y(n_1038)
);

OAI21x1_ASAP7_75t_L g1039 ( 
.A1(n_982),
.A2(n_1005),
.B(n_956),
.Y(n_1039)
);

OA21x2_ASAP7_75t_L g1040 ( 
.A1(n_1022),
.A2(n_993),
.B(n_971),
.Y(n_1040)
);

AO21x1_ASAP7_75t_L g1041 ( 
.A1(n_1023),
.A2(n_941),
.B(n_944),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_983),
.Y(n_1042)
);

CKINVDCx8_ASAP7_75t_R g1043 ( 
.A(n_983),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_L g1044 ( 
.A1(n_952),
.A2(n_930),
.B(n_944),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_954),
.A2(n_522),
.B(n_449),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_990),
.Y(n_1046)
);

NAND3xp33_ASAP7_75t_SL g1047 ( 
.A(n_957),
.B(n_915),
.C(n_893),
.Y(n_1047)
);

AOI21xp5_ASAP7_75t_L g1048 ( 
.A1(n_964),
.A2(n_522),
.B(n_449),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_967),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_1014),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_965),
.A2(n_62),
.B(n_60),
.Y(n_1051)
);

BUFx12f_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

BUFx6f_ASAP7_75t_L g1053 ( 
.A(n_1016),
.Y(n_1053)
);

OA22x2_ASAP7_75t_L g1054 ( 
.A1(n_1024),
.A2(n_915),
.B1(n_893),
.B2(n_905),
.Y(n_1054)
);

OAI22x1_ASAP7_75t_L g1055 ( 
.A1(n_1025),
.A2(n_905),
.B1(n_916),
.B2(n_887),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_955),
.Y(n_1056)
);

OAI21x1_ASAP7_75t_L g1057 ( 
.A1(n_1007),
.A2(n_64),
.B(n_63),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_1020),
.B(n_916),
.Y(n_1058)
);

AO31x2_ASAP7_75t_L g1059 ( 
.A1(n_1009),
.A2(n_522),
.A3(n_449),
.B(n_67),
.Y(n_1059)
);

OAI22xp5_ASAP7_75t_L g1060 ( 
.A1(n_987),
.A2(n_522),
.B1(n_17),
.B2(n_14),
.Y(n_1060)
);

AO21x2_ASAP7_75t_L g1061 ( 
.A1(n_979),
.A2(n_69),
.B(n_65),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_996),
.B(n_15),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_1003),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_953),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_950),
.B(n_15),
.Y(n_1065)
);

BUFx6f_ASAP7_75t_L g1066 ( 
.A(n_962),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_1026),
.B(n_18),
.Y(n_1067)
);

AOI21x1_ASAP7_75t_L g1068 ( 
.A1(n_978),
.A2(n_77),
.B(n_75),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_1010),
.A2(n_1013),
.B(n_1012),
.Y(n_1069)
);

NAND2x1p5_ASAP7_75t_L g1070 ( 
.A(n_994),
.B(n_78),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_989),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_958),
.A2(n_82),
.B(n_80),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_960),
.B(n_20),
.Y(n_1073)
);

AO31x2_ASAP7_75t_L g1074 ( 
.A1(n_966),
.A2(n_186),
.A3(n_354),
.B(n_353),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_968),
.B(n_20),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1002),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1004),
.Y(n_1077)
);

OR2x2_ASAP7_75t_L g1078 ( 
.A(n_975),
.B(n_21),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_984),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_1079)
);

AO21x2_ASAP7_75t_L g1080 ( 
.A1(n_997),
.A2(n_84),
.B(n_83),
.Y(n_1080)
);

OAI22xp5_ASAP7_75t_L g1081 ( 
.A1(n_973),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_1015),
.A2(n_86),
.B(n_85),
.Y(n_1082)
);

BUFx6f_ASAP7_75t_L g1083 ( 
.A(n_969),
.Y(n_1083)
);

OAI21x1_ASAP7_75t_L g1084 ( 
.A1(n_1001),
.A2(n_93),
.B(n_92),
.Y(n_1084)
);

OAI21xp33_ASAP7_75t_L g1085 ( 
.A1(n_959),
.A2(n_26),
.B(n_29),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1017),
.B(n_1018),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_972),
.B(n_30),
.Y(n_1087)
);

OA21x2_ASAP7_75t_L g1088 ( 
.A1(n_981),
.A2(n_95),
.B(n_94),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_985),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_974),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_1090)
);

OAI21x1_ASAP7_75t_L g1091 ( 
.A1(n_988),
.A2(n_1021),
.B(n_949),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_976),
.A2(n_97),
.B(n_96),
.Y(n_1092)
);

OR2x6_ASAP7_75t_L g1093 ( 
.A(n_980),
.B(n_1008),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_977),
.B(n_31),
.Y(n_1094)
);

INVxp67_ASAP7_75t_SL g1095 ( 
.A(n_991),
.Y(n_1095)
);

OAI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_992),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_1096)
);

CKINVDCx16_ASAP7_75t_R g1097 ( 
.A(n_1046),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1056),
.Y(n_1098)
);

INVx2_ASAP7_75t_SL g1099 ( 
.A(n_1053),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_1045),
.A2(n_999),
.B(n_998),
.Y(n_1100)
);

AOI221xp5_ASAP7_75t_L g1101 ( 
.A1(n_1047),
.A2(n_1006),
.B1(n_1000),
.B2(n_1011),
.C(n_38),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1039),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1034),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_SL g1104 ( 
.A1(n_1043),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1051),
.A2(n_102),
.B(n_98),
.Y(n_1105)
);

OAI221xp5_ASAP7_75t_L g1106 ( 
.A1(n_1085),
.A2(n_37),
.B1(n_39),
.B2(n_40),
.C(n_41),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_1034),
.Y(n_1107)
);

AO32x2_ASAP7_75t_L g1108 ( 
.A1(n_1060),
.A2(n_1081),
.A3(n_1090),
.B1(n_1050),
.B2(n_1055),
.Y(n_1108)
);

OAI21x1_ASAP7_75t_L g1109 ( 
.A1(n_1033),
.A2(n_106),
.B(n_103),
.Y(n_1109)
);

NAND2x1p5_ASAP7_75t_L g1110 ( 
.A(n_1042),
.B(n_1049),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1042),
.B(n_40),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_1030),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1064),
.Y(n_1113)
);

NAND2x1p5_ASAP7_75t_L g1114 ( 
.A(n_1049),
.B(n_109),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_1032),
.Y(n_1115)
);

AOI22x1_ASAP7_75t_L g1116 ( 
.A1(n_1092),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_1116)
);

OAI22xp5_ASAP7_75t_L g1117 ( 
.A1(n_1062),
.A2(n_42),
.B1(n_46),
.B2(n_47),
.Y(n_1117)
);

INVx1_ASAP7_75t_L g1118 ( 
.A(n_1064),
.Y(n_1118)
);

BUFx3_ASAP7_75t_L g1119 ( 
.A(n_1052),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1040),
.Y(n_1120)
);

OAI21x1_ASAP7_75t_L g1121 ( 
.A1(n_1057),
.A2(n_111),
.B(n_110),
.Y(n_1121)
);

NAND3xp33_ASAP7_75t_SL g1122 ( 
.A(n_1079),
.B(n_46),
.C(n_47),
.Y(n_1122)
);

OAI21x1_ASAP7_75t_L g1123 ( 
.A1(n_1048),
.A2(n_114),
.B(n_113),
.Y(n_1123)
);

AND2x4_ASAP7_75t_L g1124 ( 
.A(n_1093),
.B(n_356),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1040),
.Y(n_1125)
);

BUFx2_ASAP7_75t_SL g1126 ( 
.A(n_1071),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1053),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1028),
.B(n_49),
.Y(n_1128)
);

AND2x2_ASAP7_75t_L g1129 ( 
.A(n_1036),
.B(n_50),
.Y(n_1129)
);

AOI21xp5_ASAP7_75t_L g1130 ( 
.A1(n_1086),
.A2(n_116),
.B(n_115),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1068),
.A2(n_119),
.B(n_117),
.Y(n_1131)
);

AND2x4_ASAP7_75t_L g1132 ( 
.A(n_1093),
.B(n_350),
.Y(n_1132)
);

OAI21x1_ASAP7_75t_L g1133 ( 
.A1(n_1068),
.A2(n_234),
.B(n_345),
.Y(n_1133)
);

O2A1O1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1096),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_1134)
);

BUFx3_ASAP7_75t_L g1135 ( 
.A(n_1053),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1082),
.A2(n_120),
.B(n_122),
.Y(n_1136)
);

AO21x2_ASAP7_75t_L g1137 ( 
.A1(n_1038),
.A2(n_123),
.B(n_125),
.Y(n_1137)
);

BUFx6f_ASAP7_75t_L g1138 ( 
.A(n_1066),
.Y(n_1138)
);

AOI22xp33_ASAP7_75t_L g1139 ( 
.A1(n_1054),
.A2(n_126),
.B1(n_128),
.B2(n_132),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1044),
.Y(n_1140)
);

AND2x2_ASAP7_75t_SL g1141 ( 
.A(n_1031),
.B(n_133),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_1095),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_1077),
.Y(n_1143)
);

AOI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_1087),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_1144)
);

OA21x2_ASAP7_75t_L g1145 ( 
.A1(n_1037),
.A2(n_147),
.B(n_148),
.Y(n_1145)
);

BUFx3_ASAP7_75t_L g1146 ( 
.A(n_1083),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1084),
.A2(n_149),
.B(n_151),
.Y(n_1147)
);

OAI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1065),
.A2(n_152),
.B(n_154),
.Y(n_1148)
);

OAI21x1_ASAP7_75t_L g1149 ( 
.A1(n_1072),
.A2(n_1069),
.B(n_1091),
.Y(n_1149)
);

AND2x4_ASAP7_75t_L g1150 ( 
.A(n_1031),
.B(n_1063),
.Y(n_1150)
);

INVx3_ASAP7_75t_SL g1151 ( 
.A(n_1083),
.Y(n_1151)
);

OAI22xp5_ASAP7_75t_L g1152 ( 
.A1(n_1073),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1075),
.A2(n_158),
.B1(n_161),
.B2(n_164),
.Y(n_1153)
);

AND2x4_ASAP7_75t_L g1154 ( 
.A(n_1066),
.B(n_348),
.Y(n_1154)
);

OAI21x1_ASAP7_75t_L g1155 ( 
.A1(n_1088),
.A2(n_165),
.B(n_166),
.Y(n_1155)
);

OAI21x1_ASAP7_75t_L g1156 ( 
.A1(n_1088),
.A2(n_167),
.B(n_170),
.Y(n_1156)
);

NOR2xp33_ASAP7_75t_SL g1157 ( 
.A(n_1027),
.B(n_172),
.Y(n_1157)
);

CKINVDCx16_ASAP7_75t_R g1158 ( 
.A(n_1078),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1083),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1066),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1035),
.Y(n_1161)
);

INVx2_ASAP7_75t_SL g1162 ( 
.A(n_1089),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1041),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1074),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_1103),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1103),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1107),
.B(n_1118),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_1107),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1118),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1113),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1120),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1120),
.Y(n_1172)
);

AO31x2_ASAP7_75t_L g1173 ( 
.A1(n_1164),
.A2(n_1058),
.A3(n_1029),
.B(n_1067),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1161),
.B(n_1059),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1125),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1125),
.Y(n_1176)
);

OR2x2_ASAP7_75t_L g1177 ( 
.A(n_1158),
.B(n_1094),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1100),
.A2(n_1102),
.B(n_1148),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1115),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_1150),
.B(n_1074),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1112),
.Y(n_1181)
);

AO31x2_ASAP7_75t_L g1182 ( 
.A1(n_1164),
.A2(n_1076),
.A3(n_1059),
.B(n_1074),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1127),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1129),
.B(n_1076),
.Y(n_1184)
);

OAI21x1_ASAP7_75t_L g1185 ( 
.A1(n_1149),
.A2(n_1070),
.B(n_1059),
.Y(n_1185)
);

HB1xp67_ASAP7_75t_L g1186 ( 
.A(n_1126),
.Y(n_1186)
);

OAI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_1141),
.A2(n_1080),
.B1(n_1061),
.B2(n_179),
.Y(n_1187)
);

OAI22xp5_ASAP7_75t_L g1188 ( 
.A1(n_1111),
.A2(n_173),
.B1(n_174),
.B2(n_180),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1161),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1098),
.Y(n_1190)
);

OAI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_1106),
.A2(n_182),
.B1(n_185),
.B2(n_188),
.Y(n_1191)
);

AND2x2_ASAP7_75t_L g1192 ( 
.A(n_1128),
.B(n_189),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1143),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_1162),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1140),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1155),
.A2(n_191),
.B(n_196),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1124),
.A2(n_198),
.B1(n_200),
.B2(n_201),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1122),
.A2(n_202),
.B1(n_205),
.B2(n_207),
.Y(n_1198)
);

INVx2_ASAP7_75t_L g1199 ( 
.A(n_1140),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1163),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1150),
.B(n_343),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1163),
.Y(n_1202)
);

BUFx3_ASAP7_75t_L g1203 ( 
.A(n_1135),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1160),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1102),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1160),
.Y(n_1206)
);

O2A1O1Ixp33_ASAP7_75t_SL g1207 ( 
.A1(n_1134),
.A2(n_1117),
.B(n_1142),
.C(n_1153),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1145),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1138),
.Y(n_1209)
);

OAI21x1_ASAP7_75t_L g1210 ( 
.A1(n_1156),
.A2(n_208),
.B(n_209),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1138),
.Y(n_1211)
);

HB1xp67_ASAP7_75t_L g1212 ( 
.A(n_1138),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1099),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_1159),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1108),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_1146),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1108),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_1097),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_1109),
.A2(n_1133),
.B(n_1131),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1145),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1108),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_1119),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1154),
.Y(n_1223)
);

OR2x2_ASAP7_75t_L g1224 ( 
.A(n_1151),
.B(n_210),
.Y(n_1224)
);

AND2x2_ASAP7_75t_L g1225 ( 
.A(n_1124),
.B(n_211),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1132),
.B(n_213),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_1154),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1132),
.B(n_342),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1137),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1137),
.Y(n_1230)
);

OAI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1157),
.A2(n_216),
.B1(n_217),
.B2(n_219),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1110),
.B(n_220),
.Y(n_1232)
);

INVx1_ASAP7_75t_SL g1233 ( 
.A(n_1114),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1116),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1105),
.Y(n_1235)
);

HB1xp67_ASAP7_75t_L g1236 ( 
.A(n_1116),
.Y(n_1236)
);

HB1xp67_ASAP7_75t_L g1237 ( 
.A(n_1104),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1139),
.B(n_1144),
.Y(n_1238)
);

OR2x6_ASAP7_75t_L g1239 ( 
.A(n_1130),
.B(n_222),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1165),
.Y(n_1240)
);

NAND2xp33_ASAP7_75t_R g1241 ( 
.A(n_1218),
.B(n_1222),
.Y(n_1241)
);

INVxp67_ASAP7_75t_L g1242 ( 
.A(n_1214),
.Y(n_1242)
);

AND2x4_ASAP7_75t_L g1243 ( 
.A(n_1167),
.B(n_1147),
.Y(n_1243)
);

AND2x4_ASAP7_75t_L g1244 ( 
.A(n_1203),
.B(n_1136),
.Y(n_1244)
);

XNOR2xp5_ASAP7_75t_L g1245 ( 
.A(n_1218),
.B(n_1101),
.Y(n_1245)
);

NAND2xp33_ASAP7_75t_R g1246 ( 
.A(n_1222),
.B(n_223),
.Y(n_1246)
);

AND2x2_ASAP7_75t_L g1247 ( 
.A(n_1184),
.B(n_1152),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1203),
.B(n_1121),
.Y(n_1248)
);

NAND2xp33_ASAP7_75t_R g1249 ( 
.A(n_1216),
.B(n_227),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1190),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1212),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1193),
.Y(n_1252)
);

NOR2xp33_ASAP7_75t_R g1253 ( 
.A(n_1226),
.B(n_228),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_R g1254 ( 
.A(n_1225),
.B(n_236),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1189),
.B(n_1123),
.Y(n_1255)
);

XNOR2xp5_ASAP7_75t_L g1256 ( 
.A(n_1237),
.B(n_1179),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_1186),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_R g1258 ( 
.A(n_1192),
.B(n_238),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_R g1259 ( 
.A(n_1224),
.B(n_239),
.Y(n_1259)
);

BUFx3_ASAP7_75t_L g1260 ( 
.A(n_1209),
.Y(n_1260)
);

BUFx10_ASAP7_75t_L g1261 ( 
.A(n_1211),
.Y(n_1261)
);

NAND2xp33_ASAP7_75t_R g1262 ( 
.A(n_1192),
.B(n_240),
.Y(n_1262)
);

NOR2xp33_ASAP7_75t_R g1263 ( 
.A(n_1228),
.B(n_241),
.Y(n_1263)
);

AND2x4_ASAP7_75t_L g1264 ( 
.A(n_1167),
.B(n_244),
.Y(n_1264)
);

NOR2xp33_ASAP7_75t_R g1265 ( 
.A(n_1177),
.B(n_245),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1183),
.Y(n_1266)
);

BUFx3_ASAP7_75t_L g1267 ( 
.A(n_1213),
.Y(n_1267)
);

OR2x6_ASAP7_75t_L g1268 ( 
.A(n_1223),
.B(n_248),
.Y(n_1268)
);

NAND2xp33_ASAP7_75t_R g1269 ( 
.A(n_1232),
.B(n_250),
.Y(n_1269)
);

NOR2xp33_ASAP7_75t_R g1270 ( 
.A(n_1232),
.B(n_252),
.Y(n_1270)
);

HB1xp67_ASAP7_75t_L g1271 ( 
.A(n_1166),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1194),
.B(n_254),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1204),
.B(n_255),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_R g1274 ( 
.A(n_1233),
.B(n_257),
.Y(n_1274)
);

NAND2xp33_ASAP7_75t_SL g1275 ( 
.A(n_1198),
.B(n_259),
.Y(n_1275)
);

NAND2xp33_ASAP7_75t_R g1276 ( 
.A(n_1238),
.B(n_261),
.Y(n_1276)
);

AND2x4_ASAP7_75t_L g1277 ( 
.A(n_1180),
.B(n_264),
.Y(n_1277)
);

BUFx3_ASAP7_75t_L g1278 ( 
.A(n_1206),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_R g1279 ( 
.A(n_1201),
.B(n_268),
.Y(n_1279)
);

INVxp67_ASAP7_75t_L g1280 ( 
.A(n_1181),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1166),
.B(n_269),
.Y(n_1281)
);

NAND2xp33_ASAP7_75t_R g1282 ( 
.A(n_1238),
.B(n_270),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_R g1283 ( 
.A(n_1227),
.B(n_271),
.Y(n_1283)
);

OR2x6_ASAP7_75t_L g1284 ( 
.A(n_1180),
.B(n_272),
.Y(n_1284)
);

BUFx3_ASAP7_75t_L g1285 ( 
.A(n_1170),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1168),
.B(n_273),
.Y(n_1286)
);

OR2x6_ASAP7_75t_L g1287 ( 
.A(n_1180),
.B(n_1168),
.Y(n_1287)
);

NAND2xp33_ASAP7_75t_R g1288 ( 
.A(n_1215),
.B(n_274),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1170),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1169),
.Y(n_1290)
);

NOR2xp33_ASAP7_75t_R g1291 ( 
.A(n_1217),
.B(n_277),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_R g1292 ( 
.A(n_1221),
.B(n_279),
.Y(n_1292)
);

BUFx10_ASAP7_75t_L g1293 ( 
.A(n_1239),
.Y(n_1293)
);

BUFx3_ASAP7_75t_L g1294 ( 
.A(n_1169),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1173),
.B(n_283),
.Y(n_1295)
);

XOR2xp5_ASAP7_75t_L g1296 ( 
.A(n_1197),
.B(n_284),
.Y(n_1296)
);

XNOR2xp5_ASAP7_75t_L g1297 ( 
.A(n_1231),
.B(n_285),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1200),
.Y(n_1298)
);

INVxp67_ASAP7_75t_L g1299 ( 
.A(n_1202),
.Y(n_1299)
);

XNOR2xp5_ASAP7_75t_L g1300 ( 
.A(n_1231),
.B(n_286),
.Y(n_1300)
);

NOR2xp33_ASAP7_75t_R g1301 ( 
.A(n_1195),
.B(n_287),
.Y(n_1301)
);

AND2x4_ASAP7_75t_L g1302 ( 
.A(n_1173),
.B(n_289),
.Y(n_1302)
);

NAND2xp33_ASAP7_75t_R g1303 ( 
.A(n_1174),
.B(n_1239),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_SL g1304 ( 
.A(n_1187),
.B(n_290),
.Y(n_1304)
);

AND2x4_ASAP7_75t_L g1305 ( 
.A(n_1173),
.B(n_291),
.Y(n_1305)
);

AND2x4_ASAP7_75t_L g1306 ( 
.A(n_1173),
.B(n_292),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1174),
.B(n_293),
.Y(n_1307)
);

AND2x4_ASAP7_75t_L g1308 ( 
.A(n_1199),
.B(n_294),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1199),
.Y(n_1309)
);

NOR2xp33_ASAP7_75t_R g1310 ( 
.A(n_1234),
.B(n_1236),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1298),
.Y(n_1311)
);

INVx3_ASAP7_75t_L g1312 ( 
.A(n_1243),
.Y(n_1312)
);

OR2x2_ASAP7_75t_L g1313 ( 
.A(n_1240),
.B(n_1205),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1287),
.B(n_1299),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1309),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1287),
.B(n_1205),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1256),
.B(n_1188),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1290),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1289),
.Y(n_1319)
);

BUFx3_ASAP7_75t_L g1320 ( 
.A(n_1257),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1271),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1294),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1280),
.Y(n_1323)
);

BUFx2_ASAP7_75t_L g1324 ( 
.A(n_1310),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1250),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1252),
.Y(n_1326)
);

BUFx3_ASAP7_75t_L g1327 ( 
.A(n_1260),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1255),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1285),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1243),
.B(n_1171),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1305),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1305),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1247),
.B(n_1171),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1295),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1302),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1278),
.Y(n_1336)
);

INVx3_ASAP7_75t_L g1337 ( 
.A(n_1293),
.Y(n_1337)
);

AND2x4_ASAP7_75t_L g1338 ( 
.A(n_1277),
.B(n_1172),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1264),
.B(n_1172),
.Y(n_1339)
);

INVxp67_ASAP7_75t_SL g1340 ( 
.A(n_1266),
.Y(n_1340)
);

BUFx6f_ASAP7_75t_L g1341 ( 
.A(n_1284),
.Y(n_1341)
);

AND2x2_ASAP7_75t_L g1342 ( 
.A(n_1264),
.B(n_1242),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1306),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1244),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1251),
.Y(n_1345)
);

INVx2_ASAP7_75t_L g1346 ( 
.A(n_1248),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1267),
.B(n_1175),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1307),
.B(n_1175),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1277),
.B(n_1176),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_1281),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1284),
.B(n_1176),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1286),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1303),
.Y(n_1353)
);

INVx2_ASAP7_75t_L g1354 ( 
.A(n_1308),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1297),
.A2(n_1198),
.B1(n_1239),
.B2(n_1191),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1261),
.B(n_1178),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1272),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1273),
.B(n_1182),
.Y(n_1358)
);

AND2x4_ASAP7_75t_L g1359 ( 
.A(n_1268),
.B(n_1182),
.Y(n_1359)
);

INVxp67_ASAP7_75t_SL g1360 ( 
.A(n_1288),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1245),
.B(n_1182),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1291),
.B(n_1182),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1292),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1361),
.A2(n_1275),
.B1(n_1300),
.B2(n_1304),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1333),
.B(n_1312),
.Y(n_1365)
);

AND2x2_ASAP7_75t_L g1366 ( 
.A(n_1333),
.B(n_1185),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1319),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1312),
.B(n_1185),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1311),
.Y(n_1369)
);

NOR2xp33_ASAP7_75t_L g1370 ( 
.A(n_1320),
.B(n_1296),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1340),
.B(n_1301),
.Y(n_1371)
);

INVx2_ASAP7_75t_SL g1372 ( 
.A(n_1327),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1327),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1312),
.B(n_1235),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1320),
.B(n_1241),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1311),
.Y(n_1376)
);

OAI31xp33_ASAP7_75t_L g1377 ( 
.A1(n_1355),
.A2(n_1207),
.A3(n_1282),
.B(n_1276),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1330),
.B(n_1235),
.Y(n_1378)
);

AND2x2_ASAP7_75t_L g1379 ( 
.A(n_1330),
.B(n_1208),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1315),
.Y(n_1380)
);

AOI221xp5_ASAP7_75t_L g1381 ( 
.A1(n_1317),
.A2(n_1207),
.B1(n_1258),
.B2(n_1265),
.C(n_1254),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_1315),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1323),
.B(n_1253),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1319),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1318),
.Y(n_1385)
);

INVxp67_ASAP7_75t_SL g1386 ( 
.A(n_1356),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1321),
.B(n_1230),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1324),
.B(n_1270),
.Y(n_1388)
);

HB1xp67_ASAP7_75t_L g1389 ( 
.A(n_1345),
.Y(n_1389)
);

OAI222xp33_ASAP7_75t_L g1390 ( 
.A1(n_1360),
.A2(n_1363),
.B1(n_1334),
.B2(n_1353),
.C1(n_1362),
.C2(n_1358),
.Y(n_1390)
);

AND2x4_ASAP7_75t_L g1391 ( 
.A(n_1330),
.B(n_1220),
.Y(n_1391)
);

INVx2_ASAP7_75t_L g1392 ( 
.A(n_1318),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1325),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1321),
.Y(n_1394)
);

AND2x2_ASAP7_75t_L g1395 ( 
.A(n_1330),
.B(n_1220),
.Y(n_1395)
);

AND2x2_ASAP7_75t_L g1396 ( 
.A(n_1386),
.B(n_1324),
.Y(n_1396)
);

OR2x2_ASAP7_75t_L g1397 ( 
.A(n_1389),
.B(n_1323),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1387),
.Y(n_1398)
);

AND2x2_ASAP7_75t_L g1399 ( 
.A(n_1365),
.B(n_1344),
.Y(n_1399)
);

NAND2x1_ASAP7_75t_L g1400 ( 
.A(n_1372),
.B(n_1328),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1365),
.B(n_1313),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1394),
.B(n_1328),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1369),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1372),
.B(n_1344),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1369),
.Y(n_1405)
);

AND2x2_ASAP7_75t_L g1406 ( 
.A(n_1373),
.B(n_1342),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1394),
.B(n_1352),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1376),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1373),
.B(n_1346),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1376),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1380),
.B(n_1352),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1366),
.B(n_1346),
.Y(n_1412)
);

INVx2_ASAP7_75t_L g1413 ( 
.A(n_1387),
.Y(n_1413)
);

AND2x4_ASAP7_75t_L g1414 ( 
.A(n_1366),
.B(n_1314),
.Y(n_1414)
);

NOR2xp33_ASAP7_75t_SL g1415 ( 
.A(n_1377),
.B(n_1363),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1385),
.Y(n_1416)
);

AND2x2_ASAP7_75t_L g1417 ( 
.A(n_1368),
.B(n_1336),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1415),
.A2(n_1341),
.B1(n_1262),
.B2(n_1371),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1411),
.Y(n_1419)
);

NAND2x1_ASAP7_75t_L g1420 ( 
.A(n_1396),
.B(n_1375),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1396),
.B(n_1380),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1407),
.Y(n_1422)
);

NAND2xp33_ASAP7_75t_SL g1423 ( 
.A(n_1400),
.B(n_1388),
.Y(n_1423)
);

CKINVDCx5p33_ASAP7_75t_R g1424 ( 
.A(n_1397),
.Y(n_1424)
);

AO221x2_ASAP7_75t_L g1425 ( 
.A1(n_1403),
.A2(n_1390),
.B1(n_1383),
.B2(n_1377),
.C(n_1381),
.Y(n_1425)
);

OAI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1401),
.A2(n_1341),
.B1(n_1331),
.B2(n_1334),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1402),
.A2(n_1341),
.B1(n_1331),
.B2(n_1249),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1417),
.A2(n_1246),
.B1(n_1269),
.B2(n_1364),
.Y(n_1428)
);

OAI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1398),
.A2(n_1259),
.B1(n_1357),
.B2(n_1322),
.C(n_1336),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1406),
.B(n_1370),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1404),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1420),
.B(n_1431),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1419),
.B(n_1416),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1422),
.B(n_1416),
.Y(n_1434)
);

INVx1_ASAP7_75t_SL g1435 ( 
.A(n_1423),
.Y(n_1435)
);

INVx2_ASAP7_75t_SL g1436 ( 
.A(n_1424),
.Y(n_1436)
);

INVx2_ASAP7_75t_L g1437 ( 
.A(n_1421),
.Y(n_1437)
);

INVx1_ASAP7_75t_SL g1438 ( 
.A(n_1428),
.Y(n_1438)
);

AND2x2_ASAP7_75t_L g1439 ( 
.A(n_1430),
.B(n_1417),
.Y(n_1439)
);

INVx1_ASAP7_75t_SL g1440 ( 
.A(n_1425),
.Y(n_1440)
);

BUFx3_ASAP7_75t_L g1441 ( 
.A(n_1425),
.Y(n_1441)
);

INVx1_ASAP7_75t_SL g1442 ( 
.A(n_1418),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1427),
.B(n_1405),
.Y(n_1443)
);

INVxp67_ASAP7_75t_L g1444 ( 
.A(n_1429),
.Y(n_1444)
);

INVx1_ASAP7_75t_SL g1445 ( 
.A(n_1426),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1420),
.B(n_1414),
.Y(n_1446)
);

NAND2xp5_ASAP7_75t_L g1447 ( 
.A(n_1419),
.B(n_1408),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1419),
.B(n_1410),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1447),
.Y(n_1449)
);

OAI322xp33_ASAP7_75t_L g1450 ( 
.A1(n_1440),
.A2(n_1382),
.A3(n_1313),
.B1(n_1385),
.B2(n_1392),
.C1(n_1413),
.C2(n_1398),
.Y(n_1450)
);

AOI31xp33_ASAP7_75t_L g1451 ( 
.A1(n_1435),
.A2(n_1342),
.A3(n_1404),
.B(n_1414),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1448),
.Y(n_1452)
);

NOR2x1_ASAP7_75t_L g1453 ( 
.A(n_1441),
.B(n_1414),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1433),
.Y(n_1454)
);

O2A1O1Ixp33_ASAP7_75t_L g1455 ( 
.A1(n_1441),
.A2(n_1239),
.B(n_1268),
.C(n_1350),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1439),
.B(n_1399),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1434),
.Y(n_1457)
);

OAI21xp5_ASAP7_75t_L g1458 ( 
.A1(n_1444),
.A2(n_1409),
.B(n_1399),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1437),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1459),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1456),
.B(n_1432),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1453),
.A2(n_1436),
.B1(n_1438),
.B2(n_1432),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1449),
.B(n_1452),
.Y(n_1463)
);

NOR2x1_ASAP7_75t_L g1464 ( 
.A(n_1451),
.B(n_1446),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1454),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1457),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1458),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1450),
.Y(n_1468)
);

NOR2xp33_ASAP7_75t_L g1469 ( 
.A(n_1451),
.B(n_1436),
.Y(n_1469)
);

INVxp33_ASAP7_75t_SL g1470 ( 
.A(n_1462),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_L g1471 ( 
.A(n_1462),
.B(n_1437),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1460),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1467),
.B(n_1443),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1463),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1465),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1466),
.Y(n_1476)
);

OAI211xp5_ASAP7_75t_SL g1477 ( 
.A1(n_1473),
.A2(n_1464),
.B(n_1469),
.C(n_1468),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1471),
.A2(n_1470),
.B1(n_1474),
.B2(n_1472),
.C(n_1475),
.Y(n_1478)
);

NAND3xp33_ASAP7_75t_L g1479 ( 
.A(n_1476),
.B(n_1461),
.C(n_1455),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1470),
.B(n_1446),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1473),
.B(n_1445),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_L g1482 ( 
.A(n_1470),
.B(n_1442),
.Y(n_1482)
);

NAND5xp2_ASAP7_75t_L g1483 ( 
.A(n_1470),
.B(n_1368),
.C(n_1409),
.D(n_1314),
.E(n_1351),
.Y(n_1483)
);

O2A1O1Ixp33_ASAP7_75t_L g1484 ( 
.A1(n_1470),
.A2(n_1362),
.B(n_1350),
.C(n_1382),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1470),
.B(n_1412),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1480),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1477),
.A2(n_1357),
.B1(n_1341),
.B2(n_1359),
.Y(n_1487)
);

AOI21xp5_ASAP7_75t_L g1488 ( 
.A1(n_1482),
.A2(n_1392),
.B(n_1412),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1479),
.A2(n_1341),
.B1(n_1413),
.B2(n_1337),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1481),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1485),
.Y(n_1491)
);

AOI21xp5_ASAP7_75t_L g1492 ( 
.A1(n_1478),
.A2(n_1374),
.B(n_1337),
.Y(n_1492)
);

NAND4xp25_ASAP7_75t_SL g1493 ( 
.A(n_1484),
.B(n_1483),
.C(n_1332),
.D(n_1374),
.Y(n_1493)
);

NAND4xp75_ASAP7_75t_L g1494 ( 
.A(n_1486),
.B(n_1274),
.C(n_1263),
.D(n_1347),
.Y(n_1494)
);

AOI22xp5_ASAP7_75t_L g1495 ( 
.A1(n_1487),
.A2(n_1359),
.B1(n_1358),
.B2(n_1322),
.Y(n_1495)
);

NOR4xp75_ASAP7_75t_L g1496 ( 
.A(n_1489),
.B(n_1337),
.C(n_1279),
.D(n_1347),
.Y(n_1496)
);

XNOR2xp5_ASAP7_75t_L g1497 ( 
.A(n_1491),
.B(n_1490),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1493),
.B(n_1329),
.Y(n_1498)
);

XNOR2xp5_ASAP7_75t_L g1499 ( 
.A(n_1492),
.B(n_1359),
.Y(n_1499)
);

AND2x4_ASAP7_75t_L g1500 ( 
.A(n_1488),
.B(n_1378),
.Y(n_1500)
);

NAND2xp33_ASAP7_75t_SL g1501 ( 
.A(n_1497),
.B(n_1283),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1498),
.B(n_1393),
.Y(n_1502)
);

NAND3xp33_ASAP7_75t_SL g1503 ( 
.A(n_1496),
.B(n_1335),
.C(n_1343),
.Y(n_1503)
);

NOR2xp33_ASAP7_75t_R g1504 ( 
.A(n_1499),
.B(n_297),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_R g1505 ( 
.A(n_1494),
.B(n_304),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_R g1506 ( 
.A(n_1500),
.B(n_305),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1495),
.B(n_1393),
.Y(n_1507)
);

NAND2xp33_ASAP7_75t_SL g1508 ( 
.A(n_1497),
.B(n_1332),
.Y(n_1508)
);

NAND2xp33_ASAP7_75t_SL g1509 ( 
.A(n_1497),
.B(n_1343),
.Y(n_1509)
);

OAI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1502),
.A2(n_1329),
.B1(n_1348),
.B2(n_1335),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1507),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1501),
.A2(n_1196),
.B(n_1210),
.Y(n_1512)
);

AOI22xp5_ASAP7_75t_L g1513 ( 
.A1(n_1509),
.A2(n_1351),
.B1(n_1354),
.B2(n_1378),
.Y(n_1513)
);

AOI211xp5_ASAP7_75t_L g1514 ( 
.A1(n_1505),
.A2(n_1196),
.B(n_1210),
.C(n_1339),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1508),
.Y(n_1515)
);

AO22x2_ASAP7_75t_L g1516 ( 
.A1(n_1503),
.A2(n_1354),
.B1(n_1367),
.B2(n_1384),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1506),
.Y(n_1517)
);

OAI21xp33_ASAP7_75t_L g1518 ( 
.A1(n_1504),
.A2(n_1339),
.B(n_1395),
.Y(n_1518)
);

INVx2_ASAP7_75t_L g1519 ( 
.A(n_1507),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1506),
.B(n_1384),
.Y(n_1520)
);

AOI221xp5_ASAP7_75t_SL g1521 ( 
.A1(n_1515),
.A2(n_1326),
.B1(n_1325),
.B2(n_1367),
.C(n_1395),
.Y(n_1521)
);

AOI22x1_ASAP7_75t_L g1522 ( 
.A1(n_1517),
.A2(n_1349),
.B1(n_1326),
.B2(n_1338),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1511),
.B(n_1391),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1519),
.Y(n_1524)
);

AOI21xp5_ASAP7_75t_L g1525 ( 
.A1(n_1514),
.A2(n_1219),
.B(n_1391),
.Y(n_1525)
);

BUFx3_ASAP7_75t_L g1526 ( 
.A(n_1520),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1512),
.A2(n_306),
.B(n_307),
.Y(n_1527)
);

XNOR2xp5_ASAP7_75t_L g1528 ( 
.A(n_1524),
.B(n_1516),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1523),
.B(n_1510),
.Y(n_1529)
);

NOR2xp33_ASAP7_75t_L g1530 ( 
.A(n_1526),
.B(n_1518),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1525),
.A2(n_1513),
.B1(n_1391),
.B2(n_1338),
.Y(n_1531)
);

NAND3xp33_ASAP7_75t_L g1532 ( 
.A(n_1521),
.B(n_1391),
.C(n_1379),
.Y(n_1532)
);

AOI31xp33_ASAP7_75t_L g1533 ( 
.A1(n_1530),
.A2(n_1527),
.A3(n_1522),
.B(n_1349),
.Y(n_1533)
);

AOI31xp33_ASAP7_75t_L g1534 ( 
.A1(n_1528),
.A2(n_1522),
.A3(n_1338),
.B(n_316),
.Y(n_1534)
);

AOI31xp33_ASAP7_75t_L g1535 ( 
.A1(n_1529),
.A2(n_1338),
.A3(n_315),
.B(n_317),
.Y(n_1535)
);

AOI211xp5_ASAP7_75t_L g1536 ( 
.A1(n_1534),
.A2(n_1531),
.B(n_1532),
.C(n_1219),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1533),
.A2(n_1230),
.B1(n_1229),
.B2(n_1208),
.Y(n_1537)
);

OAI22x1_ASAP7_75t_L g1538 ( 
.A1(n_1536),
.A2(n_1535),
.B1(n_1316),
.B2(n_1379),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_1538),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1539),
.A2(n_1537),
.B1(n_322),
.B2(n_323),
.C(n_325),
.Y(n_1540)
);

AOI211xp5_ASAP7_75t_L g1541 ( 
.A1(n_1540),
.A2(n_313),
.B(n_330),
.C(n_331),
.Y(n_1541)
);


endmodule