module real_aes_17258_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_565;
wire n_443;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_756;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
AND2x4_ASAP7_75t_L g114 ( .A(n_0), .B(n_115), .Y(n_114) );
AOI22xp5_ASAP7_75t_L g599 ( .A1(n_1), .A2(n_4), .B1(n_216), .B2(n_600), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g153 ( .A1(n_2), .A2(n_44), .B1(n_154), .B2(n_156), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_3), .A2(n_25), .B1(n_156), .B2(n_180), .Y(n_590) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_5), .A2(n_16), .B1(n_197), .B2(n_234), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_6), .A2(n_61), .B1(n_182), .B2(n_254), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_7), .A2(n_17), .B1(n_154), .B2(n_201), .Y(n_523) );
INVx1_ASAP7_75t_L g115 ( .A(n_8), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g585 ( .A(n_9), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g270 ( .A(n_10), .Y(n_270) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_11), .A2(n_18), .B1(n_199), .B2(n_253), .Y(n_252) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_12), .A2(n_65), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_12), .Y(n_824) );
BUFx2_ASAP7_75t_L g111 ( .A(n_13), .Y(n_111) );
OR2x2_ASAP7_75t_L g135 ( .A(n_13), .B(n_39), .Y(n_135) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_14), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g237 ( .A(n_15), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g215 ( .A1(n_19), .A2(n_100), .B1(n_197), .B2(n_216), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g828 ( .A1(n_20), .A2(n_490), .B(n_829), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_21), .A2(n_40), .B1(n_230), .B2(n_231), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_22), .B(n_198), .Y(n_271) );
OAI22x1_ASAP7_75t_SL g821 ( .A1(n_23), .A2(n_822), .B1(n_823), .B2(n_826), .Y(n_821) );
CKINVDCx5p33_ASAP7_75t_R g826 ( .A(n_23), .Y(n_826) );
OAI21x1_ASAP7_75t_L g170 ( .A1(n_24), .A2(n_59), .B(n_171), .Y(n_170) );
CKINVDCx5p33_ASAP7_75t_R g223 ( .A(n_26), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g593 ( .A(n_27), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_28), .B(n_160), .Y(n_547) );
INVx4_ASAP7_75t_R g536 ( .A(n_29), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g161 ( .A1(n_30), .A2(n_48), .B1(n_162), .B2(n_164), .Y(n_161) );
AOI22xp33_ASAP7_75t_L g243 ( .A1(n_31), .A2(n_55), .B1(n_164), .B2(n_197), .Y(n_243) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_32), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_33), .B(n_230), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g206 ( .A(n_34), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_35), .B(n_156), .Y(n_554) );
INVx1_ASAP7_75t_L g602 ( .A(n_36), .Y(n_602) );
A2O1A1Ixp33_ASAP7_75t_SL g583 ( .A1(n_37), .A2(n_154), .B(n_166), .C(n_584), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_38), .A2(n_56), .B1(n_154), .B2(n_164), .Y(n_591) );
HB1xp67_ASAP7_75t_L g110 ( .A(n_39), .Y(n_110) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_41), .A2(n_88), .B1(n_154), .B2(n_179), .Y(n_178) );
OAI22xp5_ASAP7_75t_SL g138 ( .A1(n_42), .A2(n_54), .B1(n_139), .B2(n_140), .Y(n_138) );
INVx1_ASAP7_75t_L g140 ( .A(n_42), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g256 ( .A1(n_43), .A2(n_47), .B1(n_154), .B2(n_201), .Y(n_256) );
CKINVDCx5p33_ASAP7_75t_R g581 ( .A(n_45), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g218 ( .A1(n_46), .A2(n_60), .B1(n_197), .B2(n_219), .Y(n_218) );
INVx1_ASAP7_75t_L g551 ( .A(n_49), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_50), .B(n_154), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g564 ( .A(n_51), .Y(n_564) );
INVx2_ASAP7_75t_L g123 ( .A(n_52), .Y(n_123) );
BUFx3_ASAP7_75t_L g118 ( .A(n_53), .Y(n_118) );
INVx1_ASAP7_75t_L g133 ( .A(n_53), .Y(n_133) );
INVx1_ASAP7_75t_L g139 ( .A(n_54), .Y(n_139) );
CKINVDCx5p33_ASAP7_75t_R g537 ( .A(n_57), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_58), .A2(n_89), .B1(n_154), .B2(n_164), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_62), .A2(n_77), .B1(n_162), .B2(n_219), .Y(n_242) );
CKINVDCx5p33_ASAP7_75t_R g526 ( .A(n_63), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_64), .A2(n_79), .B1(n_154), .B2(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g825 ( .A(n_65), .Y(n_825) );
CKINVDCx5p33_ASAP7_75t_R g491 ( .A(n_66), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g196 ( .A1(n_67), .A2(n_99), .B1(n_197), .B2(n_199), .Y(n_196) );
AND2x4_ASAP7_75t_L g150 ( .A(n_68), .B(n_151), .Y(n_150) );
INVx1_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_70), .A2(n_91), .B1(n_162), .B2(n_164), .Y(n_598) );
AO22x1_ASAP7_75t_L g512 ( .A1(n_71), .A2(n_78), .B1(n_231), .B2(n_513), .Y(n_512) );
INVx1_ASAP7_75t_L g151 ( .A(n_72), .Y(n_151) );
AND2x2_ASAP7_75t_L g586 ( .A(n_73), .B(n_168), .Y(n_586) );
CKINVDCx14_ASAP7_75t_R g127 ( .A(n_74), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_74), .B(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_75), .B(n_182), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g579 ( .A(n_76), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_80), .B(n_156), .Y(n_565) );
INVx2_ASAP7_75t_L g160 ( .A(n_81), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_82), .B(n_168), .Y(n_544) );
CKINVDCx5p33_ASAP7_75t_R g533 ( .A(n_83), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_84), .A2(n_98), .B1(n_164), .B2(n_182), .Y(n_181) );
CKINVDCx5p33_ASAP7_75t_R g245 ( .A(n_85), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_86), .B(n_189), .Y(n_517) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_87), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_90), .B(n_168), .Y(n_276) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_92), .Y(n_258) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_93), .B(n_168), .Y(n_561) );
INVx1_ASAP7_75t_L g117 ( .A(n_94), .Y(n_117) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_94), .B(n_132), .Y(n_131) );
NAND2xp33_ASAP7_75t_L g274 ( .A(n_95), .B(n_198), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g531 ( .A1(n_96), .A2(n_182), .B(n_184), .C(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g538 ( .A(n_97), .B(n_539), .Y(n_538) );
NAND2xp33_ASAP7_75t_L g569 ( .A(n_101), .B(n_163), .Y(n_569) );
CKINVDCx5p33_ASAP7_75t_R g837 ( .A(n_102), .Y(n_837) );
AOI21xp5_ASAP7_75t_L g103 ( .A1(n_104), .A2(n_119), .B(n_836), .Y(n_103) );
BUFx3_ASAP7_75t_L g104 ( .A(n_105), .Y(n_104) );
INVx6_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx8_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g839 ( .A(n_107), .Y(n_839) );
AND2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_112), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_110), .B(n_111), .Y(n_109) );
NOR3x1_ASAP7_75t_L g112 ( .A(n_113), .B(n_116), .C(n_118), .Y(n_112) );
INVx2_ASAP7_75t_SL g113 ( .A(n_114), .Y(n_113) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx2_ASAP7_75t_L g819 ( .A(n_117), .Y(n_819) );
INVx1_ASAP7_75t_L g499 ( .A(n_118), .Y(n_499) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_118), .B(n_135), .Y(n_835) );
OR2x6_ASAP7_75t_L g119 ( .A(n_120), .B(n_493), .Y(n_119) );
NOR2x1_ASAP7_75t_L g120 ( .A(n_121), .B(n_124), .Y(n_120) );
BUFx8_ASAP7_75t_SL g121 ( .A(n_122), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx1_ASAP7_75t_L g497 ( .A(n_123), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g832 ( .A(n_123), .B(n_833), .Y(n_832) );
AND2x2_ASAP7_75t_L g124 ( .A(n_125), .B(n_485), .Y(n_124) );
NAND2xp5_ASAP7_75t_L g125 ( .A(n_126), .B(n_136), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_127), .B(n_128), .Y(n_126) );
INVx3_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
CKINVDCx8_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
INVx4_ASAP7_75t_L g489 ( .A(n_130), .Y(n_489) );
INVx5_ASAP7_75t_L g492 ( .A(n_130), .Y(n_492) );
AND2x6_ASAP7_75t_SL g130 ( .A(n_131), .B(n_134), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_134), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AOI21xp33_ASAP7_75t_SL g485 ( .A1(n_137), .A2(n_486), .B(n_490), .Y(n_485) );
XNOR2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_141), .Y(n_137) );
OAI22x1_ASAP7_75t_L g502 ( .A1(n_141), .A2(n_503), .B1(n_817), .B2(n_820), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g141 ( .A(n_142), .B(n_395), .Y(n_141) );
NAND4xp75_ASAP7_75t_L g142 ( .A(n_143), .B(n_340), .C(n_360), .D(n_376), .Y(n_142) );
NOR2x1p5_ASAP7_75t_SL g143 ( .A(n_144), .B(n_310), .Y(n_143) );
NAND4xp75_ASAP7_75t_L g144 ( .A(n_145), .B(n_246), .C(n_287), .D(n_296), .Y(n_144) );
NAND2xp5_ASAP7_75t_L g145 ( .A(n_146), .B(n_207), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_174), .Y(n_146) );
AND2x4_ASAP7_75t_L g420 ( .A(n_147), .B(n_347), .Y(n_420) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_148), .Y(n_263) );
INVx2_ASAP7_75t_L g281 ( .A(n_148), .Y(n_281) );
AND2x2_ASAP7_75t_L g304 ( .A(n_148), .B(n_266), .Y(n_304) );
OR2x2_ASAP7_75t_L g359 ( .A(n_148), .B(n_175), .Y(n_359) );
AO31x2_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_152), .A3(n_167), .B(n_172), .Y(n_148) );
INVx2_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
AO31x2_ASAP7_75t_L g227 ( .A1(n_149), .A2(n_176), .A3(n_228), .B(n_236), .Y(n_227) );
AO31x2_ASAP7_75t_L g250 ( .A1(n_149), .A2(n_193), .A3(n_251), .B(n_257), .Y(n_250) );
AO31x2_ASAP7_75t_L g521 ( .A1(n_149), .A2(n_224), .A3(n_522), .B(n_525), .Y(n_521) );
BUFx10_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g186 ( .A(n_150), .Y(n_186) );
INVx1_ASAP7_75t_L g519 ( .A(n_150), .Y(n_519) );
BUFx10_ASAP7_75t_L g556 ( .A(n_150), .Y(n_556) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B1(n_161), .B2(n_165), .Y(n_152) );
INVx1_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx4_ASAP7_75t_L g201 ( .A(n_154), .Y(n_201) );
INVx1_ASAP7_75t_L g219 ( .A(n_154), .Y(n_219) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_155), .Y(n_156) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_155), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
INVx2_ASAP7_75t_L g180 ( .A(n_155), .Y(n_180) );
INVx1_ASAP7_75t_L g182 ( .A(n_155), .Y(n_182) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_155), .Y(n_198) );
INVx1_ASAP7_75t_L g217 ( .A(n_155), .Y(n_217) );
INVx1_ASAP7_75t_L g232 ( .A(n_155), .Y(n_232) );
INVx1_ASAP7_75t_L g235 ( .A(n_155), .Y(n_235) );
INVx1_ASAP7_75t_L g255 ( .A(n_155), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_156), .B(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g214 ( .A1(n_157), .A2(n_165), .B1(n_215), .B2(n_218), .Y(n_214) );
OAI22xp5_ASAP7_75t_L g228 ( .A1(n_157), .A2(n_165), .B1(n_229), .B2(n_233), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_157), .A2(n_165), .B1(n_242), .B2(n_243), .Y(n_241) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g515 ( .A(n_158), .Y(n_515) );
BUFx3_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
INVx2_ASAP7_75t_L g567 ( .A(n_159), .Y(n_567) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx8_ASAP7_75t_L g166 ( .A(n_160), .Y(n_166) );
INVx1_ASAP7_75t_L g184 ( .A(n_160), .Y(n_184) );
INVx1_ASAP7_75t_L g550 ( .A(n_160), .Y(n_550) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
INVx1_ASAP7_75t_L g230 ( .A(n_163), .Y(n_230) );
OAI22xp33_ASAP7_75t_L g535 ( .A1(n_163), .A2(n_235), .B1(n_536), .B2(n_537), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_164), .B(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g600 ( .A(n_164), .Y(n_600) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_165), .A2(n_178), .B1(n_181), .B2(n_183), .Y(n_177) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_165), .A2(n_196), .B1(n_200), .B2(n_202), .Y(n_195) );
OAI22xp5_ASAP7_75t_L g251 ( .A1(n_165), .A2(n_202), .B1(n_252), .B2(n_256), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g272 ( .A1(n_165), .A2(n_273), .B(n_274), .Y(n_272) );
OAI22x1_ASAP7_75t_L g522 ( .A1(n_165), .A2(n_183), .B1(n_523), .B2(n_524), .Y(n_522) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_165), .A2(n_515), .B1(n_590), .B2(n_591), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g597 ( .A1(n_165), .A2(n_183), .B1(n_598), .B2(n_599), .Y(n_597) );
INVx6_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
O2A1O1Ixp5_ASAP7_75t_L g269 ( .A1(n_166), .A2(n_201), .B(n_270), .C(n_271), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_166), .A2(n_512), .B(n_514), .C(n_518), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_166), .A2(n_569), .B(n_570), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_166), .B(n_512), .Y(n_614) );
AO31x2_ASAP7_75t_L g588 ( .A1(n_167), .A2(n_556), .A3(n_589), .B(n_592), .Y(n_588) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2x1_ASAP7_75t_L g571 ( .A(n_168), .B(n_572), .Y(n_571) );
INVx4_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g172 ( .A(n_169), .B(n_173), .Y(n_172) );
BUFx3_ASAP7_75t_L g176 ( .A(n_169), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g205 ( .A(n_169), .B(n_206), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_169), .B(n_237), .Y(n_236) );
INVx2_ASAP7_75t_SL g267 ( .A(n_169), .Y(n_267) );
AND2x2_ASAP7_75t_L g555 ( .A(n_169), .B(n_556), .Y(n_555) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
AND2x2_ASAP7_75t_L g277 ( .A(n_174), .B(n_278), .Y(n_277) );
AND2x4_ASAP7_75t_L g427 ( .A(n_174), .B(n_304), .Y(n_427) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_191), .Y(n_174) );
OR2x2_ASAP7_75t_L g264 ( .A(n_175), .B(n_265), .Y(n_264) );
BUFx2_ASAP7_75t_L g295 ( .A(n_175), .Y(n_295) );
AND2x2_ASAP7_75t_L g301 ( .A(n_175), .B(n_192), .Y(n_301) );
INVx1_ASAP7_75t_L g319 ( .A(n_175), .Y(n_319) );
INVx2_ASAP7_75t_L g348 ( .A(n_175), .Y(n_348) );
AO31x2_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .A3(n_185), .B(n_187), .Y(n_175) );
INVx2_ASAP7_75t_SL g179 ( .A(n_180), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g584 ( .A(n_180), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_183), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g183 ( .A(n_184), .Y(n_183) );
INVx1_ASAP7_75t_SL g202 ( .A(n_184), .Y(n_202) );
AO31x2_ASAP7_75t_L g240 ( .A1(n_185), .A2(n_220), .A3(n_241), .B(n_244), .Y(n_240) );
AO31x2_ASAP7_75t_L g596 ( .A1(n_185), .A2(n_193), .A3(n_597), .B(n_601), .Y(n_596) );
INVx2_ASAP7_75t_SL g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_SL g275 ( .A(n_186), .Y(n_275) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_188), .B(n_190), .Y(n_187) );
INVx2_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
NOR2xp33_ASAP7_75t_SL g257 ( .A(n_188), .B(n_258), .Y(n_257) );
INVx2_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
INVx2_ASAP7_75t_L g194 ( .A(n_189), .Y(n_194) );
INVx2_ASAP7_75t_L g224 ( .A(n_189), .Y(n_224) );
OAI21xp33_ASAP7_75t_L g518 ( .A1(n_189), .A2(n_517), .B(n_519), .Y(n_518) );
INVx3_ASAP7_75t_L g324 ( .A(n_191), .Y(n_324) );
INVx2_ASAP7_75t_L g329 ( .A(n_191), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_191), .B(n_280), .Y(n_334) );
AND2x2_ASAP7_75t_L g357 ( .A(n_191), .B(n_336), .Y(n_357) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_191), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_191), .B(n_412), .Y(n_411) );
INVx3_ASAP7_75t_L g191 ( .A(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g346 ( .A(n_192), .Y(n_346) );
AND2x2_ASAP7_75t_L g394 ( .A(n_192), .B(n_348), .Y(n_394) );
AO31x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_195), .A3(n_203), .B(n_205), .Y(n_192) );
AOI21x1_ASAP7_75t_L g575 ( .A1(n_193), .A2(n_576), .B(n_586), .Y(n_575) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_194), .B(n_526), .Y(n_525) );
INVx2_ASAP7_75t_L g539 ( .A(n_194), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_194), .B(n_593), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_194), .B(n_602), .Y(n_601) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_198), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g563 ( .A1(n_201), .A2(n_564), .B(n_565), .C(n_566), .Y(n_563) );
AO31x2_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .A3(n_220), .B(n_222), .Y(n_213) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g530 ( .A1(n_204), .A2(n_531), .B(n_534), .Y(n_530) );
INVx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_209), .B(n_225), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_209), .B(n_338), .Y(n_385) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
NAND2x1p5_ASAP7_75t_L g382 ( .A(n_210), .B(n_338), .Y(n_382) );
INVx1_ASAP7_75t_L g483 ( .A(n_210), .Y(n_483) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g433 ( .A(n_211), .B(n_434), .Y(n_433) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
INVx1_ASAP7_75t_L g286 ( .A(n_212), .Y(n_286) );
OR2x2_ASAP7_75t_L g367 ( .A(n_212), .B(n_239), .Y(n_367) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
INVx2_ASAP7_75t_L g309 ( .A(n_213), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_213), .B(n_316), .Y(n_315) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_217), .B(n_581), .Y(n_580) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_220), .A2(n_530), .B(n_538), .Y(n_529) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_224), .B(n_245), .Y(n_244) );
AOI32xp33_ASAP7_75t_L g453 ( .A1(n_225), .A2(n_356), .A3(n_454), .B1(n_456), .B2(n_457), .Y(n_453) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
OR2x2_ASAP7_75t_L g402 ( .A(n_226), .B(n_403), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_227), .B(n_238), .Y(n_226) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_227), .Y(n_248) );
OR2x2_ASAP7_75t_L g284 ( .A(n_227), .B(n_240), .Y(n_284) );
INVx1_ASAP7_75t_L g299 ( .A(n_227), .Y(n_299) );
AND2x2_ASAP7_75t_L g308 ( .A(n_227), .B(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g314 ( .A(n_227), .Y(n_314) );
INVx2_ASAP7_75t_L g339 ( .A(n_227), .Y(n_339) );
AND2x2_ASAP7_75t_L g458 ( .A(n_227), .B(n_250), .Y(n_458) );
OAI21xp33_ASAP7_75t_SL g546 ( .A1(n_231), .A2(n_547), .B(n_548), .Y(n_546) );
INVx1_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_238), .B(n_291), .Y(n_378) );
INVx1_ASAP7_75t_L g238 ( .A(n_239), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g249 ( .A(n_240), .B(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g307 ( .A(n_240), .Y(n_307) );
INVx2_ASAP7_75t_L g316 ( .A(n_240), .Y(n_316) );
AND2x4_ASAP7_75t_L g338 ( .A(n_240), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_240), .Y(n_430) );
AOI22x1_ASAP7_75t_SL g246 ( .A1(n_247), .A2(n_259), .B1(n_277), .B2(n_282), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND4xp25_ASAP7_75t_L g407 ( .A(n_249), .B(n_408), .C(n_409), .D(n_410), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_249), .B(n_308), .Y(n_438) );
INVx4_ASAP7_75t_SL g291 ( .A(n_250), .Y(n_291) );
BUFx2_ASAP7_75t_L g354 ( .A(n_250), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g417 ( .A(n_250), .B(n_299), .Y(n_417) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_255), .B(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g379 ( .A(n_261), .B(n_328), .Y(n_379) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
AND2x4_ASAP7_75t_L g302 ( .A(n_265), .B(n_280), .Y(n_302) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_266), .B(n_281), .Y(n_326) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_267), .A2(n_268), .B(n_276), .Y(n_266) );
OAI21x1_ASAP7_75t_L g321 ( .A1(n_267), .A2(n_268), .B(n_276), .Y(n_321) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_272), .B(n_275), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g293 ( .A(n_278), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g344 ( .A(n_278), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g383 ( .A(n_279), .B(n_301), .Y(n_383) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g426 ( .A(n_281), .B(n_336), .Y(n_426) );
AOI221xp5_ASAP7_75t_L g398 ( .A1(n_282), .A2(n_399), .B1(n_401), .B2(n_404), .C(n_406), .Y(n_398) );
INVx2_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx2_ASAP7_75t_L g292 ( .A(n_284), .Y(n_292) );
OR2x2_ASAP7_75t_L g392 ( .A(n_284), .B(n_331), .Y(n_392) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_293), .Y(n_287) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_288), .A2(n_414), .B1(n_418), .B2(n_421), .Y(n_413) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_292), .Y(n_288) );
AND2x4_ASAP7_75t_L g337 ( .A(n_289), .B(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g449 ( .A(n_289), .B(n_367), .Y(n_449) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x4_ASAP7_75t_L g297 ( .A(n_291), .B(n_298), .Y(n_297) );
AND2x2_ASAP7_75t_L g313 ( .A(n_291), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g372 ( .A(n_291), .B(n_309), .Y(n_372) );
HB1xp67_ASAP7_75t_L g389 ( .A(n_291), .Y(n_389) );
INVx1_ASAP7_75t_L g403 ( .A(n_291), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_291), .B(n_316), .Y(n_446) );
AND2x4_ASAP7_75t_L g353 ( .A(n_292), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g351 ( .A(n_294), .Y(n_351) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_295), .B(n_336), .Y(n_335) );
NAND2x1_ASAP7_75t_L g455 ( .A(n_295), .B(n_357), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_300), .B1(n_303), .B2(n_305), .Y(n_296) );
AND2x2_ASAP7_75t_L g322 ( .A(n_297), .B(n_315), .Y(n_322) );
INVx1_ASAP7_75t_L g363 ( .A(n_297), .Y(n_363) );
AND2x2_ASAP7_75t_L g470 ( .A(n_297), .B(n_331), .Y(n_470) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x4_ASAP7_75t_SL g300 ( .A(n_301), .B(n_302), .Y(n_300) );
AND2x2_ASAP7_75t_L g303 ( .A(n_301), .B(n_304), .Y(n_303) );
INVx2_ASAP7_75t_L g443 ( .A(n_301), .Y(n_443) );
AND2x2_ASAP7_75t_L g460 ( .A(n_301), .B(n_320), .Y(n_460) );
AND2x2_ASAP7_75t_L g476 ( .A(n_301), .B(n_426), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_302), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g399 ( .A(n_302), .B(n_400), .Y(n_399) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_302), .A2(n_392), .B1(n_407), .B2(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g362 ( .A(n_304), .Y(n_362) );
AND2x2_ASAP7_75t_L g393 ( .A(n_304), .B(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_304), .B(n_400), .Y(n_422) );
AND2x2_ASAP7_75t_L g305 ( .A(n_306), .B(n_308), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g428 ( .A(n_308), .B(n_429), .Y(n_428) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_308), .A2(n_332), .B1(n_437), .B2(n_439), .Y(n_436) );
INVx3_ASAP7_75t_L g331 ( .A(n_309), .Y(n_331) );
AND2x2_ASAP7_75t_L g463 ( .A(n_309), .B(n_316), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_327), .Y(n_310) );
AOI32xp33_ASAP7_75t_L g311 ( .A1(n_312), .A2(n_317), .A3(n_320), .B1(n_322), .B2(n_323), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_315), .Y(n_312) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_314), .Y(n_409) );
INVx1_ASAP7_75t_L g434 ( .A(n_314), .Y(n_434) );
INVx3_ASAP7_75t_L g390 ( .A(n_315), .Y(n_390) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OAI221xp5_ASAP7_75t_L g465 ( .A1(n_318), .A2(n_466), .B1(n_467), .B2(n_468), .C(n_469), .Y(n_465) );
BUFx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
OR2x2_ASAP7_75t_L g442 ( .A(n_320), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g478 ( .A(n_320), .B(n_439), .Y(n_478) );
BUFx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g336 ( .A(n_321), .Y(n_336) );
NAND2x1p5_ASAP7_75t_L g350 ( .A(n_323), .B(n_351), .Y(n_350) );
AO22x1_ASAP7_75t_L g380 ( .A1(n_323), .A2(n_381), .B1(n_383), .B2(n_384), .Y(n_380) );
NAND2x1p5_ASAP7_75t_L g484 ( .A(n_323), .B(n_351), .Y(n_484) );
AND2x4_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx2_ASAP7_75t_L g400 ( .A(n_324), .Y(n_400) );
INVx1_ASAP7_75t_L g410 ( .A(n_324), .Y(n_410) );
AND2x2_ASAP7_75t_L g330 ( .A(n_325), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g325 ( .A(n_326), .Y(n_325) );
INVxp67_ASAP7_75t_SL g412 ( .A(n_326), .Y(n_412) );
INVx1_ASAP7_75t_L g452 ( .A(n_326), .Y(n_452) );
A2O1A1Ixp33_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_330), .B(n_332), .C(n_337), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NOR2x1p5_ASAP7_75t_L g439 ( .A(n_329), .B(n_359), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_330), .B(n_389), .Y(n_466) );
AOI31xp33_ASAP7_75t_L g349 ( .A1(n_331), .A2(n_350), .A3(n_352), .B(n_355), .Y(n_349) );
INVx4_ASAP7_75t_L g408 ( .A(n_331), .Y(n_408) );
OR2x2_ASAP7_75t_L g445 ( .A(n_331), .B(n_446), .Y(n_445) );
INVx2_ASAP7_75t_SL g332 ( .A(n_333), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
AND2x4_ASAP7_75t_L g347 ( .A(n_336), .B(n_348), .Y(n_347) );
HB1xp67_ASAP7_75t_L g343 ( .A(n_338), .Y(n_343) );
AND2x2_ASAP7_75t_L g374 ( .A(n_338), .B(n_372), .Y(n_374) );
NOR2xp67_ASAP7_75t_L g340 ( .A(n_341), .B(n_349), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g467 ( .A(n_344), .Y(n_467) );
INVx1_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
AND2x2_ASAP7_75t_L g404 ( .A(n_347), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_358), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
OAI322xp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_363), .A3(n_364), .B1(n_368), .B2(n_371), .C1(n_373), .C2(n_375), .Y(n_361) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
AOI211x1_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_379), .B(n_380), .C(n_386), .Y(n_376) );
INVx1_ASAP7_75t_L g481 ( .A(n_377), .Y(n_481) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g435 ( .A(n_379), .Y(n_435) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
OA21x2_ASAP7_75t_L g386 ( .A1(n_387), .A2(n_391), .B(n_393), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
INVx2_ASAP7_75t_L g456 ( .A(n_390), .Y(n_456) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
NAND2xp33_ASAP7_75t_L g451 ( .A(n_394), .B(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_396), .B(n_464), .Y(n_395) );
NOR3xp33_ASAP7_75t_L g396 ( .A(n_397), .B(n_431), .C(n_447), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_398), .B(n_413), .C(n_423), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_400), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
OAI21xp33_ASAP7_75t_L g459 ( .A1(n_404), .A2(n_460), .B(n_461), .Y(n_459) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_408), .B(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_408), .B(n_458), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_409), .B(n_483), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g418 ( .A(n_410), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
OAI21xp5_ASAP7_75t_L g469 ( .A1(n_420), .A2(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
OAI21xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_427), .B(n_428), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_432), .A2(n_435), .B(n_436), .C(n_440), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_444), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_SL g450 ( .A(n_442), .B(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
HB1xp67_ASAP7_75t_L g468 ( .A(n_446), .Y(n_468) );
OAI211xp5_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_450), .B(n_453), .C(n_459), .Y(n_447) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_458), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g479 ( .A(n_458), .Y(n_479) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g475 ( .A(n_463), .Y(n_475) );
NOR3xp33_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .C(n_480), .Y(n_464) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AOI21xp33_ASAP7_75t_SL g473 ( .A1(n_474), .A2(n_477), .B(n_479), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_475), .B(n_476), .Y(n_474) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
AOI21xp33_ASAP7_75t_R g480 ( .A1(n_481), .A2(n_482), .B(n_484), .Y(n_480) );
INVx4_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
OAI21xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_500), .B(n_828), .Y(n_493) );
CKINVDCx5p33_ASAP7_75t_R g494 ( .A(n_495), .Y(n_494) );
BUFx12f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
AND2x6_ASAP7_75t_SL g496 ( .A(n_497), .B(n_498), .Y(n_496) );
AOI22xp5_ASAP7_75t_L g500 ( .A1(n_501), .A2(n_502), .B1(n_821), .B2(n_827), .Y(n_500) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_727), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_656), .C(n_698), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_506), .B(n_630), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_540), .B1(n_605), .B2(n_616), .Y(n_506) );
INVx3_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_527), .Y(n_508) );
AOI21xp33_ASAP7_75t_L g649 ( .A1(n_509), .A2(n_650), .B(n_652), .Y(n_649) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_509), .A2(n_723), .B(n_724), .Y(n_722) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
INVx2_ASAP7_75t_L g642 ( .A(n_510), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_510), .B(n_521), .Y(n_672) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g613 ( .A(n_514), .Y(n_613) );
OAI21x1_ASAP7_75t_L g514 ( .A1(n_515), .A2(n_516), .B(n_517), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g552 ( .A1(n_515), .A2(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g615 ( .A(n_518), .Y(n_615) );
AOI21xp5_ASAP7_75t_L g576 ( .A1(n_519), .A2(n_577), .B(n_583), .Y(n_576) );
AND2x2_ASAP7_75t_L g712 ( .A(n_520), .B(n_559), .Y(n_712) );
INVx1_ASAP7_75t_L g745 ( .A(n_520), .Y(n_745) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g607 ( .A(n_521), .B(n_560), .Y(n_607) );
AND2x2_ASAP7_75t_L g638 ( .A(n_521), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_L g647 ( .A(n_521), .Y(n_647) );
OR2x2_ASAP7_75t_L g666 ( .A(n_521), .B(n_529), .Y(n_666) );
AND2x2_ASAP7_75t_L g681 ( .A(n_521), .B(n_529), .Y(n_681) );
INVx1_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_528), .B(n_680), .Y(n_723) );
OR2x2_ASAP7_75t_L g811 ( .A(n_528), .B(n_672), .Y(n_811) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx2_ASAP7_75t_L g639 ( .A(n_529), .Y(n_639) );
AND2x2_ASAP7_75t_L g648 ( .A(n_529), .B(n_611), .Y(n_648) );
AND2x2_ASAP7_75t_L g651 ( .A(n_529), .B(n_560), .Y(n_651) );
AND2x2_ASAP7_75t_L g670 ( .A(n_529), .B(n_559), .Y(n_670) );
AND2x4_ASAP7_75t_L g689 ( .A(n_529), .B(n_612), .Y(n_689) );
OAI21xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_557), .B(n_594), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_541), .B(n_684), .Y(n_787) );
CKINVDCx14_ASAP7_75t_R g541 ( .A(n_542), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_543), .B(n_604), .Y(n_603) );
INVx3_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
OR2x2_ASAP7_75t_L g628 ( .A(n_543), .B(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_543), .B(n_621), .Y(n_653) );
AND2x2_ASAP7_75t_L g678 ( .A(n_543), .B(n_596), .Y(n_678) );
AND2x2_ASAP7_75t_L g696 ( .A(n_543), .B(n_626), .Y(n_696) );
INVx1_ASAP7_75t_L g735 ( .A(n_543), .Y(n_735) );
AND2x2_ASAP7_75t_L g737 ( .A(n_543), .B(n_738), .Y(n_737) );
NAND2x1p5_ASAP7_75t_SL g756 ( .A(n_543), .B(n_677), .Y(n_756) );
AND2x4_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
OAI21xp5_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_552), .B(n_555), .Y(n_545) );
NOR2xp33_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
BUFx4f_ASAP7_75t_L g582 ( .A(n_550), .Y(n_582) );
INVx1_ASAP7_75t_L g572 ( .A(n_556), .Y(n_572) );
OAI32xp33_ASAP7_75t_L g640 ( .A1(n_557), .A2(n_632), .A3(n_641), .B1(n_643), .B2(n_645), .Y(n_640) );
OR2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_573), .Y(n_557) );
INVx1_ASAP7_75t_L g680 ( .A(n_558), .Y(n_680) );
AND2x2_ASAP7_75t_L g688 ( .A(n_558), .B(n_689), .Y(n_688) );
BUFx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
AND2x2_ASAP7_75t_L g687 ( .A(n_559), .B(n_611), .Y(n_687) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
BUFx3_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
AND2x2_ASAP7_75t_L g646 ( .A(n_560), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g752 ( .A(n_560), .Y(n_752) );
NAND2x1p5_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI21x1_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .B(n_571), .Y(n_562) );
INVx2_ASAP7_75t_SL g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g622 ( .A(n_573), .Y(n_622) );
OR2x2_ASAP7_75t_L g632 ( .A(n_573), .B(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g754 ( .A(n_573), .Y(n_754) );
OR2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_587), .Y(n_573) );
AND2x2_ASAP7_75t_L g655 ( .A(n_574), .B(n_588), .Y(n_655) );
INVx2_ASAP7_75t_L g677 ( .A(n_574), .Y(n_677) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_574), .B(n_596), .Y(n_697) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g604 ( .A(n_575), .Y(n_604) );
OAI21xp5_ASAP7_75t_L g577 ( .A1(n_578), .A2(n_580), .B(n_582), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_587), .B(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g686 ( .A(n_587), .Y(n_686) );
INVx2_ASAP7_75t_SL g587 ( .A(n_588), .Y(n_587) );
BUFx2_ASAP7_75t_L g626 ( .A(n_588), .Y(n_626) );
OR2x2_ASAP7_75t_L g692 ( .A(n_588), .B(n_596), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_588), .B(n_596), .Y(n_725) );
INVx2_ASAP7_75t_L g673 ( .A(n_594), .Y(n_673) );
OR2x2_ASAP7_75t_L g594 ( .A(n_595), .B(n_603), .Y(n_594) );
OR2x2_ASAP7_75t_L g660 ( .A(n_595), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g738 ( .A(n_595), .Y(n_738) );
INVx1_ASAP7_75t_L g621 ( .A(n_596), .Y(n_621) );
INVx1_ASAP7_75t_L g629 ( .A(n_596), .Y(n_629) );
INVx1_ASAP7_75t_L g644 ( .A(n_596), .Y(n_644) );
OR2x2_ASAP7_75t_L g748 ( .A(n_603), .B(n_725), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_604), .B(n_620), .Y(n_661) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_604), .Y(n_663) );
OR2x2_ASAP7_75t_L g762 ( .A(n_604), .B(n_686), .Y(n_762) );
INVxp67_ASAP7_75t_L g786 ( .A(n_604), .Y(n_786) );
INVx2_ASAP7_75t_SL g605 ( .A(n_606), .Y(n_605) );
NAND2x1_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_607), .B(n_648), .Y(n_715) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AND2x2_ASAP7_75t_L g664 ( .A(n_609), .B(n_665), .Y(n_664) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx1_ASAP7_75t_L g777 ( .A(n_610), .Y(n_777) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND2x2_ASAP7_75t_L g806 ( .A(n_611), .B(n_639), .Y(n_806) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
AND2x2_ASAP7_75t_L g732 ( .A(n_612), .B(n_639), .Y(n_732) );
AOI21x1_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_614), .B(n_615), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_617), .B(n_623), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_619), .B(n_622), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_619), .B(n_655), .Y(n_769) );
AND2x4_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx2_ASAP7_75t_L g633 ( .A(n_620), .Y(n_633) );
AND2x2_ASAP7_75t_L g683 ( .A(n_620), .B(n_684), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_620), .B(n_677), .Y(n_726) );
OR2x2_ASAP7_75t_L g798 ( .A(n_620), .B(n_685), .Y(n_798) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g718 ( .A(n_624), .B(n_719), .Y(n_718) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
INVx2_ASAP7_75t_L g709 ( .A(n_625), .Y(n_709) );
INVx2_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g699 ( .A(n_628), .B(n_700), .Y(n_699) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_628), .Y(n_710) );
OR2x2_ASAP7_75t_L g761 ( .A(n_628), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g816 ( .A(n_628), .Y(n_816) );
AOI211xp5_ASAP7_75t_L g630 ( .A1(n_631), .A2(n_634), .B(n_640), .C(n_649), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g705 ( .A(n_633), .B(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g753 ( .A(n_633), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g778 ( .A(n_633), .B(n_655), .Y(n_778) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_636), .B(n_681), .Y(n_703) );
NAND2x1p5_ASAP7_75t_L g720 ( .A(n_636), .B(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g788 ( .A(n_636), .B(n_789), .Y(n_788) );
INVx3_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
BUFx2_ASAP7_75t_L g731 ( .A(n_637), .Y(n_731) );
AND2x2_ASAP7_75t_L g759 ( .A(n_638), .B(n_687), .Y(n_759) );
INVx2_ASAP7_75t_L g782 ( .A(n_638), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_638), .B(n_680), .Y(n_814) );
AND2x4_ASAP7_75t_SL g768 ( .A(n_641), .B(n_646), .Y(n_768) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g721 ( .A(n_642), .B(n_647), .Y(n_721) );
OR2x2_ASAP7_75t_L g773 ( .A(n_642), .B(n_666), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_643), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g809 ( .A(n_643), .B(n_655), .Y(n_809) );
BUFx3_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g757 ( .A(n_644), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_648), .Y(n_645) );
INVx1_ASAP7_75t_L g740 ( .A(n_646), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g805 ( .A(n_646), .B(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g790 ( .A(n_647), .Y(n_790) );
BUFx2_ASAP7_75t_L g658 ( .A(n_648), .Y(n_658) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AND2x2_ASAP7_75t_L g776 ( .A(n_651), .B(n_777), .Y(n_776) );
OR2x2_ASAP7_75t_L g652 ( .A(n_653), .B(n_654), .Y(n_652) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g700 ( .A(n_655), .Y(n_700) );
HB1xp67_ASAP7_75t_L g717 ( .A(n_655), .Y(n_717) );
NAND3xp33_ASAP7_75t_SL g656 ( .A(n_657), .B(n_667), .C(n_682), .Y(n_656) );
AOI22xp33_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_664), .Y(n_657) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI222xp33_ASAP7_75t_L g770 ( .A1(n_664), .A2(n_690), .B1(n_771), .B2(n_774), .C1(n_776), .C2(n_778), .Y(n_770) );
AND2x2_ASAP7_75t_L g802 ( .A(n_665), .B(n_751), .Y(n_802) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g750 ( .A(n_666), .B(n_751), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_673), .B1(n_674), .B2(n_679), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_SL g746 ( .A(n_670), .Y(n_746) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_678), .Y(n_674) );
AND2x2_ASAP7_75t_L g733 ( .A(n_675), .B(n_734), .Y(n_733) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
OR2x2_ASAP7_75t_L g691 ( .A(n_676), .B(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g685 ( .A(n_677), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g800 ( .A(n_678), .Y(n_800) );
AND2x2_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_681), .B(n_777), .Y(n_796) );
INVx1_ASAP7_75t_L g813 ( .A(n_681), .Y(n_813) );
AOI222xp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_687), .B1(n_688), .B2(n_690), .C1(n_693), .C2(n_694), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
HB1xp67_ASAP7_75t_L g693 ( .A(n_689), .Y(n_693) );
AND2x2_ASAP7_75t_L g711 ( .A(n_689), .B(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g742 ( .A(n_689), .Y(n_742) );
INVx2_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx2_ASAP7_75t_L g706 ( .A(n_692), .Y(n_706) );
OR2x2_ASAP7_75t_L g775 ( .A(n_692), .B(n_756), .Y(n_775) );
INVx2_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B(n_704), .C(n_713), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
OAI21xp33_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_707), .B(n_711), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g791 ( .A1(n_705), .A2(n_743), .B1(n_792), .B2(n_795), .C(n_797), .Y(n_791) );
AND2x4_ASAP7_75t_L g734 ( .A(n_706), .B(n_735), .Y(n_734) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .Y(n_708) );
INVx1_ASAP7_75t_L g765 ( .A(n_712), .Y(n_765) );
AOI211x1_ASAP7_75t_L g713 ( .A1(n_714), .A2(n_716), .B(n_718), .C(n_722), .Y(n_713) );
INVxp67_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g783 ( .A(n_721), .Y(n_783) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_724), .B(n_772), .C(n_773), .Y(n_771) );
OR2x2_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
INVx1_ASAP7_75t_L g807 ( .A(n_725), .Y(n_807) );
NOR2x1_ASAP7_75t_L g727 ( .A(n_728), .B(n_779), .Y(n_727) );
NAND4xp25_ASAP7_75t_L g728 ( .A(n_729), .B(n_736), .C(n_758), .D(n_770), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g729 ( .A(n_730), .B(n_733), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
AND2x2_ASAP7_75t_L g789 ( .A(n_732), .B(n_790), .Y(n_789) );
AOI221x1_ASAP7_75t_L g758 ( .A1(n_734), .A2(n_759), .B1(n_760), .B2(n_763), .C(n_766), .Y(n_758) );
AND2x2_ASAP7_75t_L g784 ( .A(n_734), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g794 ( .A(n_735), .Y(n_794) );
AOI221xp5_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_739), .B1(n_743), .B2(n_747), .C(n_749), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_741), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_741), .B(n_765), .Y(n_764) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
OR2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_746), .A2(n_750), .B1(n_753), .B2(n_755), .Y(n_749) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g766 ( .A1(n_750), .A2(n_767), .B(n_769), .Y(n_766) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx1_ASAP7_75t_L g772 ( .A(n_752), .Y(n_772) );
OR2x2_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVxp67_ASAP7_75t_L g793 ( .A(n_762), .Y(n_793) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
OAI22xp33_ASAP7_75t_L g812 ( .A1(n_775), .A2(n_813), .B1(n_814), .B2(n_815), .Y(n_812) );
NAND3xp33_ASAP7_75t_L g779 ( .A(n_780), .B(n_791), .C(n_803), .Y(n_779) );
AOI22xp5_ASAP7_75t_L g780 ( .A1(n_781), .A2(n_784), .B1(n_787), .B2(n_788), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
INVxp67_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
OR2x2_ASAP7_75t_L g799 ( .A(n_786), .B(n_800), .Y(n_799) );
NAND2x1_ASAP7_75t_L g815 ( .A(n_786), .B(n_816), .Y(n_815) );
AND2x2_ASAP7_75t_L g792 ( .A(n_793), .B(n_794), .Y(n_792) );
INVx2_ASAP7_75t_SL g795 ( .A(n_796), .Y(n_795) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B(n_801), .Y(n_797) );
INVx1_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
AOI221xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_807), .B1(n_808), .B2(n_810), .C(n_812), .Y(n_803) );
INVx1_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
INVx3_ASAP7_75t_R g810 ( .A(n_811), .Y(n_810) );
INVx4_ASAP7_75t_L g820 ( .A(n_817), .Y(n_820) );
BUFx12f_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
CKINVDCx5p33_ASAP7_75t_R g818 ( .A(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g834 ( .A(n_819), .B(n_835), .Y(n_834) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_821), .Y(n_827) );
INVx1_ASAP7_75t_L g822 ( .A(n_823), .Y(n_822) );
INVx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g830 ( .A(n_831), .Y(n_830) );
BUFx10_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
NOR2xp33_ASAP7_75t_R g836 ( .A(n_837), .B(n_838), .Y(n_836) );
INVx2_ASAP7_75t_L g838 ( .A(n_839), .Y(n_838) );
endmodule