module fake_jpeg_15999_n_287 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_102;
wire n_99;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_273;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_176;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_100;
wire n_258;
wire n_282;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx4_ASAP7_75t_SL g43 ( 
.A(n_39),
.Y(n_43)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_43),
.Y(n_109)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_45),
.Y(n_95)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_47),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_6),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_48),
.B(n_51),
.Y(n_113)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_15),
.Y(n_49)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_49),
.Y(n_93)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_50),
.B(n_58),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_19),
.B(n_6),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_0),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_57),
.Y(n_88)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_31),
.C(n_41),
.Y(n_54)
);

A2O1A1Ixp33_ASAP7_75t_L g126 ( 
.A1(n_54),
.A2(n_37),
.B(n_35),
.C(n_33),
.Y(n_126)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_21),
.B(n_9),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_34),
.B(n_0),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_59),
.B(n_70),
.Y(n_98)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_60),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_21),
.B(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_65),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_63),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_22),
.B(n_4),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g107 ( 
.A(n_64),
.B(n_29),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g65 ( 
.A(n_17),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_39),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_66),
.B(n_76),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_67),
.Y(n_115)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_17),
.B(n_0),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_32),
.Y(n_71)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_73),
.Y(n_99)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_18),
.Y(n_74)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_74),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_24),
.Y(n_75)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_75),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_22),
.B(n_4),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_20),
.B(n_11),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_77),
.B(n_27),
.Y(n_114)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_31),
.Y(n_78)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_78),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_31),
.B1(n_40),
.B2(n_25),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_80),
.A2(n_84),
.B1(n_97),
.B2(n_127),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_36),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_81),
.B(n_110),
.Y(n_150)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx3_ASAP7_75t_SL g133 ( 
.A(n_82),
.Y(n_133)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_56),
.A2(n_41),
.B1(n_40),
.B2(n_25),
.Y(n_84)
);

BUFx10_ASAP7_75t_L g90 ( 
.A(n_55),
.Y(n_90)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_90),
.Y(n_139)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_53),
.A2(n_37),
.B1(n_35),
.B2(n_23),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_68),
.A2(n_46),
.B1(n_42),
.B2(n_47),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_104),
.A2(n_106),
.B1(n_49),
.B2(n_45),
.Y(n_137)
);

OA22x2_ASAP7_75t_L g105 ( 
.A1(n_54),
.A2(n_23),
.B1(n_33),
.B2(n_28),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_13),
.B1(n_14),
.B2(n_12),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_63),
.A2(n_27),
.B1(n_36),
.B2(n_29),
.Y(n_106)
);

NAND2xp33_ASAP7_75t_SL g167 ( 
.A(n_107),
.B(n_126),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_49),
.B(n_20),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_69),
.B(n_33),
.C(n_28),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_114),
.B(n_117),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_50),
.B(n_30),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_78),
.Y(n_118)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_118),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_30),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_120),
.B(n_123),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_43),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_30),
.Y(n_123)
);

OAI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_67),
.A2(n_37),
.B1(n_30),
.B2(n_2),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_129),
.B(n_146),
.Y(n_172)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g191 ( 
.A(n_132),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_13),
.Y(n_134)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_136),
.A2(n_137),
.B1(n_149),
.B2(n_169),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_79),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_140),
.B(n_144),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_98),
.B(n_0),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_153),
.Y(n_183)
);

AO22x2_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_69),
.B1(n_71),
.B2(n_1),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_166),
.B(n_122),
.Y(n_171)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_100),
.Y(n_143)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_91),
.B(n_3),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_145),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_124),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_147),
.B(n_152),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_103),
.A2(n_108),
.B1(n_109),
.B2(n_125),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_12),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_2),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_94),
.Y(n_154)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_105),
.B(n_2),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_164),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_85),
.B(n_71),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_156),
.B(n_157),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_124),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_94),
.Y(n_158)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_158),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_95),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_90),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_160),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_161),
.A2(n_163),
.B1(n_133),
.B2(n_138),
.Y(n_199)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_88),
.A2(n_106),
.B(n_121),
.C(n_93),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_141),
.Y(n_185)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_97),
.B(n_104),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_101),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_111),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_109),
.A2(n_99),
.B(n_119),
.Y(n_166)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_82),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_168),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_101),
.A2(n_122),
.B1(n_99),
.B2(n_119),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_171),
.A2(n_174),
.B(n_175),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_159),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_173),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_115),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_95),
.Y(n_175)
);

HAxp5_ASAP7_75t_SL g179 ( 
.A(n_142),
.B(n_83),
.CON(n_179),
.SN(n_179)
);

AND2x2_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_180),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_116),
.C(n_89),
.Y(n_180)
);

AOI32xp33_ASAP7_75t_L g181 ( 
.A1(n_167),
.A2(n_83),
.A3(n_89),
.B1(n_96),
.B2(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_186),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_153),
.A2(n_155),
.B1(n_136),
.B2(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_182),
.A2(n_165),
.B1(n_145),
.B2(n_151),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_185),
.B(n_199),
.Y(n_219)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_162),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_200),
.Y(n_216)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_154),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_150),
.B(n_140),
.Y(n_200)
);

AO22x1_ASAP7_75t_L g203 ( 
.A1(n_179),
.A2(n_138),
.B1(n_163),
.B2(n_133),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_204),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_199),
.A2(n_161),
.B1(n_164),
.B2(n_131),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_210),
.B1(n_193),
.B2(n_189),
.Y(n_229)
);

OR2x2_ASAP7_75t_L g206 ( 
.A(n_184),
.B(n_161),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_206),
.A2(n_215),
.B(n_224),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_207),
.B(n_209),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_200),
.B(n_148),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_171),
.A2(n_143),
.B1(n_130),
.B2(n_157),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_190),
.B(n_128),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_213),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_135),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_183),
.B(n_184),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_177),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_220),
.Y(n_238)
);

OA22x2_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_175),
.B1(n_170),
.B2(n_186),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_197),
.B1(n_168),
.B2(n_135),
.Y(n_230)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_221),
.B(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_198),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_130),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_223),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_180),
.B(n_158),
.Y(n_224)
);

AOI221xp5_ASAP7_75t_L g225 ( 
.A1(n_205),
.A2(n_187),
.B1(n_185),
.B2(n_174),
.C(n_175),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_225),
.A2(n_227),
.B(n_219),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_219),
.B(n_172),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_232),
.C(n_227),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_211),
.A2(n_193),
.B1(n_189),
.B2(n_195),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_229),
.B(n_235),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_214),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_201),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_239),
.B(n_241),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_218),
.A2(n_198),
.B1(n_178),
.B2(n_197),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_139),
.B1(n_178),
.B2(n_188),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_246),
.C(n_228),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_211),
.B1(n_219),
.B2(n_224),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_235),
.B1(n_241),
.B2(n_206),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_226),
.C(n_231),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_247),
.A2(n_250),
.B(n_240),
.Y(n_261)
);

OAI322xp33_ASAP7_75t_L g248 ( 
.A1(n_237),
.A2(n_206),
.A3(n_216),
.B1(n_223),
.B2(n_209),
.C1(n_215),
.C2(n_224),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_L g267 ( 
.A(n_248),
.B(n_192),
.C(n_220),
.Y(n_267)
);

OA21x2_ASAP7_75t_L g249 ( 
.A1(n_242),
.A2(n_210),
.B(n_218),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g258 ( 
.A1(n_249),
.A2(n_202),
.B(n_225),
.Y(n_258)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_243),
.B(n_211),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_230),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_254),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_236),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_233),
.A2(n_216),
.B1(n_203),
.B2(n_202),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_238),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_257),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g257 ( 
.A(n_236),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_258),
.A2(n_261),
.B(n_265),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_246),
.B(n_228),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_234),
.C(n_240),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_250),
.A2(n_238),
.B(n_234),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_267),
.B(n_252),
.Y(n_269)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_266),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_268),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_271),
.B(n_273),
.Y(n_277)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_249),
.B(n_251),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_272),
.A2(n_255),
.B1(n_247),
.B2(n_260),
.Y(n_276)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_276),
.B(n_278),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_270),
.A2(n_176),
.B(n_259),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_221),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_208),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_279),
.B(n_277),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_284),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_283),
.B(n_173),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_286),
.Y(n_287)
);


endmodule