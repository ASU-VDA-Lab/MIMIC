module real_aes_7596_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_769;
wire n_434;
wire n_505;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_756;
wire n_598;
wire n_735;
wire n_713;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_212;
wire n_575;
wire n_210;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g500 ( .A1(n_0), .A2(n_182), .B(n_501), .C(n_504), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_1), .B(n_495), .Y(n_506) );
NAND3xp33_ASAP7_75t_SL g112 ( .A(n_2), .B(n_113), .C(n_114), .Y(n_112) );
INVx1_ASAP7_75t_L g452 ( .A(n_2), .Y(n_452) );
INVx1_ASAP7_75t_L g231 ( .A(n_3), .Y(n_231) );
OAI211xp5_ASAP7_75t_L g123 ( .A1(n_4), .A2(n_124), .B(n_454), .C(n_457), .Y(n_123) );
OAI211xp5_ASAP7_75t_L g454 ( .A1(n_4), .A2(n_126), .B(n_445), .C(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_5), .B(n_170), .Y(n_529) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_6), .A2(n_479), .B(n_549), .Y(n_548) );
OAI22xp5_ASAP7_75t_SL g441 ( .A1(n_7), .A2(n_11), .B1(n_442), .B2(n_443), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g442 ( .A(n_7), .Y(n_442) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_8), .A2(n_187), .B(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g181 ( .A1(n_9), .A2(n_38), .B1(n_143), .B2(n_155), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_10), .B(n_187), .Y(n_220) );
CKINVDCx20_ASAP7_75t_R g443 ( .A(n_11), .Y(n_443) );
AOI22xp5_ASAP7_75t_L g462 ( .A1(n_11), .A2(n_128), .B1(n_443), .B2(n_444), .Y(n_462) );
AND2x6_ASAP7_75t_L g158 ( .A(n_12), .B(n_159), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g570 ( .A1(n_13), .A2(n_158), .B(n_482), .C(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g110 ( .A(n_14), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g453 ( .A(n_14), .B(n_39), .Y(n_453) );
INVx1_ASAP7_75t_L g139 ( .A(n_15), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_16), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g225 ( .A(n_17), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_18), .B(n_170), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_19), .B(n_185), .Y(n_203) );
AO32x2_ASAP7_75t_L g179 ( .A1(n_20), .A2(n_180), .A3(n_184), .B1(n_186), .B2(n_187), .Y(n_179) );
OAI22xp5_ASAP7_75t_L g764 ( .A1(n_21), .A2(n_57), .B1(n_765), .B2(n_766), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g766 ( .A(n_21), .Y(n_766) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_22), .B(n_143), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_23), .B(n_185), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g183 ( .A1(n_24), .A2(n_55), .B1(n_143), .B2(n_155), .Y(n_183) );
AOI22xp33_ASAP7_75t_SL g196 ( .A1(n_25), .A2(n_83), .B1(n_143), .B2(n_147), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_26), .B(n_143), .Y(n_173) );
A2O1A1Ixp33_ASAP7_75t_L g481 ( .A1(n_27), .A2(n_186), .B(n_482), .C(n_484), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g560 ( .A1(n_28), .A2(n_186), .B(n_482), .C(n_561), .Y(n_560) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_29), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_30), .B(n_135), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_31), .A2(n_479), .B(n_497), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_32), .B(n_135), .Y(n_177) );
INVx2_ASAP7_75t_L g145 ( .A(n_33), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g512 ( .A1(n_34), .A2(n_513), .B(n_514), .C(n_518), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_35), .B(n_143), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_36), .B(n_135), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_37), .B(n_150), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_39), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_40), .B(n_478), .Y(n_477) );
CKINVDCx20_ASAP7_75t_R g575 ( .A(n_41), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_42), .B(n_170), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_43), .B(n_479), .Y(n_559) );
A2O1A1Ixp33_ASAP7_75t_L g539 ( .A1(n_44), .A2(n_513), .B(n_518), .C(n_540), .Y(n_539) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_45), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_45), .Y(n_762) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_46), .B(n_143), .Y(n_213) );
INVx1_ASAP7_75t_L g502 ( .A(n_47), .Y(n_502) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_48), .A2(n_93), .B1(n_155), .B2(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g541 ( .A(n_49), .Y(n_541) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_50), .B(n_143), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_51), .B(n_143), .Y(n_227) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_52), .B(n_448), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_53), .B(n_479), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_54), .B(n_218), .Y(n_217) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_56), .A2(n_61), .B1(n_143), .B2(n_147), .Y(n_207) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_57), .Y(n_765) );
CKINVDCx20_ASAP7_75t_R g491 ( .A(n_58), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g142 ( .A(n_59), .B(n_143), .Y(n_142) );
NAND2xp5_ASAP7_75t_SL g244 ( .A(n_60), .B(n_143), .Y(n_244) );
INVx1_ASAP7_75t_L g159 ( .A(n_62), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_63), .B(n_479), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_64), .B(n_495), .Y(n_554) );
A2O1A1Ixp33_ASAP7_75t_L g551 ( .A1(n_65), .A2(n_218), .B(n_228), .C(n_552), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_66), .B(n_143), .Y(n_232) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_68), .Y(n_122) );
NAND2xp5_ASAP7_75t_SL g516 ( .A(n_69), .B(n_170), .Y(n_516) );
AO32x2_ASAP7_75t_L g192 ( .A1(n_70), .A2(n_186), .A3(n_187), .B1(n_193), .B2(n_197), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_71), .B(n_171), .Y(n_572) );
INVx1_ASAP7_75t_L g243 ( .A(n_72), .Y(n_243) );
INVx1_ASAP7_75t_L g168 ( .A(n_73), .Y(n_168) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_74), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_75), .B(n_486), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g104 ( .A1(n_76), .A2(n_105), .B1(n_117), .B2(n_774), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_77), .B(n_127), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_77), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g526 ( .A1(n_78), .A2(n_482), .B(n_518), .C(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_79), .B(n_147), .Y(n_169) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_80), .Y(n_550) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_82), .B(n_488), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_84), .B(n_155), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g520 ( .A(n_85), .Y(n_520) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_86), .B(n_147), .Y(n_174) );
AOI222xp33_ASAP7_75t_L g459 ( .A1(n_87), .A2(n_460), .B1(n_760), .B2(n_761), .C1(n_767), .C2(n_769), .Y(n_459) );
INVx2_ASAP7_75t_L g136 ( .A(n_88), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g533 ( .A(n_89), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g573 ( .A(n_90), .B(n_157), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_91), .B(n_147), .Y(n_214) );
INVx2_ASAP7_75t_L g113 ( .A(n_92), .Y(n_113) );
OR2x2_ASAP7_75t_L g449 ( .A(n_92), .B(n_450), .Y(n_449) );
OR2x2_ASAP7_75t_L g465 ( .A(n_92), .B(n_451), .Y(n_465) );
AOI22xp33_ASAP7_75t_L g206 ( .A1(n_94), .A2(n_103), .B1(n_147), .B2(n_148), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_95), .B(n_479), .Y(n_511) );
INVx1_ASAP7_75t_L g515 ( .A(n_96), .Y(n_515) );
INVxp67_ASAP7_75t_L g553 ( .A(n_97), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_98), .B(n_147), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g115 ( .A(n_99), .B(n_116), .Y(n_115) );
INVx1_ASAP7_75t_L g528 ( .A(n_100), .Y(n_528) );
INVx1_ASAP7_75t_L g568 ( .A(n_101), .Y(n_568) );
AND2x2_ASAP7_75t_L g543 ( .A(n_102), .B(n_135), .Y(n_543) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g774 ( .A(n_107), .Y(n_774) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g759 ( .A(n_113), .B(n_451), .Y(n_759) );
NOR2x2_ASAP7_75t_L g771 ( .A(n_113), .B(n_450), .Y(n_771) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
OA21x2_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_123), .B(n_458), .Y(n_117) );
BUFx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
CKINVDCx20_ASAP7_75t_R g119 ( .A(n_120), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g773 ( .A(n_121), .Y(n_773) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
NOR3xp33_ASAP7_75t_L g125 ( .A(n_126), .B(n_445), .C(n_448), .Y(n_125) );
INVx1_ASAP7_75t_L g447 ( .A(n_127), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_440), .B1(n_441), .B2(n_444), .Y(n_127) );
INVx1_ASAP7_75t_L g444 ( .A(n_128), .Y(n_444) );
OR2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_362), .Y(n_128) );
NAND5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_281), .C(n_296), .D(n_322), .E(n_344), .Y(n_129) );
NOR2xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_261), .Y(n_130) );
OAI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_198), .B1(n_234), .B2(n_250), .C(n_251), .Y(n_131) );
NOR2xp33_ASAP7_75t_SL g132 ( .A(n_133), .B(n_188), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_133), .B(n_311), .Y(n_310) );
INVx1_ASAP7_75t_SL g438 ( .A(n_133), .Y(n_438) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_161), .Y(n_133) );
INVx1_ASAP7_75t_L g278 ( .A(n_134), .Y(n_278) );
AND2x2_ASAP7_75t_L g280 ( .A(n_134), .B(n_179), .Y(n_280) );
AND2x2_ASAP7_75t_L g290 ( .A(n_134), .B(n_178), .Y(n_290) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_134), .Y(n_308) );
INVx1_ASAP7_75t_L g318 ( .A(n_134), .Y(n_318) );
OR2x2_ASAP7_75t_L g356 ( .A(n_134), .B(n_255), .Y(n_356) );
INVx2_ASAP7_75t_L g406 ( .A(n_134), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_134), .B(n_254), .Y(n_423) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_140), .B(n_160), .Y(n_134) );
OA21x2_ASAP7_75t_L g164 ( .A1(n_135), .A2(n_165), .B(n_177), .Y(n_164) );
INVx2_ASAP7_75t_L g197 ( .A(n_135), .Y(n_197) );
INVx1_ASAP7_75t_L g492 ( .A(n_135), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_135), .A2(n_511), .B(n_512), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_135), .A2(n_538), .B(n_539), .Y(n_537) );
AND2x2_ASAP7_75t_SL g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_L g185 ( .A(n_136), .B(n_137), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_152), .B(n_158), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_146), .B(n_149), .Y(n_141) );
INVx3_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
HB1xp67_ASAP7_75t_L g530 ( .A(n_143), .Y(n_530) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g155 ( .A(n_144), .Y(n_155) );
BUFx3_ASAP7_75t_L g195 ( .A(n_144), .Y(n_195) );
AND2x6_ASAP7_75t_L g482 ( .A(n_144), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g148 ( .A(n_145), .Y(n_148) );
INVx1_ASAP7_75t_L g219 ( .A(n_145), .Y(n_219) );
INVx2_ASAP7_75t_L g226 ( .A(n_147), .Y(n_226) );
INVx3_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_151), .Y(n_157) );
INVx3_ASAP7_75t_L g171 ( .A(n_151), .Y(n_171) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_151), .Y(n_176) );
AND2x2_ASAP7_75t_L g480 ( .A(n_151), .B(n_219), .Y(n_480) );
INVx1_ASAP7_75t_L g483 ( .A(n_151), .Y(n_483) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_154), .B(n_156), .Y(n_152) );
O2A1O1Ixp5_ASAP7_75t_L g242 ( .A1(n_156), .A2(n_230), .B(n_243), .C(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g180 ( .A1(n_157), .A2(n_181), .B1(n_182), .B2(n_183), .Y(n_180) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_157), .A2(n_171), .B1(n_194), .B2(n_196), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g205 ( .A1(n_157), .A2(n_182), .B1(n_206), .B2(n_207), .Y(n_205) );
INVx4_ASAP7_75t_L g503 ( .A(n_157), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g165 ( .A1(n_158), .A2(n_166), .B(n_172), .Y(n_165) );
BUFx3_ASAP7_75t_L g186 ( .A(n_158), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_212), .B(n_215), .Y(n_211) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_158), .A2(n_224), .B(n_229), .Y(n_223) );
AND2x4_ASAP7_75t_L g479 ( .A(n_158), .B(n_480), .Y(n_479) );
INVx4_ASAP7_75t_SL g505 ( .A(n_158), .Y(n_505) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_158), .B(n_480), .Y(n_569) );
NOR2xp67_ASAP7_75t_L g161 ( .A(n_162), .B(n_178), .Y(n_161) );
INVx1_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_163), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_163), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_163), .B(n_278), .Y(n_338) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_164), .Y(n_190) );
INVx2_ASAP7_75t_L g255 ( .A(n_164), .Y(n_255) );
OR2x2_ASAP7_75t_L g317 ( .A(n_164), .B(n_318), .Y(n_317) );
O2A1O1Ixp5_ASAP7_75t_SL g166 ( .A1(n_167), .A2(n_168), .B(n_169), .C(n_170), .Y(n_166) );
INVx2_ASAP7_75t_L g182 ( .A(n_170), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_170), .A2(n_213), .B(n_214), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_170), .A2(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_170), .B(n_553), .Y(n_552) );
INVx5_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
INVx1_ASAP7_75t_L g228 ( .A(n_175), .Y(n_228) );
INVx4_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g486 ( .A(n_176), .Y(n_486) );
AND2x2_ASAP7_75t_L g256 ( .A(n_178), .B(n_192), .Y(n_256) );
AND2x2_ASAP7_75t_L g273 ( .A(n_178), .B(n_253), .Y(n_273) );
INVx2_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
AND2x2_ASAP7_75t_L g191 ( .A(n_179), .B(n_192), .Y(n_191) );
BUFx2_ASAP7_75t_L g276 ( .A(n_179), .Y(n_276) );
AND2x2_ASAP7_75t_L g405 ( .A(n_179), .B(n_406), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_182), .A2(n_216), .B(n_217), .Y(n_215) );
O2A1O1Ixp33_ASAP7_75t_L g229 ( .A1(n_182), .A2(n_230), .B(n_231), .C(n_232), .Y(n_229) );
INVx2_ASAP7_75t_L g222 ( .A(n_184), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_184), .B(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
BUFx6f_ASAP7_75t_L g187 ( .A(n_185), .Y(n_187) );
NAND3xp33_ASAP7_75t_L g204 ( .A(n_186), .B(n_205), .C(n_208), .Y(n_204) );
OAI21xp5_ASAP7_75t_L g238 ( .A1(n_186), .A2(n_239), .B(n_242), .Y(n_238) );
INVx4_ASAP7_75t_L g208 ( .A(n_187), .Y(n_208) );
OA21x2_ASAP7_75t_L g210 ( .A1(n_187), .A2(n_211), .B(n_220), .Y(n_210) );
HB1xp67_ASAP7_75t_L g547 ( .A(n_187), .Y(n_547) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_187), .A2(n_559), .B(n_560), .Y(n_558) );
INVx1_ASAP7_75t_L g250 ( .A(n_188), .Y(n_250) );
AND2x2_ASAP7_75t_L g188 ( .A(n_189), .B(n_191), .Y(n_188) );
AND2x2_ASAP7_75t_L g368 ( .A(n_189), .B(n_256), .Y(n_368) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
AND2x2_ASAP7_75t_L g369 ( .A(n_190), .B(n_280), .Y(n_369) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_191), .A2(n_337), .B(n_339), .C(n_341), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_191), .B(n_337), .Y(n_346) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_191), .A2(n_267), .B1(n_410), .B2(n_411), .C(n_413), .Y(n_409) );
INVx1_ASAP7_75t_L g253 ( .A(n_192), .Y(n_253) );
INVx1_ASAP7_75t_L g289 ( .A(n_192), .Y(n_289) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_192), .Y(n_298) );
INVx2_ASAP7_75t_L g504 ( .A(n_195), .Y(n_504) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_195), .Y(n_517) );
INVx1_ASAP7_75t_L g489 ( .A(n_197), .Y(n_489) );
INVx1_ASAP7_75t_SL g198 ( .A(n_199), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
AND2x2_ASAP7_75t_L g315 ( .A(n_200), .B(n_260), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_200), .B(n_335), .Y(n_334) );
INVx2_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
NOR2xp33_ASAP7_75t_L g283 ( .A(n_201), .B(n_284), .Y(n_283) );
OR2x2_ASAP7_75t_L g407 ( .A(n_201), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g439 ( .A(n_201), .Y(n_439) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx3_ASAP7_75t_L g269 ( .A(n_202), .Y(n_269) );
AND2x2_ASAP7_75t_L g295 ( .A(n_202), .B(n_249), .Y(n_295) );
NOR2x1_ASAP7_75t_L g304 ( .A(n_202), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g311 ( .A(n_202), .B(n_312), .Y(n_311) );
AND2x4_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
INVx1_ASAP7_75t_L g247 ( .A(n_203), .Y(n_247) );
AO21x1_ASAP7_75t_L g246 ( .A1(n_205), .A2(n_208), .B(n_247), .Y(n_246) );
INVx3_ASAP7_75t_L g495 ( .A(n_208), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g519 ( .A(n_208), .B(n_520), .Y(n_519) );
AO21x2_ASAP7_75t_L g524 ( .A1(n_208), .A2(n_525), .B(n_532), .Y(n_524) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_208), .B(n_533), .Y(n_532) );
AO21x2_ASAP7_75t_L g566 ( .A1(n_208), .A2(n_567), .B(n_574), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_209), .B(n_351), .Y(n_386) );
INVx1_ASAP7_75t_SL g390 ( .A(n_209), .Y(n_390) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_221), .Y(n_209) );
INVx3_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
AND2x2_ASAP7_75t_L g260 ( .A(n_210), .B(n_237), .Y(n_260) );
AND2x2_ASAP7_75t_L g282 ( .A(n_210), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g327 ( .A(n_210), .B(n_321), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_210), .B(n_259), .Y(n_408) );
INVx2_ASAP7_75t_L g230 ( .A(n_218), .Y(n_230) );
INVx1_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g248 ( .A(n_221), .B(n_249), .Y(n_248) );
INVx2_ASAP7_75t_L g259 ( .A(n_221), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_221), .B(n_237), .Y(n_284) );
AND2x2_ASAP7_75t_L g320 ( .A(n_221), .B(n_321), .Y(n_320) );
OA21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_223), .B(n_233), .Y(n_221) );
OA21x2_ASAP7_75t_L g237 ( .A1(n_222), .A2(n_238), .B(n_245), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .C(n_228), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_226), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_226), .A2(n_572), .B(n_573), .Y(n_571) );
O2A1O1Ixp33_ASAP7_75t_L g527 ( .A1(n_228), .A2(n_528), .B(n_529), .C(n_530), .Y(n_527) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_230), .A2(n_485), .B(n_487), .Y(n_484) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_236), .B(n_248), .Y(n_235) );
INVx1_ASAP7_75t_L g300 ( .A(n_236), .Y(n_300) );
AND2x2_ASAP7_75t_L g342 ( .A(n_236), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g348 ( .A(n_236), .B(n_263), .Y(n_348) );
AOI21xp5_ASAP7_75t_SL g422 ( .A1(n_236), .A2(n_254), .B(n_277), .Y(n_422) );
AND2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_246), .Y(n_236) );
OR2x2_ASAP7_75t_L g265 ( .A(n_237), .B(n_246), .Y(n_265) );
AND2x2_ASAP7_75t_L g312 ( .A(n_237), .B(n_249), .Y(n_312) );
INVx2_ASAP7_75t_L g321 ( .A(n_237), .Y(n_321) );
INVx1_ASAP7_75t_L g427 ( .A(n_237), .Y(n_427) );
AND2x2_ASAP7_75t_L g351 ( .A(n_246), .B(n_321), .Y(n_351) );
INVx1_ASAP7_75t_L g376 ( .A(n_246), .Y(n_376) );
AND2x2_ASAP7_75t_L g285 ( .A(n_248), .B(n_269), .Y(n_285) );
AND2x2_ASAP7_75t_L g297 ( .A(n_248), .B(n_298), .Y(n_297) );
INVx2_ASAP7_75t_SL g415 ( .A(n_248), .Y(n_415) );
INVx2_ASAP7_75t_L g305 ( .A(n_249), .Y(n_305) );
AND2x2_ASAP7_75t_L g343 ( .A(n_249), .B(n_259), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_249), .B(n_427), .Y(n_426) );
OAI21xp33_ASAP7_75t_L g251 ( .A1(n_252), .A2(n_256), .B(n_257), .Y(n_251) );
AND2x2_ASAP7_75t_L g358 ( .A(n_252), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g412 ( .A(n_252), .Y(n_412) );
AND2x2_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
INVx1_ASAP7_75t_L g332 ( .A(n_253), .Y(n_332) );
BUFx2_ASAP7_75t_L g431 ( .A(n_253), .Y(n_431) );
BUFx2_ASAP7_75t_L g302 ( .A(n_254), .Y(n_302) );
AND2x2_ASAP7_75t_L g404 ( .A(n_254), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g387 ( .A(n_255), .Y(n_387) );
AND2x4_ASAP7_75t_L g314 ( .A(n_256), .B(n_277), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g350 ( .A(n_256), .B(n_338), .Y(n_350) );
AOI32xp33_ASAP7_75t_L g274 ( .A1(n_257), .A2(n_275), .A3(n_277), .B1(n_279), .B2(n_280), .Y(n_274) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
INVx3_ASAP7_75t_L g263 ( .A(n_258), .Y(n_263) );
OR2x2_ASAP7_75t_L g399 ( .A(n_258), .B(n_355), .Y(n_399) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g268 ( .A(n_259), .B(n_269), .Y(n_268) );
AND2x2_ASAP7_75t_L g375 ( .A(n_259), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g267 ( .A(n_260), .B(n_268), .Y(n_267) );
AND2x2_ASAP7_75t_L g279 ( .A(n_260), .B(n_269), .Y(n_279) );
INVx1_ASAP7_75t_L g400 ( .A(n_260), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_260), .B(n_375), .Y(n_433) );
A2O1A1Ixp33_ASAP7_75t_L g261 ( .A1(n_262), .A2(n_266), .B(n_270), .C(n_274), .Y(n_261) );
OAI322xp33_ASAP7_75t_L g370 ( .A1(n_262), .A2(n_307), .A3(n_371), .B1(n_373), .B2(n_377), .C1(n_378), .C2(n_382), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_264), .Y(n_262) );
INVxp67_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
INVx1_ASAP7_75t_SL g264 ( .A(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g389 ( .A(n_265), .B(n_390), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_265), .B(n_305), .Y(n_436) );
INVxp67_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx1_ASAP7_75t_L g328 ( .A(n_268), .Y(n_328) );
OR2x2_ASAP7_75t_L g414 ( .A(n_269), .B(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_272), .B(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g323 ( .A(n_273), .B(n_302), .Y(n_323) );
AND2x2_ASAP7_75t_L g394 ( .A(n_273), .B(n_307), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_273), .B(n_381), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g281 ( .A1(n_275), .A2(n_282), .B1(n_285), .B2(n_286), .C(n_291), .Y(n_281) );
OR2x2_ASAP7_75t_L g292 ( .A(n_275), .B(n_288), .Y(n_292) );
AND2x2_ASAP7_75t_L g380 ( .A(n_275), .B(n_381), .Y(n_380) );
AOI32xp33_ASAP7_75t_L g419 ( .A1(n_275), .A2(n_305), .A3(n_420), .B1(n_421), .B2(n_424), .Y(n_419) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
NAND3xp33_ASAP7_75t_L g353 ( .A(n_276), .B(n_312), .C(n_335), .Y(n_353) );
AND2x2_ASAP7_75t_L g379 ( .A(n_276), .B(n_372), .Y(n_379) );
INVxp67_ASAP7_75t_L g359 ( .A(n_277), .Y(n_359) );
BUFx3_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_SL g388 ( .A(n_280), .B(n_332), .Y(n_388) );
INVx2_ASAP7_75t_L g398 ( .A(n_280), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_280), .B(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g367 ( .A(n_283), .Y(n_367) );
OR2x2_ASAP7_75t_L g293 ( .A(n_284), .B(n_294), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_286), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_290), .Y(n_286) );
INVx1_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_289), .Y(n_372) );
AND2x2_ASAP7_75t_L g331 ( .A(n_290), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g377 ( .A(n_290), .Y(n_377) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_290), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AOI21xp33_ASAP7_75t_SL g316 ( .A1(n_292), .A2(n_317), .B(n_319), .Y(n_316) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g410 ( .A(n_295), .B(n_320), .Y(n_410) );
AOI211xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_299), .B(n_309), .C(n_316), .Y(n_296) );
AND2x2_ASAP7_75t_L g340 ( .A(n_298), .B(n_308), .Y(n_340) );
INVx2_ASAP7_75t_L g355 ( .A(n_298), .Y(n_355) );
OR2x2_ASAP7_75t_L g393 ( .A(n_298), .B(n_356), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_298), .B(n_436), .Y(n_435) );
AOI211xp5_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_301), .B(n_303), .C(n_306), .Y(n_299) );
INVxp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_302), .B(n_340), .Y(n_339) );
OAI211xp5_ASAP7_75t_L g421 ( .A1(n_303), .A2(n_398), .B(n_422), .C(n_423), .Y(n_421) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
NAND2x1p5_ASAP7_75t_L g319 ( .A(n_304), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g361 ( .A(n_305), .B(n_351), .Y(n_361) );
INVx1_ASAP7_75t_L g366 ( .A(n_305), .Y(n_366) );
INVx1_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_SL g309 ( .A(n_310), .B(n_313), .Y(n_309) );
INVxp33_ASAP7_75t_L g417 ( .A(n_311), .Y(n_417) );
AND2x2_ASAP7_75t_L g396 ( .A(n_312), .B(n_375), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g378 ( .A1(n_317), .A2(n_379), .B(n_380), .Y(n_378) );
OAI322xp33_ASAP7_75t_L g397 ( .A1(n_319), .A2(n_398), .A3(n_399), .B1(n_400), .B2(n_401), .C1(n_403), .C2(n_407), .Y(n_397) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_323), .A2(n_324), .B1(n_329), .B2(n_333), .C(n_336), .Y(n_322) );
INVx2_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
AND2x2_ASAP7_75t_L g374 ( .A(n_327), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g418 ( .A(n_331), .Y(n_418) );
INVxp67_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_334), .B(n_354), .Y(n_420) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g383 ( .A(n_343), .B(n_351), .Y(n_383) );
AOI221xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_347), .B1(n_349), .B2(n_351), .C(n_352), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI221xp5_ASAP7_75t_L g363 ( .A1(n_347), .A2(n_364), .B1(n_368), .B2(n_369), .C(n_370), .Y(n_363) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
INVxp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_351), .B(n_366), .Y(n_365) );
OAI22xp5_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_354), .B1(n_357), .B2(n_360), .Y(n_352) );
OR2x2_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx2_ASAP7_75t_SL g381 ( .A(n_356), .Y(n_381) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
NAND5xp2_ASAP7_75t_L g362 ( .A(n_363), .B(n_384), .C(n_409), .D(n_419), .E(n_429), .Y(n_362) );
NAND2xp5_ASAP7_75t_SL g364 ( .A(n_365), .B(n_367), .Y(n_364) );
NOR4xp25_ASAP7_75t_L g437 ( .A(n_366), .B(n_372), .C(n_438), .D(n_439), .Y(n_437) );
AOI221xp5_ASAP7_75t_L g429 ( .A1(n_369), .A2(n_430), .B1(n_432), .B2(n_434), .C(n_437), .Y(n_429) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g428 ( .A(n_375), .Y(n_428) );
OAI322xp33_ASAP7_75t_L g385 ( .A1(n_379), .A2(n_386), .A3(n_387), .B1(n_388), .B2(n_389), .C1(n_391), .C2(n_395), .Y(n_385) );
INVx1_ASAP7_75t_SL g382 ( .A(n_383), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g384 ( .A(n_385), .B(n_397), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g391 ( .A(n_392), .B(n_394), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g430 ( .A(n_405), .B(n_431), .Y(n_430) );
OAI22xp33_ASAP7_75t_L g413 ( .A1(n_414), .A2(n_416), .B1(n_417), .B2(n_418), .Y(n_413) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
NOR2xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_447), .Y(n_445) );
INVx1_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g456 ( .A(n_449), .Y(n_456) );
INVx2_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_453), .Y(n_451) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g458 ( .A(n_457), .B(n_459), .C(n_772), .Y(n_458) );
OAI22x1_ASAP7_75t_SL g460 ( .A1(n_461), .A2(n_463), .B1(n_466), .B2(n_757), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OAI22xp5_ASAP7_75t_SL g767 ( .A1(n_462), .A2(n_467), .B1(n_757), .B2(n_768), .Y(n_767) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx2_ASAP7_75t_L g768 ( .A(n_464), .Y(n_768) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
AND2x2_ASAP7_75t_SL g467 ( .A(n_468), .B(n_712), .Y(n_467) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_647), .Y(n_468) );
NAND4xp25_ASAP7_75t_SL g469 ( .A(n_470), .B(n_592), .C(n_616), .D(n_639), .Y(n_469) );
AOI221xp5_ASAP7_75t_L g470 ( .A1(n_471), .A2(n_534), .B1(n_564), .B2(n_576), .C(n_579), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_473), .B(n_507), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_473), .A2(n_493), .B1(n_535), .B2(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_473), .B(n_508), .Y(n_650) );
AND2x2_ASAP7_75t_L g669 ( .A(n_473), .B(n_670), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_473), .B(n_653), .Y(n_739) );
AND2x4_ASAP7_75t_L g473 ( .A(n_474), .B(n_493), .Y(n_473) );
AND2x2_ASAP7_75t_L g607 ( .A(n_474), .B(n_508), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_474), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g630 ( .A(n_474), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g635 ( .A(n_474), .B(n_494), .Y(n_635) );
INVx2_ASAP7_75t_L g667 ( .A(n_474), .Y(n_667) );
HB1xp67_ASAP7_75t_L g711 ( .A(n_474), .Y(n_711) );
AND2x2_ASAP7_75t_L g728 ( .A(n_474), .B(n_605), .Y(n_728) );
INVx5_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AND2x2_ASAP7_75t_L g646 ( .A(n_475), .B(n_605), .Y(n_646) );
AND2x4_ASAP7_75t_L g660 ( .A(n_475), .B(n_493), .Y(n_660) );
HB1xp67_ASAP7_75t_L g664 ( .A(n_475), .Y(n_664) );
AND2x2_ASAP7_75t_L g684 ( .A(n_475), .B(n_599), .Y(n_684) );
AND2x2_ASAP7_75t_L g734 ( .A(n_475), .B(n_509), .Y(n_734) );
AND2x2_ASAP7_75t_L g744 ( .A(n_475), .B(n_494), .Y(n_744) );
OR2x6_ASAP7_75t_L g475 ( .A(n_476), .B(n_490), .Y(n_475) );
AOI21xp5_ASAP7_75t_SL g476 ( .A1(n_477), .A2(n_481), .B(n_489), .Y(n_476) );
BUFx2_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVx5_ASAP7_75t_L g499 ( .A(n_482), .Y(n_499) );
INVx2_ASAP7_75t_L g488 ( .A(n_486), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_488), .A2(n_515), .B(n_516), .C(n_517), .Y(n_514) );
O2A1O1Ixp33_ASAP7_75t_L g540 ( .A1(n_488), .A2(n_517), .B(n_541), .C(n_542), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x2_ASAP7_75t_L g600 ( .A(n_493), .B(n_508), .Y(n_600) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_493), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_493), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g690 ( .A(n_493), .Y(n_690) );
INVx2_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AND2x2_ASAP7_75t_L g578 ( .A(n_494), .B(n_523), .Y(n_578) );
AND2x2_ASAP7_75t_L g605 ( .A(n_494), .B(n_524), .Y(n_605) );
OA21x2_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_496), .B(n_506), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g497 ( .A1(n_498), .A2(n_499), .B(n_500), .C(n_505), .Y(n_497) );
INVx2_ASAP7_75t_L g513 ( .A(n_499), .Y(n_513) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_499), .A2(n_505), .B(n_550), .C(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g518 ( .A(n_505), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_507), .B(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_521), .Y(n_507) );
OR2x2_ASAP7_75t_L g631 ( .A(n_508), .B(n_522), .Y(n_631) );
AND2x2_ASAP7_75t_L g668 ( .A(n_508), .B(n_578), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_508), .B(n_599), .Y(n_679) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_508), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_508), .B(n_635), .Y(n_752) );
INVx5_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g577 ( .A(n_509), .Y(n_577) );
AND2x2_ASAP7_75t_L g586 ( .A(n_509), .B(n_522), .Y(n_586) );
AND2x2_ASAP7_75t_L g702 ( .A(n_509), .B(n_597), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_509), .B(n_635), .Y(n_724) );
OR2x6_ASAP7_75t_L g509 ( .A(n_510), .B(n_519), .Y(n_509) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_522), .Y(n_670) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
HB1xp67_ASAP7_75t_L g622 ( .A(n_523), .Y(n_622) );
INVx2_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g599 ( .A(n_524), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_544), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_535), .B(n_612), .Y(n_731) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g564 ( .A(n_536), .B(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g583 ( .A(n_536), .B(n_584), .Y(n_583) );
INVx5_ASAP7_75t_SL g591 ( .A(n_536), .Y(n_591) );
OR2x2_ASAP7_75t_L g614 ( .A(n_536), .B(n_584), .Y(n_614) );
OR2x2_ASAP7_75t_L g624 ( .A(n_536), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g687 ( .A(n_536), .B(n_546), .Y(n_687) );
AND2x2_ASAP7_75t_SL g725 ( .A(n_536), .B(n_545), .Y(n_725) );
NOR4xp25_ASAP7_75t_L g746 ( .A(n_536), .B(n_667), .C(n_747), .D(n_748), .Y(n_746) );
AND2x2_ASAP7_75t_L g756 ( .A(n_536), .B(n_588), .Y(n_756) );
OR2x6_ASAP7_75t_L g536 ( .A(n_537), .B(n_543), .Y(n_536) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
AND2x2_ASAP7_75t_L g581 ( .A(n_545), .B(n_577), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_545), .B(n_583), .Y(n_750) );
AND2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_555), .Y(n_545) );
OR2x2_ASAP7_75t_L g590 ( .A(n_546), .B(n_591), .Y(n_590) );
INVx3_ASAP7_75t_L g597 ( .A(n_546), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_546), .B(n_566), .Y(n_609) );
INVxp67_ASAP7_75t_L g612 ( .A(n_546), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_546), .B(n_584), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_546), .B(n_556), .Y(n_678) );
AND2x2_ASAP7_75t_L g693 ( .A(n_546), .B(n_588), .Y(n_693) );
OR2x2_ASAP7_75t_L g722 ( .A(n_546), .B(n_556), .Y(n_722) );
OA21x2_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B(n_554), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_555), .B(n_627), .Y(n_626) );
NOR2xp33_ASAP7_75t_L g730 ( .A(n_555), .B(n_591), .Y(n_730) );
OR2x2_ASAP7_75t_L g751 ( .A(n_555), .B(n_628), .Y(n_751) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g565 ( .A(n_556), .B(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g588 ( .A(n_556), .B(n_584), .Y(n_588) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_556), .B(n_566), .Y(n_603) );
AND2x2_ASAP7_75t_L g673 ( .A(n_556), .B(n_597), .Y(n_673) );
AND2x2_ASAP7_75t_L g707 ( .A(n_556), .B(n_591), .Y(n_707) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_557), .B(n_591), .Y(n_610) );
AND2x2_ASAP7_75t_L g638 ( .A(n_557), .B(n_566), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_564), .B(n_646), .Y(n_645) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_565), .A2(n_653), .B1(n_689), .B2(n_706), .C(n_708), .Y(n_705) );
INVx5_ASAP7_75t_SL g584 ( .A(n_566), .Y(n_584) );
OAI21xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_569), .B(n_570), .Y(n_567) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
OAI33xp33_ASAP7_75t_L g604 ( .A1(n_577), .A2(n_605), .A3(n_606), .B1(n_608), .B2(n_611), .B3(n_615), .Y(n_604) );
OR2x2_ASAP7_75t_L g620 ( .A(n_577), .B(n_621), .Y(n_620) );
AOI322xp5_ASAP7_75t_L g729 ( .A1(n_577), .A2(n_646), .A3(n_653), .B1(n_730), .B2(n_731), .C1(n_732), .C2(n_735), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_577), .B(n_605), .Y(n_747) );
A2O1A1Ixp33_ASAP7_75t_SL g753 ( .A1(n_577), .A2(n_605), .B(n_754), .C(n_756), .Y(n_753) );
AOI221xp5_ASAP7_75t_L g592 ( .A1(n_578), .A2(n_593), .B1(n_598), .B2(n_601), .C(n_604), .Y(n_592) );
INVx1_ASAP7_75t_L g685 ( .A(n_578), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_578), .B(n_734), .Y(n_733) );
OAI22xp33_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B1(n_585), .B2(n_587), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g662 ( .A(n_583), .B(n_597), .Y(n_662) );
AND2x2_ASAP7_75t_L g720 ( .A(n_583), .B(n_721), .Y(n_720) );
OR2x2_ASAP7_75t_L g628 ( .A(n_584), .B(n_591), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_584), .B(n_597), .Y(n_656) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_586), .B(n_659), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_586), .B(n_664), .Y(n_718) );
OAI321xp33_ASAP7_75t_L g737 ( .A1(n_586), .A2(n_659), .A3(n_738), .B1(n_739), .B2(n_740), .C(n_741), .Y(n_737) );
INVx1_ASAP7_75t_L g704 ( .A(n_587), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_588), .B(n_589), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_588), .B(n_595), .Y(n_594) );
AND2x2_ASAP7_75t_L g643 ( .A(n_588), .B(n_591), .Y(n_643) );
AOI321xp33_ASAP7_75t_L g701 ( .A1(n_588), .A2(n_605), .A3(n_702), .B1(n_703), .B2(n_704), .C(n_705), .Y(n_701) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g618 ( .A(n_590), .B(n_603), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_591), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_591), .B(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_591), .B(n_677), .Y(n_714) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AND2x4_ASAP7_75t_L g637 ( .A(n_595), .B(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g602 ( .A(n_596), .B(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g710 ( .A(n_597), .Y(n_710) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_600), .B(n_653), .Y(n_652) );
INVx2_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g633 ( .A(n_605), .Y(n_633) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NOR2xp33_ASAP7_75t_L g691 ( .A(n_607), .B(n_642), .Y(n_691) );
OR2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
OR2x2_ASAP7_75t_L g655 ( .A(n_610), .B(n_656), .Y(n_655) );
INVx1_ASAP7_75t_SL g700 ( .A(n_610), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_611), .A2(n_658), .B1(n_661), .B2(n_663), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
INVx1_ASAP7_75t_SL g613 ( .A(n_614), .Y(n_613) );
OR2x2_ASAP7_75t_L g755 ( .A(n_614), .B(n_678), .Y(n_755) );
AOI221xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_619), .B1(n_623), .B2(n_629), .C(n_632), .Y(n_616) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
INVx2_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
BUFx2_ASAP7_75t_L g653 ( .A(n_622), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
INVx1_ASAP7_75t_SL g699 ( .A(n_625), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_627), .B(n_677), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g694 ( .A1(n_627), .A2(n_695), .B(n_697), .Y(n_694) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
OR2x2_ASAP7_75t_L g740 ( .A(n_628), .B(n_722), .Y(n_740) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx2_ASAP7_75t_SL g642 ( .A(n_631), .Y(n_642) );
AOI21xp33_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_634), .B(n_636), .Y(n_632) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx2_ASAP7_75t_SL g636 ( .A(n_637), .Y(n_636) );
AND2x2_ASAP7_75t_L g686 ( .A(n_638), .B(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_L g748 ( .A(n_638), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_644), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_642), .B(n_660), .Y(n_696) );
INVxp67_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g717 ( .A(n_646), .Y(n_717) );
NAND5xp2_ASAP7_75t_L g647 ( .A(n_648), .B(n_665), .C(n_674), .D(n_694), .E(n_701), .Y(n_647) );
O2A1O1Ixp33_ASAP7_75t_L g648 ( .A1(n_649), .A2(n_651), .B(n_654), .C(n_657), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx1_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g689 ( .A(n_653), .Y(n_689) );
CKINVDCx16_ASAP7_75t_R g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_661), .B(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g703 ( .A(n_663), .Y(n_703) );
OAI21xp5_ASAP7_75t_SL g665 ( .A1(n_666), .A2(n_669), .B(n_671), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_666), .A2(n_720), .B1(n_723), .B2(n_725), .C(n_726), .Y(n_719) );
AND2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AOI321xp33_ASAP7_75t_L g674 ( .A1(n_667), .A2(n_675), .A3(n_679), .B1(n_680), .B2(n_686), .C(n_688), .Y(n_674) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g745 ( .A(n_679), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g680 ( .A(n_681), .B(n_685), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g697 ( .A(n_682), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
NOR2xp67_ASAP7_75t_SL g709 ( .A(n_683), .B(n_690), .Y(n_709) );
AOI321xp33_ASAP7_75t_SL g741 ( .A1(n_686), .A2(n_742), .A3(n_743), .B1(n_744), .B2(n_745), .C(n_746), .Y(n_741) );
O2A1O1Ixp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_691), .C(n_692), .Y(n_688) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_699), .B(n_707), .Y(n_736) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
NAND3xp33_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_711), .Y(n_708) );
NOR3xp33_ASAP7_75t_L g712 ( .A(n_713), .B(n_737), .C(n_749), .Y(n_712) );
OAI211xp5_ASAP7_75t_SL g713 ( .A1(n_714), .A2(n_715), .B(n_719), .C(n_729), .Y(n_713) );
INVxp67_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g716 ( .A(n_717), .B(n_718), .Y(n_716) );
OAI221xp5_ASAP7_75t_L g749 ( .A1(n_718), .A2(n_750), .B1(n_751), .B2(n_752), .C(n_753), .Y(n_749) );
INVx1_ASAP7_75t_L g738 ( .A(n_720), .Y(n_738) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g742 ( .A(n_740), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
CKINVDCx14_ASAP7_75t_R g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_SL g769 ( .A(n_770), .Y(n_769) );
INVx3_ASAP7_75t_SL g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_SL g772 ( .A(n_773), .Y(n_772) );
endmodule