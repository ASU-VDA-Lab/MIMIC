module fake_jpeg_23687_n_53 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_53);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_53;

wire n_33;
wire n_45;
wire n_27;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx8_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_20),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_19),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_29),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_30),
.B(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_27),
.B(n_1),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_1),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_31),
.Y(n_34)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_30),
.A2(n_27),
.B1(n_24),
.B2(n_28),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g40 ( 
.A1(n_35),
.A2(n_36),
.B1(n_38),
.B2(n_39),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_31),
.Y(n_36)
);

NAND2xp33_ASAP7_75t_SL g37 ( 
.A(n_32),
.B(n_25),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g43 ( 
.A(n_37),
.B(n_2),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_24),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_25),
.B1(n_14),
.B2(n_4),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_41),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_43),
.A2(n_33),
.B(n_3),
.Y(n_44)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

NOR3xp33_ASAP7_75t_SL g46 ( 
.A(n_43),
.B(n_40),
.C(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_48),
.B(n_7),
.C(n_8),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_47),
.C(n_11),
.Y(n_50)
);

AOI322xp5_ASAP7_75t_L g51 ( 
.A1(n_50),
.A2(n_9),
.A3(n_12),
.B1(n_13),
.B2(n_15),
.C1(n_16),
.C2(n_17),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_51),
.Y(n_52)
);

OAI21x1_ASAP7_75t_L g53 ( 
.A1(n_52),
.A2(n_22),
.B(n_23),
.Y(n_53)
);


endmodule