module fake_jpeg_20771_n_238 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_238);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_238;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx2_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_10),
.Y(n_31)
);

BUFx24_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_4),
.B(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_8),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_44),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_39),
.B(n_31),
.Y(n_82)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_1),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_45),
.B(n_48),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_26),
.Y(n_48)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g51 ( 
.A(n_33),
.B(n_1),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_52),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_55),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_18),
.B(n_15),
.Y(n_55)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_58),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_40),
.A2(n_27),
.B1(n_30),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_31),
.B1(n_20),
.B2(n_21),
.Y(n_103)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_70),
.Y(n_92)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_46),
.Y(n_62)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_62),
.Y(n_105)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_63),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_39),
.B(n_36),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_66),
.Y(n_91)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g97 ( 
.A(n_65),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_36),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_48),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_27),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_73),
.B(n_82),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_78),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_54),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_38),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_83),
.Y(n_114)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_47),
.A2(n_30),
.B1(n_27),
.B2(n_23),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_84),
.A2(n_19),
.B1(n_29),
.B2(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g85 ( 
.A(n_43),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_85),
.B(n_89),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_51),
.B(n_17),
.Y(n_89)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_94),
.A2(n_96),
.B1(n_68),
.B2(n_3),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_73),
.B(n_56),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_95),
.B(n_99),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_57),
.A2(n_35),
.B1(n_23),
.B2(n_24),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_56),
.B(n_89),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_102),
.Y(n_139)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_77),
.A2(n_24),
.B1(n_21),
.B2(n_20),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_104),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_118),
.B1(n_90),
.B2(n_75),
.Y(n_124)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_110),
.Y(n_138)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_86),
.Y(n_111)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_61),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_80),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_7),
.Y(n_137)
);

FAx1_ASAP7_75t_L g116 ( 
.A(n_59),
.B(n_25),
.CI(n_28),
.CON(n_116),
.SN(n_116)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_60),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_25),
.B1(n_3),
.B2(n_4),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_119),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_117),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_121),
.B(n_134),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_113),
.B(n_88),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_127),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_124),
.A2(n_126),
.B1(n_135),
.B2(n_136),
.Y(n_161)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_72),
.Y(n_127)
);

AOI32xp33_ASAP7_75t_L g128 ( 
.A1(n_116),
.A2(n_72),
.A3(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

OA21x2_ASAP7_75t_L g130 ( 
.A1(n_94),
.A2(n_71),
.B(n_68),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_130),
.A2(n_98),
.B(n_106),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_108),
.B(n_16),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_2),
.B1(n_5),
.B2(n_7),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_109),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_9),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_140),
.Y(n_150)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_105),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_105),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_92),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_142),
.B(n_143),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_91),
.B(n_11),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_144),
.Y(n_166)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_147),
.A2(n_155),
.B(n_156),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_139),
.B(n_95),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_148),
.B(n_145),
.Y(n_171)
);

OR2x2_ASAP7_75t_L g153 ( 
.A(n_139),
.B(n_99),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_158),
.Y(n_170)
);

XOR2x2_ASAP7_75t_L g155 ( 
.A(n_126),
.B(n_107),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_126),
.A2(n_115),
.B(n_102),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_134),
.B(n_97),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_162),
.B(n_167),
.Y(n_179)
);

AOI22x1_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_102),
.B1(n_118),
.B2(n_97),
.Y(n_163)
);

OAI21x1_ASAP7_75t_SL g186 ( 
.A1(n_163),
.A2(n_168),
.B(n_125),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_100),
.C(n_110),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_164),
.B(n_129),
.C(n_124),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_10),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_100),
.B(n_13),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_120),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_173),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_166),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_172),
.Y(n_189)
);

OA21x2_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_130),
.B(n_135),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_175),
.B(n_182),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_132),
.C(n_119),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_164),
.C(n_153),
.Y(n_193)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_157),
.Y(n_180)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_180),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_121),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_141),
.Y(n_182)
);

NOR3xp33_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_144),
.C(n_130),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_186),
.B(n_155),
.C(n_148),
.D(n_154),
.Y(n_188)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_157),
.Y(n_184)
);

AO221x1_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_185),
.B1(n_187),
.B2(n_150),
.C(n_138),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_169),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_188),
.A2(n_198),
.B1(n_170),
.B2(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_173),
.A2(n_151),
.B1(n_154),
.B2(n_161),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_192),
.A2(n_184),
.B1(n_178),
.B2(n_138),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_193),
.B(n_140),
.C(n_14),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_174),
.A2(n_156),
.B(n_147),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_194),
.A2(n_197),
.B1(n_177),
.B2(n_170),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_174),
.A2(n_153),
.B(n_165),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_161),
.B1(n_149),
.B2(n_120),
.Y(n_198)
);

AOI322xp5_ASAP7_75t_L g199 ( 
.A1(n_186),
.A2(n_159),
.A3(n_146),
.B1(n_167),
.B2(n_158),
.C1(n_152),
.C2(n_150),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_199),
.B(n_150),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g204 ( 
.A(n_200),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_171),
.B(n_146),
.C(n_152),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_140),
.C(n_122),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_187),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_202),
.B(n_203),
.Y(n_215)
);

AO22x2_ASAP7_75t_SL g203 ( 
.A1(n_188),
.A2(n_175),
.B1(n_177),
.B2(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_179),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_205),
.B(n_209),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_206),
.A2(n_210),
.B(n_211),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_207),
.B(n_208),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_190),
.B(n_178),
.Y(n_209)
);

OA21x2_ASAP7_75t_SL g219 ( 
.A1(n_212),
.A2(n_195),
.B(n_192),
.Y(n_219)
);

NOR3xp33_ASAP7_75t_L g214 ( 
.A(n_203),
.B(n_194),
.C(n_197),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_220),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_208),
.A2(n_191),
.B(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_217),
.B(n_219),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_204),
.A2(n_191),
.B(n_190),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_216),
.B(n_196),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_193),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_211),
.C(n_196),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_213),
.B(n_200),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_215),
.B(n_201),
.CI(n_206),
.CON(n_225),
.SN(n_225)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_11),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_227),
.B(n_221),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_226),
.A2(n_213),
.B1(n_203),
.B2(n_199),
.Y(n_228)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_228),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_223),
.B(n_212),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_230),
.B(n_231),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_227),
.Y(n_235)
);

AOI321xp33_ASAP7_75t_L g237 ( 
.A1(n_235),
.A2(n_236),
.A3(n_234),
.B1(n_233),
.B2(n_222),
.C(n_225),
.Y(n_237)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_232),
.B(n_229),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_237),
.B(n_225),
.Y(n_238)
);


endmodule