module fake_jpeg_30493_n_83 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_83);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_83;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_8),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_9),
.B(n_4),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_21),
.Y(n_29)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_22),
.B(n_24),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

AOI21xp33_ASAP7_75t_SL g24 ( 
.A1(n_16),
.A2(n_0),
.B(n_1),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_2),
.Y(n_26)
);

AOI21xp5_ASAP7_75t_L g27 ( 
.A1(n_15),
.A2(n_1),
.B(n_5),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_27),
.B(n_28),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_8),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_12),
.B1(n_17),
.B2(n_18),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_31),
.A2(n_18),
.B1(n_17),
.B2(n_22),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_11),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_37),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_35),
.B(n_13),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_21),
.A2(n_12),
.B1(n_20),
.B2(n_14),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_39),
.A2(n_46),
.B1(n_30),
.B2(n_36),
.Y(n_54)
);

OAI32xp33_ASAP7_75t_L g40 ( 
.A1(n_30),
.A2(n_17),
.A3(n_20),
.B1(n_23),
.B2(n_25),
.Y(n_40)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_6),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_33),
.B(n_7),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_45),
.A2(n_48),
.B(n_49),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_47),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_34),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_7),
.Y(n_49)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_40),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_43),
.C(n_41),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_57),
.B(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_42),
.C(n_46),
.Y(n_58)
);

INVxp33_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_59),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_61),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_47),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_57),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_63),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_50),
.A2(n_54),
.B1(n_51),
.B2(n_56),
.Y(n_64)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_65),
.B(n_63),
.C(n_51),
.Y(n_68)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_68),
.A2(n_65),
.B(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_74),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_69),
.A2(n_50),
.B1(n_60),
.B2(n_52),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_70),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_72),
.B(n_59),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_66),
.Y(n_78)
);

OAI31xp33_ASAP7_75t_L g80 ( 
.A1(n_78),
.A2(n_79),
.A3(n_75),
.B(n_77),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_76),
.A2(n_66),
.B(n_52),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_80),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_52),
.C(n_55),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_55),
.Y(n_83)
);


endmodule