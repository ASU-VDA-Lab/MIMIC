module fake_aes_7922_n_13 (n_1, n_2, n_0, n_13);
input n_1;
input n_2;
input n_0;
output n_13;
wire n_11;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
NOR2x1p5_ASAP7_75t_L g3 ( .A(n_0), .B(n_1), .Y(n_3) );
INVx1_ASAP7_75t_L g4 ( .A(n_0), .Y(n_4) );
OAI221xp5_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_3), .B1(n_1), .B2(n_2), .C(n_0), .Y(n_5) );
AND2x4_ASAP7_75t_L g6 ( .A(n_3), .B(n_2), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_6), .Y(n_7) );
OAI221xp5_ASAP7_75t_SL g8 ( .A1(n_5), .A2(n_4), .B1(n_1), .B2(n_2), .C(n_0), .Y(n_8) );
INVxp67_ASAP7_75t_SL g9 ( .A(n_7), .Y(n_9) );
AOI32xp33_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_6), .A3(n_7), .B1(n_8), .B2(n_2), .Y(n_10) );
AOI211xp5_ASAP7_75t_L g11 ( .A1(n_9), .A2(n_8), .B(n_6), .C(n_1), .Y(n_11) );
AND2x2_ASAP7_75t_L g12 ( .A(n_11), .B(n_10), .Y(n_12) );
HB1xp67_ASAP7_75t_L g13 ( .A(n_12), .Y(n_13) );
endmodule