module fake_jpeg_6207_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx1_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_6),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_2),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_16),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_13),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

BUFx24_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_22),
.B(n_17),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_19),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_17),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g26 ( 
.A1(n_25),
.A2(n_15),
.B1(n_12),
.B2(n_16),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_27),
.B(n_28),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_25),
.A2(n_15),
.B1(n_12),
.B2(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_21),
.A2(n_16),
.B1(n_19),
.B2(n_10),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_31),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_24),
.A2(n_19),
.B1(n_10),
.B2(n_8),
.Y(n_31)
);

CKINVDCx10_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_19),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_20),
.Y(n_38)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_44),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g40 ( 
.A1(n_33),
.A2(n_27),
.B(n_21),
.Y(n_40)
);

AOI221xp5_ASAP7_75t_L g46 ( 
.A1(n_40),
.A2(n_41),
.B1(n_35),
.B2(n_32),
.C(n_37),
.Y(n_46)
);

XOR2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR3xp33_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_3),
.C(n_5),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_47),
.B(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_14),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_47),
.A2(n_43),
.B1(n_42),
.B2(n_41),
.Y(n_50)
);

AOI21xp5_ASAP7_75t_L g53 ( 
.A1(n_50),
.A2(n_45),
.B(n_8),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g52 ( 
.A(n_49),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_49),
.C(n_14),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_1),
.A3(n_2),
.B1(n_3),
.B2(n_5),
.C1(n_55),
.C2(n_52),
.Y(n_57)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_1),
.Y(n_58)
);

FAx1_ASAP7_75t_SL g59 ( 
.A(n_58),
.B(n_1),
.CI(n_2),
.CON(n_59),
.SN(n_59)
);


endmodule