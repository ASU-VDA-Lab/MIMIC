module real_jpeg_13470_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx10_ASAP7_75t_L g88 ( 
.A(n_0),
.Y(n_88)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_3),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_3),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_3),
.A2(n_64),
.B1(n_66),
.B2(n_69),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_69),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_3),
.A2(n_31),
.B1(n_32),
.B2(n_69),
.Y(n_111)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_6),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_36),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_6),
.A2(n_36),
.B1(n_48),
.B2(n_50),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_6),
.A2(n_36),
.B1(n_64),
.B2(n_66),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_7),
.A2(n_25),
.B1(n_26),
.B2(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_7),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g181 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_143),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_7),
.A2(n_48),
.B1(n_50),
.B2(n_143),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_7),
.A2(n_64),
.B1(n_66),
.B2(n_143),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_8),
.A2(n_25),
.B1(n_26),
.B2(n_164),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_8),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_164),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_48),
.B1(n_50),
.B2(n_164),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_8),
.A2(n_64),
.B1(n_66),
.B2(n_164),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_10),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_10),
.A2(n_24),
.B1(n_31),
.B2(n_32),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_10),
.A2(n_24),
.B1(n_48),
.B2(n_50),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_24),
.B1(n_64),
.B2(n_66),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_13),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_13),
.B(n_28),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_13),
.B(n_62),
.C(n_64),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_13),
.A2(n_48),
.B1(n_50),
.B2(n_178),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_13),
.A2(n_86),
.B1(n_89),
.B2(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_13),
.B(n_83),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_14),
.A2(n_25),
.B1(n_26),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_14),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_14),
.A2(n_31),
.B1(n_32),
.B2(n_185),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_185),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_14),
.A2(n_64),
.B1(n_66),
.B2(n_185),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_15),
.A2(n_31),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_15),
.A2(n_48),
.B1(n_50),
.B2(n_53),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_15),
.A2(n_25),
.B1(n_26),
.B2(n_53),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_15),
.A2(n_53),
.B1(n_64),
.B2(n_66),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_118),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_116),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_100),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_100),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_73),
.C(n_84),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_20),
.A2(n_21),
.B1(n_73),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_39),
.B1(n_71),
.B2(n_72),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_22),
.B(n_41),
.C(n_57),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_22),
.A2(n_71),
.B1(n_104),
.B2(n_114),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_34),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_23),
.A2(n_28),
.B1(n_97),
.B2(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_25),
.A2(n_26),
.B1(n_30),
.B2(n_33),
.Y(n_38)
);

HAxp5_ASAP7_75t_SL g177 ( 
.A(n_25),
.B(n_178),
.CON(n_177),
.SN(n_177)
);

NAND3xp33_ASAP7_75t_L g179 ( 
.A(n_25),
.B(n_31),
.C(n_33),
.Y(n_179)
);

INVx3_ASAP7_75t_SL g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_28),
.B(n_98),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_28),
.A2(n_97),
.B1(n_177),
.B2(n_184),
.Y(n_200)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_29),
.B(n_35),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_29),
.A2(n_37),
.B1(n_142),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_29),
.A2(n_37),
.B1(n_163),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_30),
.A2(n_32),
.B(n_177),
.C(n_179),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_31),
.A2(n_32),
.B1(n_45),
.B2(n_46),
.Y(n_44)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

HAxp5_ASAP7_75t_SL g236 ( 
.A(n_32),
.B(n_178),
.CON(n_236),
.SN(n_236)
);

NAND3xp33_ASAP7_75t_L g237 ( 
.A(n_32),
.B(n_46),
.C(n_50),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_37),
.A2(n_142),
.B(n_144),
.Y(n_141)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_57),
.B2(n_70),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_51),
.B(n_54),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_42),
.A2(n_110),
.B(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_42),
.A2(n_47),
.B1(n_181),
.B2(n_204),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_42),
.A2(n_47),
.B1(n_204),
.B2(n_212),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_43),
.A2(n_52),
.B1(n_81),
.B2(n_83),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_43),
.B(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_43),
.A2(n_55),
.B(n_111),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_43),
.A2(n_83),
.B1(n_213),
.B2(n_236),
.Y(n_238)
);

AND2x4_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_47),
.Y(n_43)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_45),
.Y(n_46)
);

OA22x2_ASAP7_75t_SL g47 ( 
.A1(n_45),
.A2(n_46),
.B1(n_48),
.B2(n_50),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_45),
.A2(n_48),
.B(n_236),
.C(n_237),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_47),
.B(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_47),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_47),
.A2(n_82),
.B(n_112),
.Y(n_140)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_50),
.B1(n_60),
.B2(n_62),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_48),
.B(n_260),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_57),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_57),
.A2(n_70),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_67),
.B(n_68),
.Y(n_57)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_58),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_58),
.A2(n_67),
.B1(n_94),
.B2(n_139),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_58),
.A2(n_68),
.B(n_95),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_58),
.A2(n_75),
.B(n_250),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_58),
.A2(n_67),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_58),
.A2(n_67),
.B1(n_241),
.B2(n_264),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_63),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_SL g62 ( 
.A(n_60),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.Y(n_63)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_63),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_63),
.B(n_78),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_63),
.A2(n_79),
.B1(n_240),
.B2(n_242),
.Y(n_239)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_64),
.Y(n_66)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_66),
.B(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_66),
.B(n_273),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_67),
.A2(n_77),
.B(n_139),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_67),
.B(n_178),
.Y(n_277)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_68),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_73),
.A2(n_74),
.B(n_80),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_80),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_77),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_79),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_83),
.B(n_111),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_146),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_92),
.B(n_96),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_85),
.A2(n_96),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_85),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_85),
.A2(n_93),
.B1(n_126),
.B2(n_194),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B(n_90),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_86),
.A2(n_155),
.B(n_157),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_86),
.A2(n_89),
.B1(n_267),
.B2(n_275),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_86),
.A2(n_137),
.B(n_269),
.Y(n_289)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_87),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_87),
.A2(n_88),
.B1(n_156),
.B2(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_87),
.A2(n_91),
.B(n_158),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_87),
.A2(n_88),
.B1(n_266),
.B2(n_268),
.Y(n_265)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_88),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_91),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_89),
.B(n_136),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_89),
.A2(n_134),
.B(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_89),
.B(n_178),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_124),
.Y(n_123)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_93),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g125 ( 
.A(n_96),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_98),
.B(n_99),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_102),
.B1(n_103),
.B2(n_115),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_103),
.Y(n_115)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_148),
.B(n_317),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_145),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_121),
.B(n_145),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_127),
.C(n_128),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_122),
.A2(n_123),
.B1(n_127),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_127),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_128),
.A2(n_129),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_140),
.C(n_141),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_130),
.A2(n_131),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_138),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_132),
.A2(n_133),
.B1(n_138),
.B2(n_168),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_137),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_138),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_141),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_149),
.A2(n_310),
.B(n_316),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_196),
.B(n_309),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_186),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_151),
.B(n_186),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_167),
.C(n_169),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_152),
.B(n_167),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_160),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_161),
.C(n_166),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_159),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_154),
.B(n_159),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_165),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_169),
.B(n_307),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_180),
.C(n_182),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_170),
.A2(n_171),
.B1(n_219),
.B2(n_220),
.Y(n_218)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_173),
.B1(n_176),
.B2(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_176),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_182),
.Y(n_219)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_195),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_188),
.B(n_193),
.C(n_195),
.Y(n_315)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

O2A1O1Ixp33_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_224),
.B(n_304),
.C(n_308),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_217),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_217),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.C(n_210),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_199),
.B(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_202),
.C(n_206),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_202),
.A2(n_203),
.B1(n_205),
.B2(n_206),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_207),
.A2(n_208),
.B1(n_210),
.B2(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_210),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_214),
.C(n_216),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g244 ( 
.A(n_211),
.B(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_214),
.A2(n_215),
.B1(n_216),
.B2(n_246),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_218),
.B(n_222),
.C(n_223),
.Y(n_305)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_219),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_298),
.B(n_303),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_253),
.B(n_297),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_243),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_229),
.B(n_243),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_238),
.C(n_239),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_230),
.A2(n_231),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_235),
.Y(n_248)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_238),
.B(n_239),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_242),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_247),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_244),
.B(n_249),
.C(n_251),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_251),
.B2(n_252),
.Y(n_247)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_248),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_249),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_291),
.B(n_296),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_281),
.B(n_290),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_270),
.B(n_280),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_257),
.B(n_265),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_261),
.B2(n_262),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_259),
.B(n_261),
.Y(n_282)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_276),
.B(n_279),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_274),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_278),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_289),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_285),
.B(n_288),
.C(n_289),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_295),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_295),
.Y(n_296)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_299),
.B(n_302),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_302),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_305),
.B(n_306),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_315),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_311),
.B(n_315),
.Y(n_316)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);


endmodule