module fake_jpeg_9359_n_54 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_54);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_54;

wire n_53;
wire n_33;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

AO22x1_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_9),
.B1(n_20),
.B2(n_19),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_29),
.A2(n_34),
.B1(n_16),
.B2(n_33),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_23),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_32),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_0),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_2),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_26),
.B(n_0),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_23),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_33),
.A2(n_22),
.B1(n_3),
.B2(n_4),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_26),
.A2(n_11),
.B1(n_18),
.B2(n_17),
.Y(n_34)
);

AOI21xp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_22),
.C(n_5),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_4),
.C(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

OA21x2_ASAP7_75t_L g41 ( 
.A1(n_33),
.A2(n_21),
.B(n_7),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_31),
.B(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_13),
.Y(n_43)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_43),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_50),
.C(n_46),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_48),
.C(n_39),
.Y(n_53)
);

AOI221xp5_ASAP7_75t_L g54 ( 
.A1(n_53),
.A2(n_44),
.B1(n_35),
.B2(n_45),
.C(n_40),
.Y(n_54)
);


endmodule