module real_jpeg_5917_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_173;
wire n_105;
wire n_40;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_139;
wire n_33;
wire n_188;
wire n_65;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_225;
wire n_103;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

INVx8_ASAP7_75t_L g90 ( 
.A(n_0),
.Y(n_90)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_1),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_1),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_1),
.B(n_143),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_1),
.B(n_193),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_3),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_4),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_4),
.B(n_92),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_4),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_4),
.B(n_124),
.Y(n_123)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_6),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_7),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_7),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_7),
.B(n_73),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_7),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_7),
.B(n_182),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_7),
.B(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_7),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_8),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_8),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_8),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_8),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_8),
.B(n_193),
.Y(n_221)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_9),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_9),
.Y(n_135)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g29 ( 
.A(n_11),
.B(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_13),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_13),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_13),
.B(n_133),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_13),
.B(n_184),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_13),
.B(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_13),
.B(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_14),
.B(n_53),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_14),
.B(n_109),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_14),
.B(n_139),
.Y(n_138)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_15),
.Y(n_94)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_15),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_15),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_15),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_16),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_16),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_16),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_16),
.B(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_16),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_16),
.B(n_211),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_16),
.B(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_173),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_171),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_147),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_21),
.B(n_147),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_62),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_36),
.B2(n_61),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

XNOR2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_31),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_31),
.Y(n_194)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_35),
.Y(n_220)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

XNOR2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_45),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_L g81 ( 
.A1(n_37),
.A2(n_38),
.B(n_40),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_40),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_44),
.Y(n_145)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_44),
.Y(n_159)
);

MAJx2_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_51),
.C(n_55),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_46),
.A2(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_101)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx8_ASAP7_75t_L g202 ( 
.A(n_54),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_55),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_60),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_59),
.Y(n_131)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_59),
.Y(n_166)
);

BUFx3_ASAP7_75t_L g232 ( 
.A(n_59),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_60),
.B(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_81),
.C(n_82),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_63),
.B(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_71),
.C(n_76),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_64),
.B(n_261),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_68),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_65),
.A2(n_66),
.B1(n_68),
.B2(n_69),
.Y(n_248)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_70),
.Y(n_109)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_72),
.B(n_77),
.Y(n_261)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_81),
.A2(n_82),
.B1(n_83),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_81),
.Y(n_150)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_86),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_84),
.B(n_91),
.C(n_95),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_86)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_90),
.Y(n_116)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_90),
.Y(n_125)
);

BUFx5_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_90),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_91),
.Y(n_96)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_94),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_SL g97 ( 
.A(n_98),
.B(n_121),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_102),
.C(n_110),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_99),
.A2(n_100),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_103),
.B(n_111),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_108),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_104),
.B(n_108),
.Y(n_167)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_107),
.Y(n_182)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.C(n_117),
.Y(n_111)
);

FAx1_ASAP7_75t_SL g152 ( 
.A(n_112),
.B(n_114),
.CI(n_117),
.CON(n_152),
.SN(n_152)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_120),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_136),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_126),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_132),
.Y(n_126)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_146),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_142),
.Y(n_137)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_141),
.Y(n_208)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_168),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_148),
.B(n_270),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_151),
.B(n_168),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.C(n_167),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_152),
.B(n_264),
.Y(n_263)
);

BUFx24_ASAP7_75t_SL g275 ( 
.A(n_152),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_153),
.A2(n_154),
.B1(n_167),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.Y(n_153)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_160),
.C(n_163),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_155),
.A2(n_156),
.B1(n_163),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_160),
.B(n_254),
.Y(n_253)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_163),
.Y(n_255)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

OAI21x1_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_268),
.B(n_273),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_257),
.B(n_267),
.Y(n_174)
);

OAI21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_237),
.B(n_256),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_214),
.B(n_236),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_196),
.B(n_213),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_191),
.B(n_195),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_187),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_180),
.B(n_187),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_183),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_181),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_181),
.B(n_183),
.Y(n_197)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_197),
.B(n_198),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_204),
.B2(n_205),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_199),
.B(n_207),
.C(n_209),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_201),
.B(n_203),
.Y(n_222)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_215),
.B(n_235),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_235),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_222),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.C(n_239),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_218),
.B(n_221),
.Y(n_242)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_224),
.B(n_251),
.C(n_252),
.Y(n_250)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_233),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_240),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_238),
.B(n_240),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_249),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_250),
.C(n_253),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_242),
.B(n_244),
.C(n_248),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_248),
.Y(n_243)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_253),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_266),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_263),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_262),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_262),
.C(n_272),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_263),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_271),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_271),
.Y(n_273)
);


endmodule