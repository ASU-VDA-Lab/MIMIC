module fake_netlist_1_7796_n_704 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_704);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_704;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_529;
wire n_455;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_624;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_420;
wire n_342;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
NOR2xp67_ASAP7_75t_L g78 ( .A(n_41), .B(n_35), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_50), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_46), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_6), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_16), .Y(n_82) );
CKINVDCx5p33_ASAP7_75t_R g83 ( .A(n_72), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_14), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_55), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_48), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_14), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_31), .Y(n_88) );
CKINVDCx14_ASAP7_75t_R g89 ( .A(n_26), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_10), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_51), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_34), .Y(n_92) );
INVx2_ASAP7_75t_SL g93 ( .A(n_38), .Y(n_93) );
CKINVDCx5p33_ASAP7_75t_R g94 ( .A(n_0), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_49), .Y(n_95) );
CKINVDCx20_ASAP7_75t_R g96 ( .A(n_33), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_28), .Y(n_97) );
BUFx5_ASAP7_75t_L g98 ( .A(n_64), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_61), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_11), .Y(n_100) );
INVx2_ASAP7_75t_L g101 ( .A(n_56), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_17), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_8), .Y(n_103) );
INVxp67_ASAP7_75t_L g104 ( .A(n_71), .Y(n_104) );
INVxp67_ASAP7_75t_L g105 ( .A(n_63), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_9), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_74), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_13), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_42), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_47), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_59), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_2), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_57), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_43), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_40), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_68), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_32), .Y(n_117) );
INVxp33_ASAP7_75t_L g118 ( .A(n_53), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_16), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_1), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g121 ( .A(n_52), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_39), .Y(n_122) );
NOR2xp67_ASAP7_75t_L g123 ( .A(n_58), .B(n_69), .Y(n_123) );
INVxp33_ASAP7_75t_SL g124 ( .A(n_8), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_13), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_98), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_90), .Y(n_127) );
NAND2xp33_ASAP7_75t_SL g128 ( .A(n_118), .B(n_0), .Y(n_128) );
OAI21x1_ASAP7_75t_L g129 ( .A1(n_101), .A2(n_24), .B(n_76), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_93), .B(n_1), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_90), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_122), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_122), .B(n_2), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_79), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_112), .B(n_3), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_101), .Y(n_139) );
CKINVDCx16_ASAP7_75t_R g140 ( .A(n_81), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_98), .Y(n_141) );
BUFx6f_ASAP7_75t_L g142 ( .A(n_85), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_98), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g144 ( .A(n_118), .B(n_3), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_89), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_92), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_89), .B(n_4), .Y(n_147) );
OAI22xp5_ASAP7_75t_SL g148 ( .A1(n_81), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g149 ( .A1(n_124), .A2(n_5), .B1(n_7), .B2(n_9), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_102), .Y(n_150) );
OAI22x1_ASAP7_75t_L g151 ( .A1(n_108), .A2(n_7), .B1(n_10), .B2(n_11), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_97), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_96), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_99), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_109), .Y(n_155) );
BUFx2_ASAP7_75t_L g156 ( .A(n_82), .Y(n_156) );
CKINVDCx20_ASAP7_75t_R g157 ( .A(n_84), .Y(n_157) );
CKINVDCx5p33_ASAP7_75t_R g158 ( .A(n_96), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_84), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_110), .Y(n_161) );
BUFx2_ASAP7_75t_L g162 ( .A(n_100), .Y(n_162) );
BUFx6f_ASAP7_75t_L g163 ( .A(n_114), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_119), .B(n_12), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_116), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_117), .Y(n_167) );
INVx5_ASAP7_75t_L g168 ( .A(n_98), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_156), .B(n_103), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_126), .Y(n_170) );
A2O1A1Ixp33_ASAP7_75t_L g171 ( .A1(n_137), .A2(n_125), .B(n_120), .C(n_113), .Y(n_171) );
OR2x2_ASAP7_75t_L g172 ( .A(n_156), .B(n_106), .Y(n_172) );
AOI22xp5_ASAP7_75t_L g173 ( .A1(n_147), .A2(n_121), .B1(n_111), .B2(n_86), .Y(n_173) );
BUFx3_ASAP7_75t_L g174 ( .A(n_132), .Y(n_174) );
AND2x2_ASAP7_75t_L g175 ( .A(n_162), .B(n_147), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_126), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_133), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_132), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_133), .Y(n_179) );
NAND2x1p5_ASAP7_75t_L g180 ( .A(n_134), .B(n_123), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_162), .B(n_104), .Y(n_181) );
BUFx6f_ASAP7_75t_L g182 ( .A(n_129), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_132), .Y(n_183) );
INVxp67_ASAP7_75t_L g184 ( .A(n_159), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_135), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_134), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_167), .B(n_95), .Y(n_187) );
HB1xp67_ASAP7_75t_L g188 ( .A(n_145), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_135), .Y(n_190) );
INVx3_ASAP7_75t_L g191 ( .A(n_134), .Y(n_191) );
AND2x2_ASAP7_75t_SL g192 ( .A(n_144), .B(n_121), .Y(n_192) );
BUFx4f_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
BUFx4f_ASAP7_75t_L g194 ( .A(n_142), .Y(n_194) );
BUFx10_ASAP7_75t_L g195 ( .A(n_145), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_128), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_141), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_141), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_139), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_167), .B(n_105), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_139), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_139), .Y(n_203) );
INVx3_ASAP7_75t_L g204 ( .A(n_142), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_132), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_143), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_132), .Y(n_207) );
AND2x4_ASAP7_75t_L g208 ( .A(n_136), .B(n_78), .Y(n_208) );
INVx1_ASAP7_75t_L g209 ( .A(n_143), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_168), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_142), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_137), .B(n_107), .Y(n_212) );
AND2x2_ASAP7_75t_L g213 ( .A(n_136), .B(n_98), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_146), .B(n_91), .Y(n_214) );
AND2x6_ASAP7_75t_L g215 ( .A(n_146), .B(n_111), .Y(n_215) );
BUFx10_ASAP7_75t_L g216 ( .A(n_152), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_136), .B(n_88), .Y(n_217) );
BUFx6f_ASAP7_75t_L g218 ( .A(n_129), .Y(n_218) );
AND3x4_ASAP7_75t_L g219 ( .A(n_148), .B(n_12), .C(n_15), .Y(n_219) );
INVx6_ASAP7_75t_L g220 ( .A(n_168), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_168), .Y(n_222) );
OAI21xp33_ASAP7_75t_SL g223 ( .A1(n_152), .A2(n_15), .B(n_17), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_168), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_142), .Y(n_225) );
AND2x6_ASAP7_75t_L g226 ( .A(n_154), .B(n_18), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_155), .Y(n_227) );
INVx4_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
BUFx6f_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_155), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_150), .B(n_83), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_195), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_216), .Y(n_233) );
AOI22xp33_ASAP7_75t_L g234 ( .A1(n_175), .A2(n_166), .B1(n_154), .B2(n_164), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_216), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_216), .B(n_166), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_231), .B(n_164), .Y(n_237) );
AND2x4_ASAP7_75t_L g238 ( .A(n_217), .B(n_150), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_182), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_184), .B(n_140), .Y(n_240) );
INVx2_ASAP7_75t_SL g241 ( .A(n_172), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_231), .B(n_161), .Y(n_242) );
INVx5_ASAP7_75t_L g243 ( .A(n_228), .Y(n_243) );
INVx4_ASAP7_75t_L g244 ( .A(n_228), .Y(n_244) );
BUFx12f_ASAP7_75t_L g245 ( .A(n_195), .Y(n_245) );
INVx3_ASAP7_75t_L g246 ( .A(n_186), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_173), .Y(n_247) );
HB1xp67_ASAP7_75t_L g248 ( .A(n_175), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_217), .B(n_130), .Y(n_249) );
OR2x6_ASAP7_75t_L g250 ( .A(n_196), .B(n_151), .Y(n_250) );
HB1xp67_ASAP7_75t_L g251 ( .A(n_172), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_186), .B(n_161), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_174), .Y(n_253) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_196), .A2(n_138), .B1(n_149), .B2(n_165), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_182), .A2(n_150), .B(n_155), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_174), .Y(n_256) );
AND2x4_ASAP7_75t_L g257 ( .A(n_217), .B(n_131), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_201), .B(n_131), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_186), .B(n_163), .Y(n_259) );
AND2x4_ASAP7_75t_SL g260 ( .A(n_195), .B(n_160), .Y(n_260) );
BUFx4f_ASAP7_75t_L g261 ( .A(n_226), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_178), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_191), .B(n_163), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_191), .B(n_163), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g265 ( .A(n_181), .B(n_158), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_215), .A2(n_153), .B1(n_158), .B2(n_151), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_213), .Y(n_267) );
BUFx2_ASAP7_75t_L g268 ( .A(n_215), .Y(n_268) );
AND2x2_ASAP7_75t_L g269 ( .A(n_181), .B(n_153), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_215), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_169), .B(n_80), .Y(n_271) );
BUFx6f_ASAP7_75t_L g272 ( .A(n_182), .Y(n_272) );
BUFx3_ASAP7_75t_L g273 ( .A(n_208), .Y(n_273) );
INVx8_ASAP7_75t_L g274 ( .A(n_215), .Y(n_274) );
NOR2x1_ASAP7_75t_L g275 ( .A(n_187), .B(n_127), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_191), .B(n_163), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_182), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_213), .Y(n_278) );
INVx5_ASAP7_75t_L g279 ( .A(n_228), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_212), .B(n_155), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_208), .Y(n_281) );
AND2x4_ASAP7_75t_L g282 ( .A(n_208), .B(n_127), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_208), .Y(n_283) );
BUFx3_ASAP7_75t_L g284 ( .A(n_178), .Y(n_284) );
AND2x4_ASAP7_75t_L g285 ( .A(n_188), .B(n_163), .Y(n_285) );
OR2x2_ASAP7_75t_L g286 ( .A(n_171), .B(n_157), .Y(n_286) );
NAND2xp5_ASAP7_75t_SL g287 ( .A(n_214), .B(n_180), .Y(n_287) );
NOR2x1_ASAP7_75t_L g288 ( .A(n_219), .B(n_185), .Y(n_288) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_180), .A2(n_19), .B1(n_20), .B2(n_21), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
INVx2_ASAP7_75t_SL g291 ( .A(n_180), .Y(n_291) );
OAI21xp5_ASAP7_75t_L g292 ( .A1(n_170), .A2(n_22), .B(n_23), .Y(n_292) );
INVx4_ASAP7_75t_L g293 ( .A(n_220), .Y(n_293) );
NOR2xp33_ASAP7_75t_L g294 ( .A(n_192), .B(n_25), .Y(n_294) );
AND2x2_ASAP7_75t_SL g295 ( .A(n_192), .B(n_27), .Y(n_295) );
INVx2_ASAP7_75t_L g296 ( .A(n_183), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_170), .B(n_29), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_176), .B(n_30), .Y(n_298) );
AOI22xp33_ASAP7_75t_L g299 ( .A1(n_295), .A2(n_215), .B1(n_192), .B2(n_219), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_246), .Y(n_300) );
INVxp67_ASAP7_75t_L g301 ( .A(n_251), .Y(n_301) );
AO22x1_ASAP7_75t_L g302 ( .A1(n_288), .A2(n_215), .B1(n_219), .B2(n_226), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_236), .B(n_215), .Y(n_303) );
O2A1O1Ixp33_ASAP7_75t_L g304 ( .A1(n_248), .A2(n_223), .B(n_237), .C(n_242), .Y(n_304) );
INVx2_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
INVx4_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
AND2x2_ASAP7_75t_L g307 ( .A(n_251), .B(n_223), .Y(n_307) );
CKINVDCx8_ASAP7_75t_R g308 ( .A(n_250), .Y(n_308) );
INVx3_ASAP7_75t_L g309 ( .A(n_244), .Y(n_309) );
INVx4_ASAP7_75t_L g310 ( .A(n_232), .Y(n_310) );
INVx3_ASAP7_75t_L g311 ( .A(n_244), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_236), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_241), .B(n_182), .Y(n_313) );
BUFx3_ASAP7_75t_L g314 ( .A(n_260), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_237), .B(n_197), .Y(n_315) );
INVx2_ASAP7_75t_L g316 ( .A(n_259), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_242), .B(n_197), .Y(n_317) );
OAI21xp5_ASAP7_75t_L g318 ( .A1(n_255), .A2(n_198), .B(n_177), .Y(n_318) );
AOI21xp5_ASAP7_75t_L g319 ( .A1(n_255), .A2(n_218), .B(n_209), .Y(n_319) );
INVx2_ASAP7_75t_SL g320 ( .A(n_240), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_248), .A2(n_198), .B(n_177), .C(n_176), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_269), .Y(n_322) );
CKINVDCx14_ASAP7_75t_R g323 ( .A(n_250), .Y(n_323) );
AOI21xp5_ASAP7_75t_L g324 ( .A1(n_252), .A2(n_218), .B(n_185), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_252), .A2(n_218), .B(n_190), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_265), .Y(n_326) );
O2A1O1Ixp33_ASAP7_75t_L g327 ( .A1(n_249), .A2(n_179), .B(n_206), .C(n_190), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_239), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_234), .A2(n_218), .B1(n_209), .B2(n_179), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_259), .Y(n_330) );
INVx2_ASAP7_75t_L g331 ( .A(n_263), .Y(n_331) );
AOI21xp5_ASAP7_75t_L g332 ( .A1(n_261), .A2(n_218), .B(n_206), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_243), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_239), .Y(n_334) );
OAI22x1_ASAP7_75t_L g335 ( .A1(n_266), .A2(n_226), .B1(n_227), .B2(n_211), .Y(n_335) );
AND2x6_ASAP7_75t_L g336 ( .A(n_267), .B(n_226), .Y(n_336) );
OR2x6_ASAP7_75t_L g337 ( .A(n_274), .B(n_220), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_257), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_291), .B(n_226), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_261), .A2(n_221), .B(n_210), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_263), .A2(n_221), .B(n_210), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_239), .Y(n_342) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_272), .Y(n_343) );
O2A1O1Ixp33_ASAP7_75t_L g344 ( .A1(n_286), .A2(n_224), .B(n_222), .C(n_204), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_264), .Y(n_345) );
OAI22x1_ASAP7_75t_L g346 ( .A1(n_247), .A2(n_226), .B1(n_227), .B2(n_211), .Y(n_346) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_238), .A2(n_226), .B1(n_193), .B2(n_194), .Y(n_347) );
BUFx3_ASAP7_75t_L g348 ( .A(n_285), .Y(n_348) );
A2O1A1Ixp33_ASAP7_75t_L g349 ( .A1(n_278), .A2(n_193), .B(n_194), .C(n_204), .Y(n_349) );
O2A1O1Ixp5_ASAP7_75t_SL g350 ( .A1(n_280), .A2(n_225), .B(n_204), .C(n_229), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_350), .A2(n_292), .B(n_297), .Y(n_351) );
OAI222xp33_ASAP7_75t_L g352 ( .A1(n_299), .A2(n_250), .B1(n_289), .B2(n_294), .C1(n_254), .C2(n_268), .Y(n_352) );
OAI21x1_ASAP7_75t_L g353 ( .A1(n_319), .A2(n_292), .B(n_297), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_312), .B(n_233), .Y(n_354) );
NAND2x1p5_ASAP7_75t_L g355 ( .A(n_333), .B(n_235), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g356 ( .A1(n_315), .A2(n_317), .B1(n_301), .B2(n_326), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_310), .B(n_238), .Y(n_357) );
NOR2xp33_ASAP7_75t_R g358 ( .A(n_323), .B(n_274), .Y(n_358) );
BUFx2_ASAP7_75t_L g359 ( .A(n_337), .Y(n_359) );
CKINVDCx11_ASAP7_75t_R g360 ( .A(n_306), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_319), .A2(n_298), .B(n_207), .Y(n_361) );
OAI21x1_ASAP7_75t_L g362 ( .A1(n_332), .A2(n_324), .B(n_325), .Y(n_362) );
OAI21x1_ASAP7_75t_L g363 ( .A1(n_332), .A2(n_298), .B(n_264), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_324), .A2(n_276), .B(n_275), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_320), .B(n_273), .Y(n_365) );
OAI221xp5_ASAP7_75t_L g366 ( .A1(n_322), .A2(n_281), .B1(n_283), .B2(n_287), .C(n_271), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_315), .Y(n_367) );
A2O1A1Ixp33_ASAP7_75t_L g368 ( .A1(n_304), .A2(n_276), .B(n_257), .C(n_285), .Y(n_368) );
OAI21x1_ASAP7_75t_L g369 ( .A1(n_325), .A2(n_207), .B(n_205), .Y(n_369) );
OAI21x1_ASAP7_75t_L g370 ( .A1(n_329), .A2(n_205), .B(n_272), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_329), .A2(n_289), .B(n_203), .Y(n_371) );
INVx6_ASAP7_75t_L g372 ( .A(n_310), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_307), .B(n_282), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_316), .Y(n_374) );
INVx5_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
INVx3_ASAP7_75t_L g376 ( .A(n_333), .Y(n_376) );
OA21x2_ASAP7_75t_L g377 ( .A1(n_318), .A2(n_203), .B(n_202), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_317), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_330), .Y(n_379) );
NAND3x1_ASAP7_75t_L g380 ( .A(n_308), .B(n_274), .C(n_270), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_340), .A2(n_277), .B(n_272), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_328), .Y(n_382) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_367), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_378), .B(n_331), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_356), .A2(n_348), .B1(n_282), .B2(n_338), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_378), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_367), .A2(n_314), .B1(n_313), .B2(n_303), .Y(n_387) );
AOI21xp5_ASAP7_75t_L g388 ( .A1(n_351), .A2(n_334), .B(n_343), .Y(n_388) );
AOI22xp33_ASAP7_75t_L g389 ( .A1(n_366), .A2(n_303), .B1(n_336), .B2(n_335), .Y(n_389) );
INVxp67_ASAP7_75t_L g390 ( .A(n_365), .Y(n_390) );
OAI211xp5_ASAP7_75t_L g391 ( .A1(n_373), .A2(n_304), .B(n_344), .C(n_347), .Y(n_391) );
AOI21xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_328), .B(n_334), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_379), .B(n_302), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_379), .B(n_374), .Y(n_394) );
AOI221xp5_ASAP7_75t_L g395 ( .A1(n_352), .A2(n_321), .B1(n_258), .B2(n_327), .C(n_306), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_360), .A2(n_349), .B(n_327), .C(n_225), .Y(n_396) );
AOI22xp33_ASAP7_75t_SL g397 ( .A1(n_375), .A2(n_336), .B1(n_339), .B2(n_337), .Y(n_397) );
OAI221xp5_ASAP7_75t_L g398 ( .A1(n_368), .A2(n_318), .B1(n_345), .B2(n_305), .C(n_300), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_374), .B(n_258), .Y(n_399) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_375), .A2(n_336), .B1(n_311), .B2(n_309), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_364), .Y(n_401) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_354), .A2(n_340), .B1(n_341), .B2(n_311), .C(n_309), .Y(n_402) );
OA21x2_ASAP7_75t_L g403 ( .A1(n_370), .A2(n_341), .B(n_189), .Y(n_403) );
AO21x1_ASAP7_75t_L g404 ( .A1(n_362), .A2(n_189), .B(n_199), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_362), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_364), .Y(n_406) );
AND2x2_ASAP7_75t_L g407 ( .A(n_357), .B(n_336), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_371), .B(n_346), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_371), .B(n_253), .Y(n_409) );
AND2x4_ASAP7_75t_L g410 ( .A(n_375), .B(n_343), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_383), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_394), .B(n_376), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_405), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_394), .B(n_376), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_386), .B(n_375), .Y(n_415) );
HB1xp67_ASAP7_75t_L g416 ( .A(n_401), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_386), .B(n_357), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_401), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_405), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_406), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_384), .B(n_376), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_406), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_384), .B(n_371), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_405), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_399), .B(n_376), .Y(n_425) );
AND2x4_ASAP7_75t_L g426 ( .A(n_410), .B(n_375), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_393), .B(n_377), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_393), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_403), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_404), .Y(n_430) );
NOR2x1_ASAP7_75t_L g431 ( .A(n_396), .B(n_359), .Y(n_431) );
AOI22xp33_ASAP7_75t_SL g432 ( .A1(n_391), .A2(n_359), .B1(n_375), .B2(n_358), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_403), .Y(n_433) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_403), .Y(n_434) );
NAND3xp33_ASAP7_75t_L g435 ( .A(n_395), .B(n_361), .C(n_377), .Y(n_435) );
AO21x2_ASAP7_75t_L g436 ( .A1(n_408), .A2(n_370), .B(n_353), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_409), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx3_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
INVx3_ASAP7_75t_L g441 ( .A(n_410), .Y(n_441) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_403), .Y(n_442) );
AO21x2_ASAP7_75t_L g443 ( .A1(n_408), .A2(n_353), .B(n_381), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_399), .B(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_398), .Y(n_445) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_412), .B(n_377), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_418), .Y(n_448) );
INVx5_ASAP7_75t_L g449 ( .A(n_446), .Y(n_449) );
NAND4xp25_ASAP7_75t_L g450 ( .A(n_432), .B(n_395), .C(n_385), .D(n_390), .Y(n_450) );
INVx2_ASAP7_75t_L g451 ( .A(n_413), .Y(n_451) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_411), .Y(n_452) );
INVx4_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
OAI221xp5_ASAP7_75t_L g454 ( .A1(n_432), .A2(n_387), .B1(n_389), .B2(n_398), .C(n_397), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_423), .B(n_377), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_418), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_412), .B(n_361), .Y(n_457) );
INVx4_ASAP7_75t_L g458 ( .A(n_415), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_413), .Y(n_459) );
NAND4xp25_ASAP7_75t_L g460 ( .A(n_411), .B(n_357), .C(n_402), .D(n_400), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_413), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_420), .B(n_392), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_420), .Y(n_463) );
INVx2_ASAP7_75t_L g464 ( .A(n_419), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_414), .B(n_361), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_423), .B(n_361), .Y(n_467) );
NAND4xp25_ASAP7_75t_L g468 ( .A(n_431), .B(n_357), .C(n_402), .D(n_407), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_419), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_422), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_419), .Y(n_471) );
AOI21xp5_ASAP7_75t_L g472 ( .A1(n_435), .A2(n_388), .B(n_381), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_415), .A2(n_372), .B1(n_355), .B2(n_363), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_416), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_414), .B(n_363), .Y(n_475) );
AND2x2_ASAP7_75t_L g476 ( .A(n_444), .B(n_369), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_416), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_446), .B(n_369), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_446), .B(n_382), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_428), .Y(n_481) );
INVx2_ASAP7_75t_L g482 ( .A(n_424), .Y(n_482) );
AOI33xp33_ASAP7_75t_L g483 ( .A1(n_445), .A2(n_230), .A3(n_199), .B1(n_200), .B2(n_202), .B3(n_262), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_431), .A2(n_372), .B1(n_355), .B2(n_193), .C(n_194), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_446), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_424), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_444), .B(n_382), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_421), .B(n_372), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_438), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_421), .B(n_382), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_415), .B(n_355), .Y(n_492) );
INVxp67_ASAP7_75t_L g493 ( .A(n_417), .Y(n_493) );
INVx1_ASAP7_75t_SL g494 ( .A(n_426), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_429), .Y(n_495) );
INVxp67_ASAP7_75t_SL g496 ( .A(n_429), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_427), .B(n_372), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_493), .B(n_445), .Y(n_498) );
OAI211xp5_ASAP7_75t_L g499 ( .A1(n_450), .A2(n_417), .B(n_441), .C(n_440), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_480), .B(n_438), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_475), .B(n_427), .Y(n_501) );
HB1xp67_ASAP7_75t_L g502 ( .A(n_452), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_448), .Y(n_503) );
NAND4xp25_ASAP7_75t_L g504 ( .A(n_450), .B(n_435), .C(n_425), .D(n_430), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_475), .B(n_427), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_457), .B(n_439), .Y(n_506) );
OAI221xp5_ASAP7_75t_L g507 ( .A1(n_460), .A2(n_430), .B1(n_437), .B2(n_441), .C(n_440), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_457), .B(n_439), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_465), .B(n_434), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_465), .B(n_434), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_480), .B(n_425), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_481), .B(n_440), .Y(n_513) );
INVx3_ASAP7_75t_L g514 ( .A(n_453), .Y(n_514) );
HB1xp67_ASAP7_75t_L g515 ( .A(n_497), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_482), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_474), .B(n_437), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_476), .B(n_442), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_497), .B(n_440), .Y(n_519) );
NAND3xp33_ASAP7_75t_SL g520 ( .A(n_484), .B(n_442), .C(n_433), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_476), .B(n_433), .Y(n_521) );
OAI33xp33_ASAP7_75t_L g522 ( .A1(n_481), .A2(n_200), .A3(n_230), .B1(n_443), .B2(n_436), .B3(n_380), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_490), .B(n_441), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_456), .Y(n_524) );
BUFx2_ASAP7_75t_L g525 ( .A(n_453), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_456), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_482), .Y(n_527) );
OR2x2_ASAP7_75t_L g528 ( .A(n_474), .B(n_443), .Y(n_528) );
INVx1_ASAP7_75t_SL g529 ( .A(n_494), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_463), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_463), .Y(n_531) );
NAND3xp33_ASAP7_75t_L g532 ( .A(n_460), .B(n_446), .C(n_441), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_447), .B(n_443), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_489), .B(n_426), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_466), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_490), .B(n_446), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_487), .B(n_446), .Y(n_537) );
BUFx2_ASAP7_75t_L g538 ( .A(n_453), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_487), .B(n_426), .Y(n_539) );
AND2x4_ASAP7_75t_L g540 ( .A(n_453), .B(n_443), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_466), .B(n_426), .Y(n_541) );
INVxp67_ASAP7_75t_SL g542 ( .A(n_496), .Y(n_542) );
AND2x4_ASAP7_75t_SL g543 ( .A(n_458), .B(n_328), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_447), .B(n_436), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_470), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_470), .B(n_436), .Y(n_546) );
NAND2xp33_ASAP7_75t_L g547 ( .A(n_473), .B(n_380), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_495), .B(n_436), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_477), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_449), .B(n_343), .Y(n_550) );
BUFx3_ASAP7_75t_L g551 ( .A(n_449), .Y(n_551) );
A2O1A1Ixp33_ASAP7_75t_L g552 ( .A1(n_468), .A2(n_277), .B(n_334), .C(n_342), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_477), .B(n_229), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_491), .B(n_229), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_491), .B(n_229), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_502), .B(n_467), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_547), .A2(n_468), .B1(n_454), .B2(n_458), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_501), .B(n_462), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_525), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_542), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_516), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_549), .B(n_467), .Y(n_563) );
NAND2xp33_ASAP7_75t_R g564 ( .A(n_538), .B(n_478), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_501), .B(n_462), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_503), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_505), .B(n_458), .Y(n_567) );
INVxp33_ASAP7_75t_L g568 ( .A(n_534), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_505), .B(n_458), .Y(n_569) );
HB1xp67_ASAP7_75t_L g570 ( .A(n_555), .Y(n_570) );
HB1xp67_ASAP7_75t_L g571 ( .A(n_529), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_533), .B(n_462), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_511), .Y(n_573) );
NAND2x1_ASAP7_75t_L g574 ( .A(n_514), .B(n_482), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_533), .B(n_544), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_506), .B(n_455), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_544), .B(n_462), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_518), .B(n_486), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_524), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_518), .B(n_521), .Y(n_580) );
INVx2_ASAP7_75t_SL g581 ( .A(n_551), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_526), .Y(n_582) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_512), .B(n_449), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_521), .B(n_486), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_509), .B(n_486), .Y(n_585) );
AOI21xp33_ASAP7_75t_SL g586 ( .A1(n_499), .A2(n_492), .B(n_455), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_509), .B(n_488), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_530), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_510), .B(n_488), .Y(n_589) );
NOR2xp33_ASAP7_75t_SL g590 ( .A(n_551), .B(n_449), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_514), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_531), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_506), .B(n_485), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_508), .B(n_485), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_510), .B(n_464), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_535), .Y(n_597) );
OR2x2_ASAP7_75t_L g598 ( .A(n_508), .B(n_471), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_547), .B(n_459), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_498), .B(n_464), .Y(n_600) );
AND2x4_ASAP7_75t_L g601 ( .A(n_540), .B(n_449), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_545), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_515), .B(n_461), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
BUFx2_ASAP7_75t_L g605 ( .A(n_514), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_546), .B(n_469), .Y(n_606) );
INVx1_ASAP7_75t_L g607 ( .A(n_528), .Y(n_607) );
INVx1_ASAP7_75t_SL g608 ( .A(n_543), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_558), .A2(n_504), .B1(n_532), .B2(n_541), .Y(n_609) );
INVxp67_ASAP7_75t_L g610 ( .A(n_561), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_580), .B(n_546), .Y(n_611) );
AOI222xp33_ASAP7_75t_L g612 ( .A1(n_599), .A2(n_557), .B1(n_607), .B2(n_566), .C1(n_579), .C2(n_582), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_575), .B(n_517), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_570), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_566), .Y(n_615) );
INVx1_ASAP7_75t_SL g616 ( .A(n_560), .Y(n_616) );
AND2x4_ASAP7_75t_L g617 ( .A(n_601), .B(n_540), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_589), .B(n_598), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_573), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_599), .A2(n_552), .B1(n_539), .B2(n_519), .Y(n_621) );
OAI22xp33_ASAP7_75t_L g622 ( .A1(n_590), .A2(n_520), .B1(n_449), .B2(n_507), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_579), .Y(n_623) );
OAI21xp33_ASAP7_75t_L g624 ( .A1(n_568), .A2(n_552), .B(n_540), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g625 ( .A1(n_574), .A2(n_522), .B(n_550), .Y(n_625) );
OAI322xp33_ASAP7_75t_L g626 ( .A1(n_607), .A2(n_517), .A3(n_528), .B1(n_523), .B2(n_513), .C1(n_500), .C2(n_553), .Y(n_626) );
OAI211xp5_ASAP7_75t_L g627 ( .A1(n_586), .A2(n_537), .B(n_536), .C(n_548), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_571), .A2(n_553), .B(n_483), .Y(n_628) );
AOI22xp5_ASAP7_75t_L g629 ( .A1(n_583), .A2(n_564), .B1(n_577), .B2(n_572), .Y(n_629) );
AOI221xp5_ASAP7_75t_L g630 ( .A1(n_572), .A2(n_548), .B1(n_554), .B2(n_556), .C(n_472), .Y(n_630) );
OAI221xp5_ASAP7_75t_L g631 ( .A1(n_605), .A2(n_527), .B1(n_459), .B2(n_451), .C(n_461), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_580), .B(n_478), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_575), .B(n_471), .Y(n_633) );
OAI33xp33_ASAP7_75t_L g634 ( .A1(n_593), .A2(n_469), .A3(n_451), .B1(n_550), .B2(n_478), .B3(n_479), .Y(n_634) );
AOI221xp5_ASAP7_75t_L g635 ( .A1(n_577), .A2(n_478), .B1(n_479), .B2(n_229), .C(n_543), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_582), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g637 ( .A1(n_588), .A2(n_479), .B1(n_225), .B2(n_296), .C(n_290), .Y(n_637) );
NOR2xp67_ASAP7_75t_SL g638 ( .A(n_581), .B(n_605), .Y(n_638) );
OAI22xp33_ASAP7_75t_L g639 ( .A1(n_608), .A2(n_479), .B1(n_277), .B2(n_342), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_588), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_592), .Y(n_641) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_581), .B(n_342), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_559), .A2(n_284), .B1(n_256), .B2(n_293), .Y(n_643) );
AOI22xp5_ASAP7_75t_L g644 ( .A1(n_559), .A2(n_293), .B1(n_279), .B2(n_243), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_565), .B(n_36), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_614), .Y(n_646) );
AOI22xp5_ASAP7_75t_L g647 ( .A1(n_609), .A2(n_565), .B1(n_567), .B2(n_569), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_615), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g649 ( .A1(n_629), .A2(n_576), .B1(n_591), .B2(n_598), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_618), .Y(n_650) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_612), .A2(n_622), .B(n_627), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_634), .A2(n_626), .B1(n_610), .B2(n_630), .C(n_624), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_620), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_623), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g655 ( .A1(n_612), .A2(n_594), .B1(n_587), .B2(n_596), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_636), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_616), .B(n_587), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_640), .Y(n_658) );
OAI22xp5_ASAP7_75t_L g659 ( .A1(n_616), .A2(n_591), .B1(n_589), .B2(n_574), .Y(n_659) );
OAI22xp33_ASAP7_75t_SL g660 ( .A1(n_621), .A2(n_601), .B1(n_563), .B2(n_602), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_619), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_641), .Y(n_662) );
OR2x2_ASAP7_75t_L g663 ( .A(n_613), .B(n_585), .Y(n_663) );
NAND2xp33_ASAP7_75t_SL g664 ( .A(n_638), .B(n_617), .Y(n_664) );
OA22x2_ASAP7_75t_L g665 ( .A1(n_617), .A2(n_601), .B1(n_597), .B2(n_592), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_611), .B(n_596), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_633), .B(n_585), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_632), .B(n_578), .Y(n_668) );
BUFx8_ASAP7_75t_SL g669 ( .A(n_661), .Y(n_669) );
AOI22xp5_ASAP7_75t_L g670 ( .A1(n_664), .A2(n_645), .B1(n_635), .B2(n_628), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_651), .A2(n_644), .B(n_603), .Y(n_671) );
NAND2x1_ASAP7_75t_L g672 ( .A(n_659), .B(n_625), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_655), .A2(n_642), .B1(n_578), .B2(n_584), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_652), .B(n_584), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g675 ( .A1(n_660), .A2(n_631), .B(n_639), .C(n_597), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_665), .A2(n_600), .B1(n_602), .B2(n_604), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_SL g677 ( .A1(n_659), .A2(n_643), .B(n_604), .C(n_595), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_648), .Y(n_678) );
AOI211xp5_ASAP7_75t_L g679 ( .A1(n_660), .A2(n_637), .B(n_606), .C(n_595), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_650), .Y(n_680) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_649), .A2(n_606), .B1(n_562), .B2(n_45), .C(n_54), .Y(n_681) );
XNOR2xp5_ASAP7_75t_L g682 ( .A(n_657), .B(n_562), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_676), .B(n_647), .Y(n_683) );
OAI211xp5_ASAP7_75t_L g684 ( .A1(n_672), .A2(n_646), .B(n_658), .C(n_656), .Y(n_684) );
OAI211xp5_ASAP7_75t_L g685 ( .A1(n_670), .A2(n_662), .B(n_654), .C(n_653), .Y(n_685) );
BUFx2_ASAP7_75t_L g686 ( .A(n_669), .Y(n_686) );
NOR3xp33_ASAP7_75t_L g687 ( .A(n_674), .B(n_667), .C(n_668), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_671), .A2(n_666), .B1(n_663), .B2(n_60), .Y(n_688) );
OAI22x1_ASAP7_75t_L g689 ( .A1(n_682), .A2(n_37), .B1(n_44), .B2(n_62), .Y(n_689) );
AOI21xp33_ASAP7_75t_L g690 ( .A1(n_677), .A2(n_65), .B(n_66), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_687), .B(n_673), .Y(n_691) );
OR5x1_ASAP7_75t_L g692 ( .A(n_684), .B(n_679), .C(n_675), .D(n_681), .E(n_678), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_690), .B(n_680), .C(n_70), .Y(n_693) );
NOR2xp67_ASAP7_75t_L g694 ( .A(n_685), .B(n_67), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_691), .Y(n_695) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_694), .A2(n_683), .B1(n_688), .B2(n_686), .Y(n_696) );
OAI322xp33_ASAP7_75t_L g697 ( .A1(n_692), .A2(n_689), .A3(n_75), .B1(n_77), .B2(n_73), .C1(n_224), .C2(n_222), .Y(n_697) );
AO22x2_ASAP7_75t_L g698 ( .A1(n_695), .A2(n_693), .B1(n_243), .B2(n_279), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_696), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_699), .B(n_697), .C(n_243), .Y(n_700) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_700), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g702 ( .A1(n_701), .A2(n_698), .B1(n_279), .B2(n_220), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_702), .Y(n_703) );
AO21x2_ASAP7_75t_L g704 ( .A1(n_703), .A2(n_279), .B(n_220), .Y(n_704) );
endmodule