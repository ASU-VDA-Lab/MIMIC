module fake_jpeg_14084_n_143 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_143);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVxp67_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

BUFx10_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_2),
.B(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_29),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_60),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g60 ( 
.A1(n_42),
.A2(n_0),
.B(n_1),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_64),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_45),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_40),
.B1(n_49),
.B2(n_50),
.Y(n_69)
);

AO21x1_ASAP7_75t_L g93 ( 
.A1(n_69),
.A2(n_71),
.B(n_77),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_55),
.B1(n_54),
.B2(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_41),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_73),
.B(n_7),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_20),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_51),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_SL g82 ( 
.A(n_75),
.B(n_66),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_73),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_48),
.B1(n_53),
.B2(n_46),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_62),
.A2(n_48),
.B1(n_52),
.B2(n_56),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_56),
.B1(n_39),
.B2(n_4),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_80),
.B(n_82),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_81),
.B(n_85),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_67),
.A2(n_39),
.B1(n_2),
.B2(n_4),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_10),
.B(n_11),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_77),
.B(n_0),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_86),
.B(n_89),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_70),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_87),
.B(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_67),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_88),
.A2(n_93),
.B1(n_96),
.B2(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_5),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_78),
.B(n_6),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_91),
.Y(n_100)
);

INVxp67_ASAP7_75t_SL g92 ( 
.A(n_78),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_77),
.A2(n_8),
.B(n_9),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_12),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g95 ( 
.A1(n_68),
.A2(n_10),
.B(n_11),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_68),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_24),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_38),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_101),
.B(n_108),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_15),
.B1(n_19),
.B2(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_37),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_26),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_111),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_80),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_114),
.Y(n_117)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_92),
.Y(n_113)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_113),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_14),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_106),
.A2(n_36),
.B1(n_16),
.B2(n_18),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_118),
.A2(n_126),
.B1(n_107),
.B2(n_103),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_125),
.B(n_108),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_123),
.Y(n_130)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_98),
.Y(n_124)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

FAx1_ASAP7_75t_SL g125 ( 
.A(n_110),
.B(n_23),
.CI(n_27),
.CON(n_125),
.SN(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_127),
.B(n_128),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_112),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_102),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_130),
.A2(n_122),
.B1(n_120),
.B2(n_125),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_132),
.B(n_134),
.C(n_129),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_133),
.A2(n_122),
.B1(n_121),
.B2(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_137),
.A2(n_119),
.B1(n_99),
.B2(n_116),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_138),
.A2(n_100),
.B(n_115),
.Y(n_139)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_139),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_140),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_141),
.B(n_115),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_109),
.Y(n_143)
);


endmodule