module fake_jpeg_6020_n_55 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_55);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_55;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx8_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_1),
.B(n_3),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_17),
.A2(n_18),
.B1(n_16),
.B2(n_10),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_12),
.A2(n_0),
.B1(n_6),
.B2(n_7),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_14),
.A2(n_6),
.B1(n_7),
.B2(n_13),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_14),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_21),
.B(n_22),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_9),
.Y(n_22)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_25),
.B(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_26),
.B(n_27),
.Y(n_38)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_29),
.B(n_25),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g30 ( 
.A(n_17),
.B(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_18),
.B(n_23),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_33),
.B(n_25),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_35),
.A2(n_39),
.B1(n_37),
.B2(n_40),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_15),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_27),
.Y(n_41)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_30),
.B1(n_40),
.B2(n_33),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_45),
.B1(n_41),
.B2(n_44),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_46),
.B1(n_48),
.B2(n_42),
.Y(n_52)
);

FAx1_ASAP7_75t_SL g51 ( 
.A(n_49),
.B(n_42),
.CI(n_45),
.CON(n_51),
.SN(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_51),
.B(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_52),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_51),
.Y(n_55)
);


endmodule