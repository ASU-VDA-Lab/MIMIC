module fake_jpeg_13475_n_441 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx13_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_7),
.B(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx8_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx16f_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_3),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx12_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_16),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_48),
.Y(n_121)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_28),
.Y(n_49)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_50),
.Y(n_107)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_52),
.Y(n_112)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_54),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_23),
.B(n_8),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_55),
.B(n_56),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_22),
.B(n_16),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_19),
.Y(n_57)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_57),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_29),
.Y(n_60)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_60),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_61),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_23),
.B(n_15),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_62),
.B(n_72),
.Y(n_115)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx5_ASAP7_75t_L g120 ( 
.A(n_65),
.Y(n_120)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx5_ASAP7_75t_L g124 ( 
.A(n_66),
.Y(n_124)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_68),
.Y(n_127)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_69),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_70),
.Y(n_135)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_71),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_22),
.B(n_15),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_75),
.Y(n_114)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g98 ( 
.A(n_76),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_42),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_77),
.B(n_81),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_27),
.A2(n_14),
.B(n_12),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_78),
.B(n_11),
.Y(n_96)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_79),
.B(n_80),
.Y(n_134)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_82),
.B(n_86),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_25),
.B(n_45),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_83),
.B(n_84),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_27),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_85),
.B(n_88),
.Y(n_138)
);

BUFx5_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

CKINVDCx11_ASAP7_75t_R g95 ( 
.A(n_87),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_25),
.B(n_14),
.Y(n_88)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_18),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_90),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_24),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_24),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_91),
.B(n_30),
.Y(n_117)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_24),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_92),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_41),
.B1(n_26),
.B2(n_43),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_93),
.A2(n_140),
.B1(n_73),
.B2(n_75),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_96),
.B(n_136),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_51),
.A2(n_26),
.B1(n_18),
.B2(n_32),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_101),
.A2(n_143),
.B1(n_61),
.B2(n_79),
.Y(n_151)
);

O2A1O1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_53),
.A2(n_20),
.B(n_44),
.C(n_46),
.Y(n_102)
);

OA22x2_ASAP7_75t_L g164 ( 
.A1(n_102),
.A2(n_50),
.B1(n_46),
.B2(n_17),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_67),
.A2(n_26),
.B1(n_41),
.B2(n_45),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_129),
.B1(n_111),
.B2(n_119),
.Y(n_150)
);

NAND2xp33_ASAP7_75t_R g110 ( 
.A(n_66),
.B(n_21),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_110),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_41),
.B1(n_26),
.B2(n_20),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_111),
.A2(n_119),
.B1(n_38),
.B2(n_42),
.Y(n_171)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_52),
.A2(n_74),
.B1(n_58),
.B2(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_47),
.B(n_34),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_128),
.B(n_133),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_59),
.A2(n_41),
.B1(n_44),
.B2(n_43),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_47),
.B(n_34),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_48),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_60),
.A2(n_32),
.B1(n_39),
.B2(n_37),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_71),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_142),
.B(n_61),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_69),
.A2(n_32),
.B1(n_39),
.B2(n_37),
.Y(n_143)
);

OA22x2_ASAP7_75t_L g201 ( 
.A1(n_145),
.A2(n_156),
.B1(n_161),
.B2(n_164),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_148),
.Y(n_220)
);

INVx4_ASAP7_75t_L g149 ( 
.A(n_106),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_149),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_150),
.A2(n_162),
.B1(n_171),
.B2(n_175),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_97),
.Y(n_152)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_30),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_153),
.B(n_5),
.Y(n_230)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_105),
.Y(n_154)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g155 ( 
.A(n_97),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_89),
.B1(n_57),
.B2(n_76),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_157),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_159),
.B(n_181),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_0),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_160),
.B(n_170),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_134),
.A2(n_70),
.B1(n_65),
.B2(n_37),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_46),
.B1(n_17),
.B2(n_86),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_94),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_165),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_121),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_104),
.A2(n_17),
.B1(n_87),
.B2(n_38),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_166),
.A2(n_192),
.B1(n_193),
.B2(n_123),
.Y(n_216)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_167),
.Y(n_207)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_168),
.Y(n_215)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_116),
.Y(n_169)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_116),
.B(n_1),
.Y(n_170)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_118),
.Y(n_172)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_172),
.Y(n_229)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_121),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_173),
.Y(n_211)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_118),
.Y(n_174)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_174),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_96),
.A2(n_103),
.B1(n_115),
.B2(n_122),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_2),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_177),
.B(n_4),
.Y(n_203)
);

AND2x4_ASAP7_75t_SL g178 ( 
.A(n_131),
.B(n_38),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_178),
.B(n_179),
.C(n_182),
.Y(n_210)
);

XNOR2x1_ASAP7_75t_L g179 ( 
.A(n_95),
.B(n_42),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_180),
.Y(n_226)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_108),
.Y(n_181)
);

AND2x2_ASAP7_75t_SL g182 ( 
.A(n_125),
.B(n_2),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g183 ( 
.A1(n_135),
.A2(n_38),
.B1(n_42),
.B2(n_5),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_183),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_107),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_184),
.B(n_120),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_104),
.A2(n_38),
.B1(n_42),
.B2(n_11),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_185),
.A2(n_190),
.B1(n_126),
.B2(n_112),
.Y(n_232)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_188),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_113),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_123),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_114),
.A2(n_10),
.B1(n_4),
.B2(n_5),
.Y(n_190)
);

AND2x2_ASAP7_75t_SL g191 ( 
.A(n_125),
.B(n_2),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_191),
.B(n_135),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_102),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_114),
.A2(n_127),
.B1(n_130),
.B2(n_144),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_99),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_194),
.B(n_157),
.Y(n_239)
);

BUFx12_ASAP7_75t_L g195 ( 
.A(n_107),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_195),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_203),
.B(n_191),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_195),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_205),
.B(n_222),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_146),
.A2(n_136),
.B(n_124),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_209),
.A2(n_159),
.B(n_164),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_188),
.A2(n_99),
.B1(n_132),
.B2(n_113),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_214),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_216),
.A2(n_185),
.B1(n_190),
.B2(n_178),
.Y(n_257)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_217),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_170),
.B(n_142),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_236),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_178),
.B(n_191),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_147),
.B(n_132),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_221),
.B(n_233),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g222 ( 
.A(n_167),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_145),
.A2(n_130),
.B1(n_127),
.B2(n_139),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_224),
.A2(n_216),
.B1(n_196),
.B2(n_235),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g225 ( 
.A(n_192),
.B(n_124),
.Y(n_225)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_225),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_227),
.B(n_238),
.Y(n_274)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_171),
.A2(n_126),
.B1(n_112),
.B2(n_139),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_228),
.A2(n_232),
.B1(n_211),
.B2(n_225),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_230),
.B(n_238),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_186),
.B(n_10),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_177),
.B(n_144),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_195),
.Y(n_238)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_243),
.A2(n_248),
.B(n_217),
.Y(n_279)
);

OR2x2_ASAP7_75t_L g245 ( 
.A(n_210),
.B(n_179),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_245),
.A2(n_254),
.B(n_275),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_212),
.A2(n_160),
.B1(n_158),
.B2(n_193),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g308 ( 
.A1(n_246),
.A2(n_250),
.B1(n_256),
.B2(n_258),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_247),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_164),
.B(n_173),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_263),
.Y(n_281)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_237),
.Y(n_251)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_251),
.Y(n_289)
);

BUFx3_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

INVx13_ASAP7_75t_L g313 ( 
.A(n_252),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_210),
.B(n_182),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_198),
.C(n_205),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_221),
.A2(n_182),
.B(n_164),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_196),
.Y(n_255)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_255),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_225),
.B1(n_232),
.B2(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_257),
.A2(n_262),
.B1(n_269),
.B2(n_201),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_200),
.A2(n_180),
.B1(n_169),
.B2(n_174),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_226),
.Y(n_259)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_259),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_197),
.B(n_152),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_220),
.B(n_176),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_273),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_236),
.A2(n_168),
.B1(n_172),
.B2(n_154),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_266),
.B(n_270),
.Y(n_295)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_226),
.Y(n_268)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_268),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_224),
.A2(n_194),
.B1(n_149),
.B2(n_187),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_197),
.B(n_120),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_203),
.B(n_6),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_275),
.Y(n_299)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_207),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_272),
.B(n_235),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_220),
.B(n_189),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_274),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_219),
.B(n_6),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_213),
.B(n_7),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_277),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_201),
.A2(n_7),
.B1(n_208),
.B2(n_206),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_206),
.B(n_204),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g284 ( 
.A(n_278),
.B(n_263),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_279),
.A2(n_283),
.B(n_254),
.Y(n_322)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_247),
.B(n_230),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g333 ( 
.A1(n_282),
.A2(n_305),
.B(n_283),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_243),
.A2(n_204),
.B(n_239),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_287),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_285),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_261),
.B(n_233),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g290 ( 
.A1(n_257),
.A2(n_201),
.B1(n_207),
.B2(n_202),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_290),
.A2(n_292),
.B1(n_298),
.B2(n_303),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_267),
.A2(n_201),
.B1(n_215),
.B2(n_231),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_294),
.C(n_300),
.Y(n_324)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_253),
.B(n_223),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_260),
.B(n_223),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_297),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g297 ( 
.A(n_278),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_245),
.B(n_198),
.C(n_215),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_244),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_301),
.B(n_309),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_262),
.A2(n_201),
.B1(n_199),
.B2(n_229),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_304),
.B(n_240),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_199),
.B(n_229),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_267),
.A2(n_231),
.B1(n_199),
.B2(n_234),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_307),
.B(n_269),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_260),
.B(n_234),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_266),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_258),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_245),
.B(n_240),
.C(n_270),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_312),
.B(n_242),
.C(n_249),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_316),
.B(n_300),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_290),
.A2(n_277),
.B1(n_264),
.B2(n_256),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_318),
.A2(n_322),
.B(n_333),
.Y(n_359)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_280),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_320),
.Y(n_361)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_285),
.Y(n_321)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_321),
.Y(n_345)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_323),
.Y(n_343)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_291),
.Y(n_325)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_325),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_326),
.B(n_335),
.C(n_341),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_301),
.B(n_242),
.Y(n_327)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_327),
.Y(n_353)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_291),
.Y(n_328)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_328),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_308),
.A2(n_246),
.B1(n_241),
.B2(n_250),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_329),
.A2(n_337),
.B1(n_340),
.B2(n_303),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_331),
.Y(n_347)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_306),
.Y(n_332)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_332),
.Y(n_356)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_280),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_338),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_294),
.B(n_255),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_295),
.B(n_272),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_336),
.B(n_339),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_308),
.A2(n_241),
.B1(n_264),
.B2(n_276),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_288),
.B(n_252),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_306),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_302),
.A2(n_271),
.B1(n_259),
.B2(n_268),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_294),
.B(n_251),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g342 ( 
.A1(n_279),
.A2(n_305),
.B(n_286),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_342),
.B(n_292),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_330),
.A2(n_302),
.B1(n_312),
.B2(n_284),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_346),
.A2(n_329),
.B1(n_317),
.B2(n_321),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_330),
.B1(n_318),
.B2(n_336),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_327),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_SL g368 ( 
.A(n_349),
.B(n_357),
.Y(n_368)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_351),
.A2(n_364),
.B(n_339),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_324),
.B(n_293),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_354),
.B(n_363),
.C(n_341),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_320),
.B(n_288),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_334),
.B(n_287),
.Y(n_358)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_358),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_360),
.B(n_299),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_324),
.B(n_304),
.C(n_281),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_337),
.A2(n_298),
.B1(n_297),
.B2(n_309),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_365),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_319),
.B(n_296),
.Y(n_366)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_366),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_370),
.B(n_371),
.C(n_374),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_354),
.B(n_335),
.C(n_326),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g372 ( 
.A1(n_361),
.A2(n_345),
.B1(n_351),
.B2(n_343),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_372),
.A2(n_375),
.B1(n_379),
.B2(n_384),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_362),
.B(n_316),
.C(n_322),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_344),
.Y(n_376)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_376),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_346),
.B(n_314),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_377),
.B(n_380),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g396 ( 
.A1(n_378),
.A2(n_347),
.B1(n_361),
.B2(n_359),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_353),
.A2(n_317),
.B1(n_342),
.B2(n_333),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_359),
.A2(n_315),
.B(n_282),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_344),
.Y(n_381)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_381),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_362),
.B(n_282),
.C(n_281),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_360),
.C(n_353),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_385),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_343),
.A2(n_340),
.B1(n_323),
.B2(n_325),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_363),
.B(n_299),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_386),
.B(n_366),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_389),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_368),
.Y(n_389)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_384),
.Y(n_391)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_391),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_373),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_392),
.B(n_401),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_367),
.Y(n_395)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_395),
.B(n_390),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_396),
.A2(n_355),
.B1(n_328),
.B2(n_311),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g403 ( 
.A(n_399),
.B(n_402),
.Y(n_403)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_375),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g406 ( 
.A1(n_400),
.A2(n_385),
.B(n_348),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_369),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_370),
.B(n_364),
.Y(n_402)
);

AOI321xp33_ASAP7_75t_L g404 ( 
.A1(n_394),
.A2(n_380),
.A3(n_379),
.B1(n_350),
.B2(n_382),
.C(n_374),
.Y(n_404)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_404),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_405),
.B(n_408),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_406),
.Y(n_424)
);

AO221x1_ASAP7_75t_L g408 ( 
.A1(n_393),
.A2(n_356),
.B1(n_352),
.B2(n_332),
.C(n_311),
.Y(n_408)
);

OAI322xp33_ASAP7_75t_L g409 ( 
.A1(n_388),
.A2(n_383),
.A3(n_386),
.B1(n_371),
.B2(n_365),
.C1(n_356),
.C2(n_352),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g419 ( 
.A(n_409),
.B(n_414),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_410),
.B(n_411),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_355),
.C(n_289),
.Y(n_411)
);

OAI322xp33_ASAP7_75t_L g414 ( 
.A1(n_387),
.A2(n_289),
.A3(n_307),
.B1(n_313),
.B2(n_399),
.C1(n_398),
.C2(n_402),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_413),
.A2(n_400),
.B1(n_391),
.B2(n_397),
.Y(n_415)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_415),
.Y(n_427)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_407),
.A2(n_313),
.B1(n_398),
.B2(n_412),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_416),
.B(n_404),
.Y(n_425)
);

NOR2x1_ASAP7_75t_SL g418 ( 
.A(n_411),
.B(n_313),
.Y(n_418)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_418),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_410),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g431 ( 
.A(n_420),
.B(n_423),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_403),
.B(n_405),
.Y(n_423)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_425),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_422),
.B(n_417),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_426),
.B(n_428),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_415),
.B(n_420),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_424),
.A2(n_419),
.B(n_423),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_421),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_430),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_432),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_SL g436 ( 
.A1(n_434),
.A2(n_424),
.B(n_429),
.C(n_427),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_436),
.B(n_435),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_438),
.B(n_433),
.C(n_437),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_431),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_440),
.B(n_431),
.Y(n_441)
);


endmodule