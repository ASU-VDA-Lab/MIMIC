module fake_ariane_1781_n_1261 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1261);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1261;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_423;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_319;
wire n_690;
wire n_416;
wire n_1109;
wire n_525;
wire n_187;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_524;
wire n_634;
wire n_1214;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_232;
wire n_568;
wire n_1088;
wire n_766;
wire n_377;
wire n_520;
wire n_870;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1018;
wire n_259;
wire n_953;
wire n_1224;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_200;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_868;
wire n_884;
wire n_1034;
wire n_1085;
wire n_277;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_352;
wire n_206;
wire n_899;
wire n_611;
wire n_238;
wire n_365;
wire n_1013;
wire n_334;
wire n_192;
wire n_661;
wire n_300;
wire n_533;
wire n_438;
wire n_440;
wire n_273;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_461;
wire n_1121;
wire n_209;
wire n_490;
wire n_225;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_513;
wire n_288;
wire n_179;
wire n_1178;
wire n_1026;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_746;
wire n_292;
wire n_1079;
wire n_615;
wire n_1139;
wire n_517;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1101;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1220;
wire n_356;
wire n_698;
wire n_307;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_299;
wire n_836;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_370;
wire n_706;
wire n_286;
wire n_776;
wire n_424;
wire n_466;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_855;
wire n_808;
wire n_553;
wire n_814;
wire n_578;
wire n_405;
wire n_320;
wire n_1134;
wire n_647;
wire n_600;
wire n_481;
wire n_1053;
wire n_529;
wire n_502;
wire n_218;
wire n_247;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_545;
wire n_1015;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_233;
wire n_957;
wire n_388;
wire n_1242;
wire n_1218;
wire n_321;
wire n_221;
wire n_861;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_845;
wire n_888;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_769;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_999;
wire n_456;
wire n_852;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1243;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_317;
wire n_1257;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_687;
wire n_797;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_602;
wire n_592;
wire n_854;
wire n_393;
wire n_474;
wire n_805;
wire n_295;
wire n_190;
wire n_1072;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_752;
wire n_985;
wire n_421;
wire n_906;
wire n_1180;
wire n_283;
wire n_806;
wire n_649;
wire n_374;
wire n_643;
wire n_226;
wire n_682;
wire n_819;
wire n_586;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_818;
wire n_779;
wire n_594;
wire n_1052;
wire n_272;
wire n_833;
wire n_879;
wire n_1117;
wire n_422;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_224;
wire n_894;
wire n_420;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1128;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1065;
wire n_453;
wire n_810;
wire n_181;
wire n_617;
wire n_543;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_743;
wire n_1194;
wire n_907;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_284;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_613;
wire n_1022;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_820;
wire n_872;
wire n_254;
wire n_1157;
wire n_234;
wire n_848;
wire n_280;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_223;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_213;
wire n_1014;
wire n_724;
wire n_493;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1124;
wire n_932;
wire n_1183;
wire n_981;
wire n_1110;
wire n_243;
wire n_185;
wire n_1204;
wire n_994;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1057;
wire n_191;
wire n_978;
wire n_1011;
wire n_828;
wire n_322;
wire n_558;
wire n_653;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1167;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_244;
wire n_679;
wire n_220;
wire n_663;
wire n_443;
wire n_528;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_385;
wire n_917;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1064;
wire n_633;
wire n_900;
wire n_1093;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_835;
wire n_446;
wire n_1076;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_309;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_291;
wire n_822;
wire n_1094;
wire n_840;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_240;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_188;
wire n_323;
wire n_550;
wire n_997;
wire n_635;
wire n_694;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1236;
wire n_228;
wire n_671;
wire n_1148;
wire n_654;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_658;
wire n_630;
wire n_362;
wire n_310;
wire n_709;
wire n_809;
wire n_235;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_572;
wire n_1199;
wire n_865;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_196;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1229;
wire n_415;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_195;
wire n_938;
wire n_895;
wire n_304;
wire n_583;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_265;
wire n_208;
wire n_275;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_963;
wire n_1082;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1001;
wire n_1115;
wire n_1002;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_289;
wire n_548;
wire n_523;
wire n_457;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_675;

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_158),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_160),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_5),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_117),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_107),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_59),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_60),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_12),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_159),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_125),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_74),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_39),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_62),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_150),
.Y(n_197)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_139),
.Y(n_198)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_141),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_67),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_119),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_138),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_98),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_0),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_57),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_127),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_18),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_114),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_76),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_32),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_33),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_149),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_112),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_132),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_75),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_136),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_135),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_22),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_69),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g221 ( 
.A(n_3),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_84),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_99),
.Y(n_223)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_50),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_143),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_115),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_157),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_144),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_54),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_104),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_109),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_27),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_146),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_30),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_183),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_208),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_234),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_203),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_203),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_190),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_211),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g245 ( 
.A(n_179),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_225),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_212),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_236),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_181),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_185),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_189),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_191),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_192),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_193),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_194),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_197),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_225),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_200),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_180),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_219),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_182),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_184),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_195),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_250),
.Y(n_267)
);

INVxp67_ASAP7_75t_SL g268 ( 
.A(n_247),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_237),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_262),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_238),
.Y(n_271)
);

NOR2xp67_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_201),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_244),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_239),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_262),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g278 ( 
.A(n_243),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_247),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_252),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_264),
.Y(n_282)
);

INVx3_ASAP7_75t_L g283 ( 
.A(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_259),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_266),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_254),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_245),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_245),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_255),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_245),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_245),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_245),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_246),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_248),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_240),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_249),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_257),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_260),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_241),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_241),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_263),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_237),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_237),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_259),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_261),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_261),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_250),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_262),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_261),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_277),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_270),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_279),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_267),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_282),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_284),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_312),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_316),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_312),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_312),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_312),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_270),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_283),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_283),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_282),
.Y(n_334)
);

INVxp67_ASAP7_75t_SL g335 ( 
.A(n_268),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_313),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_314),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_281),
.Y(n_340)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_299),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_306),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_308),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_314),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g345 ( 
.A(n_283),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_281),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_317),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g350 ( 
.A(n_276),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_273),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_276),
.Y(n_352)
);

INVxp67_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_271),
.Y(n_354)
);

HB1xp67_ASAP7_75t_L g355 ( 
.A(n_305),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_275),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_286),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_286),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_288),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_308),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_285),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_288),
.Y(n_362)
);

INVxp67_ASAP7_75t_SL g363 ( 
.A(n_287),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_289),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_310),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_311),
.Y(n_366)
);

INVx5_ASAP7_75t_L g367 ( 
.A(n_352),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_364),
.B(n_290),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_292),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_293),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_352),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_326),
.B(n_280),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_291),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_342),
.B(n_291),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_325),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_351),
.B(n_300),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_320),
.B(n_294),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_332),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_335),
.B(n_296),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_332),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_350),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_333),
.Y(n_383)
);

BUFx8_ASAP7_75t_SL g384 ( 
.A(n_322),
.Y(n_384)
);

AND2x4_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_296),
.Y(n_385)
);

BUFx2_ASAP7_75t_L g386 ( 
.A(n_319),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g387 ( 
.A(n_361),
.B(n_300),
.Y(n_387)
);

AND2x4_ASAP7_75t_L g388 ( 
.A(n_323),
.B(n_297),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_361),
.B(n_303),
.Y(n_390)
);

INVx5_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_333),
.Y(n_392)
);

INVx5_ASAP7_75t_L g393 ( 
.A(n_329),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_334),
.B(n_295),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_336),
.B(n_302),
.Y(n_395)
);

HB1xp67_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_330),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_331),
.Y(n_398)
);

AND2x4_ASAP7_75t_L g399 ( 
.A(n_337),
.B(n_298),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_303),
.Y(n_400)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_222),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_339),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_344),
.B(n_347),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_324),
.Y(n_404)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_348),
.Y(n_405)
);

AND2x4_ASAP7_75t_L g406 ( 
.A(n_349),
.B(n_301),
.Y(n_406)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_324),
.Y(n_407)
);

BUFx3_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_375),
.Y(n_409)
);

AND2x4_ASAP7_75t_L g410 ( 
.A(n_387),
.B(n_390),
.Y(n_410)
);

OA21x2_ASAP7_75t_L g411 ( 
.A1(n_368),
.A2(n_224),
.B(n_222),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_373),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_379),
.B(n_315),
.Y(n_413)
);

BUFx2_ASAP7_75t_L g414 ( 
.A(n_386),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_378),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_387),
.A2(n_357),
.B1(n_346),
.B2(n_362),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_380),
.Y(n_417)
);

NAND2x1p5_ASAP7_75t_L g418 ( 
.A(n_367),
.B(n_356),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_378),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_375),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_380),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_380),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_383),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_383),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_383),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_384),
.Y(n_426)
);

OAI22x1_ASAP7_75t_R g427 ( 
.A1(n_386),
.A2(n_343),
.B1(n_360),
.B2(n_362),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_373),
.B(n_327),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_379),
.B(n_315),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_373),
.B(n_322),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_375),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_375),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_387),
.B(n_365),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_379),
.B(n_274),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_375),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_390),
.B(n_366),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_374),
.B(n_390),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_392),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_397),
.Y(n_442)
);

HB1xp67_ASAP7_75t_L g443 ( 
.A(n_374),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_379),
.B(n_304),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_397),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_403),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_397),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g448 ( 
.A1(n_404),
.A2(n_405),
.B1(n_407),
.B2(n_402),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_385),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g450 ( 
.A1(n_404),
.A2(n_359),
.B1(n_338),
.B2(n_357),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_400),
.A2(n_359),
.B1(n_346),
.B2(n_340),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_375),
.Y(n_453)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_407),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_385),
.Y(n_455)
);

INVx3_ASAP7_75t_L g456 ( 
.A(n_407),
.Y(n_456)
);

BUFx3_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

AND2x4_ASAP7_75t_L g458 ( 
.A(n_406),
.B(n_358),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_385),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_376),
.A2(n_340),
.B1(n_338),
.B2(n_219),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_272),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_385),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_395),
.B(n_355),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_385),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_405),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_395),
.B(n_307),
.Y(n_466)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_406),
.A2(n_309),
.B1(n_207),
.B2(n_227),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_407),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_396),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_375),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_388),
.B(n_227),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_388),
.B(n_204),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_381),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_405),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_405),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_408),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_406),
.B(n_221),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_408),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_388),
.B(n_186),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_406),
.A2(n_186),
.B1(n_196),
.B2(n_230),
.Y(n_483)
);

AOI22x1_ASAP7_75t_SL g484 ( 
.A1(n_396),
.A2(n_235),
.B1(n_233),
.B2(n_231),
.Y(n_484)
);

AND2x4_ASAP7_75t_L g485 ( 
.A(n_406),
.B(n_206),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_388),
.B(n_399),
.Y(n_486)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_398),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_381),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_407),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_407),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_371),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_371),
.Y(n_492)
);

AND2x2_ASAP7_75t_SL g493 ( 
.A(n_407),
.B(n_402),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_372),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_377),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_372),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_371),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_372),
.B(n_198),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_381),
.Y(n_499)
);

XNOR2x2_ASAP7_75t_L g500 ( 
.A(n_370),
.B(n_218),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_381),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_371),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_371),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_426),
.Y(n_504)
);

INVx3_ASAP7_75t_L g505 ( 
.A(n_409),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_426),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_417),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_474),
.Y(n_509)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_409),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_417),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_486),
.B(n_388),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_424),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_409),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_421),
.A2(n_369),
.B(n_368),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_424),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_469),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_474),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_425),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_425),
.Y(n_520)
);

NAND2xp33_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_404),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_435),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_435),
.Y(n_523)
);

CKINVDCx16_ASAP7_75t_R g524 ( 
.A(n_427),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_436),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_416),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_436),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_422),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_441),
.B(n_399),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_423),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_440),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_415),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_419),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_442),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_442),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_409),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_445),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_445),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_452),
.B(n_399),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_447),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_447),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_484),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_460),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_450),
.B(n_399),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_465),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_420),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_420),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_414),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_494),
.Y(n_549)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_487),
.Y(n_550)
);

AND2x2_ASAP7_75t_L g551 ( 
.A(n_486),
.B(n_399),
.Y(n_551)
);

CKINVDCx20_ASAP7_75t_R g552 ( 
.A(n_487),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_475),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_496),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_476),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_446),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_451),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_496),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_449),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_430),
.Y(n_560)
);

CKINVDCx5p33_ASAP7_75t_R g561 ( 
.A(n_457),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_455),
.Y(n_562)
);

BUFx6f_ASAP7_75t_L g563 ( 
.A(n_420),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_457),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_508),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_556),
.B(n_439),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_511),
.Y(n_567)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_517),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_511),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_508),
.Y(n_570)
);

NAND3xp33_ASAP7_75t_L g571 ( 
.A(n_539),
.B(n_463),
.C(n_466),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_550),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_513),
.Y(n_573)
);

NAND3xp33_ASAP7_75t_L g574 ( 
.A(n_544),
.B(n_467),
.C(n_429),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_519),
.Y(n_575)
);

AOI21x1_ASAP7_75t_L g576 ( 
.A1(n_515),
.A2(n_411),
.B(n_448),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_554),
.B(n_458),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_558),
.B(n_458),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_519),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_520),
.Y(n_580)
);

OR2x6_ASAP7_75t_L g581 ( 
.A(n_528),
.B(n_486),
.Y(n_581)
);

AO21x2_ASAP7_75t_L g582 ( 
.A1(n_528),
.A2(n_461),
.B(n_451),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_556),
.B(n_410),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_561),
.B(n_458),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_518),
.B(n_413),
.Y(n_585)
);

OR2x2_ASAP7_75t_L g586 ( 
.A(n_517),
.B(n_443),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_520),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_513),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_516),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_514),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_522),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_522),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_525),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_560),
.B(n_410),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_525),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_538),
.Y(n_597)
);

OAI22xp33_ASAP7_75t_SL g598 ( 
.A1(n_524),
.A2(n_471),
.B1(n_412),
.B2(n_434),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_564),
.B(n_493),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_549),
.B(n_443),
.Y(n_600)
);

INVxp33_ASAP7_75t_L g601 ( 
.A(n_506),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_538),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_523),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g604 ( 
.A1(n_571),
.A2(n_526),
.B1(n_543),
.B2(n_412),
.Y(n_604)
);

AND2x6_ASAP7_75t_L g605 ( 
.A(n_565),
.B(n_510),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_565),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_581),
.B(n_518),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_595),
.B(n_600),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_568),
.B(n_478),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_570),
.Y(n_610)
);

INVxp67_ASAP7_75t_L g611 ( 
.A(n_572),
.Y(n_611)
);

AND2x2_ASAP7_75t_L g612 ( 
.A(n_568),
.B(n_478),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_581),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_574),
.B(n_514),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_577),
.B(n_428),
.Y(n_615)
);

NOR2x1p5_ASAP7_75t_L g616 ( 
.A(n_586),
.B(n_504),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g617 ( 
.A(n_586),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_578),
.B(n_548),
.Y(n_618)
);

BUFx6f_ASAP7_75t_L g619 ( 
.A(n_581),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_581),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_570),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_573),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_573),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_581),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_588),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g626 ( 
.A(n_584),
.B(n_524),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_588),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_589),
.Y(n_628)
);

BUFx6f_ASAP7_75t_SL g629 ( 
.A(n_589),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_585),
.Y(n_630)
);

NAND3xp33_ASAP7_75t_L g631 ( 
.A(n_566),
.B(n_483),
.C(n_521),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_585),
.B(n_512),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_590),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_590),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_583),
.B(n_532),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_603),
.Y(n_636)
);

OR2x2_ASAP7_75t_L g637 ( 
.A(n_603),
.B(n_532),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_598),
.B(n_514),
.Y(n_638)
);

INVx5_ASAP7_75t_L g639 ( 
.A(n_591),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_591),
.Y(n_640)
);

OR2x6_ASAP7_75t_L g641 ( 
.A(n_599),
.B(n_530),
.Y(n_641)
);

NAND2xp33_ASAP7_75t_L g642 ( 
.A(n_591),
.B(n_529),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_591),
.Y(n_643)
);

INVx4_ASAP7_75t_L g644 ( 
.A(n_582),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_587),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_587),
.Y(n_646)
);

INVxp67_ASAP7_75t_SL g647 ( 
.A(n_567),
.Y(n_647)
);

AOI22xp33_ASAP7_75t_L g648 ( 
.A1(n_582),
.A2(n_500),
.B1(n_438),
.B2(n_433),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_567),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_601),
.B(n_552),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_567),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_582),
.Y(n_652)
);

INVx1_ASAP7_75t_SL g653 ( 
.A(n_569),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_569),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_576),
.B(n_507),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_SL g657 ( 
.A(n_575),
.B(n_514),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_576),
.B(n_542),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_575),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_575),
.B(n_433),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_579),
.B(n_514),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_579),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_579),
.B(n_509),
.Y(n_663)
);

INVx3_ASAP7_75t_L g664 ( 
.A(n_580),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_580),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_580),
.Y(n_666)
);

AOI22xp33_ASAP7_75t_L g667 ( 
.A1(n_592),
.A2(n_438),
.B1(n_485),
.B2(n_498),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_592),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_592),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_593),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_593),
.Y(n_671)
);

NOR2xp33_ASAP7_75t_L g672 ( 
.A(n_593),
.B(n_512),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_SL g673 ( 
.A(n_594),
.B(n_493),
.Y(n_673)
);

BUFx10_ASAP7_75t_L g674 ( 
.A(n_594),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_594),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_596),
.B(n_602),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_596),
.B(n_530),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_596),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_597),
.Y(n_679)
);

OR2x6_ASAP7_75t_L g680 ( 
.A(n_597),
.B(n_531),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_597),
.A2(n_485),
.B1(n_444),
.B2(n_472),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_602),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_551),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_571),
.B(n_533),
.Y(n_684)
);

BUFx10_ASAP7_75t_L g685 ( 
.A(n_585),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_565),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_571),
.B(n_533),
.Y(n_687)
);

NAND2x1p5_ASAP7_75t_L g688 ( 
.A(n_654),
.B(n_613),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_606),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_625),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_610),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_617),
.B(n_515),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_621),
.Y(n_693)
);

AND2x2_ASAP7_75t_L g694 ( 
.A(n_608),
.B(n_551),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_622),
.Y(n_695)
);

XOR2xp5_ASAP7_75t_L g696 ( 
.A(n_604),
.B(n_645),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_623),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_627),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_628),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_634),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_633),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_636),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_686),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_650),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_637),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_609),
.B(n_510),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_656),
.B(n_553),
.Y(n_707)
);

INVxp33_ASAP7_75t_SL g708 ( 
.A(n_618),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_646),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_649),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_651),
.Y(n_711)
);

INVxp67_ASAP7_75t_SL g712 ( 
.A(n_647),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_605),
.Y(n_713)
);

XNOR2x2_ASAP7_75t_L g714 ( 
.A(n_604),
.B(n_531),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_665),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_684),
.B(n_553),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_629),
.B(n_555),
.Y(n_717)
);

AND2x4_ASAP7_75t_L g718 ( 
.A(n_620),
.B(n_510),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_659),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_629),
.B(n_555),
.Y(n_720)
);

INVxp33_ASAP7_75t_L g721 ( 
.A(n_663),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_685),
.B(n_536),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_662),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_666),
.Y(n_724)
);

NAND2x1p5_ASAP7_75t_L g725 ( 
.A(n_654),
.B(n_510),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_620),
.B(n_505),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_668),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_669),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_685),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_679),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_671),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_615),
.B(n_505),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_612),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_616),
.B(n_505),
.Y(n_734)
);

XOR2xp5_ASAP7_75t_L g735 ( 
.A(n_632),
.B(n_559),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_675),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_678),
.Y(n_737)
);

INVxp33_ASAP7_75t_L g738 ( 
.A(n_626),
.Y(n_738)
);

XNOR2x2_ASAP7_75t_L g739 ( 
.A(n_658),
.B(n_559),
.Y(n_739)
);

XNOR2x2_ASAP7_75t_L g740 ( 
.A(n_631),
.B(n_562),
.Y(n_740)
);

XOR2xp5_ASAP7_75t_L g741 ( 
.A(n_632),
.B(n_562),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_676),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_611),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_676),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_677),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_677),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_677),
.Y(n_747)
);

INVx2_ASAP7_75t_SL g748 ( 
.A(n_630),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_687),
.B(n_547),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_680),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_680),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_682),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_680),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_687),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_672),
.B(n_547),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_664),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_664),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_624),
.B(n_547),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_670),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_631),
.B(n_545),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_670),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_635),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_653),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_653),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_655),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_655),
.Y(n_766)
);

CKINVDCx20_ASAP7_75t_R g767 ( 
.A(n_607),
.Y(n_767)
);

NOR2xp67_ASAP7_75t_L g768 ( 
.A(n_639),
.B(n_536),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_655),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_641),
.Y(n_770)
);

INVxp33_ASAP7_75t_SL g771 ( 
.A(n_683),
.Y(n_771)
);

OR2x6_ASAP7_75t_L g772 ( 
.A(n_613),
.B(n_557),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_641),
.Y(n_773)
);

NOR2xp67_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_536),
.Y(n_774)
);

OAI221xp5_ASAP7_75t_L g775 ( 
.A1(n_717),
.A2(n_648),
.B1(n_638),
.B2(n_667),
.C(n_614),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_689),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_754),
.B(n_644),
.Y(n_777)
);

INVxp67_ASAP7_75t_L g778 ( 
.A(n_707),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_716),
.B(n_644),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_714),
.A2(n_681),
.B1(n_673),
.B2(n_641),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_708),
.B(n_0),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_716),
.B(n_652),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_692),
.B(n_652),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_707),
.B(n_605),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_743),
.Y(n_785)
);

NOR2xp33_ASAP7_75t_L g786 ( 
.A(n_721),
.B(n_1),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_733),
.B(n_624),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_690),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_701),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_706),
.B(n_607),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_749),
.B(n_605),
.Y(n_791)
);

BUFx3_ASAP7_75t_L g792 ( 
.A(n_748),
.Y(n_792)
);

INVxp67_ASAP7_75t_SL g793 ( 
.A(n_712),
.Y(n_793)
);

NOR2xp33_ASAP7_75t_L g794 ( 
.A(n_704),
.B(n_1),
.Y(n_794)
);

BUFx5_ASAP7_75t_L g795 ( 
.A(n_765),
.Y(n_795)
);

AOI22xp5_ASAP7_75t_L g796 ( 
.A1(n_717),
.A2(n_720),
.B1(n_673),
.B2(n_760),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_771),
.B(n_2),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_749),
.B(n_605),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_705),
.B(n_762),
.Y(n_799)
);

NOR2xp33_ASAP7_75t_L g800 ( 
.A(n_738),
.B(n_2),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_694),
.B(n_607),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_692),
.B(n_640),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_691),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_702),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_729),
.B(n_639),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_742),
.B(n_640),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_715),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_744),
.B(n_643),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_693),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_760),
.B(n_660),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_L g811 ( 
.A(n_729),
.B(n_643),
.Y(n_811)
);

INVx3_ASAP7_75t_L g812 ( 
.A(n_729),
.Y(n_812)
);

NAND3xp33_ASAP7_75t_L g813 ( 
.A(n_720),
.B(n_642),
.C(n_657),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_734),
.B(n_732),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_713),
.B(n_643),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_695),
.B(n_619),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_696),
.A2(n_619),
.B1(n_545),
.B2(n_515),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_697),
.B(n_698),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_L g819 ( 
.A(n_713),
.B(n_536),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_767),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_699),
.Y(n_821)
);

INVxp67_ASAP7_75t_L g822 ( 
.A(n_732),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_700),
.B(n_619),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_703),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_710),
.B(n_661),
.Y(n_825)
);

INVx4_ASAP7_75t_L g826 ( 
.A(n_726),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_755),
.B(n_674),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_726),
.B(n_758),
.Y(n_828)
);

O2A1O1Ixp5_ASAP7_75t_L g829 ( 
.A1(n_770),
.A2(n_224),
.B(n_482),
.C(n_557),
.Y(n_829)
);

OR2x6_ASAP7_75t_L g830 ( 
.A(n_772),
.B(n_536),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_773),
.B(n_674),
.Y(n_831)
);

NAND2xp33_ASAP7_75t_L g832 ( 
.A(n_688),
.B(n_546),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_758),
.B(n_515),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_712),
.B(n_411),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_711),
.Y(n_835)
);

AND2x4_ASAP7_75t_L g836 ( 
.A(n_745),
.B(n_546),
.Y(n_836)
);

INVx2_ASAP7_75t_SL g837 ( 
.A(n_766),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_719),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_718),
.B(n_546),
.Y(n_839)
);

BUFx3_ASAP7_75t_L g840 ( 
.A(n_718),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_709),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_723),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_724),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_SL g844 ( 
.A(n_735),
.B(n_205),
.C(n_202),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_SL g845 ( 
.A(n_688),
.B(n_546),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_741),
.B(n_546),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_730),
.Y(n_847)
);

AND2x2_ASAP7_75t_L g848 ( 
.A(n_769),
.B(n_563),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_727),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_722),
.B(n_3),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_778),
.B(n_756),
.Y(n_851)
);

AO22x2_ASAP7_75t_L g852 ( 
.A1(n_817),
.A2(n_747),
.B1(n_750),
.B2(n_746),
.Y(n_852)
);

AOI22xp5_ASAP7_75t_L g853 ( 
.A1(n_796),
.A2(n_753),
.B1(n_751),
.B2(n_772),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_818),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_840),
.B(n_772),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_L g856 ( 
.A(n_822),
.B(n_757),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_779),
.B(n_759),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_789),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_804),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_788),
.Y(n_860)
);

BUFx8_ASAP7_75t_L g861 ( 
.A(n_785),
.Y(n_861)
);

NAND2x1p5_ASAP7_75t_L g862 ( 
.A(n_805),
.B(n_768),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_792),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_779),
.B(n_761),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_776),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_803),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_782),
.B(n_793),
.Y(n_867)
);

INVxp67_ASAP7_75t_L g868 ( 
.A(n_799),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_814),
.Y(n_869)
);

AO22x2_ASAP7_75t_L g870 ( 
.A1(n_817),
.A2(n_731),
.B1(n_736),
.B2(n_728),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_809),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_781),
.B(n_739),
.Y(n_872)
);

AO22x2_ASAP7_75t_L g873 ( 
.A1(n_824),
.A2(n_737),
.B1(n_764),
.B2(n_763),
.Y(n_873)
);

NAND2x1p5_ASAP7_75t_L g874 ( 
.A(n_812),
.B(n_774),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_821),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_835),
.Y(n_876)
);

AND2x4_ASAP7_75t_L g877 ( 
.A(n_826),
.B(n_752),
.Y(n_877)
);

OAI221xp5_ASAP7_75t_L g878 ( 
.A1(n_794),
.A2(n_800),
.B1(n_780),
.B2(n_775),
.C(n_786),
.Y(n_878)
);

OR2x6_ASAP7_75t_L g879 ( 
.A(n_830),
.B(n_725),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_812),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_784),
.B(n_725),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_838),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_842),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_847),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_782),
.B(n_740),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_843),
.Y(n_886)
);

BUFx6f_ASAP7_75t_L g887 ( 
.A(n_848),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_849),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_806),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_826),
.B(n_563),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_806),
.Y(n_891)
);

NOR3xp33_ASAP7_75t_L g892 ( 
.A(n_813),
.B(n_850),
.C(n_844),
.Y(n_892)
);

AO22x2_ASAP7_75t_L g893 ( 
.A1(n_807),
.A2(n_527),
.B1(n_534),
.B2(n_523),
.Y(n_893)
);

BUFx6f_ASAP7_75t_SL g894 ( 
.A(n_836),
.Y(n_894)
);

NAND3xp33_ASAP7_75t_SL g895 ( 
.A(n_797),
.B(n_210),
.C(n_209),
.Y(n_895)
);

AND2x4_ASAP7_75t_L g896 ( 
.A(n_787),
.B(n_563),
.Y(n_896)
);

AO22x2_ASAP7_75t_L g897 ( 
.A1(n_841),
.A2(n_541),
.B1(n_537),
.B2(n_535),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_802),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_802),
.B(n_4),
.Y(n_899)
);

AO22x2_ASAP7_75t_L g900 ( 
.A1(n_783),
.A2(n_541),
.B1(n_537),
.B2(n_535),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_825),
.Y(n_901)
);

AO22x2_ASAP7_75t_L g902 ( 
.A1(n_783),
.A2(n_540),
.B1(n_534),
.B2(n_527),
.Y(n_902)
);

AND2x4_ASAP7_75t_L g903 ( 
.A(n_790),
.B(n_563),
.Y(n_903)
);

AO22x2_ASAP7_75t_L g904 ( 
.A1(n_777),
.A2(n_540),
.B1(n_481),
.B2(n_480),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_808),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_777),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_837),
.Y(n_907)
);

NAND2x1p5_ASAP7_75t_L g908 ( 
.A(n_839),
.B(n_845),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_808),
.Y(n_909)
);

BUFx4f_ASAP7_75t_L g910 ( 
.A(n_830),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_791),
.B(n_563),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_816),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_823),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_810),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_833),
.Y(n_915)
);

INVxp67_ASAP7_75t_L g916 ( 
.A(n_828),
.Y(n_916)
);

OR2x6_ASAP7_75t_L g917 ( 
.A(n_830),
.B(n_420),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_827),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_801),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_846),
.A2(n_477),
.B1(n_459),
.B2(n_462),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_815),
.B(n_431),
.Y(n_921)
);

AO22x2_ASAP7_75t_L g922 ( 
.A1(n_798),
.A2(n_464),
.B1(n_402),
.B2(n_490),
.Y(n_922)
);

INVxp67_ASAP7_75t_L g923 ( 
.A(n_831),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_795),
.Y(n_924)
);

BUFx6f_ASAP7_75t_SL g925 ( 
.A(n_836),
.Y(n_925)
);

BUFx8_ASAP7_75t_L g926 ( 
.A(n_820),
.Y(n_926)
);

OR2x6_ASAP7_75t_SL g927 ( 
.A(n_834),
.B(n_213),
.Y(n_927)
);

AO22x2_ASAP7_75t_L g928 ( 
.A1(n_834),
.A2(n_402),
.B1(n_502),
.B2(n_497),
.Y(n_928)
);

INVxp33_ASAP7_75t_L g929 ( 
.A(n_811),
.Y(n_929)
);

HB1xp67_ASAP7_75t_L g930 ( 
.A(n_795),
.Y(n_930)
);

OAI21xp5_ASAP7_75t_L g931 ( 
.A1(n_872),
.A2(n_829),
.B(n_832),
.Y(n_931)
);

BUFx2_ASAP7_75t_SL g932 ( 
.A(n_863),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_917),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_906),
.B(n_795),
.Y(n_934)
);

HB1xp67_ASAP7_75t_L g935 ( 
.A(n_898),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_885),
.A2(n_819),
.B(n_411),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_873),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_870),
.A2(n_795),
.B(n_492),
.Y(n_938)
);

NAND2xp33_ASAP7_75t_L g939 ( 
.A(n_892),
.B(n_795),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_889),
.B(n_891),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_926),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_907),
.B(n_4),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_929),
.B(n_431),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_878),
.A2(n_188),
.B1(n_215),
.B2(n_216),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_SL g945 ( 
.A(n_914),
.B(n_905),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_917),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_869),
.B(n_5),
.Y(n_947)
);

INVxp67_ASAP7_75t_L g948 ( 
.A(n_907),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_870),
.A2(n_492),
.B(n_491),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_861),
.Y(n_950)
);

BUFx4f_ASAP7_75t_L g951 ( 
.A(n_862),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_873),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_867),
.B(n_431),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_928),
.A2(n_497),
.B(n_491),
.Y(n_954)
);

AOI22xp5_ASAP7_75t_L g955 ( 
.A1(n_853),
.A2(n_401),
.B1(n_468),
.B2(n_456),
.Y(n_955)
);

OAI22xp5_ASAP7_75t_L g956 ( 
.A1(n_927),
.A2(n_454),
.B1(n_456),
.B2(n_468),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_909),
.B(n_6),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_915),
.B(n_6),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_858),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_928),
.A2(n_503),
.B(n_502),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_854),
.B(n_7),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_923),
.B(n_431),
.Y(n_962)
);

OAI22xp5_ASAP7_75t_L g963 ( 
.A1(n_899),
.A2(n_454),
.B1(n_489),
.B2(n_499),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_922),
.A2(n_503),
.B(n_489),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_887),
.B(n_7),
.Y(n_965)
);

INVx4_ASAP7_75t_L g966 ( 
.A(n_880),
.Y(n_966)
);

OAI21xp5_ASAP7_75t_L g967 ( 
.A1(n_895),
.A2(n_418),
.B(n_401),
.Y(n_967)
);

AND2x2_ASAP7_75t_L g968 ( 
.A(n_887),
.B(n_8),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_922),
.A2(n_437),
.B(n_432),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_904),
.A2(n_437),
.B(n_432),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_868),
.B(n_8),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_877),
.Y(n_972)
);

NOR2xp33_ASAP7_75t_L g973 ( 
.A(n_918),
.B(n_9),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_865),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_859),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_904),
.A2(n_437),
.B(n_432),
.Y(n_976)
);

BUFx4f_ASAP7_75t_L g977 ( 
.A(n_874),
.Y(n_977)
);

OAI21xp5_ASAP7_75t_L g978 ( 
.A1(n_856),
.A2(n_418),
.B(n_401),
.Y(n_978)
);

INVx5_ASAP7_75t_L g979 ( 
.A(n_879),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_910),
.A2(n_188),
.B(n_216),
.C(n_215),
.Y(n_980)
);

AOI22xp5_ASAP7_75t_L g981 ( 
.A1(n_900),
.A2(n_401),
.B1(n_215),
.B2(n_216),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_908),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_900),
.A2(n_437),
.B(n_432),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_866),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_857),
.B(n_9),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_864),
.B(n_453),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_935),
.B(n_940),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_985),
.B(n_851),
.Y(n_988)
);

NOR3xp33_ASAP7_75t_SL g989 ( 
.A(n_956),
.B(n_881),
.C(n_911),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_974),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_957),
.B(n_901),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_R g992 ( 
.A(n_950),
.B(n_871),
.Y(n_992)
);

BUFx4f_ASAP7_75t_L g993 ( 
.A(n_942),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_941),
.Y(n_994)
);

BUFx2_ASAP7_75t_L g995 ( 
.A(n_948),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_982),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_965),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_958),
.B(n_875),
.Y(n_998)
);

INVx2_ASAP7_75t_L g999 ( 
.A(n_937),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_984),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_982),
.Y(n_1001)
);

BUFx2_ASAP7_75t_L g1002 ( 
.A(n_951),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_945),
.B(n_876),
.Y(n_1003)
);

OR2x2_ASAP7_75t_L g1004 ( 
.A(n_952),
.B(n_916),
.Y(n_1004)
);

NOR3xp33_ASAP7_75t_SL g1005 ( 
.A(n_973),
.B(n_924),
.C(n_883),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_961),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_968),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_939),
.A2(n_902),
.B(n_852),
.Y(n_1008)
);

INVx6_ASAP7_75t_L g1009 ( 
.A(n_979),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_SL g1010 ( 
.A(n_951),
.B(n_912),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_944),
.A2(n_902),
.B1(n_852),
.B2(n_893),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_966),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_971),
.B(n_882),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_959),
.Y(n_1014)
);

INVx5_ASAP7_75t_L g1015 ( 
.A(n_933),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_SL g1016 ( 
.A(n_966),
.B(n_930),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_934),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_R g1018 ( 
.A(n_977),
.B(n_886),
.Y(n_1018)
);

OR2x6_ASAP7_75t_L g1019 ( 
.A(n_932),
.B(n_931),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_947),
.B(n_888),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_975),
.Y(n_1021)
);

NOR3xp33_ASAP7_75t_SL g1022 ( 
.A(n_963),
.B(n_913),
.C(n_919),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_933),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_979),
.B(n_855),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_953),
.B(n_893),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_970),
.B(n_920),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_986),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_972),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_972),
.Y(n_1029)
);

OAI22xp5_ASAP7_75t_L g1030 ( 
.A1(n_977),
.A2(n_879),
.B1(n_921),
.B2(n_896),
.Y(n_1030)
);

NOR3xp33_ASAP7_75t_SL g1031 ( 
.A(n_962),
.B(n_217),
.C(n_214),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_L g1032 ( 
.A(n_976),
.B(n_983),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_943),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_938),
.B(n_897),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_979),
.B(n_903),
.Y(n_1035)
);

AND2x2_ASAP7_75t_L g1036 ( 
.A(n_933),
.B(n_890),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_SL g1037 ( 
.A(n_969),
.B(n_223),
.C(n_220),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_SL g1038 ( 
.A(n_946),
.Y(n_1038)
);

OR2x2_ASAP7_75t_SL g1039 ( 
.A(n_946),
.B(n_860),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_946),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_981),
.Y(n_1041)
);

NOR3xp33_ASAP7_75t_SL g1042 ( 
.A(n_978),
.B(n_228),
.C(n_226),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_L g1043 ( 
.A(n_936),
.B(n_897),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_949),
.B(n_884),
.Y(n_1044)
);

HB1xp67_ASAP7_75t_L g1045 ( 
.A(n_964),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_944),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_954),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_960),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_955),
.B(n_894),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_980),
.B(n_925),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_967),
.B(n_10),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_940),
.Y(n_1052)
);

AOI33xp33_ASAP7_75t_L g1053 ( 
.A1(n_1006),
.A2(n_10),
.A3(n_11),
.B1(n_12),
.B2(n_13),
.B3(n_14),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_1052),
.B(n_11),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_R g1055 ( 
.A(n_994),
.B(n_13),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_987),
.B(n_14),
.Y(n_1056)
);

BUFx2_ASAP7_75t_SL g1057 ( 
.A(n_1002),
.Y(n_1057)
);

A2O1A1Ixp33_ASAP7_75t_L g1058 ( 
.A1(n_1008),
.A2(n_188),
.B(n_215),
.C(n_216),
.Y(n_1058)
);

OR2x6_ASAP7_75t_L g1059 ( 
.A(n_1009),
.B(n_501),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_990),
.B(n_15),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_1019),
.A2(n_215),
.B(n_188),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_1005),
.A2(n_188),
.B(n_216),
.C(n_229),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_1019),
.A2(n_470),
.B(n_453),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_1000),
.B(n_15),
.Y(n_1064)
);

BUFx6f_ASAP7_75t_L g1065 ( 
.A(n_1023),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_1039),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_1011),
.A2(n_16),
.B(n_17),
.C(n_18),
.Y(n_1067)
);

AOI221xp5_ASAP7_75t_L g1068 ( 
.A1(n_1043),
.A2(n_16),
.B1(n_17),
.B2(n_19),
.C(n_20),
.Y(n_1068)
);

NOR2xp33_ASAP7_75t_L g1069 ( 
.A(n_993),
.B(n_19),
.Y(n_1069)
);

BUFx2_ASAP7_75t_L g1070 ( 
.A(n_992),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_1001),
.B(n_20),
.Y(n_1071)
);

INVx4_ASAP7_75t_L g1072 ( 
.A(n_996),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_997),
.Y(n_1073)
);

INVxp67_ASAP7_75t_L g1074 ( 
.A(n_1038),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_1062),
.A2(n_1067),
.B(n_1058),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_1068),
.A2(n_1026),
.B1(n_1041),
.B2(n_1046),
.Y(n_1076)
);

AND2x4_ASAP7_75t_L g1077 ( 
.A(n_1070),
.B(n_996),
.Y(n_1077)
);

OAI321xp33_ASAP7_75t_L g1078 ( 
.A1(n_1069),
.A2(n_1051),
.A3(n_1034),
.B1(n_1032),
.B2(n_1050),
.C(n_1047),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_1061),
.A2(n_993),
.B(n_1045),
.Y(n_1079)
);

AOI21xp5_ASAP7_75t_L g1080 ( 
.A1(n_1056),
.A2(n_1025),
.B(n_1020),
.Y(n_1080)
);

BUFx4f_ASAP7_75t_SL g1081 ( 
.A(n_1073),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_1071),
.Y(n_1082)
);

OAI22xp33_ASAP7_75t_L g1083 ( 
.A1(n_1066),
.A2(n_1048),
.B1(n_1009),
.B2(n_1015),
.Y(n_1083)
);

OAI22xp5_ASAP7_75t_L g1084 ( 
.A1(n_1054),
.A2(n_1022),
.B1(n_989),
.B2(n_1013),
.Y(n_1084)
);

INVx2_ASAP7_75t_SL g1085 ( 
.A(n_1071),
.Y(n_1085)
);

BUFx4f_ASAP7_75t_L g1086 ( 
.A(n_1065),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_1065),
.B(n_1018),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1065),
.Y(n_1088)
);

BUFx6f_ASAP7_75t_L g1089 ( 
.A(n_1060),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_1055),
.A2(n_999),
.B1(n_1004),
.B2(n_1049),
.Y(n_1090)
);

INVx3_ASAP7_75t_L g1091 ( 
.A(n_1072),
.Y(n_1091)
);

AOI22xp33_ASAP7_75t_SL g1092 ( 
.A1(n_1057),
.A2(n_1007),
.B1(n_1038),
.B2(n_1049),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_1072),
.B(n_1015),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_1074),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1064),
.B(n_995),
.Y(n_1095)
);

BUFx6f_ASAP7_75t_L g1096 ( 
.A(n_1059),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1053),
.Y(n_1097)
);

CKINVDCx11_ASAP7_75t_R g1098 ( 
.A(n_1059),
.Y(n_1098)
);

INVx3_ASAP7_75t_L g1099 ( 
.A(n_1063),
.Y(n_1099)
);

AO21x2_ASAP7_75t_L g1100 ( 
.A1(n_1058),
.A2(n_998),
.B(n_991),
.Y(n_1100)
);

BUFx2_ASAP7_75t_SL g1101 ( 
.A(n_1077),
.Y(n_1101)
);

AOI21x1_ASAP7_75t_L g1102 ( 
.A1(n_1093),
.A2(n_1028),
.B(n_1029),
.Y(n_1102)
);

AOI21x1_ASAP7_75t_L g1103 ( 
.A1(n_1094),
.A2(n_1010),
.B(n_1033),
.Y(n_1103)
);

INVx3_ASAP7_75t_L g1104 ( 
.A(n_1082),
.Y(n_1104)
);

A2O1A1Ixp33_ASAP7_75t_L g1105 ( 
.A1(n_1080),
.A2(n_1037),
.B(n_988),
.C(n_1042),
.Y(n_1105)
);

A2O1A1Ixp33_ASAP7_75t_L g1106 ( 
.A1(n_1080),
.A2(n_1031),
.B(n_1016),
.C(n_1024),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_1089),
.Y(n_1107)
);

NAND2xp33_ASAP7_75t_L g1108 ( 
.A(n_1106),
.B(n_1085),
.Y(n_1108)
);

NAND2x1p5_ASAP7_75t_L g1109 ( 
.A(n_1104),
.B(n_1086),
.Y(n_1109)
);

OAI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_1108),
.A2(n_1079),
.B(n_1103),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_1109),
.B(n_1107),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_1111),
.B(n_1081),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1110),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1112),
.Y(n_1114)
);

CKINVDCx8_ASAP7_75t_R g1115 ( 
.A(n_1113),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_L g1116 ( 
.A1(n_1114),
.A2(n_1100),
.B1(n_1099),
.B2(n_1089),
.Y(n_1116)
);

BUFx2_ASAP7_75t_L g1117 ( 
.A(n_1115),
.Y(n_1117)
);

AND2x4_ASAP7_75t_L g1118 ( 
.A(n_1117),
.B(n_1104),
.Y(n_1118)
);

AND2x4_ASAP7_75t_L g1119 ( 
.A(n_1116),
.B(n_1077),
.Y(n_1119)
);

OR2x2_ASAP7_75t_SL g1120 ( 
.A(n_1117),
.B(n_1089),
.Y(n_1120)
);

INVxp67_ASAP7_75t_L g1121 ( 
.A(n_1118),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_1120),
.Y(n_1122)
);

AND2x4_ASAP7_75t_L g1123 ( 
.A(n_1119),
.B(n_1091),
.Y(n_1123)
);

NAND2x1_ASAP7_75t_L g1124 ( 
.A(n_1123),
.B(n_1091),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1121),
.B(n_1101),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1125),
.A2(n_1122),
.B1(n_1123),
.B2(n_1100),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1124),
.Y(n_1127)
);

NAND3xp33_ASAP7_75t_L g1128 ( 
.A(n_1127),
.B(n_1079),
.C(n_1105),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1126),
.B(n_1097),
.Y(n_1129)
);

AOI33xp33_ASAP7_75t_L g1130 ( 
.A1(n_1128),
.A2(n_1092),
.A3(n_1083),
.B1(n_1088),
.B2(n_1090),
.B3(n_1076),
.Y(n_1130)
);

AOI22xp33_ASAP7_75t_L g1131 ( 
.A1(n_1129),
.A2(n_1099),
.B1(n_1086),
.B2(n_1096),
.Y(n_1131)
);

NOR2x1_ASAP7_75t_L g1132 ( 
.A(n_1131),
.B(n_1087),
.Y(n_1132)
);

AND2x2_ASAP7_75t_SL g1133 ( 
.A(n_1130),
.B(n_1095),
.Y(n_1133)
);

NAND4xp25_ASAP7_75t_L g1134 ( 
.A(n_1132),
.B(n_1075),
.C(n_1095),
.D(n_1084),
.Y(n_1134)
);

INVx2_ASAP7_75t_SL g1135 ( 
.A(n_1133),
.Y(n_1135)
);

AOI32xp33_ASAP7_75t_L g1136 ( 
.A1(n_1135),
.A2(n_1084),
.A3(n_1078),
.B1(n_1102),
.B2(n_1098),
.Y(n_1136)
);

AND2x2_ASAP7_75t_L g1137 ( 
.A(n_1134),
.B(n_1096),
.Y(n_1137)
);

OR2x2_ASAP7_75t_L g1138 ( 
.A(n_1134),
.B(n_1096),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1137),
.B(n_1040),
.Y(n_1139)
);

NOR2xp33_ASAP7_75t_SL g1140 ( 
.A(n_1138),
.B(n_1015),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_1136),
.B(n_1040),
.Y(n_1141)
);

INVxp67_ASAP7_75t_L g1142 ( 
.A(n_1140),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_1139),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_L g1144 ( 
.A(n_1143),
.B(n_1141),
.Y(n_1144)
);

NAND4xp25_ASAP7_75t_SL g1145 ( 
.A(n_1142),
.B(n_1078),
.C(n_22),
.D(n_23),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1144),
.B(n_21),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_1145),
.B(n_21),
.Y(n_1147)
);

OAI221xp5_ASAP7_75t_L g1148 ( 
.A1(n_1147),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.C(n_26),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_1146),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1149),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1148),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_1150),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1151),
.B(n_24),
.Y(n_1153)
);

NAND2xp5_ASAP7_75t_L g1154 ( 
.A(n_1152),
.B(n_1153),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1152),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1152),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_1155),
.Y(n_1157)
);

OAI31xp33_ASAP7_75t_L g1158 ( 
.A1(n_1156),
.A2(n_25),
.A3(n_26),
.B(n_27),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_1154),
.Y(n_1159)
);

AND2x2_ASAP7_75t_L g1160 ( 
.A(n_1157),
.B(n_1023),
.Y(n_1160)
);

OR2x2_ASAP7_75t_L g1161 ( 
.A(n_1159),
.B(n_28),
.Y(n_1161)
);

OA21x2_ASAP7_75t_L g1162 ( 
.A1(n_1160),
.A2(n_1161),
.B(n_1158),
.Y(n_1162)
);

BUFx2_ASAP7_75t_L g1163 ( 
.A(n_1160),
.Y(n_1163)
);

A2O1A1Ixp33_ASAP7_75t_L g1164 ( 
.A1(n_1163),
.A2(n_1162),
.B(n_29),
.C(n_30),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1163),
.A2(n_28),
.B(n_29),
.C(n_31),
.Y(n_1165)
);

NOR3xp33_ASAP7_75t_L g1166 ( 
.A(n_1164),
.B(n_31),
.C(n_32),
.Y(n_1166)
);

OR2x2_ASAP7_75t_L g1167 ( 
.A(n_1165),
.B(n_33),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1167),
.A2(n_34),
.B(n_35),
.Y(n_1168)
);

OAI21xp33_ASAP7_75t_SL g1169 ( 
.A1(n_1166),
.A2(n_34),
.B(n_35),
.Y(n_1169)
);

NAND4xp25_ASAP7_75t_SL g1170 ( 
.A(n_1168),
.B(n_36),
.C(n_37),
.D(n_38),
.Y(n_1170)
);

INVxp67_ASAP7_75t_SL g1171 ( 
.A(n_1169),
.Y(n_1171)
);

AOI221x1_ASAP7_75t_L g1172 ( 
.A1(n_1171),
.A2(n_1023),
.B1(n_1012),
.B2(n_1024),
.C(n_370),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1170),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1171),
.Y(n_1174)
);

NAND4xp25_ASAP7_75t_L g1175 ( 
.A(n_1174),
.B(n_1012),
.C(n_41),
.D(n_42),
.Y(n_1175)
);

NAND4xp75_ASAP7_75t_L g1176 ( 
.A(n_1173),
.B(n_394),
.C(n_377),
.D(n_44),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1172),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_R g1178 ( 
.A(n_1177),
.B(n_40),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1175),
.A2(n_394),
.B(n_369),
.Y(n_1179)
);

NOR3x1_ASAP7_75t_L g1180 ( 
.A(n_1178),
.B(n_1176),
.C(n_1030),
.Y(n_1180)
);

NOR3x1_ASAP7_75t_L g1181 ( 
.A(n_1179),
.B(n_1017),
.C(n_1003),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1180),
.A2(n_1181),
.B1(n_1036),
.B2(n_1035),
.Y(n_1182)
);

NOR2x1_ASAP7_75t_L g1183 ( 
.A(n_1181),
.B(n_1021),
.Y(n_1183)
);

OAI21xp33_ASAP7_75t_SL g1184 ( 
.A1(n_1182),
.A2(n_1027),
.B(n_1014),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1183),
.A2(n_1035),
.B(n_45),
.Y(n_1185)
);

NAND2xp33_ASAP7_75t_SL g1186 ( 
.A(n_1184),
.B(n_43),
.Y(n_1186)
);

NAND3xp33_ASAP7_75t_L g1187 ( 
.A(n_1185),
.B(n_46),
.C(n_47),
.Y(n_1187)
);

INVx1_ASAP7_75t_SL g1188 ( 
.A(n_1186),
.Y(n_1188)
);

BUFx2_ASAP7_75t_L g1189 ( 
.A(n_1187),
.Y(n_1189)
);

INVx2_ASAP7_75t_L g1190 ( 
.A(n_1189),
.Y(n_1190)
);

NAND3xp33_ASAP7_75t_SL g1191 ( 
.A(n_1188),
.B(n_48),
.C(n_49),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1188),
.Y(n_1192)
);

OAI211xp5_ASAP7_75t_SL g1193 ( 
.A1(n_1190),
.A2(n_51),
.B(n_52),
.C(n_53),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1192),
.Y(n_1194)
);

NAND3xp33_ASAP7_75t_L g1195 ( 
.A(n_1191),
.B(n_55),
.C(n_56),
.Y(n_1195)
);

AOI22x1_ASAP7_75t_L g1196 ( 
.A1(n_1194),
.A2(n_58),
.B1(n_61),
.B2(n_63),
.Y(n_1196)
);

AOI22x1_ASAP7_75t_L g1197 ( 
.A1(n_1193),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1197),
.B(n_1195),
.Y(n_1198)
);

OAI22x1_ASAP7_75t_L g1199 ( 
.A1(n_1196),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1198),
.Y(n_1200)
);

HB1xp67_ASAP7_75t_L g1201 ( 
.A(n_1199),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1200),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_1201),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1203),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1202),
.Y(n_1205)
);

INVx2_ASAP7_75t_L g1206 ( 
.A(n_1204),
.Y(n_1206)
);

OR2x6_ASAP7_75t_L g1207 ( 
.A(n_1205),
.B(n_72),
.Y(n_1207)
);

NOR2x1_ASAP7_75t_L g1208 ( 
.A(n_1206),
.B(n_73),
.Y(n_1208)
);

INVx2_ASAP7_75t_SL g1209 ( 
.A(n_1207),
.Y(n_1209)
);

BUFx2_ASAP7_75t_L g1210 ( 
.A(n_1206),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_SL g1211 ( 
.A1(n_1210),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_1211)
);

OAI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1209),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_1212)
);

OAI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1208),
.A2(n_83),
.B1(n_85),
.B2(n_86),
.Y(n_1213)
);

OR3x1_ASAP7_75t_L g1214 ( 
.A(n_1212),
.B(n_87),
.C(n_88),
.Y(n_1214)
);

O2A1O1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1213),
.A2(n_89),
.B(n_90),
.C(n_92),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1214),
.B(n_1215),
.Y(n_1216)
);

XNOR2xp5_ASAP7_75t_L g1217 ( 
.A(n_1214),
.B(n_1211),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1215),
.A2(n_93),
.B(n_94),
.Y(n_1218)
);

OAI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1217),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_1219)
);

OAI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1216),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_1220)
);

AOI22xp5_ASAP7_75t_SL g1221 ( 
.A1(n_1218),
.A2(n_103),
.B1(n_105),
.B2(n_106),
.Y(n_1221)
);

NOR2xp67_ASAP7_75t_L g1222 ( 
.A(n_1219),
.B(n_108),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_1220),
.B(n_110),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1221),
.A2(n_111),
.B(n_113),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1224),
.B(n_116),
.Y(n_1225)
);

NOR2xp33_ASAP7_75t_L g1226 ( 
.A(n_1222),
.B(n_120),
.Y(n_1226)
);

AOI21xp33_ASAP7_75t_SL g1227 ( 
.A1(n_1223),
.A2(n_122),
.B(n_123),
.Y(n_1227)
);

OAI21xp33_ASAP7_75t_L g1228 ( 
.A1(n_1224),
.A2(n_126),
.B(n_128),
.Y(n_1228)
);

OAI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1224),
.A2(n_129),
.B(n_130),
.Y(n_1229)
);

OA21x2_ASAP7_75t_L g1230 ( 
.A1(n_1224),
.A2(n_131),
.B(n_134),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1224),
.B(n_137),
.Y(n_1231)
);

OAI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1224),
.A2(n_140),
.B(n_142),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_1224),
.A2(n_145),
.B(n_147),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1224),
.Y(n_1234)
);

AND2x2_ASAP7_75t_L g1235 ( 
.A(n_1224),
.B(n_148),
.Y(n_1235)
);

NAND2xp5_ASAP7_75t_L g1236 ( 
.A(n_1224),
.B(n_151),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1224),
.B(n_152),
.Y(n_1237)
);

AOI22xp5_ASAP7_75t_L g1238 ( 
.A1(n_1234),
.A2(n_1229),
.B1(n_1232),
.B2(n_1227),
.Y(n_1238)
);

AOI222xp33_ASAP7_75t_L g1239 ( 
.A1(n_1228),
.A2(n_153),
.B1(n_154),
.B2(n_155),
.C1(n_156),
.C2(n_161),
.Y(n_1239)
);

AOI222xp33_ASAP7_75t_L g1240 ( 
.A1(n_1225),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.C1(n_165),
.C2(n_166),
.Y(n_1240)
);

AOI322xp5_ASAP7_75t_L g1241 ( 
.A1(n_1231),
.A2(n_167),
.A3(n_168),
.B1(n_169),
.B2(n_171),
.C1(n_172),
.C2(n_174),
.Y(n_1241)
);

AOI222xp33_ASAP7_75t_L g1242 ( 
.A1(n_1236),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.C1(n_1044),
.C2(n_401),
.Y(n_1242)
);

AOI322xp5_ASAP7_75t_L g1243 ( 
.A1(n_1237),
.A2(n_401),
.A3(n_499),
.B1(n_488),
.B2(n_479),
.C1(n_501),
.C2(n_470),
.Y(n_1243)
);

AOI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1235),
.A2(n_401),
.B1(n_499),
.B2(n_488),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1226),
.A2(n_401),
.B1(n_501),
.B2(n_488),
.Y(n_1245)
);

AOI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1233),
.A2(n_1230),
.B1(n_401),
.B2(n_499),
.Y(n_1246)
);

AO21x2_ASAP7_75t_L g1247 ( 
.A1(n_1238),
.A2(n_1230),
.B(n_501),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1239),
.A2(n_488),
.B(n_479),
.Y(n_1248)
);

OAI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1240),
.A2(n_1241),
.B(n_1242),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1244),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1245),
.A2(n_479),
.B(n_473),
.Y(n_1251)
);

AOI22x1_ASAP7_75t_L g1252 ( 
.A1(n_1246),
.A2(n_479),
.B1(n_473),
.B2(n_470),
.Y(n_1252)
);

AOI22x1_ASAP7_75t_L g1253 ( 
.A1(n_1243),
.A2(n_473),
.B1(n_470),
.B2(n_453),
.Y(n_1253)
);

AOI221x1_ASAP7_75t_L g1254 ( 
.A1(n_1249),
.A2(n_473),
.B1(n_453),
.B2(n_367),
.C(n_391),
.Y(n_1254)
);

AOI221xp5_ASAP7_75t_L g1255 ( 
.A1(n_1247),
.A2(n_1250),
.B1(n_1248),
.B2(n_1253),
.C(n_1252),
.Y(n_1255)
);

AOI221xp5_ASAP7_75t_L g1256 ( 
.A1(n_1251),
.A2(n_367),
.B1(n_391),
.B2(n_393),
.C(n_382),
.Y(n_1256)
);

AOI221xp5_ASAP7_75t_L g1257 ( 
.A1(n_1255),
.A2(n_367),
.B1(n_391),
.B2(n_393),
.C(n_382),
.Y(n_1257)
);

AOI31xp33_ASAP7_75t_L g1258 ( 
.A1(n_1254),
.A2(n_1256),
.A3(n_367),
.B(n_391),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1258),
.A2(n_1257),
.B(n_367),
.Y(n_1259)
);

AOI211xp5_ASAP7_75t_L g1260 ( 
.A1(n_1259),
.A2(n_367),
.B(n_381),
.C(n_389),
.Y(n_1260)
);

AOI211xp5_ASAP7_75t_L g1261 ( 
.A1(n_1260),
.A2(n_367),
.B(n_381),
.C(n_389),
.Y(n_1261)
);


endmodule