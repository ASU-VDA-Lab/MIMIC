module fake_jpeg_992_n_371 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_371);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_371;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx4_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g84 ( 
.A(n_45),
.Y(n_84)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_46),
.Y(n_99)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_47),
.Y(n_96)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_48),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_49),
.B(n_59),
.Y(n_90)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_51),
.Y(n_112)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_28),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_23),
.B(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_60),
.Y(n_85)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_54),
.Y(n_108)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_55),
.Y(n_121)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_28),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_56),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_18),
.B(n_22),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_23),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_62),
.Y(n_116)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_18),
.Y(n_63)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

BUFx8_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

INVx8_ASAP7_75t_L g118 ( 
.A(n_64),
.Y(n_118)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_37),
.B(n_13),
.Y(n_67)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_68),
.Y(n_82)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_31),
.Y(n_69)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_18),
.Y(n_70)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_70),
.Y(n_104)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_73),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_35),
.B(n_13),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_74),
.B(n_75),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_38),
.B(n_12),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_40),
.Y(n_76)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_76),
.Y(n_105)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_60),
.B(n_33),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_77),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_64),
.A2(n_29),
.B1(n_33),
.B2(n_43),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_80),
.A2(n_87),
.B1(n_88),
.B2(n_97),
.Y(n_129)
);

AND2x4_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_42),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_83),
.B(n_111),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_64),
.A2(n_29),
.B1(n_33),
.B2(n_43),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_63),
.A2(n_70),
.B1(n_76),
.B2(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_44),
.A2(n_62),
.B1(n_51),
.B2(n_72),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_54),
.A2(n_40),
.B1(n_38),
.B2(n_43),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_98),
.A2(n_34),
.B1(n_24),
.B2(n_25),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_39),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_100),
.B(n_120),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_50),
.A2(n_40),
.B1(n_39),
.B2(n_20),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_103),
.A2(n_107),
.B1(n_24),
.B2(n_25),
.Y(n_139)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_45),
.Y(n_106)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_46),
.A2(n_40),
.B1(n_34),
.B2(n_26),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_20),
.B1(n_19),
.B2(n_32),
.Y(n_111)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_115),
.Y(n_125)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_52),
.Y(n_117)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_117),
.Y(n_162)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_119),
.B(n_12),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_69),
.B(n_41),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_42),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_122),
.B(n_68),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_123),
.B(n_128),
.Y(n_178)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_83),
.A2(n_56),
.B(n_41),
.C(n_71),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_124),
.A2(n_25),
.B(n_2),
.Y(n_182)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_78),
.Y(n_126)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_126),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_34),
.C(n_26),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_142),
.C(n_87),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_114),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_84),
.Y(n_130)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx13_ASAP7_75t_L g131 ( 
.A(n_118),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_107),
.A2(n_34),
.B1(n_32),
.B2(n_19),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_132),
.A2(n_94),
.B1(n_116),
.B2(n_79),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_133),
.A2(n_145),
.B1(n_3),
.B2(n_4),
.Y(n_196)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_134),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_137),
.Y(n_188)
);

AO22x1_ASAP7_75t_SL g138 ( 
.A1(n_83),
.A2(n_104),
.B1(n_95),
.B2(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_138),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_139),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_197)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_140),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_85),
.B(n_0),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_141),
.B(n_143),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_81),
.B(n_24),
.C(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_92),
.B(n_0),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_121),
.Y(n_144)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_110),
.A2(n_30),
.B1(n_11),
.B2(n_9),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_91),
.B(n_1),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_154),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_99),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_151),
.Y(n_193)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_149),
.Y(n_167)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_94),
.Y(n_150)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_93),
.B(n_11),
.Y(n_151)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_105),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_90),
.B(n_1),
.Y(n_154)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_102),
.Y(n_156)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_156),
.Y(n_199)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_116),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_157),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_86),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_158),
.B(n_160),
.Y(n_183)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_89),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_159),
.B(n_163),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_86),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_96),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_161),
.B(n_1),
.Y(n_187)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_112),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_166),
.B1(n_172),
.B2(n_176),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_129),
.A2(n_97),
.B1(n_108),
.B2(n_88),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_79),
.B1(n_109),
.B2(n_101),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_168),
.A2(n_173),
.B1(n_197),
.B2(n_130),
.Y(n_228)
);

XNOR2x1_ASAP7_75t_L g214 ( 
.A(n_170),
.B(n_140),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_153),
.A2(n_80),
.B1(n_112),
.B2(n_113),
.Y(n_172)
);

OAI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_133),
.A2(n_109),
.B1(n_101),
.B2(n_82),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_108),
.B1(n_113),
.B2(n_82),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_123),
.B(n_30),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_194),
.C(n_124),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_182),
.A2(n_149),
.B(n_134),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_153),
.A2(n_30),
.B1(n_9),
.B2(n_8),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_186),
.A2(n_190),
.B1(n_196),
.B2(n_198),
.Y(n_205)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_187),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_8),
.B1(n_2),
.B2(n_3),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_147),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_191),
.B(n_195),
.Y(n_225)
);

AND2x2_ASAP7_75t_SL g194 ( 
.A(n_127),
.B(n_1),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_146),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_135),
.A2(n_142),
.B1(n_141),
.B2(n_143),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_201),
.A2(n_154),
.B1(n_138),
.B2(n_156),
.Y(n_206)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_206),
.B(n_209),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_162),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_207),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_183),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_208),
.B(n_215),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_181),
.B(n_138),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_210),
.Y(n_242)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_211),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_180),
.Y(n_238)
);

AO22x1_ASAP7_75t_SL g213 ( 
.A1(n_184),
.A2(n_126),
.B1(n_152),
.B2(n_163),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_221),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_214),
.B(n_164),
.C(n_179),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_200),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_169),
.Y(n_216)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_216),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_193),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_178),
.B(n_161),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_184),
.A2(n_144),
.B1(n_157),
.B2(n_150),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_219),
.A2(n_229),
.B1(n_176),
.B2(n_199),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_191),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_220),
.Y(n_254)
);

OR2x6_ASAP7_75t_L g221 ( 
.A(n_170),
.B(n_194),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_185),
.Y(n_222)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_177),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_223),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_181),
.B(n_125),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_227),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_225),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_228),
.B(n_165),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_194),
.B(n_125),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_172),
.A2(n_155),
.B1(n_159),
.B2(n_148),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_187),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_230),
.B(n_231),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g231 ( 
.A(n_182),
.Y(n_231)
);

INVx13_ASAP7_75t_L g232 ( 
.A(n_171),
.Y(n_232)
);

HAxp5_ASAP7_75t_SL g252 ( 
.A(n_232),
.B(n_234),
.CON(n_252),
.SN(n_252)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_167),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g262 ( 
.A(n_233),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_177),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_169),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_235),
.A2(n_199),
.B1(n_189),
.B2(n_192),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_238),
.B(n_247),
.C(n_216),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_240),
.A2(n_249),
.B(n_260),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_226),
.A2(n_164),
.B(n_166),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_179),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_255),
.B(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g256 ( 
.A(n_212),
.B(n_190),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_258),
.Y(n_275)
);

A2O1A1O1Ixp25_ASAP7_75t_L g260 ( 
.A1(n_221),
.A2(n_186),
.B(n_192),
.C(n_198),
.D(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_230),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_263),
.B(n_267),
.Y(n_301)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_237),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_264),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_238),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_265),
.B(n_271),
.C(n_284),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_251),
.B(n_202),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_237),
.Y(n_268)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_269),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_208),
.Y(n_270)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_247),
.B(n_221),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_204),
.B1(n_209),
.B2(n_202),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_272),
.A2(n_274),
.B1(n_276),
.B2(n_278),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_254),
.A2(n_204),
.B1(n_206),
.B2(n_215),
.Y(n_274)
);

OAI21xp33_ASAP7_75t_L g276 ( 
.A1(n_259),
.A2(n_224),
.B(n_227),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_242),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_244),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_250),
.A2(n_221),
.B1(n_210),
.B2(n_203),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g293 ( 
.A1(n_280),
.A2(n_250),
.B(n_240),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g281 ( 
.A(n_259),
.B(n_229),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_281),
.Y(n_300)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_282),
.B(n_257),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_213),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_283),
.A2(n_260),
.B(n_261),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_248),
.A2(n_221),
.B1(n_205),
.B2(n_219),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_285),
.A2(n_258),
.B1(n_261),
.B2(n_243),
.Y(n_296)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_287),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_272),
.A2(n_250),
.B1(n_248),
.B2(n_253),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_288),
.A2(n_296),
.B1(n_298),
.B2(n_273),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_284),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_292),
.B(n_299),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_303),
.B(n_266),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_297),
.B(n_273),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_275),
.A2(n_246),
.B1(n_245),
.B2(n_239),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_256),
.Y(n_299)
);

A2O1A1O1Ixp25_ASAP7_75t_L g303 ( 
.A1(n_263),
.A2(n_246),
.B(n_262),
.C(n_205),
.D(n_243),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_236),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_280),
.C(n_266),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_279),
.B(n_267),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_285),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_309),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_310),
.A2(n_299),
.B(n_304),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_311),
.A2(n_312),
.B1(n_320),
.B2(n_296),
.Y(n_326)
);

AND2x6_ASAP7_75t_L g312 ( 
.A(n_293),
.B(n_281),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_290),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_313),
.B(n_315),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_292),
.B(n_275),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_283),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_291),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_316),
.B(n_317),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_302),
.B(n_278),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_318),
.A2(n_303),
.B(n_295),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_277),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_321),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_301),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_298),
.B(n_268),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_264),
.Y(n_333)
);

A2O1A1Ixp33_ASAP7_75t_SL g324 ( 
.A1(n_312),
.A2(n_288),
.B(n_300),
.C(n_297),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_324),
.A2(n_328),
.B(n_306),
.Y(n_340)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_325),
.Y(n_337)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_326),
.Y(n_339)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_310),
.A2(n_294),
.B(n_287),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_329),
.A2(n_331),
.B1(n_309),
.B2(n_252),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_308),
.A2(n_286),
.B1(n_289),
.B2(n_294),
.Y(n_331)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_333),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_315),
.B(n_239),
.C(n_235),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_314),
.C(n_319),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_338),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_334),
.B(n_327),
.C(n_307),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_340),
.A2(n_342),
.B1(n_325),
.B2(n_324),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_341),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_335),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_330),
.B(n_223),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_343),
.B(n_167),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_332),
.B(n_324),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g349 ( 
.A(n_344),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_346),
.B(n_347),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_339),
.A2(n_324),
.B1(n_323),
.B2(n_228),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_350),
.B(n_352),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_342),
.B(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_337),
.B(n_307),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_353),
.B(n_354),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_338),
.B(n_336),
.C(n_340),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_354),
.B(n_344),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_SL g363 ( 
.A(n_356),
.B(n_358),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_351),
.B(n_345),
.C(n_222),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_167),
.Y(n_360)
);

AOI21xp5_ASAP7_75t_L g362 ( 
.A1(n_360),
.A2(n_350),
.B(n_211),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_SL g361 ( 
.A1(n_359),
.A2(n_349),
.B(n_348),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_361),
.B(n_362),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_359),
.B(n_174),
.Y(n_364)
);

AO21x1_ASAP7_75t_L g366 ( 
.A1(n_364),
.A2(n_357),
.B(n_355),
.Y(n_366)
);

AOI21xp5_ASAP7_75t_L g367 ( 
.A1(n_366),
.A2(n_363),
.B(n_213),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_367),
.B(n_365),
.Y(n_368)
);

AOI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_368),
.A2(n_174),
.B(n_232),
.Y(n_369)
);

OAI321xp33_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_131),
.A3(n_171),
.B1(n_7),
.B2(n_5),
.C(n_6),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_370),
.B(n_7),
.Y(n_371)
);


endmodule