module real_jpeg_27171_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_215;
wire n_176;
wire n_166;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_200;
wire n_56;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_216;
wire n_213;
wire n_167;
wire n_179;
wire n_202;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_0),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_0),
.A2(n_36),
.B1(n_43),
.B2(n_44),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_0),
.A2(n_36),
.B1(n_76),
.B2(n_78),
.Y(n_97)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_1),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_2),
.A2(n_72),
.B1(n_73),
.B2(n_82),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_2),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_2),
.A2(n_76),
.B1(n_78),
.B2(n_82),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_2),
.A2(n_43),
.B1(n_44),
.B2(n_82),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_2),
.A2(n_28),
.B1(n_29),
.B2(n_82),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_3),
.A2(n_72),
.B1(n_73),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_3),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_3),
.A2(n_76),
.B1(n_78),
.B2(n_114),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_114),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_114),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_4),
.Y(n_71)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_5),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_5),
.B(n_78),
.Y(n_145)
);

AOI21xp33_ASAP7_75t_L g149 ( 
.A1(n_5),
.A2(n_78),
.B(n_145),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_5),
.B(n_75),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_5),
.A2(n_43),
.B1(n_44),
.B2(n_103),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_5),
.A2(n_29),
.B(n_48),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_5),
.B(n_183),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_5),
.A2(n_57),
.B1(n_200),
.B2(n_201),
.Y(n_203)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_72),
.B1(n_73),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_7),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_7),
.A2(n_76),
.B1(n_78),
.B2(n_80),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_7),
.A2(n_43),
.B1(n_44),
.B2(n_80),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_7),
.A2(n_28),
.B1(n_29),
.B2(n_80),
.Y(n_192)
);

INVx13_ASAP7_75t_L g73 ( 
.A(n_8),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_9),
.A2(n_28),
.B1(n_29),
.B2(n_50),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_10),
.A2(n_39),
.B1(n_76),
.B2(n_78),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_39),
.B1(n_43),
.B2(n_44),
.Y(n_125)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_11),
.A2(n_43),
.B1(n_44),
.B2(n_46),
.Y(n_42)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_12),
.A2(n_43),
.B1(n_44),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_12),
.A2(n_28),
.B1(n_29),
.B2(n_52),
.Y(n_58)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_13),
.Y(n_77)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_14),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_14),
.Y(n_91)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_116),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_116),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_98),
.B2(n_115),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_53),
.B2(n_54),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_40),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_37),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_26),
.A2(n_33),
.B(n_105),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_34),
.Y(n_26)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_27),
.A2(n_38),
.B(n_60),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_27),
.A2(n_32),
.B1(n_191),
.B2(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.Y(n_27)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_28),
.A2(n_29),
.B1(n_46),
.B2(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_28),
.B(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx4f_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_38),
.Y(n_37)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_33),
.B(n_35),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_33),
.A2(n_57),
.B1(n_58),
.B2(n_105),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_37),
.A2(n_57),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B1(n_49),
.B2(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_41),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_41),
.A2(n_47),
.B1(n_153),
.B2(n_154),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_SL g167 ( 
.A1(n_41),
.A2(n_154),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_41),
.A2(n_47),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_41),
.A2(n_47),
.B1(n_153),
.B2(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_47),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_43),
.A2(n_44),
.B1(n_90),
.B2(n_93),
.Y(n_92)
);

AOI32xp33_ASAP7_75t_L g143 ( 
.A1(n_43),
.A2(n_76),
.A3(n_144),
.B1(n_145),
.B2(n_146),
.Y(n_143)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

NAND2xp33_ASAP7_75t_SL g146 ( 
.A(n_44),
.B(n_89),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_L g177 ( 
.A1(n_44),
.A2(n_46),
.B(n_103),
.C(n_178),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_46),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_49),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_47),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_47),
.B(n_103),
.Y(n_198)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_56),
.B(n_61),
.Y(n_55)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_61),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B(n_59),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_57),
.A2(n_192),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_64),
.B(n_127),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_84),
.B2(n_85),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_79),
.B1(n_81),
.B2(n_83),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_68),
.A2(n_79),
.B1(n_83),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_69),
.A2(n_75),
.B1(n_102),
.B2(n_113),
.Y(n_131)
);

O2A1O1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_72),
.B(n_74),
.C(n_75),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_70),
.B(n_72),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_70),
.A2(n_71),
.B1(n_76),
.B2(n_78),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_70),
.B(n_78),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g70 ( 
.A(n_71),
.Y(n_70)
);

HAxp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_103),
.CON(n_102),
.SN(n_102)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_74),
.A2(n_76),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_78),
.B1(n_89),
.B2(n_91),
.Y(n_88)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_94),
.B(n_96),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_107),
.B(n_109),
.Y(n_106)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_87),
.A2(n_92),
.B1(n_108),
.B2(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_87),
.A2(n_92),
.B1(n_149),
.B2(n_150),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_87),
.A2(n_92),
.B1(n_130),
.B2(n_150),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_89),
.Y(n_144)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_91),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_97),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_92),
.B(n_95),
.Y(n_109)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_92),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_106),
.C(n_110),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_SL g117 ( 
.A(n_99),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_100),
.B(n_104),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_103),
.B(n_201),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_110),
.B1(n_111),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_120),
.C(n_121),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_117),
.B(n_232),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_120),
.B(n_121),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_128),
.C(n_131),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_122),
.A2(n_123),
.B1(n_128),
.B2(n_129),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_125),
.B(n_127),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_131),
.B(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_233),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_136),
.B(n_229),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_216),
.B(n_228),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_169),
.B(n_215),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_155),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_139),
.B(n_155),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_147),
.C(n_151),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_140),
.A2(n_141),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_142),
.B(n_143),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_164),
.B2(n_165),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_156),
.B(n_166),
.C(n_167),
.Y(n_217)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_158),
.B(n_160),
.C(n_163),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_170),
.A2(n_209),
.B(n_214),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_188),
.B(n_208),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_179),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_172),
.B(n_179),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_177),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_173),
.A2(n_174),
.B1(n_177),
.B2(n_195),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_186),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_184),
.B2(n_185),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_181),
.B(n_185),
.C(n_186),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_187),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_196),
.B(n_207),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_190),
.B(n_194),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_197),
.A2(n_202),
.B(n_206),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_198),
.B(n_199),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_211),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_210),
.B(n_211),
.Y(n_214)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_217),
.B(n_218),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_219),
.A2(n_224),
.B1(n_225),
.B2(n_227),
.Y(n_218)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_219),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_221),
.B1(n_222),
.B2(n_223),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_223),
.C(n_224),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_231),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_234),
.Y(n_233)
);


endmodule