module real_aes_12925_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_852;
wire n_766;
wire n_132;
wire n_857;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_746;
wire n_532;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_860;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_874;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_867;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_827;
wire n_809;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_249;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
OA21x2_ASAP7_75t_L g135 ( .A1(n_0), .A2(n_50), .B(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g173 ( .A(n_0), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_1), .B(n_167), .Y(n_209) );
AND2x2_ASAP7_75t_L g548 ( .A(n_2), .B(n_161), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_3), .B(n_294), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_4), .A2(n_96), .B1(n_140), .B2(n_212), .C(n_226), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_5), .B(n_233), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_6), .B(n_233), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_7), .B(n_134), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_8), .B(n_169), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_9), .B(n_212), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_10), .B(n_169), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_11), .B(n_148), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_12), .B(n_208), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_13), .Y(n_275) );
INVx1_ASAP7_75t_L g142 ( .A(n_14), .Y(n_142) );
BUFx3_ASAP7_75t_L g146 ( .A(n_14), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_15), .B(n_153), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_16), .B(n_526), .Y(n_553) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_17), .Y(n_289) );
CKINVDCx5p33_ASAP7_75t_R g599 ( .A(n_18), .Y(n_599) );
BUFx10_ASAP7_75t_L g114 ( .A(n_19), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g139 ( .A(n_20), .B(n_140), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_21), .B(n_567), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_22), .B(n_528), .Y(n_596) );
OAI21xp33_ASAP7_75t_L g697 ( .A1(n_22), .A2(n_71), .B(n_286), .Y(n_697) );
CKINVDCx5p33_ASAP7_75t_R g269 ( .A(n_23), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_24), .B(n_167), .Y(n_223) );
O2A1O1Ixp5_ASAP7_75t_L g630 ( .A1(n_25), .A2(n_164), .B(n_248), .C(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_SL g151 ( .A(n_26), .B(n_140), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_27), .B(n_153), .Y(n_186) );
NAND2xp33_ASAP7_75t_L g213 ( .A(n_28), .B(n_145), .Y(n_213) );
INVx1_ASAP7_75t_L g158 ( .A(n_29), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g265 ( .A1(n_30), .A2(n_189), .B(n_266), .C(n_268), .Y(n_265) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_31), .B(n_168), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_32), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_33), .B(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_34), .B(n_231), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_35), .B(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g507 ( .A(n_36), .Y(n_507) );
AND3x2_ASAP7_75t_L g851 ( .A(n_36), .B(n_109), .C(n_111), .Y(n_851) );
AO221x1_ASAP7_75t_L g160 ( .A1(n_37), .A2(n_87), .B1(n_140), .B2(n_148), .C(n_161), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_38), .B(n_185), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_39), .B(n_526), .Y(n_525) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_40), .A2(n_88), .B1(n_866), .B2(n_867), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_40), .Y(n_866) );
AND2x4_ASAP7_75t_L g157 ( .A(n_41), .B(n_158), .Y(n_157) );
NAND2x1_ASAP7_75t_L g543 ( .A(n_42), .B(n_161), .Y(n_543) );
CKINVDCx5p33_ASAP7_75t_R g602 ( .A(n_43), .Y(n_602) );
INVx1_ASAP7_75t_L g539 ( .A(n_44), .Y(n_539) );
NAND3xp33_ASAP7_75t_L g191 ( .A(n_45), .B(n_189), .C(n_192), .Y(n_191) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_46), .Y(n_615) );
AND2x2_ASAP7_75t_L g547 ( .A(n_47), .B(n_192), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_48), .B(n_231), .Y(n_584) );
AOI22xp33_ASAP7_75t_L g118 ( .A1(n_49), .A2(n_61), .B1(n_119), .B2(n_120), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_49), .Y(n_120) );
INVx1_ASAP7_75t_L g174 ( .A(n_50), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_51), .B(n_134), .Y(n_624) );
INVx1_ASAP7_75t_L g136 ( .A(n_52), .Y(n_136) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_53), .A2(n_240), .B(n_242), .C(n_244), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g273 ( .A(n_54), .Y(n_273) );
CKINVDCx5p33_ASAP7_75t_R g847 ( .A(n_55), .Y(n_847) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_56), .B(n_192), .Y(n_552) );
INVx2_ASAP7_75t_L g243 ( .A(n_57), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_58), .B(n_134), .Y(n_297) );
AND2x4_ASAP7_75t_L g882 ( .A(n_59), .B(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_60), .B(n_528), .Y(n_592) );
INVx1_ASAP7_75t_L g119 ( .A(n_61), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_62), .B(n_167), .Y(n_542) );
NOR2xp67_ASAP7_75t_L g110 ( .A(n_63), .B(n_80), .Y(n_110) );
HB1xp67_ASAP7_75t_L g887 ( .A(n_63), .Y(n_887) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_64), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g522 ( .A(n_65), .B(n_231), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_66), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g883 ( .A(n_67), .Y(n_883) );
AND2x2_ASAP7_75t_L g550 ( .A(n_68), .B(n_134), .Y(n_550) );
AND2x2_ASAP7_75t_L g236 ( .A(n_69), .B(n_134), .Y(n_236) );
INVx1_ASAP7_75t_L g177 ( .A(n_70), .Y(n_177) );
CKINVDCx5p33_ASAP7_75t_R g634 ( .A(n_71), .Y(n_634) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_72), .B(n_248), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_73), .B(n_169), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_74), .B(n_231), .Y(n_617) );
CKINVDCx5p33_ASAP7_75t_R g632 ( .A(n_75), .Y(n_632) );
INVx2_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g880 ( .A(n_76), .B(n_506), .C(n_881), .Y(n_880) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_77), .B(n_290), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g166 ( .A1(n_78), .A2(n_82), .B1(n_167), .B2(n_169), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_79), .B(n_189), .Y(n_188) );
HB1xp67_ASAP7_75t_L g886 ( .A(n_80), .Y(n_886) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_81), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_83), .B(n_252), .Y(n_561) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_84), .B(n_192), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g603 ( .A(n_85), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_86), .B(n_567), .Y(n_590) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_88), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_89), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g251 ( .A(n_90), .B(n_252), .Y(n_251) );
BUFx3_ASAP7_75t_L g149 ( .A(n_91), .Y(n_149) );
INVx1_ASAP7_75t_L g165 ( .A(n_91), .Y(n_165) );
INVx1_ASAP7_75t_L g227 ( .A(n_91), .Y(n_227) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_92), .A2(n_102), .B1(n_874), .B2(n_888), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g131 ( .A(n_93), .B(n_132), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_94), .B(n_277), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_95), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_97), .B(n_134), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_98), .B(n_623), .Y(n_622) );
CKINVDCx5p33_ASAP7_75t_R g873 ( .A(n_99), .Y(n_873) );
CKINVDCx5p33_ASAP7_75t_R g198 ( .A(n_100), .Y(n_198) );
OR2x2_ASAP7_75t_L g102 ( .A(n_103), .B(n_870), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_104), .B(n_852), .Y(n_103) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_115), .B(n_846), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
BUFx8_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
OR2x6_ASAP7_75t_L g107 ( .A(n_108), .B(n_113), .Y(n_107) );
AND2x2_ASAP7_75t_L g108 ( .A(n_109), .B(n_111), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g863 ( .A(n_110), .B(n_507), .Y(n_863) );
BUFx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
INVx1_ASAP7_75t_L g862 ( .A(n_112), .Y(n_862) );
BUFx3_ASAP7_75t_L g854 ( .A(n_113), .Y(n_854) );
INVx3_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_114), .B(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
XNOR2xp5_ASAP7_75t_L g116 ( .A(n_117), .B(n_121), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
OAI22xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_503), .B1(n_508), .B2(n_845), .Y(n_121) );
INVx2_ASAP7_75t_SL g868 ( .A(n_122), .Y(n_868) );
NOR2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_433), .Y(n_122) );
NAND4xp25_ASAP7_75t_L g123 ( .A(n_124), .B(n_340), .C(n_376), .D(n_401), .Y(n_123) );
NOR3xp33_ASAP7_75t_L g124 ( .A(n_125), .B(n_307), .C(n_323), .Y(n_124) );
OAI221xp5_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_216), .B1(n_278), .B2(n_283), .C(n_298), .Y(n_125) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_179), .Y(n_127) );
INVx2_ASAP7_75t_L g392 ( .A(n_128), .Y(n_392) );
AND2x4_ASAP7_75t_L g424 ( .A(n_128), .B(n_346), .Y(n_424) );
AND2x2_ASAP7_75t_L g502 ( .A(n_128), .B(n_368), .Y(n_502) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_159), .Y(n_128) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_129), .B(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g366 ( .A(n_129), .Y(n_366) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
NOR2xp33_ASAP7_75t_L g300 ( .A(n_130), .B(n_202), .Y(n_300) );
AND2x2_ASAP7_75t_L g326 ( .A(n_130), .B(n_280), .Y(n_326) );
HB1xp67_ASAP7_75t_L g344 ( .A(n_130), .Y(n_344) );
OR2x2_ASAP7_75t_L g348 ( .A(n_130), .B(n_159), .Y(n_348) );
AND2x2_ASAP7_75t_L g361 ( .A(n_130), .B(n_202), .Y(n_361) );
AND2x4_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .Y(n_130) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
INVxp67_ASAP7_75t_SL g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g155 ( .A(n_134), .B(n_156), .Y(n_155) );
INVx2_ASAP7_75t_L g196 ( .A(n_134), .Y(n_196) );
INVx1_ASAP7_75t_L g204 ( .A(n_134), .Y(n_204) );
INVxp33_ASAP7_75t_L g556 ( .A(n_134), .Y(n_556) );
BUFx6f_ASAP7_75t_L g581 ( .A(n_134), .Y(n_581) );
INVx1_ASAP7_75t_L g635 ( .A(n_134), .Y(n_635) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
BUFx2_ASAP7_75t_L g200 ( .A(n_135), .Y(n_200) );
INVx1_ASAP7_75t_L g253 ( .A(n_135), .Y(n_253) );
INVx1_ASAP7_75t_L g175 ( .A(n_136), .Y(n_175) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_150), .B(n_155), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g138 ( .A1(n_139), .A2(n_143), .B(n_147), .Y(n_138) );
INVx2_ASAP7_75t_L g567 ( .A(n_140), .Y(n_567) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
INVx2_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_142), .Y(n_193) );
INVx2_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
INVx3_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
INVx2_ASAP7_75t_L g233 ( .A(n_145), .Y(n_233) );
INVx2_ASAP7_75t_L g526 ( .A(n_145), .Y(n_526) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx2_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g271 ( .A1(n_147), .A2(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g154 ( .A(n_149), .Y(n_154) );
INVx2_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g538 ( .A(n_149), .B(n_539), .Y(n_538) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_154), .Y(n_150) );
INVx1_ASAP7_75t_L g536 ( .A(n_153), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_154), .A2(n_184), .B(n_186), .Y(n_183) );
O2A1O1Ixp5_ASAP7_75t_L g288 ( .A1(n_154), .A2(n_289), .B(n_290), .C(n_291), .Y(n_288) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_154), .A2(n_225), .B(n_599), .C(n_600), .Y(n_598) );
NOR2xp33_ASAP7_75t_R g171 ( .A(n_156), .B(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g195 ( .A(n_156), .Y(n_195) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_156), .B(n_629), .C(n_630), .Y(n_628) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx2_ASAP7_75t_L g263 ( .A(n_157), .Y(n_263) );
BUFx6f_ASAP7_75t_SL g296 ( .A(n_157), .Y(n_296) );
INVx1_ASAP7_75t_L g606 ( .A(n_157), .Y(n_606) );
OR2x2_ASAP7_75t_L g279 ( .A(n_159), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g301 ( .A(n_159), .B(n_282), .Y(n_301) );
BUFx3_ASAP7_75t_L g314 ( .A(n_159), .Y(n_314) );
INVx2_ASAP7_75t_SL g334 ( .A(n_159), .Y(n_334) );
AND2x2_ASAP7_75t_L g375 ( .A(n_159), .B(n_366), .Y(n_375) );
AND2x2_ASAP7_75t_L g398 ( .A(n_159), .B(n_310), .Y(n_398) );
AO31x2_ASAP7_75t_L g159 ( .A1(n_160), .A2(n_162), .A3(n_171), .B(n_176), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_163), .B(n_166), .Y(n_162) );
AOI21x1_ASAP7_75t_L g541 ( .A1(n_163), .A2(n_542), .B(n_543), .Y(n_541) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_163), .A2(n_569), .B(n_570), .Y(n_568) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_164), .A2(n_207), .B(n_209), .Y(n_206) );
INVx2_ASAP7_75t_L g587 ( .A(n_164), .Y(n_587) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
BUFx3_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
INVx1_ASAP7_75t_L g586 ( .A(n_167), .Y(n_586) );
INVx2_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
INVx2_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
INVx2_ASAP7_75t_L g231 ( .A(n_168), .Y(n_231) );
INVx1_ASAP7_75t_L g565 ( .A(n_168), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_169), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx2_ASAP7_75t_L g208 ( .A(n_170), .Y(n_208) );
INVx1_ASAP7_75t_L g612 ( .A(n_170), .Y(n_612) );
INVx2_ASAP7_75t_L g621 ( .A(n_170), .Y(n_621) );
NAND2xp5_ASAP7_75t_SL g631 ( .A(n_170), .B(n_632), .Y(n_631) );
INVx2_ASAP7_75t_L g178 ( .A(n_172), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_172), .B(n_606), .Y(n_605) );
AOI21x1_ASAP7_75t_L g172 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_172) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_173), .A2(n_174), .B(n_175), .Y(n_261) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
HB1xp67_ASAP7_75t_L g699 ( .A(n_178), .Y(n_699) );
AND2x2_ASAP7_75t_L g343 ( .A(n_179), .B(n_344), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_179), .B(n_365), .Y(n_405) );
AND2x2_ASAP7_75t_L g459 ( .A(n_179), .B(n_334), .Y(n_459) );
AND2x2_ASAP7_75t_L g473 ( .A(n_179), .B(n_474), .Y(n_473) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
OR2x2_ASAP7_75t_L g439 ( .A(n_180), .B(n_348), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_181), .B(n_201), .Y(n_180) );
INVx2_ASAP7_75t_L g282 ( .A(n_181), .Y(n_282) );
BUFx2_ASAP7_75t_SL g322 ( .A(n_181), .Y(n_322) );
AND2x2_ASAP7_75t_L g346 ( .A(n_181), .B(n_202), .Y(n_346) );
INVx1_ASAP7_75t_L g368 ( .A(n_181), .Y(n_368) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
O2A1O1Ixp5_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_187), .B(n_194), .C(n_197), .Y(n_182) );
INVx2_ASAP7_75t_SL g225 ( .A(n_185), .Y(n_225) );
OAI21xp5_ASAP7_75t_L g187 ( .A1(n_188), .A2(n_190), .B(n_191), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_189), .A2(n_524), .B(n_525), .Y(n_523) );
INVx2_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
INVx1_ASAP7_75t_L g241 ( .A(n_193), .Y(n_241) );
INVx2_ASAP7_75t_L g248 ( .A(n_193), .Y(n_248) );
INVx2_ASAP7_75t_L g294 ( .A(n_193), .Y(n_294) );
INVx1_ASAP7_75t_L g540 ( .A(n_193), .Y(n_540) );
NAND2x1_ASAP7_75t_L g221 ( .A(n_194), .B(n_222), .Y(n_221) );
AOI21x1_ASAP7_75t_L g228 ( .A1(n_194), .A2(n_229), .B(n_236), .Y(n_228) );
AND2x4_ASAP7_75t_L g194 ( .A(n_195), .B(n_196), .Y(n_194) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_195), .A2(n_206), .B(n_210), .Y(n_205) );
AOI21xp33_ASAP7_75t_L g254 ( .A1(n_195), .A2(n_199), .B(n_251), .Y(n_254) );
AOI21xp33_ASAP7_75t_L g555 ( .A1(n_195), .A2(n_550), .B(n_556), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g197 ( .A(n_198), .B(n_199), .Y(n_197) );
INVxp67_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
BUFx3_ASAP7_75t_L g286 ( .A(n_200), .Y(n_286) );
INVx1_ASAP7_75t_L g518 ( .A(n_200), .Y(n_518) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g280 ( .A(n_202), .Y(n_280) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_202), .Y(n_311) );
INVx1_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
OA21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_205), .B(n_215), .Y(n_202) );
OAI21x1_ASAP7_75t_L g532 ( .A1(n_203), .A2(n_533), .B(n_544), .Y(n_532) );
INVx1_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OAI221xp5_ASAP7_75t_L g601 ( .A1(n_208), .A2(n_294), .B1(n_602), .B2(n_603), .C(n_604), .Y(n_601) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_213), .B(n_214), .Y(n_210) );
INVx2_ASAP7_75t_L g267 ( .A(n_212), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_212), .B(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g290 ( .A(n_212), .Y(n_290) );
INVx1_ASAP7_75t_L g244 ( .A(n_214), .Y(n_244) );
INVx2_ASAP7_75t_L g554 ( .A(n_214), .Y(n_554) );
OR2x2_ASAP7_75t_L g216 ( .A(n_217), .B(n_255), .Y(n_216) );
OR2x2_ASAP7_75t_L g315 ( .A(n_217), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g471 ( .A(n_217), .Y(n_471) );
OR2x2_ASAP7_75t_L g495 ( .A(n_217), .B(n_356), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_237), .Y(n_217) );
AND2x2_ASAP7_75t_L g306 ( .A(n_218), .B(n_238), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_218), .B(n_256), .Y(n_388) );
OR2x2_ASAP7_75t_L g417 ( .A(n_218), .B(n_330), .Y(n_417) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g339 ( .A(n_219), .B(n_238), .Y(n_339) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
AND2x2_ASAP7_75t_L g284 ( .A(n_220), .B(n_285), .Y(n_284) );
INVx1_ASAP7_75t_L g320 ( .A(n_220), .Y(n_320) );
AND2x2_ASAP7_75t_L g400 ( .A(n_220), .B(n_331), .Y(n_400) );
OR2x2_ASAP7_75t_L g453 ( .A(n_220), .B(n_238), .Y(n_453) );
NAND2x1p5_ASAP7_75t_L g220 ( .A(n_221), .B(n_228), .Y(n_220) );
AOI21xp5_ASAP7_75t_SL g222 ( .A1(n_223), .A2(n_224), .B(n_226), .Y(n_222) );
INVx1_ASAP7_75t_L g604 ( .A(n_226), .Y(n_604) );
OAI22xp5_ASAP7_75t_L g610 ( .A1(n_226), .A2(n_611), .B1(n_613), .B2(n_617), .Y(n_610) );
INVx2_ASAP7_75t_SL g616 ( .A(n_226), .Y(n_616) );
BUFx3_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g235 ( .A(n_227), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_232), .B(n_234), .Y(n_229) );
INVx1_ASAP7_75t_L g250 ( .A(n_234), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_234), .A2(n_293), .B(n_295), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_234), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_234), .A2(n_564), .B(n_566), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_234), .A2(n_589), .B(n_590), .Y(n_588) );
AOI21xp5_ASAP7_75t_L g618 ( .A1(n_234), .A2(n_619), .B(n_622), .Y(n_618) );
BUFx10_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g329 ( .A(n_237), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g354 ( .A(n_238), .Y(n_354) );
INVx2_ASAP7_75t_L g380 ( .A(n_238), .Y(n_380) );
AND2x2_ASAP7_75t_L g407 ( .A(n_238), .B(n_257), .Y(n_407) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_245), .B(n_254), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g242 ( .A(n_240), .B(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g240 ( .A(n_241), .Y(n_240) );
NOR2xp33_ASAP7_75t_L g272 ( .A(n_241), .B(n_273), .Y(n_272) );
OAI21xp5_ASAP7_75t_L g546 ( .A1(n_244), .A2(n_547), .B(n_548), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_250), .B(n_251), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_247), .B(n_249), .Y(n_246) );
BUFx6f_ASAP7_75t_L g528 ( .A(n_252), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_252), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
BUFx2_ASAP7_75t_SL g255 ( .A(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g316 ( .A(n_256), .Y(n_316) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g371 ( .A(n_257), .B(n_372), .Y(n_371) );
OR2x2_ASAP7_75t_L g416 ( .A(n_257), .B(n_380), .Y(n_416) );
INVx3_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_258), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g422 ( .A(n_258), .B(n_330), .Y(n_422) );
AO21x2_ASAP7_75t_L g258 ( .A1(n_259), .A2(n_264), .B(n_270), .Y(n_258) );
AO21x1_ASAP7_75t_SL g305 ( .A1(n_259), .A2(n_264), .B(n_270), .Y(n_305) );
INVxp67_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OAI21x1_ASAP7_75t_SL g270 ( .A1(n_260), .A2(n_271), .B(n_276), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
INVx2_ASAP7_75t_L g277 ( .A(n_261), .Y(n_277) );
AO21x2_ASAP7_75t_L g627 ( .A1(n_261), .A2(n_628), .B(n_633), .Y(n_627) );
OAI21x1_ASAP7_75t_L g609 ( .A1(n_262), .A2(n_610), .B(n_618), .Y(n_609) );
INVx2_ASAP7_75t_SL g262 ( .A(n_263), .Y(n_262) );
INVx1_ASAP7_75t_L g591 ( .A(n_263), .Y(n_591) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
OR2x2_ASAP7_75t_L g321 ( .A(n_279), .B(n_322), .Y(n_321) );
NOR2x1_ASAP7_75t_SL g442 ( .A(n_279), .B(n_322), .Y(n_442) );
INVx2_ASAP7_75t_L g385 ( .A(n_281), .Y(n_385) );
INVx2_ASAP7_75t_L g310 ( .A(n_282), .Y(n_310) );
INVx6_ASAP7_75t_L g359 ( .A(n_283), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_283), .B(n_499), .Y(n_498) );
INVx4_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x2_ASAP7_75t_L g406 ( .A(n_284), .B(n_407), .Y(n_406) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_284), .Y(n_475) );
INVx2_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
INVxp33_ASAP7_75t_L g372 ( .A(n_285), .Y(n_372) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_286), .A2(n_287), .B(n_297), .Y(n_285) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_292), .B(n_296), .Y(n_287) );
INVx2_ASAP7_75t_L g623 ( .A(n_294), .Y(n_623) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_296), .A2(n_520), .B(n_523), .Y(n_519) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_296), .A2(n_534), .B(n_541), .Y(n_533) );
INVx1_ASAP7_75t_L g572 ( .A(n_296), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_302), .Y(n_298) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
INVxp67_ASAP7_75t_L g418 ( .A(n_300), .Y(n_418) );
AND2x4_ASAP7_75t_L g325 ( .A(n_301), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g363 ( .A(n_302), .Y(n_363) );
AND2x2_ASAP7_75t_L g302 ( .A(n_303), .B(n_306), .Y(n_302) );
NAND2x1_ASAP7_75t_L g358 ( .A(n_303), .B(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g444 ( .A(n_303), .Y(n_444) );
AND2x2_ASAP7_75t_L g451 ( .A(n_303), .B(n_452), .Y(n_451) );
AND2x4_ASAP7_75t_L g487 ( .A(n_303), .B(n_488), .Y(n_487) );
INVx5_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g378 ( .A(n_304), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g432 ( .A(n_304), .B(n_339), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_304), .B(n_437), .Y(n_436) );
AND2x2_ASAP7_75t_L g458 ( .A(n_304), .B(n_452), .Y(n_458) );
AND2x4_ASAP7_75t_SL g464 ( .A(n_304), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_304), .B(n_492), .Y(n_491) );
BUFx6f_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g318 ( .A(n_305), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_315), .B1(n_317), .B2(n_321), .Y(n_307) );
OR2x2_ASAP7_75t_L g308 ( .A(n_309), .B(n_312), .Y(n_308) );
OR2x2_ASAP7_75t_L g426 ( .A(n_309), .B(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
INVx1_ASAP7_75t_L g430 ( .A(n_310), .Y(n_430) );
AND2x2_ASAP7_75t_L g493 ( .A(n_310), .B(n_360), .Y(n_493) );
AND2x2_ASAP7_75t_L g411 ( .A(n_311), .B(n_412), .Y(n_411) );
INVxp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g409 ( .A(n_313), .B(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx2_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_314), .Y(n_382) );
INVx1_ASAP7_75t_L g427 ( .A(n_314), .Y(n_427) );
AND2x4_ASAP7_75t_L g423 ( .A(n_316), .B(n_339), .Y(n_423) );
OR2x2_ASAP7_75t_L g448 ( .A(n_316), .B(n_399), .Y(n_448) );
OR2x2_ASAP7_75t_L g327 ( .A(n_317), .B(n_328), .Y(n_327) );
NAND2x1p5_ASAP7_75t_L g317 ( .A(n_318), .B(n_319), .Y(n_317) );
AND2x4_ASAP7_75t_L g414 ( .A(n_319), .B(n_329), .Y(n_414) );
INVx1_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
INVx3_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g492 ( .A(n_320), .B(n_338), .Y(n_492) );
AND2x2_ASAP7_75t_L g478 ( .A(n_322), .B(n_361), .Y(n_478) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_324), .A2(n_327), .B1(n_332), .B2(n_335), .Y(n_323) );
INVx4_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
AOI21xp5_ASAP7_75t_L g468 ( .A1(n_325), .A2(n_464), .B(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g397 ( .A(n_326), .B(n_398), .Y(n_397) );
NAND2x1_ASAP7_75t_L g497 ( .A(n_326), .B(n_430), .Y(n_497) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
OR2x2_ASAP7_75t_L g379 ( .A(n_330), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g338 ( .A(n_331), .Y(n_338) );
INVx1_ASAP7_75t_L g356 ( .A(n_331), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
INVx2_ASAP7_75t_L g384 ( .A(n_333), .Y(n_384) );
AOI211x1_ASAP7_75t_L g460 ( .A1(n_333), .A2(n_461), .B(n_466), .C(n_472), .Y(n_460) );
AND2x4_ASAP7_75t_SL g360 ( .A(n_334), .B(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g474 ( .A(n_334), .B(n_366), .Y(n_474) );
INVx2_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AO22x1_ASAP7_75t_L g500 ( .A1(n_336), .A2(n_423), .B1(n_501), .B2(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
OR2x2_ASAP7_75t_L g445 ( .A(n_337), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g463 ( .A(n_337), .Y(n_463) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
OR2x2_ASAP7_75t_L g467 ( .A(n_338), .B(n_453), .Y(n_467) );
INVx1_ASAP7_75t_L g446 ( .A(n_339), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_349), .B1(n_357), .B2(n_360), .C(n_362), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_342), .B(n_345), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AOI221xp5_ASAP7_75t_SL g376 ( .A1(n_343), .A2(n_377), .B1(n_381), .B2(n_386), .C(n_391), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NOR2x1_ASAP7_75t_L g455 ( .A(n_348), .B(n_368), .Y(n_455) );
INVx2_ASAP7_75t_L g465 ( .A(n_348), .Y(n_465) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g350 ( .A(n_351), .B(n_355), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_353), .Y(n_395) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AND2x4_ASAP7_75t_SL g488 ( .A(n_356), .B(n_482), .Y(n_488) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g449 ( .A(n_360), .Y(n_449) );
AND2x2_ASAP7_75t_L g403 ( .A(n_361), .B(n_368), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_364), .B1(n_370), .B2(n_373), .Y(n_362) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_367), .Y(n_364) );
INVx1_ASAP7_75t_L g441 ( .A(n_365), .Y(n_441) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g412 ( .A(n_366), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_368), .B(n_369), .Y(n_367) );
INVx2_ASAP7_75t_L g374 ( .A(n_368), .Y(n_374) );
AND2x2_ASAP7_75t_L g501 ( .A(n_368), .B(n_465), .Y(n_501) );
INVx1_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g477 ( .A(n_371), .B(n_452), .Y(n_477) );
AND2x2_ASAP7_75t_L g390 ( .A(n_372), .B(n_380), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_374), .B(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g469 ( .A(n_374), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_374), .B(n_375), .Y(n_486) );
AND2x2_ASAP7_75t_L g429 ( .A(n_375), .B(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NOR2x1_ASAP7_75t_L g457 ( .A(n_379), .B(n_388), .Y(n_457) );
NAND2xp33_ASAP7_75t_L g480 ( .A(n_379), .B(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g421 ( .A(n_380), .Y(n_421) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_383), .Y(n_381) );
AND2x4_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2xp5_ASAP7_75t_SL g386 ( .A(n_387), .B(n_389), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g435 ( .A1(n_389), .A2(n_436), .B(n_439), .C(n_440), .Y(n_435) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_393), .B(n_396), .C(n_399), .Y(n_391) );
INVx1_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NOR3xp33_ASAP7_75t_L g401 ( .A(n_402), .B(n_408), .C(n_425), .Y(n_401) );
OA21x2_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_404), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g496 ( .A(n_403), .Y(n_496) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g476 ( .A(n_407), .Y(n_476) );
OAI221xp5_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_413), .B1(n_415), .B2(n_418), .C(n_419), .Y(n_408) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
OR2x2_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g499 ( .A(n_416), .Y(n_499) );
OAI21xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_423), .B(n_424), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_421), .B(n_422), .Y(n_420) );
AOI21xp5_ASAP7_75t_L g425 ( .A1(n_426), .A2(n_428), .B(n_431), .Y(n_425) );
INVx1_ASAP7_75t_L g485 ( .A(n_427), .Y(n_485) );
INVx1_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
NAND4xp75_ASAP7_75t_L g433 ( .A(n_434), .B(n_460), .C(n_479), .D(n_489), .Y(n_433) );
AOI21xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_443), .B(n_447), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_439), .B(n_444), .C(n_445), .Y(n_443) );
OAI22xp33_ASAP7_75t_L g466 ( .A1(n_440), .A2(n_467), .B1(n_468), .B2(n_470), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OAI221xp5_ASAP7_75t_SL g447 ( .A1(n_448), .A2(n_449), .B1(n_450), .B2(n_454), .C(n_456), .Y(n_447) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx2_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g482 ( .A(n_453), .Y(n_482) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_455), .A2(n_457), .B1(n_458), .B2(n_459), .Y(n_456) );
AND2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_464), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
AO32x1_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_475), .A3(n_476), .B1(n_477), .B2(n_478), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_478), .B(n_485), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_483), .B1(n_486), .B2(n_487), .Y(n_479) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AOI211xp5_ASAP7_75t_L g489 ( .A1(n_490), .A2(n_493), .B(n_494), .C(n_500), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
OAI22xp33_ASAP7_75t_SL g494 ( .A1(n_495), .A2(n_496), .B1(n_497), .B2(n_498), .Y(n_494) );
INVxp67_ASAP7_75t_SL g845 ( .A(n_503), .Y(n_845) );
BUFx8_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
NOR2x1_ASAP7_75t_L g508 ( .A(n_509), .B(n_771), .Y(n_508) );
NAND4xp25_ASAP7_75t_L g509 ( .A(n_510), .B(n_681), .C(n_720), .D(n_753), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_511), .B(n_656), .Y(n_510) );
OAI222xp33_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_576), .B1(n_625), .B2(n_639), .C1(n_644), .C2(n_651), .Y(n_511) );
NOR2xp67_ASAP7_75t_SL g512 ( .A(n_513), .B(n_557), .Y(n_512) );
AND2x2_ASAP7_75t_L g754 ( .A(n_513), .B(n_755), .Y(n_754) );
AND2x2_ASAP7_75t_L g513 ( .A(n_514), .B(n_529), .Y(n_513) );
AND2x2_ASAP7_75t_L g690 ( .A(n_514), .B(n_560), .Y(n_690) );
HB1xp67_ASAP7_75t_L g705 ( .A(n_514), .Y(n_705) );
INVx1_ASAP7_75t_L g726 ( .A(n_514), .Y(n_726) );
INVx1_ASAP7_75t_L g775 ( .A(n_514), .Y(n_775) );
AND2x2_ASAP7_75t_L g815 ( .A(n_514), .B(n_746), .Y(n_815) );
INVx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND2x2_ASAP7_75t_L g574 ( .A(n_515), .B(n_575), .Y(n_574) );
AND2x2_ASAP7_75t_L g718 ( .A(n_515), .B(n_531), .Y(n_718) );
AND2x2_ASAP7_75t_L g789 ( .A(n_515), .B(n_643), .Y(n_789) );
BUFx3_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g678 ( .A(n_516), .Y(n_678) );
OAI21x1_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_519), .B(n_527), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g689 ( .A(n_529), .B(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g706 ( .A(n_529), .B(n_677), .Y(n_706) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx1_ASAP7_75t_L g779 ( .A(n_530), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_545), .Y(n_530) );
INVx2_ASAP7_75t_L g575 ( .A(n_531), .Y(n_575) );
AND2x4_ASAP7_75t_SL g655 ( .A(n_531), .B(n_573), .Y(n_655) );
HB1xp67_ASAP7_75t_L g666 ( .A(n_531), .Y(n_666) );
INVx1_ASAP7_75t_L g680 ( .A(n_531), .Y(n_680) );
INVxp67_ASAP7_75t_L g747 ( .A(n_531), .Y(n_747) );
INVx1_ASAP7_75t_L g764 ( .A(n_531), .Y(n_764) );
BUFx6f_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
OAI21xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_536), .B(n_537), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
INVx2_ASAP7_75t_L g573 ( .A(n_545), .Y(n_573) );
INVx1_ASAP7_75t_L g643 ( .A(n_545), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_545), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g733 ( .A(n_545), .B(n_642), .Y(n_733) );
OR2x2_ASAP7_75t_L g768 ( .A(n_545), .B(n_560), .Y(n_768) );
AO21x2_ASAP7_75t_L g545 ( .A1(n_546), .A2(n_549), .B(n_555), .Y(n_545) );
NOR2xp67_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_552), .A2(n_553), .B(n_554), .Y(n_551) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_574), .Y(n_558) );
AND2x2_ASAP7_75t_L g715 ( .A(n_559), .B(n_716), .Y(n_715) );
BUFx3_ASAP7_75t_L g736 ( .A(n_559), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_559), .B(n_726), .Y(n_817) );
AND2x2_ASAP7_75t_L g559 ( .A(n_560), .B(n_573), .Y(n_559) );
INVx3_ASAP7_75t_L g642 ( .A(n_560), .Y(n_642) );
INVx1_ASAP7_75t_L g653 ( .A(n_560), .Y(n_653) );
AND2x2_ASAP7_75t_L g746 ( .A(n_560), .B(n_747), .Y(n_746) );
HB1xp67_ASAP7_75t_L g752 ( .A(n_560), .Y(n_752) );
INVx1_ASAP7_75t_L g813 ( .A(n_560), .Y(n_813) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_562), .Y(n_560) );
OAI21xp5_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_568), .B(n_571), .Y(n_562) );
BUFx2_ASAP7_75t_L g704 ( .A(n_573), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_574), .B(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g798 ( .A(n_574), .Y(n_798) );
AND2x2_ASAP7_75t_L g843 ( .A(n_574), .B(n_813), .Y(n_843) );
AND2x2_ASAP7_75t_L g786 ( .A(n_575), .B(n_678), .Y(n_786) );
NAND2xp5_ASAP7_75t_SL g576 ( .A(n_577), .B(n_593), .Y(n_576) );
INVx2_ASAP7_75t_L g659 ( .A(n_577), .Y(n_659) );
AND2x2_ASAP7_75t_L g719 ( .A(n_577), .B(n_669), .Y(n_719) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AND2x2_ASAP7_75t_L g702 ( .A(n_578), .B(n_650), .Y(n_702) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g708 ( .A(n_579), .B(n_627), .Y(n_708) );
OAI21xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_582), .B(n_592), .Y(n_579) );
OAI21x1_ASAP7_75t_L g608 ( .A1(n_580), .A2(n_609), .B(n_624), .Y(n_608) );
OAI21x1_ASAP7_75t_L g648 ( .A1(n_580), .A2(n_609), .B(n_624), .Y(n_648) );
OAI21x1_ASAP7_75t_L g673 ( .A1(n_580), .A2(n_582), .B(n_592), .Y(n_673) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OAI21x1_ASAP7_75t_L g582 ( .A1(n_583), .A2(n_588), .B(n_591), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_585), .B(n_587), .Y(n_583) );
AND2x2_ASAP7_75t_L g765 ( .A(n_593), .B(n_708), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_593), .B(n_659), .Y(n_776) );
AND2x2_ASAP7_75t_L g781 ( .A(n_593), .B(n_677), .Y(n_781) );
AND2x2_ASAP7_75t_L g795 ( .A(n_593), .B(n_702), .Y(n_795) );
AND2x2_ASAP7_75t_L g825 ( .A(n_593), .B(n_826), .Y(n_825) );
AND2x4_ASAP7_75t_L g593 ( .A(n_594), .B(n_607), .Y(n_593) );
INVx1_ASAP7_75t_L g809 ( .A(n_594), .Y(n_809) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g638 ( .A(n_595), .Y(n_638) );
INVx2_ASAP7_75t_L g661 ( .A(n_595), .Y(n_661) );
AND2x2_ASAP7_75t_L g669 ( .A(n_595), .B(n_608), .Y(n_669) );
AND2x2_ASAP7_75t_L g807 ( .A(n_595), .B(n_647), .Y(n_807) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND3xp33_ASAP7_75t_L g696 ( .A(n_597), .B(n_697), .C(n_698), .Y(n_696) );
NAND3xp33_ASAP7_75t_L g597 ( .A(n_598), .B(n_601), .C(n_605), .Y(n_597) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g660 ( .A(n_608), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_616), .Y(n_613) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx2_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_636), .Y(n_625) );
AND2x2_ASAP7_75t_L g662 ( .A(n_626), .B(n_646), .Y(n_662) );
HB1xp67_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
INVx2_ASAP7_75t_L g650 ( .A(n_627), .Y(n_650) );
AND2x2_ASAP7_75t_L g671 ( .A(n_627), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g783 ( .A(n_627), .Y(n_783) );
NAND2xp33_ASAP7_75t_L g698 ( .A(n_628), .B(n_699), .Y(n_698) );
NOR2xp33_ASAP7_75t_R g633 ( .A(n_634), .B(n_635), .Y(n_633) );
INVx2_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_637), .Y(n_722) );
AND2x2_ASAP7_75t_L g796 ( .A(n_637), .B(n_671), .Y(n_796) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
AND2x2_ASAP7_75t_L g649 ( .A(n_638), .B(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g663 ( .A(n_640), .B(n_664), .Y(n_663) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_649), .Y(n_644) );
AND2x2_ASAP7_75t_L g670 ( .A(n_645), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g701 ( .A(n_646), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g804 ( .A(n_646), .Y(n_804) );
BUFx3_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
BUFx3_ASAP7_75t_L g687 ( .A(n_648), .Y(n_687) );
AND2x4_ASAP7_75t_L g826 ( .A(n_650), .B(n_742), .Y(n_826) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_L g755 ( .A(n_652), .Y(n_755) );
AOI32xp33_ASAP7_75t_L g780 ( .A1(n_652), .A2(n_781), .A3(n_782), .B1(n_784), .B2(n_785), .Y(n_780) );
AND2x4_ASAP7_75t_L g822 ( .A(n_652), .B(n_779), .Y(n_822) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OR2x2_ASAP7_75t_L g763 ( .A(n_653), .B(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g729 ( .A(n_654), .Y(n_729) );
INVx2_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_L g684 ( .A(n_655), .B(n_677), .Y(n_684) );
AND2x2_ASAP7_75t_L g713 ( .A(n_655), .B(n_676), .Y(n_713) );
AND2x2_ASAP7_75t_L g751 ( .A(n_655), .B(n_752), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_667), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_658), .A2(n_662), .B(n_663), .Y(n_657) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AND2x2_ASAP7_75t_L g668 ( .A(n_659), .B(n_669), .Y(n_668) );
OR2x2_ASAP7_75t_L g838 ( .A(n_659), .B(n_770), .Y(n_838) );
AND2x2_ASAP7_75t_L g711 ( .A(n_660), .B(n_708), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g714 ( .A1(n_660), .A2(n_690), .B1(n_715), .B2(n_719), .Y(n_714) );
AND2x2_ASAP7_75t_L g784 ( .A(n_660), .B(n_671), .Y(n_784) );
AND2x2_ASAP7_75t_L g792 ( .A(n_660), .B(n_702), .Y(n_792) );
AND2x4_ASAP7_75t_SL g844 ( .A(n_660), .B(n_826), .Y(n_844) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVxp67_ASAP7_75t_L g732 ( .A(n_666), .Y(n_732) );
OAI21xp5_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_670), .B(n_674), .Y(n_667) );
AND2x2_ASAP7_75t_L g738 ( .A(n_669), .B(n_708), .Y(n_738) );
INVx1_ASAP7_75t_L g756 ( .A(n_669), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_671), .B(n_686), .Y(n_685) );
INVx2_ASAP7_75t_L g742 ( .A(n_672), .Y(n_742) );
INVx2_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVxp67_ASAP7_75t_L g694 ( .A(n_673), .Y(n_694) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OR2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AND2x2_ASAP7_75t_L g840 ( .A(n_677), .B(n_733), .Y(n_840) );
INVx2_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OR2x2_ASAP7_75t_L g774 ( .A(n_679), .B(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_709), .Y(n_681) );
OAI221xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B1(n_688), .B2(n_691), .C(n_700), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g707 ( .A(n_686), .B(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g744 ( .A(n_687), .Y(n_744) );
OR2x2_ASAP7_75t_L g770 ( .A(n_687), .B(n_696), .Y(n_770) );
INVx2_ASAP7_75t_SL g688 ( .A(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_695), .Y(n_692) );
INVx1_ASAP7_75t_L g757 ( .A(n_693), .Y(n_757) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
AND2x2_ASAP7_75t_L g749 ( .A(n_694), .B(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
OR2x2_ASAP7_75t_L g743 ( .A(n_696), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g750 ( .A(n_696), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B1(n_706), .B2(n_707), .Y(n_700) );
AND2x2_ASAP7_75t_L g721 ( .A(n_701), .B(n_722), .Y(n_721) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx1_ASAP7_75t_L g760 ( .A(n_704), .Y(n_760) );
AND2x2_ASAP7_75t_L g785 ( .A(n_704), .B(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g761 ( .A(n_705), .Y(n_761) );
AND2x2_ASAP7_75t_L g808 ( .A(n_708), .B(n_809), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_708), .B(n_830), .Y(n_829) );
AND2x2_ASAP7_75t_L g835 ( .A(n_708), .B(n_807), .Y(n_835) );
OAI21xp5_ASAP7_75t_SL g709 ( .A1(n_710), .A2(n_712), .B(n_714), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_713), .B(n_755), .Y(n_802) );
INVx2_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g812 ( .A(n_718), .B(n_813), .Y(n_812) );
AOI21xp5_ASAP7_75t_L g720 ( .A1(n_721), .A2(n_723), .B(n_734), .Y(n_720) );
NAND3xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .C(n_730), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_725), .Y(n_724) );
AND2x2_ASAP7_75t_L g766 ( .A(n_725), .B(n_767), .Y(n_766) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
HB1xp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g730 ( .A(n_731), .Y(n_730) );
AND2x2_ASAP7_75t_L g731 ( .A(n_732), .B(n_733), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_737), .B1(n_739), .B2(n_745), .C(n_748), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_740), .B(n_778), .Y(n_777) );
NOR2x1p5_ASAP7_75t_SL g740 ( .A(n_741), .B(n_743), .Y(n_740) );
AND2x2_ASAP7_75t_L g806 ( .A(n_741), .B(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_SL g820 ( .A(n_741), .B(n_781), .Y(n_820) );
INVx2_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
OAI21xp5_ASAP7_75t_L g827 ( .A1(n_749), .A2(n_828), .B(n_831), .Y(n_827) );
AOI322xp5_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_756), .A3(n_757), .B1(n_758), .B2(n_765), .C1(n_766), .C2(n_769), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_762), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
INVx1_ASAP7_75t_L g790 ( .A(n_762), .Y(n_790) );
BUFx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g794 ( .A(n_768), .Y(n_794) );
INVx1_ASAP7_75t_L g799 ( .A(n_768), .Y(n_799) );
INVx2_ASAP7_75t_L g832 ( .A(n_768), .Y(n_832) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_768), .B(n_786), .Y(n_837) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NOR2xp33_ASAP7_75t_L g816 ( .A(n_770), .B(n_817), .Y(n_816) );
NAND3xp33_ASAP7_75t_L g771 ( .A(n_772), .B(n_800), .C(n_818), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_773), .B(n_787), .Y(n_772) );
OAI211xp5_ASAP7_75t_L g773 ( .A1(n_774), .A2(n_776), .B(n_777), .C(n_780), .Y(n_773) );
INVx2_ASAP7_75t_L g842 ( .A(n_774), .Y(n_842) );
BUFx3_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
AOI221x1_ASAP7_75t_L g805 ( .A1(n_785), .A2(n_806), .B1(n_808), .B2(n_810), .C(n_816), .Y(n_805) );
AND2x2_ASAP7_75t_L g831 ( .A(n_786), .B(n_832), .Y(n_831) );
OAI21xp33_ASAP7_75t_SL g787 ( .A1(n_788), .A2(n_791), .B(n_793), .Y(n_787) );
NOR2xp33_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .Y(n_788) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_795), .B1(n_796), .B2(n_797), .Y(n_793) );
NAND2x1p5_ASAP7_75t_L g803 ( .A(n_796), .B(n_804), .Y(n_803) );
NOR2x1_ASAP7_75t_L g797 ( .A(n_798), .B(n_799), .Y(n_797) );
OA21x2_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B(n_805), .Y(n_800) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AOI21xp33_ASAP7_75t_SL g819 ( .A1(n_803), .A2(n_820), .B(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g830 ( .A(n_809), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_811), .B(n_814), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_812), .B(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g814 ( .A(n_815), .Y(n_814) );
NOR3xp33_ASAP7_75t_SL g818 ( .A(n_819), .B(n_823), .C(n_833), .Y(n_818) );
INVx1_ASAP7_75t_L g821 ( .A(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g823 ( .A(n_824), .B(n_827), .Y(n_823) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
OAI221xp5_ASAP7_75t_L g833 ( .A1(n_834), .A2(n_836), .B1(n_838), .B2(n_839), .C(n_841), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVxp67_ASAP7_75t_SL g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
OAI21xp33_ASAP7_75t_L g841 ( .A1(n_842), .A2(n_843), .B(n_844), .Y(n_841) );
NOR2xp33_ASAP7_75t_R g846 ( .A(n_847), .B(n_848), .Y(n_846) );
BUFx6f_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
BUFx6f_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_855), .Y(n_852) );
BUFx3_ASAP7_75t_L g853 ( .A(n_854), .Y(n_853) );
NAND2xp5_ASAP7_75t_SL g855 ( .A(n_856), .B(n_869), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_864), .Y(n_856) );
BUFx3_ASAP7_75t_L g857 ( .A(n_858), .Y(n_857) );
BUFx3_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
BUFx3_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx2_ASAP7_75t_L g860 ( .A(n_861), .Y(n_860) );
INVx2_ASAP7_75t_SL g872 ( .A(n_861), .Y(n_872) );
NOR2x1p5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
XNOR2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_868), .Y(n_864) );
INVxp67_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
NOR2xp67_ASAP7_75t_SL g870 ( .A(n_871), .B(n_873), .Y(n_870) );
BUFx2_ASAP7_75t_SL g871 ( .A(n_872), .Y(n_871) );
BUFx8_ASAP7_75t_SL g874 ( .A(n_875), .Y(n_874) );
BUFx6f_ASAP7_75t_SL g875 ( .A(n_876), .Y(n_875) );
BUFx4f_ASAP7_75t_L g890 ( .A(n_876), .Y(n_890) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
NAND2x1p5_ASAP7_75t_L g877 ( .A(n_878), .B(n_884), .Y(n_877) );
INVx1_ASAP7_75t_L g878 ( .A(n_879), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVxp67_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_886), .B(n_887), .Y(n_885) );
BUFx2_ASAP7_75t_L g888 ( .A(n_889), .Y(n_888) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_890), .Y(n_889) );
endmodule