module fake_jpeg_11241_n_553 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_553);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_553;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx8_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_12),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_1),
.B(n_8),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_3),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_14),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_15),
.Y(n_57)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_27),
.Y(n_58)
);

INVx1_ASAP7_75t_SL g209 ( 
.A(n_58),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_60),
.Y(n_126)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_63),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx5_ASAP7_75t_L g200 ( 
.A(n_64),
.Y(n_200)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_27),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g150 ( 
.A(n_65),
.Y(n_150)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_66),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

BUFx4f_ASAP7_75t_L g69 ( 
.A(n_27),
.Y(n_69)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_69),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_18),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_70),
.B(n_94),
.Y(n_127)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_40),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_73),
.B(n_82),
.Y(n_148)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_74),
.Y(n_166)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_75),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_78),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_19),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_79),
.Y(n_174)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_80),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_19),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_81),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_40),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_83),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_43),
.Y(n_85)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_32),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_86),
.B(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_87),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_88),
.Y(n_163)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_35),
.Y(n_89)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_89),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_40),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_91),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_92),
.Y(n_201)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_56),
.Y(n_93)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_93),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_52),
.B(n_18),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_95),
.Y(n_172)
);

BUFx8_ASAP7_75t_L g96 ( 
.A(n_37),
.Y(n_96)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_18),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_125),
.Y(n_138)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_43),
.Y(n_98)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_98),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_55),
.B(n_35),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_99),
.B(n_109),
.Y(n_136)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_100),
.Y(n_154)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_32),
.Y(n_101)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_102),
.Y(n_155)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_57),
.Y(n_103)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_103),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_31),
.Y(n_104)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_104),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx3_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_106),
.B(n_112),
.Y(n_161)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_34),
.Y(n_107)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_44),
.Y(n_108)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_108),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_55),
.B(n_17),
.Y(n_109)
);

INVx8_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_110),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_31),
.Y(n_111)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_40),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_113),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_34),
.Y(n_114)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_114),
.Y(n_192)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_28),
.Y(n_116)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_44),
.B(n_17),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_117),
.B(n_124),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_34),
.Y(n_118)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_118),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_23),
.Y(n_119)
);

NAND2xp33_ASAP7_75t_SL g193 ( 
.A(n_119),
.B(n_123),
.Y(n_193)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_39),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_122),
.Y(n_169)
);

INVx11_ASAP7_75t_L g121 ( 
.A(n_32),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_121),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_23),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_23),
.Y(n_123)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_30),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_30),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_24),
.B1(n_48),
.B2(n_42),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_128),
.A2(n_132),
.B1(n_134),
.B2(n_145),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_86),
.A2(n_30),
.B1(n_49),
.B2(n_45),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_101),
.A2(n_39),
.B1(n_48),
.B2(n_42),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_101),
.A2(n_39),
.B1(n_41),
.B2(n_53),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_137),
.A2(n_141),
.B1(n_167),
.B2(n_198),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_20),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_139),
.B(n_153),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_78),
.B(n_39),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_140),
.B(n_171),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_98),
.A2(n_53),
.B1(n_41),
.B2(n_24),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_36),
.C(n_49),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_144),
.B(n_182),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_111),
.A2(n_51),
.B1(n_45),
.B2(n_38),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_72),
.A2(n_51),
.B1(n_38),
.B2(n_36),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_149),
.A2(n_175),
.B1(n_186),
.B2(n_207),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_33),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_80),
.B(n_22),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_157),
.B(n_170),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_74),
.A2(n_67),
.B1(n_61),
.B2(n_110),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_165),
.A2(n_177),
.B1(n_203),
.B2(n_58),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_92),
.A2(n_33),
.B1(n_29),
.B2(n_22),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_95),
.B(n_29),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_60),
.B(n_20),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_83),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_76),
.A2(n_16),
.B1(n_15),
.B2(n_5),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_120),
.B(n_3),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_66),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_78),
.B(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_191),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_88),
.B(n_6),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_88),
.B(n_8),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_194),
.B(n_196),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_77),
.B(n_9),
.Y(n_195)
);

NAND3xp33_ASAP7_75t_L g242 ( 
.A(n_195),
.B(n_65),
.C(n_63),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_105),
.B(n_9),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_64),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_198)
);

OAI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_79),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_81),
.A2(n_10),
.B1(n_11),
.B2(n_125),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_124),
.A2(n_10),
.B1(n_11),
.B2(n_106),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g229 ( 
.A1(n_208),
.A2(n_105),
.B1(n_106),
.B2(n_63),
.Y(n_229)
);

INVx11_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_213),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_148),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_214),
.B(n_220),
.Y(n_293)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx4_ASAP7_75t_L g320 ( 
.A(n_215),
.Y(n_320)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_180),
.Y(n_216)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_176),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g331 ( 
.A(n_217),
.Y(n_331)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_147),
.Y(n_218)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_218),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_219),
.A2(n_222),
.B1(n_229),
.B2(n_236),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_126),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_164),
.Y(n_221)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_221),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_167),
.A2(n_119),
.B1(n_84),
.B2(n_118),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_138),
.B(n_114),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_223),
.B(n_246),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g224 ( 
.A(n_150),
.Y(n_224)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_155),
.Y(n_227)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_227),
.Y(n_294)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_143),
.Y(n_231)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_231),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_232),
.B(n_233),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_169),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_131),
.Y(n_235)
);

INVx6_ASAP7_75t_L g324 ( 
.A(n_235),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_L g236 ( 
.A1(n_167),
.A2(n_107),
.B1(n_122),
.B2(n_69),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_151),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_237),
.B(n_242),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_136),
.B(n_122),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_239),
.B(n_248),
.Y(n_308)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_159),
.Y(n_240)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_240),
.Y(n_330)
);

INVx11_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_241),
.Y(n_327)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_178),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_243),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_128),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_244),
.B(n_250),
.Y(n_318)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_192),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_245),
.B(n_247),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_152),
.B(n_127),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_212),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_173),
.B(n_179),
.Y(n_248)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_149),
.A2(n_203),
.B1(n_145),
.B2(n_134),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_249),
.A2(n_252),
.B1(n_276),
.B2(n_283),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_130),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_187),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_253),
.Y(n_321)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_208),
.A2(n_186),
.B1(n_175),
.B2(n_183),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_150),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_130),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_255),
.B(n_258),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_184),
.B(n_181),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_257),
.B(n_261),
.Y(n_326)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_183),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_202),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_259),
.B(n_262),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_172),
.A2(n_166),
.B1(n_205),
.B2(n_201),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_260),
.A2(n_266),
.B1(n_277),
.B2(n_278),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_197),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_205),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_263),
.Y(n_288)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_L g266 ( 
.A1(n_146),
.A2(n_185),
.B1(n_154),
.B2(n_189),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_210),
.B(n_172),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_267),
.B(n_270),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_156),
.B(n_163),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_268),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_202),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g306 ( 
.A(n_269),
.B(n_271),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_158),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_156),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_133),
.B(n_158),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_272),
.B(n_273),
.Y(n_334)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_133),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_163),
.B(n_190),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_274),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_142),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_275),
.Y(n_335)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_200),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_166),
.A2(n_201),
.B1(n_142),
.B2(n_189),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_168),
.A2(n_174),
.B1(n_206),
.B2(n_162),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_168),
.Y(n_279)
);

NAND2x1_ASAP7_75t_SL g302 ( 
.A(n_279),
.B(n_280),
.Y(n_302)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_206),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_190),
.Y(n_281)
);

NAND2x1_ASAP7_75t_SL g332 ( 
.A(n_281),
.B(n_284),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_174),
.Y(n_283)
);

INVx4_ASAP7_75t_L g284 ( 
.A(n_160),
.Y(n_284)
);

MAJx2_ASAP7_75t_L g287 ( 
.A(n_246),
.B(n_129),
.C(n_200),
.Y(n_287)
);

MAJx2_ASAP7_75t_L g370 ( 
.A(n_287),
.B(n_315),
.C(n_322),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_219),
.A2(n_254),
.B1(n_244),
.B2(n_223),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_313),
.B1(n_235),
.B2(n_303),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_256),
.A2(n_199),
.B1(n_204),
.B2(n_129),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_296),
.A2(n_304),
.B1(n_309),
.B2(n_338),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_234),
.B(n_199),
.C(n_131),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_301),
.B(n_314),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_282),
.A2(n_204),
.B1(n_270),
.B2(n_254),
.Y(n_304)
);

OA22x2_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_260),
.B1(n_232),
.B2(n_277),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_305),
.B(n_297),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_267),
.A2(n_272),
.B1(n_279),
.B2(n_243),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_225),
.A2(n_253),
.B(n_264),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_228),
.A2(n_226),
.B1(n_238),
.B2(n_231),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_220),
.B(n_214),
.C(n_227),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_273),
.B(n_247),
.C(n_240),
.Y(n_315)
);

OAI32xp33_ASAP7_75t_L g319 ( 
.A1(n_265),
.A2(n_280),
.A3(n_216),
.B1(n_258),
.B2(n_213),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_319),
.B(n_276),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g322 ( 
.A1(n_245),
.A2(n_218),
.B(n_281),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_241),
.A2(n_259),
.B(n_224),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g348 ( 
.A(n_323),
.Y(n_348)
);

FAx1_ASAP7_75t_L g337 ( 
.A(n_221),
.B(n_230),
.CI(n_284),
.CON(n_337),
.SN(n_337)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_337),
.B(n_217),
.Y(n_340)
);

AOI22x1_ASAP7_75t_L g338 ( 
.A1(n_263),
.A2(n_283),
.B1(n_255),
.B2(n_250),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_339),
.A2(n_340),
.B(n_345),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_304),
.A2(n_275),
.B1(n_215),
.B2(n_235),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_341),
.A2(n_342),
.B1(n_349),
.B2(n_362),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_317),
.A2(n_235),
.B1(n_328),
.B2(n_295),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_344),
.B(n_347),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_326),
.B(n_312),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_317),
.A2(n_328),
.B1(n_291),
.B2(n_309),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_297),
.A2(n_334),
.B1(n_337),
.B2(n_291),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_350),
.A2(n_363),
.B1(n_378),
.B2(n_333),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_334),
.B(n_314),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_351),
.B(n_359),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_312),
.Y(n_352)
);

CKINVDCx14_ASAP7_75t_R g407 ( 
.A(n_352),
.Y(n_407)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_324),
.Y(n_353)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_353),
.Y(n_380)
);

BUFx24_ASAP7_75t_SL g354 ( 
.A(n_293),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_354),
.B(n_355),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_331),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_298),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_356),
.B(n_358),
.Y(n_409)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_316),
.Y(n_357)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_357),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_292),
.B(n_308),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_292),
.B(n_299),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_316),
.Y(n_360)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_294),
.Y(n_361)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_361),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g362 ( 
.A1(n_318),
.A2(n_337),
.B1(n_310),
.B2(n_301),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_337),
.A2(n_305),
.B1(n_313),
.B2(n_319),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_305),
.A2(n_287),
.B1(n_300),
.B2(n_306),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_364),
.A2(n_371),
.B1(n_373),
.B2(n_290),
.Y(n_403)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_320),
.Y(n_365)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_365),
.Y(n_396)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_294),
.Y(n_366)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_366),
.Y(n_397)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_298),
.Y(n_367)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_321),
.B(n_336),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_289),
.B(n_306),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_369),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_305),
.A2(n_338),
.B1(n_329),
.B2(n_315),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_298),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_L g392 ( 
.A1(n_372),
.A2(n_375),
.B(n_376),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_338),
.A2(n_329),
.B1(n_325),
.B2(n_335),
.Y(n_373)
);

BUFx24_ASAP7_75t_SL g374 ( 
.A(n_289),
.Y(n_374)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_322),
.B(n_333),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_302),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_302),
.B(n_332),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_377),
.B(n_332),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_311),
.A2(n_335),
.B1(n_285),
.B2(n_302),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_340),
.A2(n_323),
.B(n_332),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_SL g424 ( 
.A1(n_381),
.A2(n_403),
.B(n_377),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_382),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g425 ( 
.A1(n_383),
.A2(n_400),
.B1(n_408),
.B2(n_343),
.Y(n_425)
);

MAJx2_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_285),
.C(n_330),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_386),
.B(n_393),
.Y(n_416)
);

XOR2xp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_330),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_389),
.B(n_364),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_379),
.B(n_288),
.C(n_311),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_370),
.B(n_288),
.C(n_307),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_394),
.B(n_395),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_370),
.B(n_307),
.C(n_286),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_370),
.B(n_286),
.C(n_327),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_399),
.B(n_362),
.Y(n_434)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_345),
.A2(n_320),
.B1(n_290),
.B2(n_327),
.Y(n_400)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_357),
.Y(n_402)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_402),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_346),
.A2(n_324),
.B1(n_341),
.B2(n_373),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_406),
.A2(n_371),
.B1(n_343),
.B2(n_342),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g408 ( 
.A1(n_350),
.A2(n_363),
.B1(n_344),
.B2(n_339),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_360),
.Y(n_410)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_410),
.Y(n_418)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_411),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_349),
.Y(n_414)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_414),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_415),
.B(n_389),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_419),
.A2(n_437),
.B(n_380),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_409),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_420),
.B(n_421),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_405),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_424),
.A2(n_381),
.B(n_392),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_425),
.A2(n_441),
.B1(n_397),
.B2(n_402),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_359),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_426),
.Y(n_447)
);

OR2x2_ASAP7_75t_L g427 ( 
.A(n_387),
.B(n_375),
.Y(n_427)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_427),
.Y(n_456)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_429),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_413),
.B(n_376),
.Y(n_430)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_430),
.Y(n_461)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_384),
.Y(n_431)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_431),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_412),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_432),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g433 ( 
.A(n_388),
.B(n_347),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g444 ( 
.A(n_433),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_434),
.B(n_393),
.C(n_399),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g435 ( 
.A(n_391),
.B(n_352),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_435),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g436 ( 
.A1(n_404),
.A2(n_348),
.B1(n_378),
.B2(n_356),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_436),
.A2(n_439),
.B1(n_380),
.B2(n_396),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_408),
.A2(n_348),
.B1(n_372),
.B2(n_367),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_385),
.Y(n_438)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_438),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_403),
.A2(n_368),
.B1(n_366),
.B2(n_355),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_391),
.B(n_365),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g462 ( 
.A(n_440),
.B(n_410),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_398),
.B(n_353),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_SL g442 ( 
.A(n_398),
.B(n_392),
.Y(n_442)
);

NOR2xp67_ASAP7_75t_L g457 ( 
.A(n_442),
.B(n_411),
.Y(n_457)
);

XOR2xp5_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_446),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g446 ( 
.A(n_416),
.B(n_395),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_448),
.B(n_465),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_394),
.C(n_386),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_449),
.B(n_458),
.C(n_427),
.Y(n_476)
);

OAI22x1_ASAP7_75t_L g451 ( 
.A1(n_425),
.A2(n_404),
.B1(n_387),
.B2(n_383),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g472 ( 
.A1(n_451),
.A2(n_455),
.B1(n_468),
.B2(n_419),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g479 ( 
.A(n_452),
.B(n_463),
.Y(n_479)
);

XOR2x2_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_382),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_454),
.B(n_422),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_439),
.A2(n_400),
.B1(n_385),
.B2(n_390),
.Y(n_455)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_457),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_423),
.B(n_390),
.C(n_397),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g473 ( 
.A1(n_460),
.A2(n_436),
.B1(n_442),
.B2(n_432),
.Y(n_473)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_462),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_416),
.B(n_434),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_466),
.B(n_421),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_475),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_481),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g493 ( 
.A1(n_473),
.A2(n_468),
.B1(n_445),
.B2(n_456),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_446),
.B(n_437),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_474),
.B(n_476),
.C(n_488),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g475 ( 
.A(n_444),
.B(n_426),
.Y(n_475)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_461),
.Y(n_477)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_477),
.Y(n_490)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_461),
.Y(n_478)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_478),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_450),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_480),
.B(n_482),
.Y(n_503)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_453),
.A2(n_420),
.B1(n_414),
.B2(n_427),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_464),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_464),
.Y(n_483)
);

BUFx12_ASAP7_75t_L g491 ( 
.A(n_483),
.Y(n_491)
);

BUFx12f_ASAP7_75t_SL g502 ( 
.A(n_484),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_L g485 ( 
.A1(n_444),
.A2(n_430),
.B1(n_440),
.B2(n_417),
.Y(n_485)
);

INVxp33_ASAP7_75t_SL g497 ( 
.A(n_485),
.Y(n_497)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_448),
.B(n_424),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_447),
.B(n_458),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_489),
.A2(n_449),
.B(n_452),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_493),
.A2(n_496),
.B1(n_504),
.B2(n_505),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_494),
.B(n_499),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_473),
.A2(n_456),
.B1(n_445),
.B2(n_455),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_487),
.B(n_465),
.C(n_443),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g500 ( 
.A(n_487),
.B(n_462),
.C(n_463),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_500),
.B(n_486),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_469),
.A2(n_451),
.B1(n_422),
.B2(n_467),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_469),
.A2(n_477),
.B1(n_478),
.B2(n_471),
.Y(n_505)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_492),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_SL g520 ( 
.A(n_506),
.B(n_502),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_494),
.A2(n_476),
.B(n_479),
.Y(n_508)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_508),
.A2(n_510),
.B(n_516),
.Y(n_524)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_498),
.A2(n_482),
.B1(n_483),
.B2(n_467),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_509),
.B(n_512),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_498),
.A2(n_479),
.B(n_471),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_503),
.Y(n_511)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_511),
.B(n_513),
.Y(n_519)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_501),
.Y(n_513)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_497),
.A2(n_479),
.B1(n_474),
.B2(n_459),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_514),
.B(n_518),
.Y(n_526)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_499),
.B(n_486),
.Y(n_515)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_515),
.B(n_454),
.Y(n_529)
);

OAI21xp5_ASAP7_75t_L g516 ( 
.A1(n_496),
.A2(n_441),
.B(n_459),
.Y(n_516)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_493),
.A2(n_505),
.B1(n_504),
.B2(n_490),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_522),
.Y(n_534)
);

XOR2xp5_ASAP7_75t_L g522 ( 
.A(n_514),
.B(n_500),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_495),
.C(n_488),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_523),
.B(n_525),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_507),
.B(n_401),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g527 ( 
.A(n_517),
.B(n_401),
.Y(n_527)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_527),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_510),
.B(n_495),
.C(n_501),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_528),
.A2(n_517),
.B(n_516),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_429),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_530),
.B(n_532),
.Y(n_539)
);

OAI22xp5_ASAP7_75t_SL g532 ( 
.A1(n_526),
.A2(n_518),
.B1(n_502),
.B2(n_418),
.Y(n_532)
);

MAJx2_ASAP7_75t_L g533 ( 
.A(n_528),
.B(n_491),
.C(n_417),
.Y(n_533)
);

XNOR2xp5_ASAP7_75t_L g542 ( 
.A(n_533),
.B(n_537),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_521),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_535),
.B(n_418),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g538 ( 
.A(n_531),
.B(n_523),
.Y(n_538)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_538),
.A2(n_540),
.B(n_541),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_534),
.B(n_522),
.C(n_524),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_535),
.B(n_519),
.C(n_529),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g545 ( 
.A1(n_543),
.A2(n_536),
.B(n_428),
.Y(n_545)
);

HAxp5_ASAP7_75t_SL g544 ( 
.A(n_539),
.B(n_533),
.CON(n_544),
.SN(n_544)
);

OAI21xp33_ASAP7_75t_SL g549 ( 
.A1(n_544),
.A2(n_542),
.B(n_491),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g548 ( 
.A1(n_545),
.A2(n_547),
.B(n_431),
.Y(n_548)
);

OAI21xp5_ASAP7_75t_L g547 ( 
.A1(n_543),
.A2(n_491),
.B(n_428),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g550 ( 
.A1(n_548),
.A2(n_549),
.B(n_546),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_550),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_551),
.B(n_438),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_552),
.B(n_396),
.Y(n_553)
);


endmodule