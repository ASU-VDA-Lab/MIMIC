module real_jpeg_4550_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_1),
.A2(n_52),
.B1(n_113),
.B2(n_116),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_1),
.A2(n_52),
.B1(n_194),
.B2(n_197),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_1),
.B(n_67),
.Y(n_291)
);

O2A1O1Ixp33_ASAP7_75t_L g348 ( 
.A1(n_1),
.A2(n_70),
.B(n_349),
.C(n_351),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_1),
.B(n_99),
.C(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_1),
.B(n_21),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_1),
.B(n_192),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_1),
.B(n_101),
.Y(n_413)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_2),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_2),
.Y(n_108)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_2),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_3),
.A2(n_233),
.B1(n_234),
.B2(n_235),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_3),
.Y(n_234)
);

OAI22xp33_ASAP7_75t_SL g255 ( 
.A1(n_3),
.A2(n_234),
.B1(n_256),
.B2(n_258),
.Y(n_255)
);

OAI22xp33_ASAP7_75t_SL g360 ( 
.A1(n_3),
.A2(n_234),
.B1(n_361),
.B2(n_363),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_3),
.A2(n_234),
.B1(n_384),
.B2(n_386),
.Y(n_383)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_5),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_5),
.Y(n_192)
);

INVx8_ASAP7_75t_L g297 ( 
.A(n_5),
.Y(n_297)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_6),
.Y(n_269)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_8),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_9),
.Y(n_66)
);

BUFx5_ASAP7_75t_L g79 ( 
.A(n_9),
.Y(n_79)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_9),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g141 ( 
.A(n_9),
.Y(n_141)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_9),
.Y(n_237)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_10),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_10),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_11),
.A2(n_78),
.B1(n_80),
.B2(n_82),
.Y(n_77)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_11),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_11),
.A2(n_82),
.B1(n_145),
.B2(n_149),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_11),
.A2(n_82),
.B1(n_116),
.B2(n_200),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_11),
.A2(n_82),
.B1(n_282),
.B2(n_284),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_12),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_13),
.A2(n_59),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_13),
.A2(n_71),
.B1(n_85),
.B2(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_13),
.A2(n_85),
.B1(n_175),
.B2(n_177),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_13),
.A2(n_85),
.B1(n_107),
.B2(n_224),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_446),
.B(n_449),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_156),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_154),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_129),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_18),
.B(n_129),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_54),
.B1(n_55),
.B2(n_87),
.Y(n_19)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_20),
.A2(n_87),
.B1(n_320),
.B2(n_321),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_34),
.B(n_49),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_21),
.B(n_123),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_21),
.A2(n_121),
.B(n_144),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_21),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_22),
.B(n_36),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_22),
.B(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_27),
.B1(n_29),
.B2(n_32),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g350 ( 
.A(n_25),
.Y(n_350)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_26),
.Y(n_40)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_26),
.Y(n_353)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_28),
.Y(n_31)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_28),
.Y(n_178)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_28),
.Y(n_362)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_30),
.Y(n_373)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_31),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_31),
.Y(n_176)
);

INVx6_ASAP7_75t_L g365 ( 
.A(n_31),
.Y(n_365)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_34),
.A2(n_144),
.B(n_152),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_34),
.B(n_49),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_34),
.B(n_255),
.Y(n_289)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_35),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_41),
.B1(n_44),
.B2(n_47),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_43),
.Y(n_148)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_48),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_48),
.Y(n_266)
);

INVxp67_ASAP7_75t_SL g120 ( 
.A(n_49),
.Y(n_120)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_50),
.Y(n_53)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx6_ASAP7_75t_L g277 ( 
.A(n_51),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_52),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_52),
.B(n_141),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_L g351 ( 
.A1(n_52),
.A2(n_352),
.B(n_354),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_77),
.B(n_83),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_56),
.A2(n_127),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_57),
.B(n_84),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_57),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_57),
.B(n_232),
.Y(n_231)
);

NOR2x1_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_67),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_62),
.B2(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_61),
.Y(n_63)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_67),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_67),
.B(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_67),
.B(n_232),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_72),
.B2(n_75),
.Y(n_67)
);

INVx6_ASAP7_75t_L g279 ( 
.A(n_68),
.Y(n_279)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_77),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_81),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_83),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_83),
.B(n_231),
.Y(n_309)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_86),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_87),
.B(n_318),
.C(n_320),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_118),
.C(n_125),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_89),
.A2(n_118),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_89),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_89),
.A2(n_135),
.B1(n_143),
.B2(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_89),
.A2(n_135),
.B1(n_252),
.B2(n_259),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_89),
.B(n_249),
.C(n_252),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_110),
.B(n_111),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_90),
.A2(n_199),
.B(n_203),
.Y(n_198)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_91),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_91),
.B(n_112),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_91),
.B(n_360),
.Y(n_359)
);

NOR2x1_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_101),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx4_ASAP7_75t_SL g109 ( 
.A(n_99),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_101),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_101),
.B(n_174),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g378 ( 
.A(n_101),
.B(n_360),
.Y(n_378)
);

AO22x1_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_104),
.B1(n_107),
.B2(n_109),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx3_ASAP7_75t_SL g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_106),
.Y(n_186)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_106),
.Y(n_286)
);

INVx3_ASAP7_75t_L g376 ( 
.A(n_106),
.Y(n_376)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_108),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_110),
.B(n_111),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_110),
.A2(n_173),
.B(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_114),
.Y(n_202)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_115),
.Y(n_355)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_121),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g311 ( 
.A(n_119),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_121),
.Y(n_253)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_125),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_128),
.B(n_250),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_136),
.C(n_142),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_130),
.A2(n_131),
.B1(n_136),
.B2(n_164),
.Y(n_240)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_135),
.B(n_136),
.C(n_143),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_164),
.B1(n_165),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_137),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_138),
.Y(n_206)
);

INVxp33_ASAP7_75t_L g272 ( 
.A(n_140),
.Y(n_272)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_141),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_142),
.B(n_240),
.Y(n_239)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx5_ASAP7_75t_L g257 ( 
.A(n_151),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_153),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_153),
.B(n_289),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_242),
.B(n_442),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_238),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_207),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_160),
.B(n_207),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_180),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_162),
.A2(n_163),
.B1(n_168),
.B2(n_169),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_163),
.B(n_168),
.C(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_169),
.A2(n_170),
.B(n_179),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_170),
.B(n_179),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_171),
.Y(n_358)
);

INVxp67_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_173),
.B(n_378),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_204),
.B(n_205),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_181),
.A2(n_182),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_198),
.Y(n_182)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_183),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_183),
.A2(n_204),
.B1(n_205),
.B2(n_211),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_183),
.A2(n_198),
.B1(n_204),
.B2(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_183),
.B(n_348),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g424 ( 
.A1(n_183),
.A2(n_204),
.B1(n_348),
.B2(n_425),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_189),
.B(n_193),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_184),
.B(n_193),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_184),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_184),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_187),
.Y(n_184)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_188),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_190),
.A2(n_222),
.B(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_194),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g283 ( 
.A(n_195),
.Y(n_283)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g385 ( 
.A(n_196),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_198),
.Y(n_330)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AND2x2_ASAP7_75t_SL g304 ( 
.A(n_203),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_203),
.B(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_205),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_214),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_208),
.A2(n_212),
.B1(n_213),
.B2(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_208),
.Y(n_334)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_214),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_227),
.C(n_229),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_215),
.A2(n_216),
.B1(n_327),
.B2(n_328),
.Y(n_326)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_226),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_217),
.B(n_226),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_221),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_218),
.B(n_381),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_220),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_221),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_223),
.B(n_295),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_225),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_227),
.B(n_229),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_228),
.B(n_254),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_238),
.A2(n_444),
.B(n_445),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_239),
.B(n_241),
.Y(n_445)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_434),
.Y(n_243)
);

NAND3xp33_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_323),
.C(n_338),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_312),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_298),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_247),
.B(n_298),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_260),
.C(n_287),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_248),
.B(n_341),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_251),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_252),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_254),
.Y(n_252)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_256),
.Y(n_258)
);

INVx6_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_260),
.A2(n_261),
.B1(n_287),
.B2(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_280),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_262),
.B(n_280),
.Y(n_307)
);

AOI32xp33_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_267),
.A3(n_270),
.B1(n_272),
.B2(n_273),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx4_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx5_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp33_ASAP7_75t_SL g273 ( 
.A(n_274),
.B(n_278),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_294),
.B(n_303),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_284),
.Y(n_386)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_287),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_288),
.B(n_345),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_311),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_346),
.Y(n_345)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_292),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_293),
.B(n_398),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_294),
.B(n_382),
.Y(n_412)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_297),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_306),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_301),
.C(n_306),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_304),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_378),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_309),
.C(n_310),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g436 ( 
.A1(n_312),
.A2(n_437),
.B(n_438),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_322),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_313),
.B(n_322),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_314),
.B(n_316),
.C(n_317),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_319),
.Y(n_317)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_320),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_335),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_324),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_332),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_325),
.B(n_332),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_329),
.C(n_331),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_329),
.CI(n_331),
.CON(n_336),
.SN(n_336)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_335),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_336),
.B(n_337),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_336),
.B(n_337),
.Y(n_439)
);

BUFx24_ASAP7_75t_SL g452 ( 
.A(n_336),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_339),
.A2(n_366),
.B(n_433),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_340),
.B(n_343),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_340),
.B(n_343),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_347),
.C(n_356),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_344),
.B(n_429),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_347),
.A2(n_356),
.B1(n_357),
.B2(n_430),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_347),
.Y(n_430)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_348),
.Y(n_425)
);

INVx8_ASAP7_75t_L g349 ( 
.A(n_350),
.Y(n_349)
);

INVx6_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_359),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_367),
.A2(n_427),
.B(n_432),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_368),
.A2(n_417),
.B(n_426),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g368 ( 
.A1(n_369),
.A2(n_392),
.B(n_416),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_379),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_370),
.B(n_379),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_377),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_371),
.A2(n_372),
.B1(n_377),
.B2(n_395),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_372),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_374),
.Y(n_372)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_377),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_387),
.Y(n_379)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_383),
.B(n_399),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_388),
.A2(n_389),
.B1(n_390),
.B2(n_391),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_388),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_389),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_390),
.C(n_419),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_393),
.A2(n_401),
.B(n_415),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_396),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_396),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g401 ( 
.A1(n_402),
.A2(n_411),
.B(n_414),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_410),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_404),
.B(n_409),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_412),
.B(n_413),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_420),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_418),
.B(n_420),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_422),
.B(n_423),
.C(n_424),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_428),
.B(n_431),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_431),
.Y(n_432)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g434 ( 
.A1(n_435),
.A2(n_436),
.B(n_439),
.C(n_440),
.D(n_441),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

BUFx4f_ASAP7_75t_SL g446 ( 
.A(n_447),
.Y(n_446)
);

INVx13_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx8_ASAP7_75t_L g450 ( 
.A(n_448),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);


endmodule