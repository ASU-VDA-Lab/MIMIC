module fake_jpeg_18473_n_328 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_328);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_328;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_13),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

CKINVDCx9p33_ASAP7_75t_R g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_27),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_38),
.Y(n_44)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_30),
.C(n_19),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_42),
.Y(n_79)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_55),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_25),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_51),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_59),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_56),
.A2(n_22),
.B(n_20),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_61),
.A2(n_25),
.B(n_17),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_15),
.B1(n_28),
.B2(n_18),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_50),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_63),
.B(n_77),
.Y(n_113)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_64),
.B(n_70),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_43),
.A2(n_39),
.B1(n_18),
.B2(n_30),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_65),
.A2(n_73),
.B1(n_79),
.B2(n_85),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_32),
.B1(n_18),
.B2(n_31),
.Y(n_67)
);

OAI22x1_ASAP7_75t_L g95 ( 
.A1(n_67),
.A2(n_41),
.B1(n_38),
.B2(n_27),
.Y(n_95)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_54),
.Y(n_69)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_69),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g70 ( 
.A(n_49),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_71),
.B(n_21),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_39),
.B1(n_42),
.B2(n_40),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_83),
.Y(n_93)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_78),
.Y(n_90)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_48),
.Y(n_80)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_38),
.B1(n_42),
.B2(n_40),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_81),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_82),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_37),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_52),
.A2(n_42),
.B1(n_40),
.B2(n_37),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_37),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_41),
.Y(n_118)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_57),
.A2(n_15),
.B(n_28),
.C(n_27),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_40),
.Y(n_99)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_99),
.B(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_77),
.B1(n_76),
.B2(n_33),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_98),
.B(n_102),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_118),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_60),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_106),
.A2(n_109),
.B1(n_85),
.B2(n_73),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_107),
.Y(n_122)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_62),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_74),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_110),
.Y(n_123)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_87),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_111),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_112),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_32),
.B1(n_33),
.B2(n_15),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_93),
.B(n_79),
.C(n_66),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_135),
.Y(n_153)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_104),
.A2(n_79),
.B1(n_61),
.B2(n_81),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_125),
.A2(n_126),
.B1(n_140),
.B2(n_109),
.Y(n_158)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_132),
.A2(n_105),
.B(n_41),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_133),
.A2(n_137),
.B1(n_141),
.B2(n_147),
.Y(n_174)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_117),
.Y(n_134)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_93),
.B(n_65),
.C(n_64),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_84),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_136),
.B(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_94),
.A2(n_63),
.B1(n_89),
.B2(n_88),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_21),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_146),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_101),
.B(n_69),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_139),
.B(n_147),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_104),
.A2(n_35),
.B1(n_41),
.B2(n_28),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_94),
.A2(n_35),
.B1(n_33),
.B2(n_32),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_72),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_100),
.B(n_72),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_35),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_148),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_132),
.A2(n_92),
.B(n_112),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_149),
.A2(n_154),
.B(n_160),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_95),
.B(n_96),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_118),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_156),
.B(n_177),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_158),
.A2(n_122),
.B1(n_129),
.B2(n_141),
.Y(n_183)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_159),
.B(n_165),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_144),
.A2(n_96),
.B(n_114),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_103),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_162),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_128),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_133),
.A2(n_103),
.B1(n_110),
.B2(n_108),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_163),
.A2(n_174),
.B1(n_17),
.B2(n_20),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_137),
.A2(n_100),
.B(n_111),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_164),
.A2(n_168),
.B(n_23),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_128),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_105),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_169),
.B(n_170),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_120),
.B(n_106),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g172 ( 
.A(n_125),
.B(n_27),
.C(n_91),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_172),
.B(n_123),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_135),
.B(n_59),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_173),
.B(n_176),
.Y(n_205)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_138),
.B(n_31),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_27),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g178 ( 
.A(n_124),
.Y(n_178)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_131),
.Y(n_179)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_179),
.Y(n_201)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_134),
.Y(n_180)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_180),
.Y(n_204)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g196 ( 
.A(n_181),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_202),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_189),
.B1(n_200),
.B2(n_161),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_122),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_184),
.B(n_186),
.Y(n_232)
);

OAI32xp33_ASAP7_75t_L g185 ( 
.A1(n_181),
.A2(n_127),
.A3(n_123),
.B1(n_17),
.B2(n_23),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_185),
.B(n_198),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_153),
.B(n_148),
.C(n_130),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_187),
.B(n_208),
.C(n_209),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g216 ( 
.A1(n_190),
.A2(n_172),
.B(n_157),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_191),
.A2(n_195),
.B1(n_199),
.B2(n_175),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_174),
.A2(n_22),
.B1(n_26),
.B2(n_24),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_171),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_170),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_150),
.A2(n_25),
.B1(n_26),
.B2(n_24),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_154),
.A2(n_21),
.B(n_27),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_164),
.A2(n_7),
.B(n_14),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_203),
.B(n_206),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_7),
.B(n_14),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_156),
.B(n_19),
.C(n_8),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_173),
.B(n_19),
.C(n_6),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_210),
.Y(n_214)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_178),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_212),
.B(n_152),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_0),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_213),
.A2(n_166),
.B(n_167),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_235),
.B(n_207),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_217),
.A2(n_218),
.B1(n_236),
.B2(n_207),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_196),
.A2(n_150),
.B1(n_169),
.B2(n_171),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_192),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_220),
.B(n_221),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_201),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_222),
.B(n_224),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_223),
.A2(n_189),
.B1(n_200),
.B2(n_213),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_225),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_177),
.Y(n_226)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_229),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_187),
.B(n_155),
.C(n_179),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_6),
.C(n_13),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_180),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_233),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_199),
.B(n_166),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_234),
.B(n_237),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_167),
.B1(n_178),
.B2(n_2),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_193),
.B(n_6),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_238),
.B(n_208),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_232),
.B(n_184),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_240),
.B(n_242),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_241),
.A2(n_248),
.B1(n_215),
.B2(n_217),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_232),
.B(n_193),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_197),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_245),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_219),
.B(n_197),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_247),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_216),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_215),
.A2(n_213),
.B1(n_191),
.B2(n_185),
.Y(n_248)
);

NOR3xp33_ASAP7_75t_SL g250 ( 
.A(n_231),
.B(n_195),
.C(n_198),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_250),
.B(n_252),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_251),
.A2(n_214),
.B1(n_224),
.B2(n_222),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_254),
.B(n_257),
.C(n_229),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_219),
.B(n_13),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_260),
.Y(n_279)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_261),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_263),
.B(n_268),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_249),
.Y(n_264)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_264),
.Y(n_289)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_256),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_266),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_237),
.C(n_233),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_269),
.C(n_245),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_255),
.A2(n_220),
.B(n_227),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_240),
.C(n_242),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_273),
.B1(n_225),
.B2(n_272),
.Y(n_290)
);

FAx1_ASAP7_75t_SL g273 ( 
.A(n_247),
.B(n_218),
.CI(n_221),
.CON(n_273),
.SN(n_273)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_274),
.Y(n_286)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_259),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_275),
.B(n_276),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_214),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_254),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_277),
.Y(n_278)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_278),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_262),
.A2(n_244),
.B1(n_236),
.B2(n_235),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_281),
.A2(n_9),
.B1(n_1),
.B2(n_2),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_272),
.C(n_265),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_257),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_287),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_226),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_292),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_291),
.B(n_263),
.Y(n_294)
);

FAx1_ASAP7_75t_SL g292 ( 
.A(n_267),
.B(n_14),
.CI(n_12),
.CON(n_292),
.SN(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_269),
.C(n_265),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_297),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_294),
.A2(n_304),
.B(n_289),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_282),
.B(n_273),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_303),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_296),
.B(n_299),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_12),
.C(n_11),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_285),
.B(n_9),
.C(n_1),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_302),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_284),
.B(n_9),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_280),
.B(n_0),
.Y(n_304)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_293),
.B(n_279),
.Y(n_306)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_306),
.Y(n_315)
);

A2O1A1Ixp33_ASAP7_75t_SL g307 ( 
.A1(n_301),
.A2(n_278),
.B(n_286),
.C(n_290),
.Y(n_307)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_307),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_288),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_308),
.B(n_309),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_310),
.B(n_292),
.Y(n_316)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_313),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g322 ( 
.A1(n_318),
.A2(n_319),
.B(n_307),
.Y(n_322)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_300),
.C(n_299),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_317),
.A2(n_315),
.B1(n_312),
.B2(n_314),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_321),
.B(n_322),
.Y(n_323)
);

AOI21x1_ASAP7_75t_L g324 ( 
.A1(n_323),
.A2(n_320),
.B(n_2),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_324),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_4),
.C(n_5),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_326),
.A2(n_4),
.B1(n_5),
.B2(n_284),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_327),
.B(n_5),
.Y(n_328)
);


endmodule