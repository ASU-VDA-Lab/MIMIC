module fake_jpeg_5376_n_78 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_78);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_78;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_48;
wire n_35;
wire n_46;
wire n_36;
wire n_62;
wire n_43;

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_SL g37 ( 
.A(n_14),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_23),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g42 ( 
.A(n_29),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

BUFx8_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_13),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_39),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_50),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_49),
.B(n_52),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_41),
.B(n_1),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_2),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_51),
.B(n_53),
.Y(n_54)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_50),
.A2(n_43),
.B1(n_46),
.B2(n_34),
.Y(n_55)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_59),
.B(n_6),
.C(n_15),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_52),
.A2(n_36),
.B1(n_33),
.B2(n_8),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_16),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_52),
.A2(n_38),
.B1(n_35),
.B2(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_4),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g62 ( 
.A(n_60),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_58),
.A2(n_47),
.B(n_9),
.C(n_10),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_64),
.Y(n_68)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

BUFx4f_ASAP7_75t_SL g65 ( 
.A(n_62),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_54),
.B1(n_56),
.B2(n_20),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_69),
.B(n_66),
.C(n_68),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_71),
.B(n_70),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_72),
.B(n_17),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_19),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_24),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_75),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_76),
.B(n_25),
.C(n_26),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_28),
.Y(n_78)
);


endmodule