module fake_jpeg_28566_n_122 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_122);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_122;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_12),
.Y(n_13)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx10_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

INVx2_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g47 ( 
.A1(n_29),
.A2(n_26),
.B(n_21),
.Y(n_47)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_23),
.B(n_0),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_35),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_20),
.Y(n_34)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_13),
.B(n_6),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_36),
.B(n_17),
.Y(n_41)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_37),
.Y(n_46)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_38),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_39),
.B(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_51),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_38),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_18),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_35),
.A2(n_21),
.B1(n_26),
.B2(n_25),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_52),
.B1(n_31),
.B2(n_38),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_38),
.Y(n_59)
);

NAND3xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_13),
.C(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_35),
.A2(n_25),
.B1(n_24),
.B2(n_27),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_32),
.B(n_25),
.C(n_19),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_16),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_59),
.Y(n_81)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_49),
.Y(n_56)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_34),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_58),
.B(n_61),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_43),
.B(n_19),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_60),
.B(n_64),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_40),
.B(n_34),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

INVx6_ASAP7_75t_SL g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_18),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_65),
.B(n_10),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_66),
.A2(n_29),
.B1(n_37),
.B2(n_44),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_40),
.B(n_28),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_67),
.B(n_69),
.C(n_70),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_16),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_71),
.A2(n_74),
.B1(n_79),
.B2(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_63),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_80),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_58),
.A2(n_48),
.B1(n_50),
.B2(n_44),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_68),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_76),
.B(n_78),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_61),
.A2(n_50),
.B1(n_54),
.B2(n_49),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_69),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_70),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_90),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_85),
.B(n_86),
.Y(n_100)
);

NOR3xp33_ASAP7_75t_L g86 ( 
.A(n_75),
.B(n_67),
.C(n_59),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_89),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_81),
.A2(n_59),
.B(n_29),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_91),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_83),
.B(n_16),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_82),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_83),
.B(n_16),
.Y(n_94)
);

A2O1A1O1Ixp25_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_77),
.B(n_81),
.C(n_79),
.D(n_74),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_87),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g104 ( 
.A(n_96),
.B(n_88),
.C(n_22),
.Y(n_104)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_94),
.Y(n_97)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_97),
.Y(n_106)
);

A2O1A1O1Ixp25_ASAP7_75t_L g107 ( 
.A1(n_99),
.A2(n_71),
.B(n_22),
.C(n_3),
.D(n_5),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_100),
.A2(n_81),
.B(n_90),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_103),
.B(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_104),
.B(n_105),
.Y(n_111)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_101),
.A2(n_89),
.B(n_84),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_95),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_102),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_106),
.B(n_102),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_112),
.Y(n_115)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_113),
.B(n_8),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g114 ( 
.A1(n_110),
.A2(n_98),
.B(n_99),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_114),
.A2(n_116),
.B(n_115),
.Y(n_117)
);

AOI21xp33_ASAP7_75t_L g116 ( 
.A1(n_109),
.A2(n_108),
.B(n_98),
.Y(n_116)
);

OAI221xp5_ASAP7_75t_SL g120 ( 
.A1(n_117),
.A2(n_118),
.B1(n_119),
.B2(n_9),
.C(n_10),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_114),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_119)
);

OAI21x1_ASAP7_75t_L g121 ( 
.A1(n_120),
.A2(n_0),
.B(n_1),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_121),
.B(n_22),
.Y(n_122)
);


endmodule