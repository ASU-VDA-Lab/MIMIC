module real_jpeg_24591_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_131;
wire n_47;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_202;
wire n_128;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_89;
wire n_16;

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_0),
.A2(n_56),
.B1(n_106),
.B2(n_107),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_0),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_0),
.A2(n_58),
.B1(n_60),
.B2(n_106),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_0),
.A2(n_33),
.B1(n_37),
.B2(n_106),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_0),
.A2(n_22),
.B1(n_23),
.B2(n_106),
.Y(n_217)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_1),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_5),
.A2(n_33),
.B1(n_37),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_5),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_5),
.A2(n_40),
.B1(n_58),
.B2(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_5),
.A2(n_22),
.B1(n_23),
.B2(n_40),
.Y(n_119)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_6),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_33),
.B1(n_37),
.B2(n_43),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_7),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_7),
.A2(n_43),
.B1(n_58),
.B2(n_60),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_7),
.A2(n_22),
.B1(n_23),
.B2(n_43),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_43),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_8),
.A2(n_28),
.B1(n_51),
.B2(n_52),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_8),
.A2(n_28),
.B1(n_33),
.B2(n_37),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_8),
.A2(n_28),
.B1(n_58),
.B2(n_60),
.Y(n_100)
);

O2A1O1Ixp33_ASAP7_75t_L g164 ( 
.A1(n_8),
.A2(n_54),
.B(n_55),
.C(n_165),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_8),
.B(n_57),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g187 ( 
.A1(n_8),
.A2(n_60),
.B(n_77),
.C(n_188),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_8),
.B(n_22),
.C(n_36),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_8),
.B(n_75),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_8),
.B(n_223),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_8),
.B(n_38),
.Y(n_233)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_134),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_132),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_109),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_109),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_85),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_17),
.A2(n_18),
.B1(n_64),
.B2(n_65),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_44),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_20),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_20),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_20),
.A2(n_29),
.B1(n_45),
.B2(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_20),
.B(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_20),
.A2(n_45),
.B1(n_187),
.B2(n_245),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B(n_27),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_21),
.B(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_21),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_21),
.B(n_27),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_21),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_22),
.A2(n_23),
.B1(n_35),
.B2(n_36),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_22),
.B(n_229),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_25),
.B(n_93),
.Y(n_121)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_25),
.Y(n_223)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

OAI21xp33_ASAP7_75t_L g165 ( 
.A1(n_28),
.A2(n_53),
.B(n_60),
.Y(n_165)
);

OAI21xp33_ASAP7_75t_L g188 ( 
.A1(n_28),
.A2(n_37),
.B(n_79),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_29),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_39),
.B(n_41),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_30),
.A2(n_68),
.B(n_70),
.Y(n_146)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_31),
.B(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_31),
.B(n_69),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_31),
.B(n_192),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_38),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_32)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_33),
.A2(n_37),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_33),
.B(n_205),
.Y(n_204)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_38),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_38),
.B(n_192),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_39),
.A2(n_70),
.B(n_72),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_41),
.B(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_41),
.B(n_191),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_48),
.A2(n_61),
.B(n_62),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_49),
.B(n_129),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_49),
.B(n_63),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_57),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_50)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_51),
.Y(n_131)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx8_ASAP7_75t_L g108 ( 
.A(n_52),
.Y(n_108)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_53),
.A2(n_54),
.B1(n_58),
.B2(n_60),
.Y(n_57)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_57),
.B(n_63),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_57),
.B(n_105),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_57),
.B(n_129),
.Y(n_160)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_58),
.A2(n_60),
.B1(n_77),
.B2(n_79),
.Y(n_82)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_65),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_73),
.B(n_84),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_71),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_67),
.B(n_190),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_72),
.B(n_202),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_80),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_75),
.B(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_76),
.B(n_83),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_76),
.A2(n_81),
.B(n_125),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_76),
.B(n_125),
.Y(n_158)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_80),
.B(n_148),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_81),
.B(n_157),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_95),
.C(n_101),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_94),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_87),
.B(n_94),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_92),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_88),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_91),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_92),
.B(n_119),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_92),
.B(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_95),
.A2(n_101),
.B1(n_102),
.B2(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_96),
.B(n_156),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_98),
.B(n_149),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_99),
.B(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_104),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_104),
.B(n_160),
.Y(n_159)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_113),
.C(n_115),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_110),
.B(n_113),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_115),
.B(n_271),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_124),
.C(n_126),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_116),
.A2(n_117),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_121),
.B(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_121),
.B(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_123),
.B(n_202),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_124),
.A2(n_126),
.B1(n_262),
.B2(n_263),
.Y(n_261)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_124),
.Y(n_262)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_126),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_127),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_268),
.B(n_272),
.Y(n_134)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_180),
.B(n_254),
.C(n_267),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_168),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_137),
.B(n_168),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_153),
.B2(n_167),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_151),
.B2(n_152),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_140),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_140),
.B(n_152),
.C(n_167),
.Y(n_255)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_147),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_142),
.A2(n_143),
.B1(n_171),
.B2(n_172),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_145),
.A2(n_146),
.B1(n_147),
.B2(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_147),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g157 ( 
.A(n_150),
.Y(n_157)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_163),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_159),
.B1(n_161),
.B2(n_162),
.Y(n_154)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_155),
.B(n_162),
.C(n_163),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_158),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_159),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_174),
.C(n_175),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_170),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_175),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_177),
.C(n_178),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_185),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_178),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_179),
.B(n_231),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_253),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_196),
.B(n_252),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_183),
.B(n_193),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.C(n_189),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_184),
.B(n_250),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_186),
.B(n_189),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

INVxp33_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_247),
.B(n_251),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_198),
.A2(n_238),
.B(n_246),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_219),
.B(n_237),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_206),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_200),
.B(n_206),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_201),
.A2(n_203),
.B1(n_204),
.B2(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_201),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_208),
.B1(n_213),
.B2(n_218),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_210),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_212),
.C(n_218),
.Y(n_239)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_210),
.Y(n_212)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_217),
.B(n_223),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_220),
.A2(n_226),
.B(n_236),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_224),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_221),
.B(n_224),
.Y(n_236)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_222),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_232),
.B(n_235),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_233),
.B(n_234),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_239),
.B(n_240),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_244),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_243),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_243),
.C(n_244),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_248),
.B(n_249),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_256),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_266),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_259),
.B1(n_264),
.B2(n_265),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_265),
.C(n_266),
.Y(n_269)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_269),
.B(n_270),
.Y(n_272)
);


endmodule