module fake_ibex_1451_n_842 (n_151, n_147, n_85, n_128, n_84, n_64, n_3, n_73, n_152, n_145, n_65, n_103, n_95, n_139, n_55, n_130, n_63, n_98, n_129, n_29, n_143, n_106, n_148, n_2, n_76, n_8, n_118, n_67, n_9, n_38, n_124, n_37, n_110, n_47, n_108, n_10, n_82, n_21, n_27, n_16, n_78, n_60, n_86, n_70, n_7, n_20, n_87, n_69, n_75, n_109, n_121, n_127, n_137, n_48, n_57, n_59, n_28, n_125, n_39, n_5, n_62, n_71, n_153, n_120, n_93, n_155, n_13, n_122, n_116, n_61, n_14, n_0, n_94, n_134, n_12, n_42, n_77, n_112, n_150, n_88, n_133, n_44, n_142, n_51, n_46, n_80, n_49, n_40, n_66, n_17, n_74, n_90, n_58, n_43, n_140, n_22, n_136, n_4, n_119, n_33, n_30, n_6, n_100, n_72, n_26, n_114, n_34, n_97, n_102, n_15, n_131, n_123, n_24, n_52, n_99, n_135, n_105, n_156, n_126, n_1, n_154, n_111, n_25, n_36, n_104, n_41, n_45, n_141, n_18, n_89, n_83, n_32, n_53, n_107, n_115, n_149, n_50, n_11, n_92, n_144, n_101, n_113, n_138, n_96, n_68, n_117, n_79, n_81, n_35, n_132, n_157, n_31, n_56, n_23, n_146, n_91, n_54, n_19, n_842);

input n_151;
input n_147;
input n_85;
input n_128;
input n_84;
input n_64;
input n_3;
input n_73;
input n_152;
input n_145;
input n_65;
input n_103;
input n_95;
input n_139;
input n_55;
input n_130;
input n_63;
input n_98;
input n_129;
input n_29;
input n_143;
input n_106;
input n_148;
input n_2;
input n_76;
input n_8;
input n_118;
input n_67;
input n_9;
input n_38;
input n_124;
input n_37;
input n_110;
input n_47;
input n_108;
input n_10;
input n_82;
input n_21;
input n_27;
input n_16;
input n_78;
input n_60;
input n_86;
input n_70;
input n_7;
input n_20;
input n_87;
input n_69;
input n_75;
input n_109;
input n_121;
input n_127;
input n_137;
input n_48;
input n_57;
input n_59;
input n_28;
input n_125;
input n_39;
input n_5;
input n_62;
input n_71;
input n_153;
input n_120;
input n_93;
input n_155;
input n_13;
input n_122;
input n_116;
input n_61;
input n_14;
input n_0;
input n_94;
input n_134;
input n_12;
input n_42;
input n_77;
input n_112;
input n_150;
input n_88;
input n_133;
input n_44;
input n_142;
input n_51;
input n_46;
input n_80;
input n_49;
input n_40;
input n_66;
input n_17;
input n_74;
input n_90;
input n_58;
input n_43;
input n_140;
input n_22;
input n_136;
input n_4;
input n_119;
input n_33;
input n_30;
input n_6;
input n_100;
input n_72;
input n_26;
input n_114;
input n_34;
input n_97;
input n_102;
input n_15;
input n_131;
input n_123;
input n_24;
input n_52;
input n_99;
input n_135;
input n_105;
input n_156;
input n_126;
input n_1;
input n_154;
input n_111;
input n_25;
input n_36;
input n_104;
input n_41;
input n_45;
input n_141;
input n_18;
input n_89;
input n_83;
input n_32;
input n_53;
input n_107;
input n_115;
input n_149;
input n_50;
input n_11;
input n_92;
input n_144;
input n_101;
input n_113;
input n_138;
input n_96;
input n_68;
input n_117;
input n_79;
input n_81;
input n_35;
input n_132;
input n_157;
input n_31;
input n_56;
input n_23;
input n_146;
input n_91;
input n_54;
input n_19;

output n_842;

wire n_599;
wire n_778;
wire n_822;
wire n_507;
wire n_743;
wire n_540;
wire n_754;
wire n_395;
wire n_171;
wire n_756;
wire n_529;
wire n_389;
wire n_204;
wire n_626;
wire n_274;
wire n_387;
wire n_766;
wire n_688;
wire n_177;
wire n_707;
wire n_273;
wire n_330;
wire n_309;
wire n_328;
wire n_293;
wire n_372;
wire n_341;
wire n_256;
wire n_418;
wire n_193;
wire n_510;
wire n_446;
wire n_350;
wire n_601;
wire n_621;
wire n_610;
wire n_165;
wire n_790;
wire n_452;
wire n_664;
wire n_255;
wire n_175;
wire n_586;
wire n_773;
wire n_638;
wire n_398;
wire n_304;
wire n_821;
wire n_191;
wire n_593;
wire n_545;
wire n_583;
wire n_678;
wire n_663;
wire n_194;
wire n_249;
wire n_334;
wire n_634;
wire n_733;
wire n_312;
wire n_622;
wire n_578;
wire n_478;
wire n_239;
wire n_432;
wire n_371;
wire n_403;
wire n_423;
wire n_608;
wire n_357;
wire n_412;
wire n_457;
wire n_494;
wire n_226;
wire n_336;
wire n_258;
wire n_449;
wire n_547;
wire n_176;
wire n_727;
wire n_216;
wire n_652;
wire n_781;
wire n_421;
wire n_828;
wire n_738;
wire n_475;
wire n_802;
wire n_166;
wire n_163;
wire n_753;
wire n_645;
wire n_500;
wire n_747;
wire n_542;
wire n_236;
wire n_376;
wire n_377;
wire n_584;
wire n_531;
wire n_647;
wire n_761;
wire n_556;
wire n_748;
wire n_189;
wire n_498;
wire n_708;
wire n_280;
wire n_317;
wire n_375;
wire n_340;
wire n_698;
wire n_187;
wire n_667;
wire n_682;
wire n_182;
wire n_196;
wire n_326;
wire n_327;
wire n_723;
wire n_170;
wire n_270;
wire n_346;
wire n_383;
wire n_840;
wire n_561;
wire n_417;
wire n_471;
wire n_739;
wire n_755;
wire n_265;
wire n_504;
wire n_158;
wire n_259;
wire n_276;
wire n_339;
wire n_470;
wire n_770;
wire n_210;
wire n_348;
wire n_220;
wire n_674;
wire n_481;
wire n_287;
wire n_243;
wire n_497;
wire n_711;
wire n_228;
wire n_671;
wire n_552;
wire n_384;
wire n_251;
wire n_632;
wire n_373;
wire n_458;
wire n_244;
wire n_343;
wire n_310;
wire n_714;
wire n_703;
wire n_426;
wire n_323;
wire n_469;
wire n_829;
wire n_598;
wire n_825;
wire n_740;
wire n_386;
wire n_549;
wire n_224;
wire n_183;
wire n_533;
wire n_508;
wire n_453;
wire n_591;
wire n_655;
wire n_333;
wire n_306;
wire n_400;
wire n_550;
wire n_736;
wire n_169;
wire n_732;
wire n_798;
wire n_673;
wire n_832;
wire n_242;
wire n_278;
wire n_316;
wire n_404;
wire n_557;
wire n_641;
wire n_527;
wire n_590;
wire n_465;
wire n_325;
wire n_301;
wire n_496;
wire n_617;
wire n_434;
wire n_296;
wire n_690;
wire n_835;
wire n_168;
wire n_526;
wire n_785;
wire n_824;
wire n_315;
wire n_441;
wire n_604;
wire n_637;
wire n_523;
wire n_787;
wire n_694;
wire n_614;
wire n_370;
wire n_431;
wire n_719;
wire n_574;
wire n_289;
wire n_716;
wire n_515;
wire n_642;
wire n_286;
wire n_321;
wire n_569;
wire n_600;
wire n_215;
wire n_279;
wire n_374;
wire n_235;
wire n_464;
wire n_538;
wire n_669;
wire n_838;
wire n_750;
wire n_746;
wire n_261;
wire n_742;
wire n_521;
wire n_665;
wire n_459;
wire n_518;
wire n_367;
wire n_221;
wire n_789;
wire n_654;
wire n_656;
wire n_724;
wire n_437;
wire n_731;
wire n_602;
wire n_355;
wire n_767;
wire n_474;
wire n_758;
wire n_594;
wire n_636;
wire n_720;
wire n_710;
wire n_407;
wire n_490;
wire n_568;
wire n_813;
wire n_448;
wire n_646;
wire n_595;
wire n_466;
wire n_269;
wire n_570;
wire n_623;
wire n_585;
wire n_715;
wire n_791;
wire n_530;
wire n_356;
wire n_420;
wire n_483;
wire n_543;
wire n_580;
wire n_487;
wire n_769;
wire n_222;
wire n_660;
wire n_186;
wire n_524;
wire n_349;
wire n_765;
wire n_454;
wire n_777;
wire n_295;
wire n_730;
wire n_331;
wire n_576;
wire n_230;
wire n_759;
wire n_185;
wire n_388;
wire n_625;
wire n_619;
wire n_536;
wire n_611;
wire n_352;
wire n_290;
wire n_558;
wire n_666;
wire n_174;
wire n_467;
wire n_427;
wire n_607;
wire n_827;
wire n_219;
wire n_246;
wire n_442;
wire n_207;
wire n_438;
wire n_689;
wire n_793;
wire n_167;
wire n_676;
wire n_253;
wire n_208;
wire n_234;
wire n_300;
wire n_358;
wire n_771;
wire n_205;
wire n_618;
wire n_488;
wire n_514;
wire n_705;
wire n_429;
wire n_560;
wire n_275;
wire n_541;
wire n_613;
wire n_659;
wire n_267;
wire n_662;
wire n_635;
wire n_245;
wire n_589;
wire n_571;
wire n_229;
wire n_209;
wire n_472;
wire n_648;
wire n_783;
wire n_347;
wire n_830;
wire n_473;
wire n_445;
wire n_629;
wire n_335;
wire n_413;
wire n_263;
wire n_573;
wire n_353;
wire n_359;
wire n_826;
wire n_299;
wire n_262;
wire n_439;
wire n_433;
wire n_704;
wire n_643;
wire n_679;
wire n_841;
wire n_772;
wire n_810;
wire n_768;
wire n_839;
wire n_338;
wire n_173;
wire n_696;
wire n_796;
wire n_797;
wire n_837;
wire n_477;
wire n_640;
wire n_363;
wire n_402;
wire n_725;
wire n_180;
wire n_369;
wire n_596;
wire n_201;
wire n_699;
wire n_351;
wire n_368;
wire n_456;
wire n_834;
wire n_257;
wire n_718;
wire n_801;
wire n_672;
wire n_722;
wire n_401;
wire n_553;
wire n_554;
wire n_735;
wire n_305;
wire n_713;
wire n_307;
wire n_192;
wire n_804;
wire n_484;
wire n_566;
wire n_480;
wire n_416;
wire n_581;
wire n_721;
wire n_365;
wire n_651;
wire n_814;
wire n_605;
wire n_539;
wire n_179;
wire n_354;
wire n_206;
wire n_392;
wire n_630;
wire n_516;
wire n_548;
wire n_567;
wire n_763;
wire n_745;
wire n_329;
wire n_447;
wire n_188;
wire n_200;
wire n_444;
wire n_506;
wire n_562;
wire n_564;
wire n_546;
wire n_199;
wire n_788;
wire n_795;
wire n_592;
wire n_495;
wire n_762;
wire n_410;
wire n_308;
wire n_800;
wire n_675;
wire n_463;
wire n_624;
wire n_706;
wire n_411;
wire n_520;
wire n_784;
wire n_684;
wire n_775;
wire n_658;
wire n_512;
wire n_615;
wire n_685;
wire n_283;
wire n_366;
wire n_397;
wire n_803;
wire n_692;
wire n_627;
wire n_709;
wire n_322;
wire n_227;
wire n_499;
wire n_757;
wire n_248;
wire n_702;
wire n_451;
wire n_712;
wire n_190;
wire n_650;
wire n_776;
wire n_409;
wire n_582;
wire n_818;
wire n_653;
wire n_238;
wire n_214;
wire n_579;
wire n_332;
wire n_799;
wire n_517;
wire n_211;
wire n_744;
wire n_817;
wire n_218;
wire n_314;
wire n_691;
wire n_563;
wire n_277;
wire n_555;
wire n_337;
wire n_522;
wire n_700;
wire n_479;
wire n_534;
wire n_225;
wire n_360;
wire n_272;
wire n_511;
wire n_734;
wire n_468;
wire n_223;
wire n_381;
wire n_525;
wire n_815;
wire n_780;
wire n_535;
wire n_382;
wire n_502;
wire n_681;
wire n_633;
wire n_532;
wire n_726;
wire n_405;
wire n_415;
wire n_597;
wire n_285;
wire n_288;
wire n_247;
wire n_320;
wire n_379;
wire n_551;
wire n_612;
wire n_318;
wire n_291;
wire n_819;
wire n_161;
wire n_237;
wire n_203;
wire n_268;
wire n_440;
wire n_342;
wire n_233;
wire n_385;
wire n_414;
wire n_430;
wire n_729;
wire n_741;
wire n_603;
wire n_378;
wire n_486;
wire n_422;
wire n_164;
wire n_264;
wire n_198;
wire n_616;
wire n_782;
wire n_833;
wire n_217;
wire n_324;
wire n_391;
wire n_831;
wire n_537;
wire n_728;
wire n_805;
wire n_670;
wire n_820;
wire n_390;
wire n_544;
wire n_178;
wire n_509;
wire n_695;
wire n_786;
wire n_639;
wire n_303;
wire n_362;
wire n_717;
wire n_505;
wire n_162;
wire n_482;
wire n_240;
wire n_282;
wire n_680;
wire n_501;
wire n_809;
wire n_752;
wire n_668;
wire n_779;
wire n_266;
wire n_294;
wire n_485;
wire n_284;
wire n_811;
wire n_808;
wire n_172;
wire n_250;
wire n_493;
wire n_460;
wire n_609;
wire n_476;
wire n_792;
wire n_461;
wire n_575;
wire n_313;
wire n_519;
wire n_345;
wire n_408;
wire n_361;
wire n_455;
wire n_419;
wire n_774;
wire n_319;
wire n_195;
wire n_513;
wire n_212;
wire n_588;
wire n_693;
wire n_311;
wire n_661;
wire n_406;
wire n_606;
wire n_737;
wire n_197;
wire n_528;
wire n_181;
wire n_683;
wire n_631;
wire n_260;
wire n_620;
wire n_794;
wire n_836;
wire n_462;
wire n_302;
wire n_450;
wire n_443;
wire n_686;
wire n_572;
wire n_644;
wire n_577;
wire n_344;
wire n_393;
wire n_436;
wire n_428;
wire n_491;
wire n_297;
wire n_435;
wire n_628;
wire n_252;
wire n_396;
wire n_816;
wire n_697;
wire n_489;
wire n_677;
wire n_399;
wire n_254;
wire n_213;
wire n_424;
wire n_565;
wire n_823;
wire n_701;
wire n_271;
wire n_241;
wire n_503;
wire n_292;
wire n_807;
wire n_394;
wire n_364;
wire n_687;
wire n_159;
wire n_298;
wire n_202;
wire n_231;
wire n_587;
wire n_760;
wire n_751;
wire n_806;
wire n_160;
wire n_657;
wire n_764;
wire n_184;
wire n_492;
wire n_649;
wire n_812;
wire n_232;
wire n_380;
wire n_749;
wire n_281;
wire n_559;
wire n_425;

INVx1_ASAP7_75t_L g158 ( 
.A(n_36),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_84),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_73),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_76),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_28),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_80),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_38),
.Y(n_169)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_83),
.Y(n_170)
);

CKINVDCx14_ASAP7_75t_R g171 ( 
.A(n_60),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_53),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_93),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_95),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_61),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_6),
.Y(n_176)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_50),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_101),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_68),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_48),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_132),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_90),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_59),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_111),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_107),
.Y(n_188)
);

NOR2xp67_ASAP7_75t_L g189 ( 
.A(n_104),
.B(n_20),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_140),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_49),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_131),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_2),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_86),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_114),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_142),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_98),
.Y(n_198)
);

BUFx10_ASAP7_75t_L g199 ( 
.A(n_139),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_64),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_12),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_129),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_133),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_70),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_134),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_141),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_20),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_100),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_43),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_28),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

NOR2xp67_ASAP7_75t_L g213 ( 
.A(n_37),
.B(n_35),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_117),
.Y(n_214)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_33),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_46),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_67),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_92),
.Y(n_219)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_77),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_123),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_62),
.Y(n_222)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_157),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_54),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_116),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_148),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_42),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_27),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_10),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_125),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_85),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_88),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_15),
.Y(n_233)
);

INVxp33_ASAP7_75t_SL g234 ( 
.A(n_57),
.Y(n_234)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_108),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_110),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_130),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_3),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_120),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_122),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_26),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_2),
.Y(n_242)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_32),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_66),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_82),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_5),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_15),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_74),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_14),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_41),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_78),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_127),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_128),
.Y(n_253)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_65),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_10),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_47),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_79),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_12),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_33),
.Y(n_259)
);

INVx4_ASAP7_75t_R g260 ( 
.A(n_5),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_87),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_11),
.Y(n_262)
);

OAI22x1_ASAP7_75t_R g263 ( 
.A1(n_233),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_170),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_170),
.Y(n_265)
);

AND2x6_ASAP7_75t_L g266 ( 
.A(n_223),
.B(n_34),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_201),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_1),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g269 ( 
.A(n_186),
.Y(n_269)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_207),
.B(n_4),
.Y(n_271)
);

OAI22x1_ASAP7_75t_L g272 ( 
.A1(n_194),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_174),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_207),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_174),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_235),
.Y(n_276)
);

INVx5_ASAP7_75t_L g277 ( 
.A(n_174),
.Y(n_277)
);

AND2x4_ASAP7_75t_L g278 ( 
.A(n_201),
.B(n_7),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_246),
.B(n_8),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_187),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_173),
.Y(n_281)
);

BUFx8_ASAP7_75t_L g282 ( 
.A(n_220),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_176),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_175),
.Y(n_285)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_175),
.A2(n_91),
.B(n_156),
.Y(n_286)
);

BUFx12f_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_194),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_187),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_216),
.Y(n_290)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_200),
.A2(n_89),
.B(n_155),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_246),
.A2(n_9),
.B1(n_11),
.B2(n_13),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_241),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_171),
.B(n_9),
.Y(n_294)
);

OAI22x1_ASAP7_75t_L g295 ( 
.A1(n_242),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_295)
);

OA21x2_ASAP7_75t_L g296 ( 
.A1(n_203),
.A2(n_96),
.B(n_153),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_208),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_203),
.B(n_16),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_230),
.B(n_17),
.Y(n_299)
);

AOI22x1_ASAP7_75t_SL g300 ( 
.A1(n_243),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_230),
.Y(n_301)
);

AND2x4_ASAP7_75t_L g302 ( 
.A(n_239),
.B(n_252),
.Y(n_302)
);

OA21x2_ASAP7_75t_L g303 ( 
.A1(n_239),
.A2(n_97),
.B(n_152),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_247),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_187),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_228),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g307 ( 
.A(n_171),
.B(n_18),
.Y(n_307)
);

NOR2x1_ASAP7_75t_L g308 ( 
.A(n_258),
.B(n_39),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_188),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_177),
.B(n_19),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g311 ( 
.A(n_196),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g312 ( 
.A(n_259),
.B(n_21),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_196),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_229),
.Y(n_314)
);

OA21x2_ASAP7_75t_L g315 ( 
.A1(n_158),
.A2(n_99),
.B(n_151),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_183),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_227),
.B(n_22),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_159),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_160),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_162),
.Y(n_320)
);

BUFx8_ASAP7_75t_L g321 ( 
.A(n_163),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_188),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_164),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_215),
.Y(n_324)
);

OA21x2_ASAP7_75t_L g325 ( 
.A1(n_166),
.A2(n_94),
.B(n_150),
.Y(n_325)
);

HB1xp67_ASAP7_75t_L g326 ( 
.A(n_238),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_169),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_215),
.Y(n_328)
);

INVxp33_ASAP7_75t_L g329 ( 
.A(n_297),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g330 ( 
.A(n_266),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_274),
.B(n_245),
.Y(n_331)
);

HB1xp67_ASAP7_75t_SL g332 ( 
.A(n_282),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_305),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_305),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_267),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_305),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_L g338 ( 
.A1(n_298),
.A2(n_234),
.B1(n_237),
.B2(n_212),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g339 ( 
.A(n_306),
.Y(n_339)
);

NOR2x1p5_ASAP7_75t_L g340 ( 
.A(n_269),
.B(n_249),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

INVx3_ASAP7_75t_L g342 ( 
.A(n_299),
.Y(n_342)
);

OAI22x1_ASAP7_75t_SL g343 ( 
.A1(n_263),
.A2(n_262),
.B1(n_255),
.B2(n_257),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_299),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_299),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_278),
.Y(n_347)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_276),
.B(n_199),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_278),
.Y(n_349)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_273),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_270),
.B(n_165),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_273),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_209),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_312),
.Y(n_354)
);

INVx8_ASAP7_75t_L g355 ( 
.A(n_287),
.Y(n_355)
);

NAND2xp33_ASAP7_75t_L g356 ( 
.A(n_266),
.B(n_168),
.Y(n_356)
);

BUFx6f_ASAP7_75t_SL g357 ( 
.A(n_312),
.Y(n_357)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_314),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_275),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_267),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_268),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_326),
.B(n_211),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_268),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g366 ( 
.A(n_279),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_282),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_302),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_283),
.B(n_261),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_275),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_316),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_264),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_265),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_284),
.B(n_178),
.Y(n_374)
);

NAND3xp33_ASAP7_75t_L g375 ( 
.A(n_271),
.B(n_181),
.C(n_180),
.Y(n_375)
);

BUFx2_ASAP7_75t_L g376 ( 
.A(n_282),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_281),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_287),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_L g379 ( 
.A(n_294),
.B(n_172),
.Y(n_379)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_311),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_318),
.B(n_184),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_281),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_318),
.B(n_185),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_293),
.B(n_179),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_319),
.B(n_182),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_285),
.Y(n_386)
);

HB1xp67_ASAP7_75t_L g387 ( 
.A(n_279),
.Y(n_387)
);

OR2x6_ASAP7_75t_L g388 ( 
.A(n_311),
.B(n_292),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_301),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_301),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_280),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_290),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_307),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_304),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_321),
.Y(n_395)
);

INVxp33_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

OAI22xp33_ASAP7_75t_L g397 ( 
.A1(n_295),
.A2(n_161),
.B1(n_205),
.B2(n_210),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_288),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_310),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_319),
.B(n_191),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_277),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_317),
.B(n_192),
.Y(n_402)
);

NAND2xp33_ASAP7_75t_L g403 ( 
.A(n_320),
.B(n_195),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_277),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_317),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_323),
.Y(n_407)
);

NAND2xp33_ASAP7_75t_L g408 ( 
.A(n_327),
.B(n_204),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_327),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_321),
.A2(n_224),
.B1(n_214),
.B2(n_236),
.Y(n_410)
);

OAI22xp33_ASAP7_75t_L g411 ( 
.A1(n_295),
.A2(n_189),
.B1(n_190),
.B2(n_256),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_289),
.Y(n_412)
);

BUFx10_ASAP7_75t_L g413 ( 
.A(n_289),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_277),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_289),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

BUFx6f_ASAP7_75t_SL g417 ( 
.A(n_378),
.Y(n_417)
);

INVx2_ASAP7_75t_SL g418 ( 
.A(n_355),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_366),
.B(n_308),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_366),
.B(n_286),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g421 ( 
.A(n_330),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_354),
.B(n_286),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_339),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_362),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_331),
.B(n_202),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_329),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_368),
.Y(n_427)
);

BUFx6f_ASAP7_75t_SL g428 ( 
.A(n_380),
.Y(n_428)
);

NAND2x1p5_ASAP7_75t_L g429 ( 
.A(n_376),
.B(n_291),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_342),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_342),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_345),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_336),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_L g434 ( 
.A1(n_363),
.A2(n_272),
.B1(n_296),
.B2(n_303),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_369),
.B(n_222),
.Y(n_435)
);

INVxp33_ASAP7_75t_L g436 ( 
.A(n_329),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_365),
.A2(n_272),
.B1(n_296),
.B2(n_303),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_399),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_367),
.B(n_226),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_399),
.B(n_303),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_369),
.B(n_231),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_346),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_348),
.B(n_240),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_395),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_347),
.A2(n_193),
.B1(n_244),
.B2(n_197),
.Y(n_446)
);

NOR2xp67_ASAP7_75t_L g447 ( 
.A(n_380),
.B(n_22),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_384),
.B(n_248),
.Y(n_448)
);

INVxp67_ASAP7_75t_L g449 ( 
.A(n_332),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_358),
.B(n_198),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_406),
.Y(n_451)
);

INVx2_ASAP7_75t_SL g452 ( 
.A(n_355),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_338),
.B(n_206),
.Y(n_453)
);

OAI22xp33_ASAP7_75t_L g454 ( 
.A1(n_396),
.A2(n_300),
.B1(n_232),
.B2(n_217),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_407),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_392),
.B(n_218),
.Y(n_456)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_387),
.B(n_219),
.Y(n_457)
);

INVxp67_ASAP7_75t_SL g458 ( 
.A(n_387),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_338),
.B(n_221),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g460 ( 
.A(n_393),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_394),
.B(n_374),
.Y(n_462)
);

NOR2xp67_ASAP7_75t_L g463 ( 
.A(n_375),
.B(n_23),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_374),
.B(n_250),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_396),
.B(n_251),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_402),
.B(n_253),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_349),
.B(n_213),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_360),
.A2(n_325),
.B1(n_315),
.B2(n_225),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_371),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_389),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_385),
.B(n_400),
.Y(n_472)
);

OAI22xp33_ASAP7_75t_L g473 ( 
.A1(n_405),
.A2(n_260),
.B1(n_325),
.B2(n_225),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_372),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_353),
.B(n_215),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_373),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_377),
.Y(n_479)
);

NOR2xp67_ASAP7_75t_L g480 ( 
.A(n_410),
.B(n_23),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

OR2x2_ASAP7_75t_L g482 ( 
.A(n_405),
.B(n_24),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_351),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_382),
.A2(n_328),
.B(n_324),
.C(n_322),
.Y(n_484)
);

BUFx2_ASAP7_75t_L g485 ( 
.A(n_388),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_357),
.B(n_40),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

O2A1O1Ixp33_ASAP7_75t_L g488 ( 
.A1(n_411),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_488)
);

INVx8_ASAP7_75t_L g489 ( 
.A(n_388),
.Y(n_489)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_390),
.Y(n_490)
);

AOI22x1_ASAP7_75t_L g491 ( 
.A1(n_401),
.A2(n_328),
.B1(n_324),
.B2(n_322),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_438),
.B(n_379),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_422),
.A2(n_356),
.B(n_403),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_422),
.A2(n_408),
.B(n_383),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_423),
.A2(n_388),
.B1(n_397),
.B2(n_383),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_490),
.B(n_381),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_426),
.B(n_397),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_464),
.A2(n_381),
.B1(n_340),
.B2(n_414),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_462),
.B(n_25),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_27),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_430),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_431),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g503 ( 
.A1(n_450),
.A2(n_343),
.B1(n_413),
.B2(n_309),
.Y(n_503)
);

AOI21xp5_ASAP7_75t_L g504 ( 
.A1(n_420),
.A2(n_415),
.B(n_412),
.Y(n_504)
);

NOR2x1_ASAP7_75t_R g505 ( 
.A(n_445),
.B(n_29),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_458),
.B(n_29),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_432),
.Y(n_507)
);

BUFx2_ASAP7_75t_L g508 ( 
.A(n_418),
.Y(n_508)
);

BUFx8_ASAP7_75t_SL g509 ( 
.A(n_428),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_472),
.B(n_30),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_419),
.B(n_466),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_452),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_457),
.B(n_31),
.Y(n_514)
);

AOI33xp33_ASAP7_75t_L g515 ( 
.A1(n_454),
.A2(n_333),
.A3(n_334),
.B1(n_335),
.B2(n_337),
.B3(n_370),
.Y(n_515)
);

AND2x4_ASAP7_75t_L g516 ( 
.A(n_460),
.B(n_31),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_478),
.Y(n_517)
);

INVxp33_ASAP7_75t_SL g518 ( 
.A(n_439),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_419),
.B(n_32),
.Y(n_519)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_440),
.A2(n_391),
.B(n_341),
.Y(n_520)
);

A2O1A1Ixp33_ASAP7_75t_L g521 ( 
.A1(n_442),
.A2(n_309),
.B(n_322),
.C(n_324),
.Y(n_521)
);

NAND2x1p5_ASAP7_75t_L g522 ( 
.A(n_485),
.B(n_324),
.Y(n_522)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_469),
.A2(n_429),
.B(n_434),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_482),
.A2(n_328),
.B1(n_337),
.B2(n_370),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_443),
.B(n_425),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_427),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_474),
.Y(n_527)
);

BUFx4f_ASAP7_75t_L g528 ( 
.A(n_489),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_453),
.B(n_44),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_424),
.Y(n_530)
);

O2A1O1Ixp33_ASAP7_75t_L g531 ( 
.A1(n_459),
.A2(n_352),
.B(n_350),
.C(n_344),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_477),
.Y(n_532)
);

NOR2x1_ASAP7_75t_L g533 ( 
.A(n_447),
.B(n_352),
.Y(n_533)
);

O2A1O1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_467),
.A2(n_45),
.B(n_51),
.C(n_52),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_446),
.B(n_55),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_465),
.B(n_451),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_455),
.B(n_56),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_R g538 ( 
.A(n_417),
.B(n_58),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_461),
.B(n_63),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_L g540 ( 
.A1(n_475),
.A2(n_359),
.B(n_69),
.Y(n_540)
);

INVx4_ASAP7_75t_L g541 ( 
.A(n_428),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_478),
.Y(n_542)
);

BUFx2_ASAP7_75t_L g543 ( 
.A(n_449),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_470),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_487),
.A2(n_71),
.B1(n_72),
.B2(n_75),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_478),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_479),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_444),
.B(n_102),
.Y(n_548)
);

A2O1A1Ixp33_ASAP7_75t_L g549 ( 
.A1(n_476),
.A2(n_103),
.B(n_105),
.C(n_106),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g550 ( 
.A1(n_456),
.A2(n_441),
.B1(n_435),
.B2(n_489),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_417),
.B(n_126),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_489),
.A2(n_448),
.B1(n_480),
.B2(n_471),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_433),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g554 ( 
.A1(n_463),
.A2(n_135),
.B1(n_136),
.B2(n_138),
.Y(n_554)
);

AND2x4_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_144),
.Y(n_555)
);

AND2x4_ASAP7_75t_L g556 ( 
.A(n_416),
.B(n_149),
.Y(n_556)
);

O2A1O1Ixp33_ASAP7_75t_L g557 ( 
.A1(n_488),
.A2(n_145),
.B(n_146),
.C(n_147),
.Y(n_557)
);

AOI221x1_ASAP7_75t_L g558 ( 
.A1(n_540),
.A2(n_484),
.B1(n_486),
.B2(n_481),
.C(n_491),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_526),
.B(n_421),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_536),
.B(n_514),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_510),
.A2(n_499),
.B1(n_550),
.B2(n_519),
.Y(n_561)
);

INVx3_ASAP7_75t_L g562 ( 
.A(n_542),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_544),
.B(n_547),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_532),
.Y(n_564)
);

AND2x4_ASAP7_75t_L g565 ( 
.A(n_541),
.B(n_530),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_528),
.B(n_542),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_494),
.A2(n_520),
.B(n_504),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g568 ( 
.A(n_513),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_516),
.B(n_527),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_516),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_492),
.B(n_497),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_528),
.B(n_508),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_501),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_502),
.Y(n_574)
);

AO32x2_ASAP7_75t_L g575 ( 
.A1(n_552),
.A2(n_495),
.A3(n_524),
.B1(n_498),
.B2(n_545),
.Y(n_575)
);

O2A1O1Ixp33_ASAP7_75t_L g576 ( 
.A1(n_506),
.A2(n_500),
.B(n_557),
.C(n_496),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_507),
.Y(n_577)
);

OR2x2_ASAP7_75t_L g578 ( 
.A(n_512),
.B(n_541),
.Y(n_578)
);

NOR2x1_ASAP7_75t_R g579 ( 
.A(n_509),
.B(n_543),
.Y(n_579)
);

BUFx3_ASAP7_75t_L g580 ( 
.A(n_518),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_556),
.A2(n_535),
.B1(n_537),
.B2(n_539),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_553),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_542),
.B(n_538),
.Y(n_583)
);

INVx2_ASAP7_75t_SL g584 ( 
.A(n_548),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_555),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_L g586 ( 
.A1(n_556),
.A2(n_554),
.B1(n_529),
.B2(n_522),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_517),
.B(n_546),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_505),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_533),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_551),
.Y(n_590)
);

OAI21xp5_ASAP7_75t_L g591 ( 
.A1(n_549),
.A2(n_531),
.B(n_521),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_546),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_536),
.A2(n_420),
.B1(n_366),
.B2(n_511),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_509),
.Y(n_594)
);

OAI21xp5_ASAP7_75t_L g595 ( 
.A1(n_523),
.A2(n_520),
.B(n_493),
.Y(n_595)
);

AOI21xp33_ASAP7_75t_L g596 ( 
.A1(n_557),
.A2(n_550),
.B(n_525),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_511),
.B(n_399),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_511),
.B(n_399),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_511),
.B(n_399),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_544),
.Y(n_600)
);

CKINVDCx6p67_ASAP7_75t_R g601 ( 
.A(n_541),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_497),
.B(n_423),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_542),
.Y(n_603)
);

AND2x4_ASAP7_75t_L g604 ( 
.A(n_526),
.B(n_445),
.Y(n_604)
);

AO21x1_ASAP7_75t_L g605 ( 
.A1(n_523),
.A2(n_473),
.B(n_534),
.Y(n_605)
);

AOI21xp5_ASAP7_75t_L g606 ( 
.A1(n_523),
.A2(n_422),
.B(n_420),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_523),
.A2(n_520),
.B(n_493),
.Y(n_607)
);

BUFx4f_ASAP7_75t_SL g608 ( 
.A(n_541),
.Y(n_608)
);

AND2x2_ASAP7_75t_L g609 ( 
.A(n_497),
.B(n_423),
.Y(n_609)
);

AOI21xp5_ASAP7_75t_L g610 ( 
.A1(n_523),
.A2(n_422),
.B(n_420),
.Y(n_610)
);

HB1xp67_ASAP7_75t_L g611 ( 
.A(n_513),
.Y(n_611)
);

HB1xp67_ASAP7_75t_L g612 ( 
.A(n_513),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_497),
.B(n_423),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_511),
.B(n_399),
.Y(n_614)
);

HB1xp67_ASAP7_75t_L g615 ( 
.A(n_513),
.Y(n_615)
);

OAI21xp5_ASAP7_75t_L g616 ( 
.A1(n_523),
.A2(n_520),
.B(n_493),
.Y(n_616)
);

NAND2x1p5_ASAP7_75t_L g617 ( 
.A(n_528),
.B(n_542),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_541),
.B(n_423),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_523),
.A2(n_422),
.B(n_420),
.Y(n_619)
);

INVx3_ASAP7_75t_L g620 ( 
.A(n_542),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_542),
.Y(n_621)
);

NAND3xp33_ASAP7_75t_L g622 ( 
.A(n_515),
.B(n_437),
.C(n_434),
.Y(n_622)
);

OAI22xp5_ASAP7_75t_L g623 ( 
.A1(n_536),
.A2(n_420),
.B1(n_366),
.B2(n_511),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_542),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_515),
.B(n_437),
.C(n_434),
.Y(n_625)
);

AOI21xp33_ASAP7_75t_L g626 ( 
.A1(n_557),
.A2(n_550),
.B(n_525),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_600),
.Y(n_627)
);

CKINVDCx8_ASAP7_75t_R g628 ( 
.A(n_565),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_602),
.B(n_609),
.Y(n_629)
);

BUFx4_ASAP7_75t_SL g630 ( 
.A(n_594),
.Y(n_630)
);

AO21x2_ASAP7_75t_L g631 ( 
.A1(n_595),
.A2(n_607),
.B(n_616),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_565),
.B(n_572),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_593),
.B(n_623),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_582),
.Y(n_634)
);

AO32x2_ASAP7_75t_L g635 ( 
.A1(n_561),
.A2(n_593),
.A3(n_623),
.B1(n_586),
.B2(n_581),
.Y(n_635)
);

NOR2x1p5_ASAP7_75t_L g636 ( 
.A(n_601),
.B(n_580),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_573),
.Y(n_637)
);

NAND2x1p5_ASAP7_75t_L g638 ( 
.A(n_562),
.B(n_603),
.Y(n_638)
);

OA21x2_ASAP7_75t_L g639 ( 
.A1(n_606),
.A2(n_610),
.B(n_619),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_574),
.Y(n_640)
);

O2A1O1Ixp33_ASAP7_75t_L g641 ( 
.A1(n_596),
.A2(n_626),
.B(n_561),
.C(n_571),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_613),
.A2(n_560),
.B1(n_596),
.B2(n_626),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_597),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_564),
.Y(n_644)
);

CKINVDCx20_ASAP7_75t_R g645 ( 
.A(n_608),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_577),
.Y(n_646)
);

CKINVDCx11_ASAP7_75t_R g647 ( 
.A(n_588),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_563),
.Y(n_648)
);

OAI21xp5_ASAP7_75t_L g649 ( 
.A1(n_622),
.A2(n_625),
.B(n_567),
.Y(n_649)
);

AND2x2_ASAP7_75t_L g650 ( 
.A(n_598),
.B(n_614),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_590),
.A2(n_570),
.B1(n_599),
.B2(n_569),
.Y(n_651)
);

HB1xp67_ASAP7_75t_L g652 ( 
.A(n_592),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_566),
.Y(n_653)
);

NOR2xp67_ASAP7_75t_L g654 ( 
.A(n_618),
.B(n_624),
.Y(n_654)
);

OA21x2_ASAP7_75t_L g655 ( 
.A1(n_591),
.A2(n_605),
.B(n_558),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_559),
.B(n_584),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_568),
.Y(n_657)
);

NAND2x1p5_ASAP7_75t_L g658 ( 
.A(n_562),
.B(n_624),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_566),
.Y(n_659)
);

AND2x2_ASAP7_75t_L g660 ( 
.A(n_604),
.B(n_615),
.Y(n_660)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_611),
.Y(n_661)
);

OAI21x1_ASAP7_75t_L g662 ( 
.A1(n_587),
.A2(n_591),
.B(n_589),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_617),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_612),
.Y(n_664)
);

BUFx3_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

NAND2x1p5_ASAP7_75t_L g666 ( 
.A(n_620),
.B(n_621),
.Y(n_666)
);

AOI21x1_ASAP7_75t_L g667 ( 
.A1(n_583),
.A2(n_575),
.B(n_604),
.Y(n_667)
);

AOI21xp5_ASAP7_75t_L g668 ( 
.A1(n_621),
.A2(n_620),
.B(n_575),
.Y(n_668)
);

NAND2x1p5_ASAP7_75t_L g669 ( 
.A(n_578),
.B(n_579),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_593),
.A2(n_623),
.B1(n_560),
.B2(n_561),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_566),
.B(n_489),
.Y(n_671)
);

OAI22xp33_ASAP7_75t_L g672 ( 
.A1(n_593),
.A2(n_623),
.B1(n_560),
.B2(n_585),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_566),
.B(n_489),
.Y(n_673)
);

INVx3_ASAP7_75t_L g674 ( 
.A(n_566),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_596),
.A2(n_626),
.B(n_576),
.C(n_561),
.Y(n_675)
);

OA21x2_ASAP7_75t_L g676 ( 
.A1(n_595),
.A2(n_616),
.B(n_607),
.Y(n_676)
);

AO21x2_ASAP7_75t_L g677 ( 
.A1(n_595),
.A2(n_616),
.B(n_607),
.Y(n_677)
);

AOI22xp33_ASAP7_75t_L g678 ( 
.A1(n_602),
.A2(n_609),
.B1(n_613),
.B2(n_571),
.Y(n_678)
);

INVxp67_ASAP7_75t_SL g679 ( 
.A(n_593),
.Y(n_679)
);

OA21x2_ASAP7_75t_L g680 ( 
.A1(n_595),
.A2(n_616),
.B(n_607),
.Y(n_680)
);

OR2x6_ASAP7_75t_L g681 ( 
.A(n_566),
.B(n_489),
.Y(n_681)
);

OA21x2_ASAP7_75t_L g682 ( 
.A1(n_595),
.A2(n_616),
.B(n_607),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_602),
.B(n_399),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_644),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_662),
.B(n_667),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_639),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_637),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_628),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_678),
.B(n_648),
.Y(n_689)
);

INVx3_ASAP7_75t_L g690 ( 
.A(n_663),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_645),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_640),
.Y(n_692)
);

BUFx4f_ASAP7_75t_SL g693 ( 
.A(n_645),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_646),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_629),
.B(n_632),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_678),
.B(n_627),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_634),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_683),
.B(n_629),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_630),
.Y(n_699)
);

INVxp33_ASAP7_75t_L g700 ( 
.A(n_652),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_663),
.Y(n_701)
);

NOR2xp33_ASAP7_75t_L g702 ( 
.A(n_632),
.B(n_660),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_630),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_665),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_653),
.Y(n_705)
);

NAND2x1p5_ASAP7_75t_L g706 ( 
.A(n_665),
.B(n_674),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_668),
.B(n_631),
.Y(n_707)
);

HB1xp67_ASAP7_75t_L g708 ( 
.A(n_652),
.Y(n_708)
);

BUFx2_ASAP7_75t_L g709 ( 
.A(n_635),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_635),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_650),
.B(n_643),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_674),
.Y(n_712)
);

AND2x4_ASAP7_75t_L g713 ( 
.A(n_631),
.B(n_677),
.Y(n_713)
);

INVx3_ASAP7_75t_L g714 ( 
.A(n_638),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_SL g715 ( 
.A1(n_670),
.A2(n_633),
.B(n_679),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_641),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_641),
.Y(n_717)
);

INVx2_ASAP7_75t_SL g718 ( 
.A(n_636),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_642),
.B(n_635),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_686),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_700),
.B(n_647),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_719),
.B(n_635),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_713),
.B(n_677),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_719),
.B(n_682),
.Y(n_724)
);

INVx5_ASAP7_75t_L g725 ( 
.A(n_714),
.Y(n_725)
);

NOR2x1_ASAP7_75t_SL g726 ( 
.A(n_684),
.B(n_670),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_713),
.B(n_676),
.Y(n_727)
);

OR2x2_ASAP7_75t_L g728 ( 
.A(n_689),
.B(n_676),
.Y(n_728)
);

BUFx2_ASAP7_75t_L g729 ( 
.A(n_704),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_685),
.Y(n_730)
);

BUFx2_ASAP7_75t_L g731 ( 
.A(n_704),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_689),
.B(n_696),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_696),
.B(n_680),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_707),
.B(n_649),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_716),
.B(n_642),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_708),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_695),
.A2(n_672),
.B1(n_679),
.B2(n_633),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_707),
.B(n_655),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_707),
.B(n_655),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_687),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_724),
.B(n_707),
.Y(n_741)
);

OAI22xp5_ASAP7_75t_L g742 ( 
.A1(n_737),
.A2(n_711),
.B1(n_698),
.B2(n_705),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_720),
.Y(n_743)
);

OR2x2_ASAP7_75t_L g744 ( 
.A(n_728),
.B(n_709),
.Y(n_744)
);

AND2x4_ASAP7_75t_L g745 ( 
.A(n_738),
.B(n_685),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_724),
.B(n_709),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_728),
.B(n_710),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_721),
.B(n_647),
.Y(n_748)
);

AND2x2_ASAP7_75t_L g749 ( 
.A(n_733),
.B(n_710),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_733),
.B(n_715),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_732),
.B(n_715),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_740),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_729),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_732),
.B(n_716),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_736),
.B(n_687),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_736),
.B(n_692),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_734),
.B(n_717),
.Y(n_757)
);

BUFx2_ASAP7_75t_L g758 ( 
.A(n_729),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_738),
.B(n_685),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_741),
.B(n_723),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_741),
.B(n_723),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_755),
.Y(n_762)
);

AND2x4_ASAP7_75t_L g763 ( 
.A(n_745),
.B(n_730),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_754),
.B(n_746),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_750),
.B(n_723),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_756),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_743),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_752),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_754),
.B(n_727),
.Y(n_769)
);

OR2x2_ASAP7_75t_L g770 ( 
.A(n_744),
.B(n_727),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_750),
.B(n_738),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_746),
.B(n_722),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_757),
.B(n_739),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_752),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_743),
.Y(n_775)
);

OR2x2_ASAP7_75t_L g776 ( 
.A(n_744),
.B(n_727),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_757),
.B(n_739),
.Y(n_777)
);

INVxp67_ASAP7_75t_SL g778 ( 
.A(n_767),
.Y(n_778)
);

BUFx2_ASAP7_75t_L g779 ( 
.A(n_763),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_764),
.B(n_769),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_769),
.B(n_747),
.Y(n_781)
);

AOI22xp33_ASAP7_75t_L g782 ( 
.A1(n_763),
.A2(n_751),
.B1(n_759),
.B2(n_745),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_768),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_774),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_767),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_760),
.B(n_749),
.Y(n_786)
);

A2O1A1Ixp33_ASAP7_75t_L g787 ( 
.A1(n_763),
.A2(n_742),
.B(n_718),
.C(n_688),
.Y(n_787)
);

OAI222xp33_ASAP7_75t_L g788 ( 
.A1(n_770),
.A2(n_753),
.B1(n_758),
.B2(n_747),
.C1(n_731),
.C2(n_759),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_762),
.B(n_722),
.Y(n_789)
);

OR2x2_ASAP7_75t_L g790 ( 
.A(n_770),
.B(n_776),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_775),
.Y(n_791)
);

OR2x2_ASAP7_75t_L g792 ( 
.A(n_781),
.B(n_776),
.Y(n_792)
);

AOI32xp33_ASAP7_75t_L g793 ( 
.A1(n_779),
.A2(n_771),
.A3(n_765),
.B1(n_761),
.B2(n_760),
.Y(n_793)
);

AOI21xp5_ASAP7_75t_L g794 ( 
.A1(n_787),
.A2(n_788),
.B(n_726),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_790),
.Y(n_795)
);

INVx1_ASAP7_75t_SL g796 ( 
.A(n_780),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_785),
.Y(n_797)
);

OAI21xp5_ASAP7_75t_L g798 ( 
.A1(n_787),
.A2(n_748),
.B(n_718),
.Y(n_798)
);

OAI322xp33_ASAP7_75t_L g799 ( 
.A1(n_781),
.A2(n_780),
.A3(n_766),
.B1(n_789),
.B2(n_772),
.C1(n_783),
.C2(n_784),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_778),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_785),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_791),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_792),
.Y(n_803)
);

AOI322xp5_ASAP7_75t_L g804 ( 
.A1(n_796),
.A2(n_786),
.A3(n_782),
.B1(n_773),
.B2(n_777),
.C1(n_765),
.C2(n_771),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_795),
.B(n_786),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_794),
.B(n_699),
.Y(n_806)
);

AOI21xp5_ASAP7_75t_L g807 ( 
.A1(n_806),
.A2(n_794),
.B(n_798),
.Y(n_807)
);

AOI222xp33_ASAP7_75t_L g808 ( 
.A1(n_803),
.A2(n_800),
.B1(n_801),
.B2(n_802),
.C1(n_797),
.C2(n_664),
.Y(n_808)
);

OAI211xp5_ASAP7_75t_SL g809 ( 
.A1(n_804),
.A2(n_793),
.B(n_675),
.C(n_735),
.Y(n_809)
);

INVxp67_ASAP7_75t_L g810 ( 
.A(n_807),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_SL g811 ( 
.A(n_808),
.B(n_703),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_810),
.B(n_809),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_811),
.B(n_805),
.Y(n_813)
);

AND2x4_ASAP7_75t_L g814 ( 
.A(n_813),
.B(n_691),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_812),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_814),
.Y(n_816)
);

NAND4xp75_ASAP7_75t_L g817 ( 
.A(n_815),
.B(n_693),
.C(n_654),
.D(n_814),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_816),
.A2(n_669),
.B1(n_797),
.B2(n_735),
.Y(n_818)
);

AO211x2_ASAP7_75t_L g819 ( 
.A1(n_817),
.A2(n_661),
.B(n_657),
.C(n_669),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_816),
.Y(n_820)
);

OR5x1_ASAP7_75t_L g821 ( 
.A(n_820),
.B(n_799),
.C(n_673),
.D(n_681),
.E(n_671),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_818),
.Y(n_822)
);

AOI22x1_ASAP7_75t_L g823 ( 
.A1(n_819),
.A2(n_659),
.B1(n_706),
.B2(n_666),
.Y(n_823)
);

XNOR2xp5_ASAP7_75t_L g824 ( 
.A(n_819),
.B(n_671),
.Y(n_824)
);

AOI22xp5_ASAP7_75t_L g825 ( 
.A1(n_819),
.A2(n_671),
.B1(n_673),
.B2(n_681),
.Y(n_825)
);

OAI22xp33_ASAP7_75t_L g826 ( 
.A1(n_822),
.A2(n_673),
.B1(n_681),
.B2(n_725),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_824),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_825),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_823),
.A2(n_643),
.B(n_656),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_821),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_822),
.Y(n_831)
);

INVx2_ASAP7_75t_L g832 ( 
.A(n_823),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_830),
.A2(n_702),
.B1(n_712),
.B2(n_651),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_L g834 ( 
.A1(n_831),
.A2(n_651),
.B1(n_706),
.B2(n_717),
.Y(n_834)
);

OAI22xp5_ASAP7_75t_L g835 ( 
.A1(n_832),
.A2(n_706),
.B1(n_694),
.B2(n_697),
.Y(n_835)
);

XNOR2xp5_ASAP7_75t_L g836 ( 
.A(n_826),
.B(n_658),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_R g837 ( 
.A(n_836),
.B(n_827),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_835),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_834),
.B(n_828),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_SL g840 ( 
.A1(n_838),
.A2(n_833),
.B(n_829),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_840),
.B(n_839),
.Y(n_841)
);

AOI22xp33_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_837),
.B1(n_701),
.B2(n_690),
.Y(n_842)
);


endmodule