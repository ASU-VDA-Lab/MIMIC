module fake_jpeg_22943_n_318 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_0),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx11_ASAP7_75t_SL g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx8_ASAP7_75t_SL g26 ( 
.A(n_12),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_3),
.B(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

INVx4_ASAP7_75t_SL g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_36),
.Y(n_42)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_19),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_39),
.C(n_24),
.Y(n_55)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g74 ( 
.A(n_41),
.Y(n_74)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_37),
.B(n_25),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_47),
.B(n_55),
.Y(n_64)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_33),
.Y(n_48)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_51),
.Y(n_84)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_50),
.A2(n_20),
.B1(n_40),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_57),
.A2(n_60),
.B1(n_65),
.B2(n_66),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_47),
.B(n_27),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g86 ( 
.A(n_58),
.B(n_73),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_59),
.B(n_61),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_52),
.A2(n_20),
.B1(n_40),
.B2(n_30),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_62),
.B(n_67),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_55),
.B(n_37),
.Y(n_63)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_63),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_71),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_41),
.A2(n_39),
.B(n_27),
.C(n_26),
.Y(n_73)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_40),
.B1(n_39),
.B2(n_20),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_79),
.B(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_43),
.B(n_27),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_80),
.Y(n_112)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_81),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_82),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_88),
.B(n_90),
.Y(n_123)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_68),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_91),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_96),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_26),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_93),
.A2(n_95),
.B(n_36),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_26),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_97),
.B(n_98),
.Y(n_133)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_71),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_100),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_76),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_40),
.B1(n_20),
.B2(n_34),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_102),
.A2(n_83),
.B1(n_84),
.B2(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

INVx2_ASAP7_75t_SL g107 ( 
.A(n_74),
.Y(n_107)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_72),
.A2(n_34),
.B1(n_54),
.B2(n_49),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_110),
.A2(n_45),
.B1(n_83),
.B2(n_74),
.Y(n_116)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_96),
.A2(n_59),
.B(n_64),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_114),
.A2(n_129),
.B(n_130),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_89),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_100),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_116),
.A2(n_117),
.B1(n_134),
.B2(n_139),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_64),
.B1(n_72),
.B2(n_82),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_54),
.B1(n_48),
.B2(n_45),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_121),
.A2(n_127),
.B1(n_131),
.B2(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_78),
.C(n_76),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_132),
.C(n_91),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_95),
.B(n_24),
.C(n_23),
.Y(n_128)
);

MAJx2_ASAP7_75t_L g167 ( 
.A(n_128),
.B(n_23),
.C(n_32),
.Y(n_167)
);

NAND2xp33_ASAP7_75t_SL g130 ( 
.A(n_95),
.B(n_19),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_38),
.B1(n_33),
.B2(n_84),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_103),
.B(n_78),
.C(n_33),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_111),
.A2(n_36),
.B1(n_83),
.B2(n_70),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_86),
.A2(n_17),
.B(n_18),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_18),
.B(n_17),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_111),
.A2(n_81),
.B1(n_75),
.B2(n_38),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_36),
.B1(n_34),
.B2(n_38),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_105),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_141),
.A2(n_107),
.B1(n_106),
.B2(n_34),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_93),
.B(n_112),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_142),
.A2(n_29),
.B(n_21),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_151),
.B1(n_160),
.B2(n_162),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_135),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_145),
.Y(n_178)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_121),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_153),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_148),
.B(n_157),
.C(n_128),
.Y(n_182)
);

AO21x2_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_93),
.B(n_107),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_149),
.A2(n_159),
.B1(n_32),
.B2(n_25),
.Y(n_190)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_136),
.A2(n_109),
.B1(n_94),
.B2(n_90),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_170),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_127),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g154 ( 
.A(n_118),
.B(n_92),
.CI(n_101),
.CON(n_154),
.SN(n_154)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_154),
.B(n_155),
.Y(n_185)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_133),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_104),
.Y(n_156)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_156),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_118),
.B(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_123),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_158),
.B(n_161),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_134),
.A2(n_85),
.B1(n_94),
.B2(n_36),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_138),
.A2(n_85),
.B1(n_113),
.B2(n_34),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_137),
.B(n_99),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_136),
.A2(n_135),
.B1(n_126),
.B2(n_124),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_163),
.B(n_164),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_119),
.B(n_99),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_131),
.A2(n_87),
.B1(n_23),
.B2(n_56),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_165),
.A2(n_168),
.B1(n_160),
.B2(n_143),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_149),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_117),
.A2(n_87),
.B1(n_17),
.B2(n_18),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_141),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_169),
.B(n_172),
.Y(n_206)
);

OAI32xp33_ASAP7_75t_L g170 ( 
.A1(n_114),
.A2(n_128),
.A3(n_130),
.B1(n_139),
.B2(n_119),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_124),
.B(n_29),
.Y(n_171)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_171),
.Y(n_184)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_120),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_32),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_19),
.Y(n_174)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_174),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_183),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_156),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_180),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_195),
.C(n_200),
.Y(n_221)
);

AOI322xp5_ASAP7_75t_L g183 ( 
.A1(n_166),
.A2(n_126),
.A3(n_140),
.B1(n_125),
.B2(n_32),
.C1(n_31),
.C2(n_15),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_144),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_187),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_140),
.Y(n_187)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_189),
.Y(n_226)
);

OAI21xp33_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_192),
.B(n_205),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g191 ( 
.A(n_154),
.B(n_19),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_191),
.B(n_170),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_157),
.B(n_32),
.C(n_19),
.Y(n_195)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_149),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_202),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_174),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_198),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_25),
.B1(n_31),
.B2(n_22),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_201),
.B1(n_203),
.B2(n_159),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_172),
.B(n_32),
.C(n_19),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_146),
.A2(n_31),
.B1(n_22),
.B2(n_16),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_149),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_22),
.B1(n_16),
.B2(n_15),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_148),
.B(n_16),
.C(n_15),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_204),
.B(n_152),
.C(n_147),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_207),
.B(n_208),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_177),
.A2(n_202),
.B(n_175),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_178),
.B(n_173),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_214),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_212),
.A2(n_213),
.B1(n_223),
.B2(n_225),
.Y(n_234)
);

OA22x2_ASAP7_75t_L g213 ( 
.A1(n_196),
.A2(n_143),
.B1(n_142),
.B2(n_165),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_206),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_176),
.B(n_147),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_228),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g218 ( 
.A(n_188),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_218),
.B(n_227),
.Y(n_243)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_189),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_222),
.B(n_191),
.C(n_195),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_177),
.A2(n_167),
.B1(n_168),
.B2(n_154),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g244 ( 
.A(n_224),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_205),
.A2(n_21),
.B(n_29),
.Y(n_225)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_28),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_199),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_231),
.B1(n_180),
.B2(n_192),
.Y(n_233)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_232),
.B(n_238),
.C(n_239),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_213),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_185),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_245),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_219),
.A2(n_181),
.B1(n_193),
.B2(n_198),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_236),
.A2(n_241),
.B1(n_247),
.B2(n_213),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_200),
.C(n_197),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_197),
.C(n_193),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_214),
.A2(n_190),
.B1(n_178),
.B2(n_184),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_217),
.B(n_204),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_242),
.B(n_249),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_228),
.B(n_230),
.C(n_222),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_211),
.A2(n_201),
.B1(n_179),
.B2(n_28),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_209),
.A2(n_179),
.B1(n_14),
.B2(n_13),
.Y(n_248)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_226),
.B(n_1),
.C(n_2),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_216),
.B(n_1),
.C(n_2),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_212),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_250),
.B(n_227),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_257),
.Y(n_269)
);

XNOR2x1_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_208),
.Y(n_253)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_253),
.B(n_242),
.Y(n_271)
);

NAND3xp33_ASAP7_75t_L g254 ( 
.A(n_237),
.B(n_223),
.C(n_225),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_236),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_256),
.B(n_258),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_243),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_251),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_260),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_215),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_262),
.B(n_265),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_263),
.A2(n_234),
.B1(n_244),
.B2(n_238),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_215),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_264),
.B(n_268),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_246),
.B(n_220),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_249),
.B(n_213),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_266),
.A2(n_11),
.B(n_4),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_240),
.B(n_14),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_271),
.B(n_268),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g273 ( 
.A(n_259),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_262),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_275),
.B(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_239),
.C(n_232),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_261),
.A2(n_235),
.B1(n_14),
.B2(n_12),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_277),
.A2(n_282),
.B1(n_5),
.B2(n_6),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_265),
.B(n_2),
.C(n_3),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_279),
.B(n_281),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_256),
.B(n_12),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_280),
.B(n_255),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_269),
.B(n_255),
.Y(n_283)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_283),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_271),
.A2(n_253),
.B1(n_254),
.B2(n_279),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_284),
.A2(n_294),
.B(n_6),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_285),
.B(n_286),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_292),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_11),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_293),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_278),
.B(n_3),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_272),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_290),
.A2(n_278),
.B1(n_272),
.B2(n_8),
.Y(n_295)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_295),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_289),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_284),
.A2(n_6),
.B(n_7),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g306 ( 
.A(n_300),
.B(n_303),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_7),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_288),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_302),
.B(n_9),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_306),
.A2(n_307),
.B(n_299),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_8),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_308),
.B(n_297),
.Y(n_311)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_309),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_310),
.C(n_302),
.Y(n_314)
);

AOI31xp33_ASAP7_75t_L g315 ( 
.A1(n_314),
.A2(n_297),
.A3(n_304),
.B(n_9),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_9),
.C(n_10),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_316),
.B(n_10),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_10),
.Y(n_318)
);


endmodule