module fake_aes_4464_n_33 (n_11, n_1, n_2, n_12, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_33);
input n_11;
input n_1;
input n_2;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_33;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_32;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
XOR2xp5_ASAP7_75t_L g14 ( .A(n_4), .B(n_9), .Y(n_14) );
INVxp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_4), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_7), .Y(n_17) );
CKINVDCx5p33_ASAP7_75t_R g18 ( .A(n_12), .Y(n_18) );
OAI21xp5_ASAP7_75t_L g19 ( .A1(n_13), .A2(n_6), .B(n_10), .Y(n_19) );
INVxp67_ASAP7_75t_SL g20 ( .A(n_15), .Y(n_20) );
INVxp67_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
OAI21xp5_ASAP7_75t_L g22 ( .A1(n_19), .A2(n_17), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
NAND3xp33_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .C(n_19), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
OAI22xp5_ASAP7_75t_L g26 ( .A1(n_24), .A2(n_16), .B1(n_14), .B2(n_2), .Y(n_26) );
AOI211x1_ASAP7_75t_SL g27 ( .A1(n_26), .A2(n_16), .B(n_1), .C(n_2), .Y(n_27) );
INVxp67_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
AOI211xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_0), .B(n_1), .C(n_3), .Y(n_29) );
BUFx2_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
NAND2xp5_ASAP7_75t_L g31 ( .A(n_30), .B(n_27), .Y(n_31) );
OAI21x1_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B(n_11), .Y(n_32) );
AOI21xp33_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_0), .B(n_3), .Y(n_33) );
endmodule