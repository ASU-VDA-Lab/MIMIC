module fake_jpeg_8319_n_192 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx16f_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

BUFx5_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_3),
.B(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_21),
.Y(n_25)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

NAND2xp33_ASAP7_75t_SL g39 ( 
.A(n_27),
.B(n_29),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx4_ASAP7_75t_SL g38 ( 
.A(n_28),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g29 ( 
.A1(n_14),
.A2(n_0),
.B(n_1),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_33),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_33),
.B1(n_19),
.B2(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_43),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_20),
.Y(n_42)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_29),
.B(n_20),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_24),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_24),
.Y(n_46)
);

AO22x1_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_14),
.B1(n_15),
.B2(n_30),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_51),
.B1(n_58),
.B2(n_35),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_33),
.B1(n_26),
.B2(n_17),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_49),
.A2(n_54),
.B1(n_36),
.B2(n_38),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_22),
.B1(n_19),
.B2(n_12),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_52),
.A2(n_59),
.B1(n_38),
.B2(n_36),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_14),
.B1(n_27),
.B2(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_18),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_60),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx24_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_43),
.A2(n_14),
.B1(n_22),
.B2(n_23),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_36),
.A2(n_22),
.B1(n_12),
.B2(n_23),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_62),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_37),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_45),
.B(n_46),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_65),
.Y(n_82)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_66),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_67),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_68),
.A2(n_61),
.B1(n_62),
.B2(n_53),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_50),
.B(n_46),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_70),
.B(n_30),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_48),
.A2(n_42),
.B(n_41),
.C(n_45),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_71),
.B(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_47),
.B(n_0),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_72),
.B(n_18),
.C(n_16),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

OA22x2_ASAP7_75t_L g85 ( 
.A1(n_74),
.A2(n_44),
.B1(n_60),
.B2(n_13),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_54),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_78),
.Y(n_96)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_58),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_80),
.A2(n_38),
.B1(n_13),
.B2(n_25),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_84),
.B(n_86),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_85),
.A2(n_91),
.B1(n_69),
.B2(n_73),
.Y(n_98)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_48),
.B1(n_53),
.B2(n_37),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_87),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_37),
.B1(n_44),
.B2(n_41),
.Y(n_90)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_37),
.B1(n_30),
.B2(n_28),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_63),
.B(n_66),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_95),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_98),
.A2(n_108),
.B1(n_107),
.B2(n_109),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_64),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_99),
.Y(n_123)
);

INVx13_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_88),
.A2(n_72),
.B(n_79),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_102),
.A2(n_108),
.B(n_111),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_94),
.B(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_106),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_97),
.B(n_71),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_89),
.A2(n_72),
.B(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_87),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_109),
.B(n_90),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_93),
.B(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_113),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_83),
.B(n_10),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_84),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_112),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_83),
.B(n_96),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g115 ( 
.A(n_102),
.B(n_104),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_124),
.C(n_131),
.Y(n_135)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_114),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_116),
.B(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_117),
.B(n_24),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_82),
.B1(n_91),
.B2(n_85),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_119),
.A2(n_103),
.B1(n_111),
.B2(n_69),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_101),
.A2(n_91),
.B1(n_86),
.B2(n_85),
.Y(n_120)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_120),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_81),
.C(n_92),
.Y(n_124)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_113),
.Y(n_126)
);

OAI22x1_ASAP7_75t_L g127 ( 
.A1(n_98),
.A2(n_85),
.B1(n_91),
.B2(n_76),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_127),
.A2(n_129),
.B(n_40),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_21),
.Y(n_130)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_99),
.B(n_25),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_115),
.B(n_110),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_137),
.C(n_144),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_125),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_134),
.A2(n_118),
.B(n_130),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_124),
.B(n_105),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_136),
.B(n_142),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_103),
.C(n_100),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_140),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_141),
.A2(n_143),
.B1(n_119),
.B2(n_121),
.Y(n_152)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_125),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_32),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_135),
.B(n_128),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_137),
.C(n_144),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_135),
.B(n_128),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g160 ( 
.A(n_148),
.B(n_151),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_24),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_133),
.B(n_118),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_6),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_139),
.A2(n_120),
.B1(n_122),
.B2(n_117),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_154),
.A2(n_139),
.B1(n_132),
.B2(n_145),
.Y(n_158)
);

XOR2x1_ASAP7_75t_SL g155 ( 
.A(n_141),
.B(n_24),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_24),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_161),
.C(n_148),
.Y(n_171)
);

INVxp33_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g159 ( 
.A(n_156),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_162),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_153),
.B(n_76),
.C(n_32),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_163),
.A2(n_165),
.B(n_76),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_147),
.A2(n_38),
.B1(n_76),
.B2(n_2),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_164),
.A2(n_155),
.B(n_154),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_160),
.A2(n_153),
.B(n_149),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_168),
.A2(n_6),
.B(n_1),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_169),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_170),
.B(n_162),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_171),
.B(n_172),
.C(n_5),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_146),
.C(n_151),
.Y(n_172)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_173),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_176),
.C(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_166),
.B(n_40),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_167),
.B(n_56),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_177),
.A2(n_2),
.B(n_3),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_0),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_180),
.A2(n_10),
.B(n_5),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_175),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_181),
.B(n_183),
.C(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_10),
.B(n_7),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_180),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_188),
.A2(n_179),
.B(n_7),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_187),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_7),
.C(n_8),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_8),
.Y(n_192)
);


endmodule