module real_aes_1472_n_382 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_379, n_374, n_26, n_235, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_382);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_379;
input n_374;
input n_26;
input n_235;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_382;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_977;
wire n_503;
wire n_905;
wire n_386;
wire n_635;
wire n_673;
wire n_518;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_1004;
wire n_577;
wire n_580;
wire n_469;
wire n_987;
wire n_759;
wire n_979;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_974;
wire n_919;
wire n_857;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_1034;
wire n_549;
wire n_694;
wire n_491;
wire n_923;
wire n_571;
wire n_894;
wire n_952;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_989;
wire n_773;
wire n_401;
wire n_538;
wire n_431;
wire n_1044;
wire n_963;
wire n_865;
wire n_537;
wire n_551;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_955;
wire n_889;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1021;
wire n_677;
wire n_958;
wire n_1046;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_961;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_578;
wire n_994;
wire n_528;
wire n_495;
wire n_892;
wire n_384;
wire n_744;
wire n_938;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_951;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_976;
wire n_1049;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_693;
wire n_496;
wire n_962;
wire n_468;
wire n_746;
wire n_755;
wire n_1025;
wire n_532;
wire n_656;
wire n_409;
wire n_748;
wire n_860;
wire n_909;
wire n_523;
wire n_781;
wire n_996;
wire n_439;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_455;
wire n_725;
wire n_960;
wire n_671;
wire n_973;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_885;
wire n_1059;
wire n_950;
wire n_993;
wire n_493;
wire n_664;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_936;
wire n_610;
wire n_1035;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_940;
wire n_770;
wire n_808;
wire n_722;
wire n_745;
wire n_867;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_1006;
wire n_690;
wire n_629;
wire n_1053;
wire n_499;
wire n_508;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_769;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_733;
wire n_602;
wire n_617;
wire n_402;
wire n_552;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1037;
wire n_1031;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_869;
wire n_613;
wire n_642;
wire n_387;
wire n_957;
wire n_995;
wire n_702;
wire n_954;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_464;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_713;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_756;
wire n_997;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_727;
wire n_1014;
wire n_397;
wire n_749;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_1001;
wire n_494;
wire n_711;
wire n_864;
wire n_1027;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_845;
wire n_850;
wire n_1043;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_653;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_789;
wire n_544;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_787;
wire n_1052;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_456;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_719;
wire n_1045;
wire n_465;
wire n_473;
wire n_566;
wire n_837;
wire n_967;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_597;
wire n_640;
wire n_483;
wire n_611;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_1040;
wire n_393;
wire n_703;
wire n_652;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_1039;
wire n_574;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp33_ASAP7_75t_L g585 ( .A1(n_0), .A2(n_329), .B1(n_586), .B2(n_587), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g623 ( .A1(n_1), .A2(n_219), .B1(n_592), .B2(n_624), .Y(n_623) );
AOI22xp33_ASAP7_75t_SL g907 ( .A1(n_2), .A2(n_281), .B1(n_608), .B2(n_686), .Y(n_907) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_3), .A2(n_116), .B1(n_485), .B2(n_684), .Y(n_1016) );
AOI22xp33_ASAP7_75t_L g901 ( .A1(n_4), .A2(n_125), .B1(n_693), .B2(n_694), .Y(n_901) );
CKINVDCx20_ASAP7_75t_R g915 ( .A(n_5), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1055 ( .A1(n_6), .A2(n_187), .B1(n_690), .B2(n_693), .Y(n_1055) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_7), .A2(n_81), .B1(n_501), .B2(n_697), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_8), .B(n_574), .Y(n_573) );
AOI22xp33_ASAP7_75t_SL g648 ( .A1(n_9), .A2(n_256), .B1(n_586), .B2(n_587), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g782 ( .A1(n_10), .A2(n_92), .B1(n_533), .B2(n_578), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_11), .A2(n_288), .B1(n_689), .B2(n_690), .Y(n_688) );
AOI22xp33_ASAP7_75t_L g786 ( .A1(n_12), .A2(n_238), .B1(n_787), .B2(n_789), .Y(n_786) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_13), .A2(n_204), .B1(n_594), .B2(n_595), .Y(n_930) );
AOI22xp33_ASAP7_75t_SL g944 ( .A1(n_14), .A2(n_79), .B1(n_581), .B2(n_582), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_15), .A2(n_141), .B1(n_424), .B2(n_609), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g1050 ( .A1(n_16), .A2(n_169), .B1(n_681), .B2(n_682), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g905 ( .A1(n_17), .A2(n_194), .B1(n_524), .B2(n_684), .Y(n_905) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_18), .A2(n_244), .B1(n_481), .B2(n_484), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g945 ( .A1(n_19), .A2(n_220), .B1(n_579), .B2(n_643), .Y(n_945) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_20), .A2(n_180), .B1(n_557), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_SL g652 ( .A1(n_21), .A2(n_177), .B1(n_592), .B2(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g764 ( .A1(n_22), .A2(n_152), .B1(n_612), .B2(n_682), .Y(n_764) );
XOR2x2_ASAP7_75t_L g732 ( .A(n_23), .B(n_733), .Y(n_732) );
AO222x2_ASAP7_75t_L g918 ( .A1(n_24), .A2(n_147), .B1(n_240), .B2(n_395), .C1(n_415), .C2(n_919), .Y(n_918) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_25), .A2(n_191), .B1(n_557), .B2(n_771), .Y(n_1052) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_26), .A2(n_139), .B1(n_694), .B2(n_708), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g922 ( .A1(n_27), .A2(n_338), .B1(n_643), .B2(n_923), .Y(n_922) );
INVx1_ASAP7_75t_SL g400 ( .A(n_28), .Y(n_400) );
NOR2xp33_ASAP7_75t_L g999 ( .A(n_28), .B(n_40), .Y(n_999) );
CKINVDCx20_ASAP7_75t_R g940 ( .A(n_29), .Y(n_940) );
OA22x2_ASAP7_75t_L g800 ( .A1(n_30), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g801 ( .A(n_30), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_31), .A2(n_174), .B1(n_716), .B2(n_771), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_32), .A2(n_377), .B1(n_693), .B2(n_743), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g423 ( .A1(n_33), .A2(n_136), .B1(n_424), .B2(n_428), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g593 ( .A1(n_34), .A2(n_296), .B1(n_594), .B2(n_595), .Y(n_593) );
AOI22x1_ASAP7_75t_L g951 ( .A1(n_35), .A2(n_199), .B1(n_452), .B2(n_594), .Y(n_951) );
AOI22xp33_ASAP7_75t_L g974 ( .A1(n_36), .A2(n_115), .B1(n_643), .B2(n_923), .Y(n_974) );
AOI22xp33_ASAP7_75t_L g712 ( .A1(n_37), .A2(n_217), .B1(n_498), .B2(n_713), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g814 ( .A1(n_38), .A2(n_367), .B1(n_682), .B2(n_815), .Y(n_814) );
AO21x1_ASAP7_75t_SL g1000 ( .A1(n_39), .A2(n_1001), .B(n_1009), .Y(n_1000) );
AO22x2_ASAP7_75t_L g402 ( .A1(n_40), .A2(n_357), .B1(n_399), .B2(n_403), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g463 ( .A1(n_41), .A2(n_173), .B1(n_464), .B2(n_467), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g851 ( .A1(n_42), .A2(n_212), .B1(n_690), .B2(n_741), .Y(n_851) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_43), .A2(n_55), .B1(n_608), .B2(n_686), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_44), .A2(n_112), .B1(n_693), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g742 ( .A1(n_45), .A2(n_366), .B1(n_708), .B2(n_743), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_46), .A2(n_153), .B1(n_492), .B2(n_494), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_47), .A2(n_183), .B1(n_485), .B2(n_602), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g1053 ( .A1(n_48), .A2(n_80), .B1(n_444), .B2(n_498), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g852 ( .A1(n_49), .A2(n_289), .B1(n_460), .B2(n_708), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g965 ( .A1(n_50), .A2(n_342), .B1(n_444), .B2(n_769), .Y(n_965) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_51), .B(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g401 ( .A(n_52), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g654 ( .A1(n_53), .A2(n_311), .B1(n_591), .B2(n_595), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g963 ( .A1(n_54), .A2(n_245), .B1(n_708), .B2(n_716), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_56), .A2(n_235), .B1(n_496), .B2(n_498), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_57), .A2(n_308), .B1(n_594), .B2(n_650), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g747 ( .A1(n_58), .A2(n_131), .B1(n_748), .B2(n_749), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_59), .A2(n_354), .B1(n_457), .B2(n_617), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g822 ( .A1(n_60), .A2(n_249), .B1(n_684), .B2(n_823), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_61), .A2(n_214), .B1(n_837), .B2(n_838), .Y(n_836) );
AOI22xp5_ASAP7_75t_L g1010 ( .A1(n_62), .A2(n_1011), .B1(n_1012), .B2(n_1034), .Y(n_1010) );
CKINVDCx20_ASAP7_75t_R g1034 ( .A(n_62), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1030 ( .A1(n_63), .A2(n_347), .B1(n_444), .B2(n_447), .Y(n_1030) );
AO22x2_ASAP7_75t_L g409 ( .A1(n_64), .A2(n_196), .B1(n_399), .B2(n_410), .Y(n_409) );
AOI22xp33_ASAP7_75t_L g774 ( .A1(n_65), .A2(n_312), .B1(n_690), .B2(n_696), .Y(n_774) );
AOI22xp33_ASAP7_75t_L g793 ( .A1(n_66), .A2(n_84), .B1(n_549), .B2(n_794), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g1029 ( .A1(n_67), .A2(n_201), .B1(n_549), .B2(n_696), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_68), .A2(n_143), .B1(n_595), .B2(n_662), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_69), .A2(n_237), .B1(n_444), .B2(n_498), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_70), .A2(n_106), .B1(n_413), .B2(n_419), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g580 ( .A1(n_71), .A2(n_163), .B1(n_581), .B2(n_582), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_72), .A2(n_295), .B1(n_450), .B2(n_694), .Y(n_879) );
AOI22xp33_ASAP7_75t_L g449 ( .A1(n_73), .A2(n_325), .B1(n_450), .B2(n_452), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g952 ( .A1(n_74), .A2(n_167), .B1(n_595), .B2(n_650), .Y(n_952) );
AOI22xp5_ASAP7_75t_L g834 ( .A1(n_75), .A2(n_202), .B1(n_494), .B2(n_708), .Y(n_834) );
AOI22xp5_ASAP7_75t_L g588 ( .A1(n_76), .A2(n_157), .B1(n_452), .B2(n_464), .Y(n_588) );
AOI22xp33_ASAP7_75t_SL g926 ( .A1(n_77), .A2(n_114), .B1(n_586), .B2(n_587), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g983 ( .A1(n_78), .A2(n_293), .B1(n_650), .B2(n_653), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_82), .A2(n_257), .B1(n_536), .B2(n_538), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_83), .A2(n_253), .B1(n_415), .B2(n_419), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_85), .A2(n_99), .B1(n_457), .B2(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_86), .A2(n_368), .B1(n_485), .B2(n_684), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_87), .A2(n_228), .B1(n_447), .B2(n_713), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g858 ( .A1(n_88), .A2(n_306), .B1(n_538), .B2(n_815), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g767 ( .A1(n_89), .A2(n_285), .B1(n_768), .B2(n_769), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g839 ( .A1(n_90), .A2(n_137), .B1(n_554), .B2(n_840), .Y(n_839) );
AO222x2_ASAP7_75t_L g640 ( .A1(n_91), .A2(n_211), .B1(n_360), .B2(n_395), .C1(n_579), .C2(n_582), .Y(n_640) );
AOI22xp33_ASAP7_75t_SL g894 ( .A1(n_93), .A2(n_127), .B1(n_895), .B2(n_897), .Y(n_894) );
AOI22xp5_ASAP7_75t_L g577 ( .A1(n_94), .A2(n_233), .B1(n_578), .B2(n_579), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g645 ( .A1(n_95), .A2(n_259), .B1(n_415), .B2(n_419), .Y(n_645) );
CKINVDCx20_ASAP7_75t_R g558 ( .A(n_96), .Y(n_558) );
AOI222xp33_ASAP7_75t_L g859 ( .A1(n_97), .A2(n_175), .B1(n_345), .B2(n_485), .C1(n_759), .C2(n_860), .Y(n_859) );
OA22x2_ASAP7_75t_L g512 ( .A1(n_98), .A2(n_513), .B1(n_514), .B2(n_515), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_98), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g959 ( .A1(n_100), .A2(n_144), .B1(n_279), .B2(n_612), .C1(n_759), .C2(n_830), .Y(n_959) );
AOI22xp33_ASAP7_75t_L g975 ( .A1(n_101), .A2(n_158), .B1(n_582), .B2(n_644), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g783 ( .A1(n_102), .A2(n_275), .B1(n_722), .B2(n_784), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_103), .A2(n_236), .B1(n_748), .B2(n_749), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g874 ( .A1(n_104), .A2(n_197), .B1(n_875), .B2(n_877), .Y(n_874) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_105), .A2(n_126), .B1(n_504), .B2(n_746), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_107), .A2(n_336), .B1(n_457), .B2(n_460), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_108), .B(n_474), .Y(n_473) );
CKINVDCx20_ASAP7_75t_R g541 ( .A(n_109), .Y(n_541) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_110), .A2(n_239), .B1(n_444), .B2(n_447), .Y(n_808) );
AO22x2_ASAP7_75t_L g406 ( .A1(n_111), .A2(n_292), .B1(n_399), .B2(n_407), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_113), .A2(n_305), .B1(n_681), .B2(n_682), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g908 ( .A1(n_117), .A2(n_155), .B1(n_681), .B2(n_830), .Y(n_908) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_118), .A2(n_376), .B1(n_457), .B2(n_716), .Y(n_715) );
AO21x2_ASAP7_75t_L g868 ( .A1(n_119), .A2(n_869), .B(n_885), .Y(n_868) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_119), .B(n_871), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_120), .A2(n_271), .B1(n_693), .B2(n_694), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_121), .A2(n_122), .B1(n_523), .B2(n_526), .Y(n_883) );
AOI22xp5_ASAP7_75t_L g1033 ( .A1(n_123), .A2(n_146), .B1(n_689), .B2(n_716), .Y(n_1033) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_124), .A2(n_269), .B1(n_488), .B2(n_489), .Y(n_487) );
INVx1_ASAP7_75t_L g861 ( .A(n_128), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g978 ( .A1(n_129), .A2(n_352), .B1(n_587), .B2(n_979), .Y(n_978) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_130), .Y(n_543) );
AOI22xp33_ASAP7_75t_L g982 ( .A1(n_132), .A2(n_206), .B1(n_592), .B2(n_624), .Y(n_982) );
AOI22xp5_ASAP7_75t_L g522 ( .A1(n_133), .A2(n_333), .B1(n_523), .B2(n_526), .Y(n_522) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_134), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_135), .B(n_475), .Y(n_1017) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_138), .A2(n_232), .B1(n_424), .B2(n_686), .Y(n_961) );
CKINVDCx20_ASAP7_75t_R g596 ( .A(n_140), .Y(n_596) );
OA22x2_ASAP7_75t_L g469 ( .A1(n_142), .A2(n_470), .B1(n_471), .B2(n_506), .Y(n_469) );
CKINVDCx20_ASAP7_75t_R g470 ( .A(n_142), .Y(n_470) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_145), .A2(n_327), .B1(n_716), .B2(n_741), .Y(n_740) );
AOI22xp5_ASAP7_75t_L g829 ( .A1(n_148), .A2(n_171), .B1(n_612), .B2(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_149), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g927 ( .A1(n_150), .A2(n_156), .B1(n_650), .B2(n_653), .Y(n_927) );
AOI22xp5_ASAP7_75t_L g824 ( .A1(n_151), .A2(n_332), .B1(n_428), .B2(n_825), .Y(n_824) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_154), .A2(n_176), .B1(n_536), .B2(n_538), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_159), .B(n_605), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_160), .A2(n_241), .B1(n_689), .B2(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_161), .A2(n_294), .B1(n_447), .B2(n_497), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g669 ( .A1(n_162), .A2(n_364), .B1(n_433), .B2(n_538), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_164), .B(n_519), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_165), .A2(n_189), .B1(n_450), .B2(n_504), .Y(n_503) );
AOI22xp33_ASAP7_75t_SL g443 ( .A1(n_166), .A2(n_324), .B1(n_444), .B2(n_446), .Y(n_443) );
AOI222xp33_ASAP7_75t_L g1057 ( .A1(n_168), .A2(n_181), .B1(n_225), .B2(n_475), .C1(n_485), .C2(n_684), .Y(n_1057) );
AOI22xp33_ASAP7_75t_L g736 ( .A1(n_170), .A2(n_348), .B1(n_479), .B2(n_612), .Y(n_736) );
OA22x2_ASAP7_75t_L g954 ( .A1(n_172), .A2(n_955), .B1(n_956), .B2(n_957), .Y(n_954) );
INVx1_ASAP7_75t_L g955 ( .A(n_172), .Y(n_955) );
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_178), .A2(n_230), .B1(n_424), .B2(n_686), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_179), .A2(n_346), .B1(n_452), .B2(n_621), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g724 ( .A1(n_182), .A2(n_378), .B1(n_484), .B2(n_526), .Y(n_724) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_184), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_185), .A2(n_209), .B1(n_428), .B2(n_608), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_186), .A2(n_302), .B1(n_530), .B2(n_533), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_188), .A2(n_261), .B1(n_608), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_190), .A2(n_365), .B1(n_485), .B2(n_684), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g792 ( .A1(n_192), .A2(n_380), .B1(n_557), .B2(n_771), .Y(n_792) );
AOI22xp33_ASAP7_75t_SL g899 ( .A1(n_193), .A2(n_313), .B1(n_696), .B2(n_900), .Y(n_899) );
AOI22xp33_ASAP7_75t_L g721 ( .A1(n_195), .A2(n_254), .B1(n_613), .B2(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g998 ( .A(n_196), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g980 ( .A1(n_198), .A2(n_231), .B1(n_594), .B2(n_595), .Y(n_980) );
AOI22xp33_ASAP7_75t_L g948 ( .A1(n_200), .A2(n_262), .B1(n_586), .B2(n_587), .Y(n_948) );
XNOR2xp5_ASAP7_75t_L g935 ( .A(n_203), .B(n_936), .Y(n_935) );
AOI22xp5_ASAP7_75t_L g607 ( .A1(n_205), .A2(n_358), .B1(n_608), .B2(n_609), .Y(n_607) );
INVx1_ASAP7_75t_L g904 ( .A(n_207), .Y(n_904) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_208), .A2(n_323), .B1(n_643), .B2(n_644), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g565 ( .A(n_210), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_213), .A2(n_272), .B1(n_684), .B2(n_813), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_215), .A2(n_284), .B1(n_707), .B2(n_709), .Y(n_706) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_216), .A2(n_315), .B1(n_450), .B2(n_504), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g960 ( .A1(n_218), .A2(n_372), .B1(n_684), .B2(n_813), .Y(n_960) );
INVx2_ASAP7_75t_L g1006 ( .A(n_221), .Y(n_1006) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_222), .A2(n_369), .B1(n_591), .B2(n_592), .Y(n_929) );
OA22x2_ASAP7_75t_L g818 ( .A1(n_223), .A2(n_819), .B1(n_842), .B2(n_843), .Y(n_818) );
CKINVDCx20_ASAP7_75t_R g842 ( .A(n_223), .Y(n_842) );
AOI22xp33_ASAP7_75t_SL g773 ( .A1(n_224), .A2(n_276), .B1(n_549), .B2(n_693), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_226), .A2(n_246), .B1(n_467), .B2(n_837), .Y(n_855) );
INVx1_ASAP7_75t_L g1041 ( .A(n_227), .Y(n_1041) );
AOI22xp5_ASAP7_75t_L g1044 ( .A1(n_227), .A2(n_1041), .B1(n_1045), .B2(n_1058), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g668 ( .A1(n_229), .A2(n_255), .B1(n_424), .B2(n_428), .Y(n_668) );
AOI22xp5_ASAP7_75t_L g964 ( .A1(n_234), .A2(n_320), .B1(n_690), .B2(n_771), .Y(n_964) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_242), .A2(n_287), .B1(n_497), .B2(n_769), .Y(n_833) );
AOI22xp5_ASAP7_75t_L g1047 ( .A1(n_243), .A2(n_316), .B1(n_424), .B2(n_1048), .Y(n_1047) );
CKINVDCx16_ASAP7_75t_R g984 ( .A(n_247), .Y(n_984) );
AOI22xp5_ASAP7_75t_L g888 ( .A1(n_248), .A2(n_889), .B1(n_890), .B2(n_909), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_248), .Y(n_889) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_250), .A2(n_637), .B1(n_638), .B2(n_655), .Y(n_636) );
INVx1_ASAP7_75t_L g655 ( .A(n_250), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_251), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_252), .A2(n_344), .B1(n_433), .B2(n_437), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g972 ( .A1(n_258), .A2(n_339), .B1(n_415), .B2(n_919), .Y(n_972) );
CKINVDCx20_ASAP7_75t_R g939 ( .A(n_260), .Y(n_939) );
AOI22xp5_ASAP7_75t_L g761 ( .A1(n_263), .A2(n_273), .B1(n_485), .B2(n_684), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_264), .A2(n_321), .B1(n_433), .B2(n_479), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g921 ( .A1(n_265), .A2(n_290), .B1(n_582), .B2(n_644), .Y(n_921) );
AOI22xp33_ASAP7_75t_L g949 ( .A1(n_266), .A2(n_381), .B1(n_592), .B2(n_624), .Y(n_949) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_267), .A2(n_351), .B1(n_622), .B2(n_708), .Y(n_807) );
NAND2xp5_ASAP7_75t_L g881 ( .A(n_268), .B(n_605), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g601 ( .A1(n_270), .A2(n_304), .B1(n_485), .B2(n_602), .Y(n_601) );
XNOR2x1_ASAP7_75t_L g754 ( .A(n_274), .B(n_755), .Y(n_754) );
CKINVDCx20_ASAP7_75t_R g1019 ( .A(n_277), .Y(n_1019) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_278), .A2(n_356), .B1(n_621), .B2(n_622), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_280), .A2(n_353), .B1(n_446), .B2(n_497), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_282), .B(n_475), .Y(n_735) );
OA22x2_ASAP7_75t_L g701 ( .A1(n_283), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_283), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_286), .Y(n_547) );
AOI22xp33_ASAP7_75t_SL g893 ( .A1(n_291), .A2(n_331), .B1(n_689), .B2(n_716), .Y(n_893) );
NOR2xp33_ASAP7_75t_L g996 ( .A(n_292), .B(n_997), .Y(n_996) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_297), .A2(n_343), .B1(n_591), .B2(n_592), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_298), .B(n_475), .Y(n_827) );
CKINVDCx20_ASAP7_75t_R g1026 ( .A(n_299), .Y(n_1026) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_300), .A2(n_379), .B1(n_444), .B2(n_446), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g941 ( .A(n_301), .Y(n_941) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_303), .A2(n_335), .B1(n_530), .B2(n_533), .Y(n_884) );
CKINVDCx20_ASAP7_75t_R g760 ( .A(n_307), .Y(n_760) );
AOI22xp33_ASAP7_75t_L g966 ( .A1(n_309), .A2(n_330), .B1(n_693), .B2(n_810), .Y(n_966) );
INVx3_ASAP7_75t_L g399 ( .A(n_310), .Y(n_399) );
AOI22xp33_ASAP7_75t_L g590 ( .A1(n_314), .A2(n_326), .B1(n_591), .B2(n_592), .Y(n_590) );
AOI222xp33_ASAP7_75t_L g795 ( .A1(n_317), .A2(n_355), .B1(n_363), .B2(n_475), .C1(n_523), .C2(n_526), .Y(n_795) );
OAI22x1_ASAP7_75t_L g676 ( .A1(n_318), .A2(n_677), .B1(n_698), .B2(n_699), .Y(n_676) );
INVx1_ASAP7_75t_L g699 ( .A(n_318), .Y(n_699) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_319), .Y(n_521) );
CKINVDCx20_ASAP7_75t_R g1024 ( .A(n_322), .Y(n_1024) );
CKINVDCx20_ASAP7_75t_R g625 ( .A(n_328), .Y(n_625) );
AOI22xp5_ASAP7_75t_L g723 ( .A1(n_334), .A2(n_361), .B1(n_530), .B2(n_609), .Y(n_723) );
XNOR2x1_ASAP7_75t_L g657 ( .A(n_337), .B(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_340), .B(n_759), .Y(n_817) );
CKINVDCx20_ASAP7_75t_R g411 ( .A(n_341), .Y(n_411) );
INVx1_ASAP7_75t_L g390 ( .A(n_349), .Y(n_390) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_350), .A2(n_375), .B1(n_612), .B2(n_613), .Y(n_611) );
INVx1_ASAP7_75t_L g993 ( .A(n_359), .Y(n_993) );
AND2x4_ASAP7_75t_L g1008 ( .A(n_359), .B(n_994), .Y(n_1008) );
AO21x1_ASAP7_75t_L g1039 ( .A1(n_359), .A2(n_1004), .B(n_1040), .Y(n_1039) );
INVx1_ASAP7_75t_L g994 ( .A(n_362), .Y(n_994) );
AND2x2_ASAP7_75t_R g1036 ( .A(n_362), .B(n_993), .Y(n_1036) );
INVxp67_ASAP7_75t_L g1005 ( .A(n_370), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g971 ( .A(n_371), .B(n_395), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_373), .B(n_605), .Y(n_667) );
CKINVDCx20_ASAP7_75t_R g1021 ( .A(n_374), .Y(n_1021) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_776), .B(n_989), .C(n_1000), .Y(n_382) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_383), .A2(n_776), .B(n_990), .Y(n_989) );
XNOR2x1_ASAP7_75t_L g383 ( .A(n_384), .B(n_630), .Y(n_383) );
OAI21x1_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_508), .B(n_629), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_385), .B(n_510), .Y(n_629) );
AO22x1_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_387), .B1(n_469), .B2(n_507), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_389), .Y(n_388) );
XNOR2x1_ASAP7_75t_L g389 ( .A(n_390), .B(n_391), .Y(n_389) );
NAND2x1_ASAP7_75t_L g391 ( .A(n_392), .B(n_441), .Y(n_391) );
NOR2xp67_ASAP7_75t_L g392 ( .A(n_393), .B(n_422), .Y(n_392) );
OAI21xp5_ASAP7_75t_SL g393 ( .A1(n_394), .A2(n_411), .B(n_412), .Y(n_393) );
OAI222xp33_ASAP7_75t_L g938 ( .A1(n_394), .A2(n_414), .B1(n_939), .B2(n_940), .C1(n_941), .C2(n_942), .Y(n_938) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AND2x4_ASAP7_75t_L g395 ( .A(n_396), .B(n_404), .Y(n_395) );
AND2x4_ASAP7_75t_L g429 ( .A(n_396), .B(n_430), .Y(n_429) );
AND2x4_ASAP7_75t_L g439 ( .A(n_396), .B(n_440), .Y(n_439) );
AND2x2_ASAP7_75t_L g477 ( .A(n_396), .B(n_404), .Y(n_477) );
AND2x2_ASAP7_75t_L g579 ( .A(n_396), .B(n_430), .Y(n_579) );
AND2x2_ASAP7_75t_L g582 ( .A(n_396), .B(n_440), .Y(n_582) );
AND2x2_ASAP7_75t_L g923 ( .A(n_396), .B(n_430), .Y(n_923) );
AND2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_402), .Y(n_396) );
AND2x2_ASAP7_75t_L g417 ( .A(n_397), .B(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
INVx2_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
OAI22x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B1(n_400), .B2(n_401), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g403 ( .A(n_399), .Y(n_403) );
INVx2_ASAP7_75t_L g407 ( .A(n_399), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_399), .Y(n_410) );
INVx2_ASAP7_75t_L g418 ( .A(n_402), .Y(n_418) );
AND2x2_ASAP7_75t_L g435 ( .A(n_402), .B(n_436), .Y(n_435) );
BUFx2_ASAP7_75t_L g448 ( .A(n_402), .Y(n_448) );
AND2x4_ASAP7_75t_L g451 ( .A(n_404), .B(n_417), .Y(n_451) );
AND2x2_ASAP7_75t_L g459 ( .A(n_404), .B(n_435), .Y(n_459) );
AND2x4_ASAP7_75t_L g466 ( .A(n_404), .B(n_454), .Y(n_466) );
AND2x2_ASAP7_75t_L g591 ( .A(n_404), .B(n_417), .Y(n_591) );
AND2x6_ASAP7_75t_L g594 ( .A(n_404), .B(n_435), .Y(n_594) );
AND2x2_ASAP7_75t_L g624 ( .A(n_404), .B(n_417), .Y(n_624) );
AND2x2_ASAP7_75t_L g650 ( .A(n_404), .B(n_454), .Y(n_650) );
AND2x4_ASAP7_75t_L g404 ( .A(n_405), .B(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AND2x4_ASAP7_75t_L g416 ( .A(n_406), .B(n_408), .Y(n_416) );
AND2x2_ASAP7_75t_L g421 ( .A(n_406), .B(n_409), .Y(n_421) );
INVx1_ASAP7_75t_L g427 ( .A(n_406), .Y(n_427) );
INVxp67_ASAP7_75t_L g440 ( .A(n_408), .Y(n_440) );
INVx2_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
AND2x2_ASAP7_75t_L g426 ( .A(n_409), .B(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
AND2x4_ASAP7_75t_L g434 ( .A(n_416), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g453 ( .A(n_416), .B(n_454), .Y(n_453) );
AND2x2_ASAP7_75t_L g483 ( .A(n_416), .B(n_417), .Y(n_483) );
AND2x2_ASAP7_75t_L g581 ( .A(n_416), .B(n_435), .Y(n_581) );
AND2x2_ASAP7_75t_L g644 ( .A(n_416), .B(n_435), .Y(n_644) );
AND2x2_ASAP7_75t_L g653 ( .A(n_416), .B(n_454), .Y(n_653) );
AND2x2_ASAP7_75t_L g425 ( .A(n_417), .B(n_426), .Y(n_425) );
AND2x4_ASAP7_75t_L g643 ( .A(n_417), .B(n_426), .Y(n_643) );
AND2x4_ASAP7_75t_L g454 ( .A(n_418), .B(n_436), .Y(n_454) );
INVxp67_ASAP7_75t_L g942 ( .A(n_419), .Y(n_942) );
AND2x2_ASAP7_75t_SL g419 ( .A(n_420), .B(n_421), .Y(n_419) );
AND2x2_ASAP7_75t_L g486 ( .A(n_420), .B(n_421), .Y(n_486) );
AND2x2_ASAP7_75t_SL g919 ( .A(n_420), .B(n_421), .Y(n_919) );
AND2x4_ASAP7_75t_L g447 ( .A(n_421), .B(n_448), .Y(n_447) );
AND2x4_ASAP7_75t_L g468 ( .A(n_421), .B(n_454), .Y(n_468) );
AND2x4_ASAP7_75t_L g587 ( .A(n_421), .B(n_448), .Y(n_587) );
AND2x4_ASAP7_75t_L g592 ( .A(n_421), .B(n_454), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_432), .Y(n_422) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_424), .Y(n_488) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx3_ASAP7_75t_L g532 ( .A(n_425), .Y(n_532) );
BUFx6f_ASAP7_75t_L g608 ( .A(n_425), .Y(n_608) );
AND2x2_ASAP7_75t_L g445 ( .A(n_426), .B(n_435), .Y(n_445) );
AND2x4_ASAP7_75t_L g462 ( .A(n_426), .B(n_454), .Y(n_462) );
AND2x2_ASAP7_75t_SL g586 ( .A(n_426), .B(n_435), .Y(n_586) );
AND2x6_ASAP7_75t_L g595 ( .A(n_426), .B(n_454), .Y(n_595) );
AND2x2_ASAP7_75t_L g979 ( .A(n_426), .B(n_435), .Y(n_979) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_427), .Y(n_431) );
BUFx2_ASAP7_75t_SL g489 ( .A(n_428), .Y(n_489) );
BUFx6f_ASAP7_75t_SL g428 ( .A(n_429), .Y(n_428) );
BUFx3_ASAP7_75t_L g534 ( .A(n_429), .Y(n_534) );
INVx2_ASAP7_75t_L g610 ( .A(n_429), .Y(n_610) );
BUFx4f_ASAP7_75t_L g686 ( .A(n_429), .Y(n_686) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx6f_ASAP7_75t_L g537 ( .A(n_434), .Y(n_537) );
BUFx3_ASAP7_75t_L g612 ( .A(n_434), .Y(n_612) );
BUFx2_ASAP7_75t_L g815 ( .A(n_434), .Y(n_815) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g479 ( .A(n_438), .Y(n_479) );
INVx2_ASAP7_75t_L g538 ( .A(n_438), .Y(n_538) );
INVx2_ASAP7_75t_L g613 ( .A(n_438), .Y(n_613) );
INVx2_ASAP7_75t_SL g682 ( .A(n_438), .Y(n_682) );
INVx2_ASAP7_75t_L g784 ( .A(n_438), .Y(n_784) );
INVx2_ASAP7_75t_SL g830 ( .A(n_438), .Y(n_830) );
OAI22xp5_ASAP7_75t_L g1023 ( .A1(n_438), .A2(n_1024), .B1(n_1025), .B2(n_1026), .Y(n_1023) );
INVx6_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g441 ( .A(n_442), .B(n_455), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_443), .B(n_449), .Y(n_442) );
BUFx6f_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
BUFx3_ASAP7_75t_L g497 ( .A(n_445), .Y(n_497) );
INVx2_ASAP7_75t_L g564 ( .A(n_445), .Y(n_564) );
BUFx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx5_ASAP7_75t_SL g499 ( .A(n_447), .Y(n_499) );
BUFx2_ASAP7_75t_L g749 ( .A(n_447), .Y(n_749) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx6_ASAP7_75t_L g542 ( .A(n_451), .Y(n_542) );
INVx2_ASAP7_75t_L g502 ( .A(n_452), .Y(n_502) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_452), .Y(n_789) );
BUFx6f_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_453), .Y(n_622) );
BUFx3_ASAP7_75t_L g690 ( .A(n_453), .Y(n_690) );
INVx2_ASAP7_75t_L g841 ( .A(n_453), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_463), .Y(n_455) );
INVx3_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx2_ASAP7_75t_L g554 ( .A(n_458), .Y(n_554) );
INVx2_ASAP7_75t_SL g689 ( .A(n_458), .Y(n_689) );
INVx2_ASAP7_75t_L g741 ( .A(n_458), .Y(n_741) );
INVx2_ASAP7_75t_SL g771 ( .A(n_458), .Y(n_771) );
INVx3_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
BUFx2_ASAP7_75t_L g876 ( .A(n_459), .Y(n_876) );
INVx2_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g494 ( .A(n_461), .Y(n_494) );
INVx2_ASAP7_75t_L g557 ( .A(n_461), .Y(n_557) );
INVx2_ASAP7_75t_SL g617 ( .A(n_461), .Y(n_617) );
INVx2_ASAP7_75t_SL g716 ( .A(n_461), .Y(n_716) );
INVx1_ASAP7_75t_SL g806 ( .A(n_461), .Y(n_806) );
INVx2_ASAP7_75t_L g877 ( .A(n_461), .Y(n_877) );
INVx8_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx3_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_SL g493 ( .A(n_465), .Y(n_493) );
INVx2_ASAP7_75t_L g621 ( .A(n_465), .Y(n_621) );
INVx4_ASAP7_75t_L g697 ( .A(n_465), .Y(n_697) );
INVx2_ASAP7_75t_SL g708 ( .A(n_465), .Y(n_708) );
INVx8_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
BUFx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g505 ( .A(n_468), .Y(n_505) );
BUFx2_ASAP7_75t_SL g549 ( .A(n_468), .Y(n_549) );
BUFx2_ASAP7_75t_SL g694 ( .A(n_468), .Y(n_694) );
BUFx3_ASAP7_75t_L g838 ( .A(n_468), .Y(n_838) );
INVx1_ASAP7_75t_L g507 ( .A(n_469), .Y(n_507) );
INVx1_ASAP7_75t_L g506 ( .A(n_471), .Y(n_506) );
OR2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_490), .Y(n_471) );
NAND4xp25_ASAP7_75t_SL g472 ( .A(n_473), .B(n_478), .C(n_480), .D(n_487), .Y(n_472) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx3_ASAP7_75t_SL g520 ( .A(n_476), .Y(n_520) );
INVx4_ASAP7_75t_SL g574 ( .A(n_476), .Y(n_574) );
INVx3_ASAP7_75t_L g605 ( .A(n_476), .Y(n_605) );
INVx4_ASAP7_75t_SL g759 ( .A(n_476), .Y(n_759) );
INVx6_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx6f_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx3_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g527 ( .A(n_483), .Y(n_527) );
INVx2_ASAP7_75t_L g603 ( .A(n_483), .Y(n_603) );
BUFx5_ASAP7_75t_L g684 ( .A(n_483), .Y(n_684) );
BUFx3_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
BUFx12f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g525 ( .A(n_486), .Y(n_525) );
NAND4xp25_ASAP7_75t_L g490 ( .A(n_491), .B(n_495), .C(n_500), .D(n_503), .Y(n_490) );
INVx1_ASAP7_75t_L g546 ( .A(n_492), .Y(n_546) );
BUFx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
BUFx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
OAI22xp33_ASAP7_75t_SL g559 ( .A1(n_499), .A2(n_560), .B1(n_565), .B2(n_566), .Y(n_559) );
INVx3_ASAP7_75t_L g769 ( .A(n_499), .Y(n_769) );
INVx2_ASAP7_75t_L g897 ( .A(n_499), .Y(n_897) );
INVx2_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_502), .A2(n_541), .B1(n_542), .B2(n_543), .Y(n_540) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
INVx2_ASAP7_75t_SL g810 ( .A(n_505), .Y(n_810) );
INVx2_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
OAI22x1_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_567), .B1(n_568), .B2(n_628), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVx1_ASAP7_75t_L g628 ( .A(n_512), .Y(n_628) );
INVx1_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
AND3x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_539), .C(n_550), .Y(n_515) );
NOR2xp67_ASAP7_75t_SL g516 ( .A(n_517), .B(n_528), .Y(n_516) );
OAI21xp5_ASAP7_75t_SL g517 ( .A1(n_518), .A2(n_521), .B(n_522), .Y(n_517) );
OAI21xp33_ASAP7_75t_L g903 ( .A1(n_518), .A2(n_904), .B(n_905), .Y(n_903) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g720 ( .A(n_520), .Y(n_720) );
BUFx6f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx3_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx2_ASAP7_75t_L g813 ( .A(n_525), .Y(n_813) );
INVx2_ASAP7_75t_L g823 ( .A(n_525), .Y(n_823) );
BUFx6f_ASAP7_75t_SL g526 ( .A(n_527), .Y(n_526) );
NAND2xp5_ASAP7_75t_SL g528 ( .A(n_529), .B(n_535), .Y(n_528) );
BUFx3_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx4_ASAP7_75t_L g578 ( .A(n_532), .Y(n_578) );
INVx2_ASAP7_75t_L g825 ( .A(n_532), .Y(n_825) );
BUFx6f_ASAP7_75t_SL g533 ( .A(n_534), .Y(n_533) );
BUFx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
BUFx4f_ASAP7_75t_SL g681 ( .A(n_537), .Y(n_681) );
BUFx2_ASAP7_75t_L g722 ( .A(n_537), .Y(n_722) );
INVx1_ASAP7_75t_L g1025 ( .A(n_537), .Y(n_1025) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_540), .B(n_544), .Y(n_539) );
INVx2_ASAP7_75t_L g693 ( .A(n_542), .Y(n_693) );
INVx3_ASAP7_75t_L g746 ( .A(n_542), .Y(n_746) );
INVx2_ASAP7_75t_L g794 ( .A(n_542), .Y(n_794) );
INVx2_ASAP7_75t_L g837 ( .A(n_542), .Y(n_837) );
OAI22xp33_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_546), .B1(n_547), .B2(n_548), .Y(n_544) );
INVx1_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
NOR2xp33_ASAP7_75t_L g550 ( .A(n_551), .B(n_559), .Y(n_550) );
OAI22xp33_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_555), .B1(n_556), .B2(n_558), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
BUFx2_ASAP7_75t_L g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g768 ( .A(n_562), .Y(n_768) );
INVx1_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_563), .Y(n_748) );
INVx1_ASAP7_75t_L g896 ( .A(n_563), .Y(n_896) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g714 ( .A(n_564), .Y(n_714) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AO22x2_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_597), .B1(n_626), .B2(n_627), .Y(n_568) );
INVx1_ASAP7_75t_SL g627 ( .A(n_569), .Y(n_627) );
INVx1_ASAP7_75t_L g672 ( .A(n_569), .Y(n_672) );
XOR2x2_ASAP7_75t_L g569 ( .A(n_570), .B(n_596), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g570 ( .A(n_571), .B(n_583), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_576), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_580), .Y(n_576) );
INVx2_ASAP7_75t_SL g1020 ( .A(n_578), .Y(n_1020) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_588), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_593), .Y(n_589) );
INVx1_ASAP7_75t_L g663 ( .A(n_594), .Y(n_663) );
INVx2_ASAP7_75t_L g626 ( .A(n_597), .Y(n_626) );
XOR2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_625), .Y(n_597) );
NAND2x1p5_ASAP7_75t_L g598 ( .A(n_599), .B(n_614), .Y(n_598) );
NOR2x1_ASAP7_75t_L g599 ( .A(n_600), .B(n_606), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_601), .B(n_604), .Y(n_600) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
INVx1_ASAP7_75t_L g860 ( .A(n_603), .Y(n_860) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_607), .B(n_611), .Y(n_606) );
INVx2_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g1049 ( .A(n_610), .Y(n_1049) );
NOR2x1_ASAP7_75t_L g614 ( .A(n_615), .B(n_619), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_616), .B(n_618), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_620), .B(n_623), .Y(n_619) );
INVx1_ASAP7_75t_L g744 ( .A(n_622), .Y(n_744) );
XOR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_726), .Y(n_630) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B1(n_671), .B2(n_725), .Y(n_631) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
OA22x2_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_636), .B1(n_656), .B2(n_657), .Y(n_634) );
AO22x2_ASAP7_75t_L g730 ( .A1(n_635), .A2(n_731), .B1(n_732), .B2(n_750), .Y(n_730) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
BUFx2_ASAP7_75t_L g750 ( .A(n_636), .Y(n_750) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g638 ( .A(n_639), .B(n_646), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_645), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_647), .B(n_651), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
NOR2x1_ASAP7_75t_L g658 ( .A(n_659), .B(n_666), .Y(n_658) );
NAND4xp25_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .C(n_664), .D(n_665), .Y(n_659) );
INVx1_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
NAND4xp25_ASAP7_75t_SL g666 ( .A(n_667), .B(n_668), .C(n_669), .D(n_670), .Y(n_666) );
INVx1_ASAP7_75t_L g725 ( .A(n_671), .Y(n_725) );
XNOR2xp5_ASAP7_75t_L g671 ( .A(n_672), .B(n_673), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g673 ( .A1(n_674), .A2(n_675), .B1(n_700), .B2(n_701), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g698 ( .A(n_677), .Y(n_698) );
OR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_687), .Y(n_677) );
NAND4xp25_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .C(n_683), .D(n_685), .Y(n_678) );
INVxp67_ASAP7_75t_L g1022 ( .A(n_686), .Y(n_1022) );
NAND4xp25_ASAP7_75t_L g687 ( .A(n_688), .B(n_691), .C(n_692), .D(n_695), .Y(n_687) );
BUFx2_ASAP7_75t_L g709 ( .A(n_690), .Y(n_709) );
BUFx6f_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g788 ( .A(n_697), .Y(n_788) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NOR3x1_ASAP7_75t_SL g704 ( .A(n_705), .B(n_711), .C(n_717), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_706), .B(n_710), .Y(n_705) );
BUFx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_712), .B(n_715), .Y(n_711) );
BUFx6f_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
NAND4xp25_ASAP7_75t_SL g717 ( .A(n_718), .B(n_721), .C(n_723), .D(n_724), .Y(n_717) );
INVx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI22xp5_ASAP7_75t_SL g728 ( .A1(n_729), .A2(n_730), .B1(n_751), .B2(n_775), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp67_ASAP7_75t_L g733 ( .A(n_734), .B(n_739), .Y(n_733) );
NAND4xp25_ASAP7_75t_SL g734 ( .A(n_735), .B(n_736), .C(n_737), .D(n_738), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .C(n_745), .D(n_747), .Y(n_739) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g775 ( .A(n_753), .Y(n_775) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
AND2x4_ASAP7_75t_L g755 ( .A(n_756), .B(n_765), .Y(n_755) );
NOR2xp67_ASAP7_75t_L g756 ( .A(n_757), .B(n_762), .Y(n_756) );
OAI21xp5_ASAP7_75t_SL g757 ( .A1(n_758), .A2(n_760), .B(n_761), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NOR2x1_ASAP7_75t_L g765 ( .A(n_766), .B(n_772), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g766 ( .A(n_767), .B(n_770), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_773), .B(n_774), .Y(n_772) );
OAI22xp5_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_864), .B1(n_865), .B2(n_988), .Y(n_776) );
INVx1_ASAP7_75t_L g988 ( .A(n_777), .Y(n_988) );
AOI22xp33_ASAP7_75t_SL g777 ( .A1(n_778), .A2(n_797), .B1(n_862), .B2(n_863), .Y(n_777) );
INVx2_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
HB1xp67_ASAP7_75t_L g862 ( .A(n_779), .Y(n_862) );
XNOR2x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_796), .Y(n_779) );
NAND4xp75_ASAP7_75t_L g780 ( .A(n_781), .B(n_785), .C(n_791), .D(n_795), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_782), .B(n_783), .Y(n_781) );
AND2x2_ASAP7_75t_L g785 ( .A(n_786), .B(n_790), .Y(n_785) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
AND2x2_ASAP7_75t_L g791 ( .A(n_792), .B(n_793), .Y(n_791) );
INVx2_ASAP7_75t_SL g863 ( .A(n_797), .Y(n_863) );
OA22x2_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_799), .B1(n_847), .B2(n_848), .Y(n_797) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
AOI22xp5_ASAP7_75t_L g799 ( .A1(n_800), .A2(n_818), .B1(n_845), .B2(n_846), .Y(n_799) );
INVx1_ASAP7_75t_L g845 ( .A(n_800), .Y(n_845) );
INVx1_ASAP7_75t_L g802 ( .A(n_803), .Y(n_802) );
NOR2x1_ASAP7_75t_L g803 ( .A(n_804), .B(n_811), .Y(n_803) );
NAND4xp25_ASAP7_75t_L g804 ( .A(n_805), .B(n_807), .C(n_808), .D(n_809), .Y(n_804) );
NAND4xp25_ASAP7_75t_L g811 ( .A(n_812), .B(n_814), .C(n_816), .D(n_817), .Y(n_811) );
INVx2_ASAP7_75t_L g846 ( .A(n_818), .Y(n_846) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_831), .Y(n_819) );
NOR3xp33_ASAP7_75t_L g820 ( .A(n_821), .B(n_826), .C(n_828), .Y(n_820) );
NOR4xp25_ASAP7_75t_L g843 ( .A(n_821), .B(n_832), .C(n_835), .D(n_844), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .Y(n_821) );
INVxp67_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_827), .B(n_829), .Y(n_844) );
INVxp67_ASAP7_75t_SL g828 ( .A(n_829), .Y(n_828) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_832), .B(n_835), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_833), .B(n_834), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g835 ( .A(n_836), .B(n_839), .Y(n_835) );
INVx2_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx1_ASAP7_75t_L g900 ( .A(n_841), .Y(n_900) );
INVx3_ASAP7_75t_L g847 ( .A(n_848), .Y(n_847) );
XOR2x2_ASAP7_75t_L g848 ( .A(n_849), .B(n_861), .Y(n_848) );
NAND4xp75_ASAP7_75t_L g849 ( .A(n_850), .B(n_853), .C(n_856), .D(n_859), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
AND2x2_ASAP7_75t_L g853 ( .A(n_854), .B(n_855), .Y(n_853) );
AND2x2_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
XNOR2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_911), .Y(n_865) );
AO22x1_ASAP7_75t_L g866 ( .A1(n_867), .A2(n_868), .B1(n_886), .B2(n_910), .Y(n_866) );
INVx2_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
INVx1_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
NOR2xp33_ASAP7_75t_L g871 ( .A(n_872), .B(n_880), .Y(n_871) );
NAND4xp25_ASAP7_75t_SL g872 ( .A(n_873), .B(n_874), .C(n_878), .D(n_879), .Y(n_872) );
BUFx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND4xp25_ASAP7_75t_SL g880 ( .A(n_881), .B(n_882), .C(n_883), .D(n_884), .Y(n_880) );
INVx2_ASAP7_75t_L g910 ( .A(n_886), .Y(n_910) );
BUFx3_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVxp33_ASAP7_75t_SL g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_SL g909 ( .A(n_890), .Y(n_909) );
AND2x2_ASAP7_75t_L g890 ( .A(n_891), .B(n_902), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_898), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
INVx1_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_899), .B(n_901), .Y(n_898) );
NOR2xp33_ASAP7_75t_L g902 ( .A(n_903), .B(n_906), .Y(n_902) );
NAND2xp5_ASAP7_75t_L g906 ( .A(n_907), .B(n_908), .Y(n_906) );
OAI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_931), .B1(n_986), .B2(n_987), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
HB1xp67_ASAP7_75t_L g986 ( .A(n_913), .Y(n_986) );
INVx2_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
XNOR2x1_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
AND2x2_ASAP7_75t_L g916 ( .A(n_917), .B(n_924), .Y(n_916) );
NOR2xp33_ASAP7_75t_L g917 ( .A(n_918), .B(n_920), .Y(n_917) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_921), .B(n_922), .Y(n_920) );
NOR2xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_928), .Y(n_924) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_929), .B(n_930), .Y(n_928) );
INVx1_ASAP7_75t_L g987 ( .A(n_931), .Y(n_987) );
OAI22x1_ASAP7_75t_SL g931 ( .A1(n_932), .A2(n_933), .B1(n_953), .B2(n_985), .Y(n_931) );
INVx2_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
HB1xp67_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
NAND2x1p5_ASAP7_75t_L g936 ( .A(n_937), .B(n_946), .Y(n_936) );
NOR2x1_ASAP7_75t_L g937 ( .A(n_938), .B(n_943), .Y(n_937) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_945), .Y(n_943) );
NOR2x1_ASAP7_75t_L g946 ( .A(n_947), .B(n_950), .Y(n_946) );
NAND2xp5_ASAP7_75t_L g947 ( .A(n_948), .B(n_949), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g950 ( .A(n_951), .B(n_952), .Y(n_950) );
INVx2_ASAP7_75t_L g985 ( .A(n_953), .Y(n_985) );
XNOR2x1_ASAP7_75t_L g953 ( .A(n_954), .B(n_967), .Y(n_953) );
INVx1_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
NOR2x1_ASAP7_75t_L g957 ( .A(n_958), .B(n_962), .Y(n_957) );
NAND3xp33_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .C(n_961), .Y(n_958) );
NAND4xp25_ASAP7_75t_L g962 ( .A(n_963), .B(n_964), .C(n_965), .D(n_966), .Y(n_962) );
XOR2x2_ASAP7_75t_L g967 ( .A(n_968), .B(n_984), .Y(n_967) );
NAND2x1p5_ASAP7_75t_L g968 ( .A(n_969), .B(n_976), .Y(n_968) );
NOR2x1_ASAP7_75t_L g969 ( .A(n_970), .B(n_973), .Y(n_969) );
NAND2xp5_ASAP7_75t_L g970 ( .A(n_971), .B(n_972), .Y(n_970) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_974), .B(n_975), .Y(n_973) );
NOR2x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_981), .Y(n_976) );
NAND2xp5_ASAP7_75t_L g977 ( .A(n_978), .B(n_980), .Y(n_977) );
NAND2xp5_ASAP7_75t_L g981 ( .A(n_982), .B(n_983), .Y(n_981) );
INVx2_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
AND2x2_ASAP7_75t_L g991 ( .A(n_992), .B(n_995), .Y(n_991) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_992), .B(n_996), .Y(n_1061) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_993), .B(n_994), .Y(n_992) );
INVx1_ASAP7_75t_L g1040 ( .A(n_994), .Y(n_1040) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
CKINVDCx20_ASAP7_75t_R g1001 ( .A(n_1002), .Y(n_1001) );
OR2x2_ASAP7_75t_L g1002 ( .A(n_1003), .B(n_1007), .Y(n_1002) );
INVx1_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NOR2xp33_ASAP7_75t_L g1004 ( .A(n_1005), .B(n_1006), .Y(n_1004) );
INVxp67_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OAI222xp33_ASAP7_75t_L g1009 ( .A1(n_1010), .A2(n_1035), .B1(n_1037), .B2(n_1041), .C1(n_1042), .C2(n_1059), .Y(n_1009) );
CKINVDCx16_ASAP7_75t_R g1011 ( .A(n_1012), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
NAND2xp5_ASAP7_75t_L g1013 ( .A(n_1014), .B(n_1027), .Y(n_1013) );
NOR3xp33_ASAP7_75t_L g1014 ( .A(n_1015), .B(n_1018), .C(n_1023), .Y(n_1014) );
NAND2xp5_ASAP7_75t_SL g1015 ( .A(n_1016), .B(n_1017), .Y(n_1015) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_1019), .A2(n_1020), .B1(n_1021), .B2(n_1022), .Y(n_1018) );
NOR2xp33_ASAP7_75t_L g1027 ( .A(n_1028), .B(n_1031), .Y(n_1027) );
NAND2xp5_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
NAND2xp5_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
INVx1_ASAP7_75t_SL g1035 ( .A(n_1036), .Y(n_1035) );
CKINVDCx20_ASAP7_75t_R g1037 ( .A(n_1038), .Y(n_1037) );
CKINVDCx20_ASAP7_75t_R g1038 ( .A(n_1039), .Y(n_1038) );
BUFx2_ASAP7_75t_L g1042 ( .A(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_SL g1043 ( .A(n_1044), .Y(n_1043) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1045), .Y(n_1058) );
NAND4xp75_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1051), .C(n_1054), .D(n_1057), .Y(n_1045) );
AND2x2_ASAP7_75t_L g1046 ( .A(n_1047), .B(n_1050), .Y(n_1046) );
INVx3_ASAP7_75t_L g1048 ( .A(n_1049), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1051 ( .A(n_1052), .B(n_1053), .Y(n_1051) );
AND2x2_ASAP7_75t_L g1054 ( .A(n_1055), .B(n_1056), .Y(n_1054) );
INVx1_ASAP7_75t_SL g1059 ( .A(n_1060), .Y(n_1059) );
CKINVDCx6p67_ASAP7_75t_R g1060 ( .A(n_1061), .Y(n_1060) );
endmodule