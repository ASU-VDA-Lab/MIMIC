module fake_ariane_2367_n_790 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_790);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_790;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_616;
wire n_617;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

OR2x2_ASAP7_75t_L g162 ( 
.A(n_148),
.B(n_24),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_62),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_153),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_11),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_8),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_113),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_45),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_96),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_140),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_66),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_26),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_122),
.Y(n_176)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_111),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_141),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_27),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_33),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_59),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_151),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_81),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_52),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_121),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_29),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_38),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_134),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g189 ( 
.A(n_150),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_76),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_152),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_16),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_3),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_131),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_42),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_31),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_60),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_104),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_112),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_71),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_130),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_54),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_44),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_124),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_123),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_4),
.Y(n_208)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_135),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_103),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_48),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_19),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_32),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_102),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_154),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_127),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_72),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_146),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_93),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_170),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_165),
.B(n_0),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_180),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_180),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx4_ASAP7_75t_L g225 ( 
.A(n_170),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

AND2x6_ASAP7_75t_L g227 ( 
.A(n_177),
.B(n_18),
.Y(n_227)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_202),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_202),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_165),
.Y(n_230)
);

BUFx12f_ASAP7_75t_L g231 ( 
.A(n_169),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_189),
.Y(n_232)
);

AND2x4_ASAP7_75t_L g233 ( 
.A(n_189),
.B(n_0),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_161),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_163),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_177),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_209),
.B(n_1),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_167),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_184),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_194),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_210),
.Y(n_243)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_172),
.Y(n_244)
);

AND2x2_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_202),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_217),
.B(n_5),
.Y(n_246)
);

OA21x2_ASAP7_75t_L g247 ( 
.A1(n_175),
.A2(n_6),
.B(n_7),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_212),
.Y(n_248)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_212),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_178),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_185),
.B(n_6),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_197),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_20),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_200),
.Y(n_255)
);

AND2x4_ASAP7_75t_L g256 ( 
.A(n_204),
.B(n_7),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_214),
.Y(n_257)
);

INVx5_ASAP7_75t_L g258 ( 
.A(n_162),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_8),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_218),
.Y(n_260)
);

INVx4_ASAP7_75t_L g261 ( 
.A(n_164),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_166),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_220),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_243),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_260),
.Y(n_267)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_220),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_225),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_181),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_205),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g272 ( 
.A(n_230),
.B(n_193),
.Y(n_272)
);

BUFx6f_ASAP7_75t_SL g273 ( 
.A(n_233),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_208),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_220),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_260),
.Y(n_277)
);

INVx8_ASAP7_75t_L g278 ( 
.A(n_258),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_224),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_243),
.B(n_168),
.Y(n_280)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_224),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_238),
.B(n_171),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_224),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_224),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_226),
.Y(n_285)
);

OR2x2_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_9),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_226),
.Y(n_287)
);

BUFx6f_ASAP7_75t_SL g288 ( 
.A(n_233),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_238),
.B(n_173),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_231),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_226),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_191),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_255),
.B(n_174),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_260),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_260),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_229),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_233),
.B(n_176),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_261),
.B(n_179),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_229),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_229),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_242),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_242),
.Y(n_304)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_221),
.Y(n_305)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_225),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_222),
.Y(n_307)
);

NAND2xp33_ASAP7_75t_SL g308 ( 
.A(n_246),
.B(n_182),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_235),
.A2(n_216),
.B1(n_215),
.B2(n_213),
.Y(n_309)
);

AND2x6_ASAP7_75t_L g310 ( 
.A(n_246),
.B(n_21),
.Y(n_310)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_225),
.Y(n_311)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_228),
.Y(n_312)
);

INVx3_ASAP7_75t_L g313 ( 
.A(n_228),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_242),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_183),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_270),
.B(n_258),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_305),
.B(n_256),
.Y(n_317)
);

INVxp33_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_293),
.Y(n_320)
);

NOR3xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_251),
.C(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_271),
.B(n_258),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_269),
.B(n_258),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_267),
.Y(n_324)
);

AOI221xp5_ASAP7_75t_L g325 ( 
.A1(n_305),
.A2(n_246),
.B1(n_259),
.B2(n_256),
.C(n_221),
.Y(n_325)
);

NAND2x1p5_ASAP7_75t_L g326 ( 
.A(n_265),
.B(n_237),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g327 ( 
.A(n_279),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_269),
.B(n_245),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_266),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_231),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_294),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_269),
.B(n_306),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_L g333 ( 
.A(n_310),
.B(n_227),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_274),
.B(n_236),
.Y(n_334)
);

NOR3xp33_ASAP7_75t_L g335 ( 
.A(n_308),
.B(n_259),
.C(n_256),
.Y(n_335)
);

BUFx6f_ASAP7_75t_SL g336 ( 
.A(n_310),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_286),
.B(n_236),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_274),
.B(n_262),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_277),
.Y(n_339)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_296),
.Y(n_340)
);

NAND2xp33_ASAP7_75t_L g341 ( 
.A(n_310),
.B(n_227),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_306),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_306),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_311),
.B(n_245),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_279),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_311),
.B(n_259),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_311),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_222),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_223),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_312),
.B(n_223),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_300),
.B(n_232),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_313),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_313),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_313),
.B(n_232),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_294),
.B(n_239),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_228),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_272),
.B(n_239),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_291),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_272),
.B(n_244),
.Y(n_359)
);

BUFx5_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_299),
.B(n_237),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_282),
.B(n_244),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_290),
.B(n_237),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g364 ( 
.A(n_286),
.B(n_280),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

NOR2xp67_ASAP7_75t_L g366 ( 
.A(n_264),
.B(n_249),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_310),
.B(n_257),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_310),
.B(n_257),
.Y(n_369)
);

AND2x4_ASAP7_75t_L g370 ( 
.A(n_309),
.B(n_241),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_278),
.B(n_257),
.Y(n_371)
);

NAND2xp33_ASAP7_75t_L g372 ( 
.A(n_278),
.B(n_227),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_273),
.B(n_186),
.Y(n_373)
);

NOR2x1_ASAP7_75t_L g374 ( 
.A(n_268),
.B(n_257),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_273),
.B(n_188),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_278),
.B(n_268),
.Y(n_376)
);

NAND2xp33_ASAP7_75t_L g377 ( 
.A(n_278),
.B(n_227),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_273),
.B(n_288),
.Y(n_378)
);

BUFx5_ASAP7_75t_L g379 ( 
.A(n_288),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_275),
.B(n_249),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_275),
.B(n_276),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_276),
.B(n_249),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_332),
.A2(n_356),
.B(n_346),
.Y(n_383)
);

O2A1O1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_325),
.A2(n_247),
.B(n_304),
.C(n_303),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_351),
.B(n_190),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g386 ( 
.A1(n_317),
.A2(n_288),
.B1(n_247),
.B2(n_196),
.Y(n_386)
);

A2O1A1Ixp33_ASAP7_75t_L g387 ( 
.A1(n_335),
.A2(n_314),
.B(n_304),
.C(n_303),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_362),
.B(n_192),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_338),
.B(n_195),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_334),
.B(n_198),
.Y(n_390)
);

NAND2x1p5_ASAP7_75t_L g391 ( 
.A(n_334),
.B(n_247),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_323),
.A2(n_314),
.B(n_302),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_333),
.A2(n_227),
.B(n_254),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_331),
.A2(n_199),
.B1(n_201),
.B2(n_203),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g395 ( 
.A1(n_364),
.A2(n_206),
.B1(n_207),
.B2(n_298),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_321),
.A2(n_254),
.B1(n_301),
.B2(n_298),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_L g398 ( 
.A1(n_341),
.A2(n_302),
.B(n_301),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_328),
.B(n_281),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_344),
.A2(n_295),
.B(n_292),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_360),
.B(n_279),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_342),
.Y(n_402)
);

AO21x1_ASAP7_75t_L g403 ( 
.A1(n_367),
.A2(n_295),
.B(n_292),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_343),
.A2(n_287),
.B(n_285),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_347),
.A2(n_287),
.B(n_285),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_318),
.B(n_9),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_10),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_329),
.B(n_281),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_369),
.A2(n_353),
.B(n_352),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_355),
.B(n_283),
.Y(n_410)
);

A2O1A1Ixp33_ASAP7_75t_L g411 ( 
.A1(n_378),
.A2(n_284),
.B(n_283),
.C(n_289),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_357),
.B(n_284),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_319),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_359),
.B(n_254),
.Y(n_414)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_348),
.A2(n_254),
.B(n_249),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_337),
.B(n_254),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g417 ( 
.A(n_360),
.B(n_279),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_349),
.A2(n_249),
.B(n_279),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_360),
.B(n_289),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_336),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_316),
.B(n_242),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

AOI21x1_ASAP7_75t_L g423 ( 
.A1(n_380),
.A2(n_289),
.B(n_252),
.Y(n_423)
);

NAND2x1p5_ASAP7_75t_L g424 ( 
.A(n_330),
.B(n_289),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_326),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_370),
.B(n_248),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_327),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_350),
.A2(n_289),
.B(n_85),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_373),
.B(n_12),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g430 ( 
.A1(n_354),
.A2(n_252),
.B(n_248),
.Y(n_430)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_361),
.B(n_13),
.Y(n_431)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_379),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_376),
.A2(n_252),
.B(n_248),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g435 ( 
.A1(n_372),
.A2(n_252),
.B(n_248),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_327),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_377),
.A2(n_84),
.B(n_159),
.Y(n_437)
);

NOR2xp67_ASAP7_75t_L g438 ( 
.A(n_322),
.B(n_22),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_327),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_379),
.B(n_13),
.Y(n_440)
);

INVx3_ASAP7_75t_L g441 ( 
.A(n_345),
.Y(n_441)
);

INVx3_ASAP7_75t_L g442 ( 
.A(n_345),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_363),
.A2(n_86),
.B(n_158),
.Y(n_443)
);

O2A1O1Ixp33_ASAP7_75t_L g444 ( 
.A1(n_375),
.A2(n_14),
.B(n_15),
.C(n_16),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_379),
.B(n_15),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_365),
.B(n_370),
.Y(n_446)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_371),
.A2(n_87),
.B(n_23),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_374),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_379),
.B(n_17),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_381),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_360),
.B(n_17),
.Y(n_451)
);

AO31x2_ASAP7_75t_L g452 ( 
.A1(n_403),
.A2(n_368),
.A3(n_382),
.B(n_360),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_429),
.A2(n_336),
.B1(n_379),
.B2(n_358),
.Y(n_453)
);

NOR2x1_ASAP7_75t_SL g454 ( 
.A(n_432),
.B(n_345),
.Y(n_454)
);

OAI21x1_ASAP7_75t_L g455 ( 
.A1(n_398),
.A2(n_366),
.B(n_28),
.Y(n_455)
);

AOI21xp5_ASAP7_75t_L g456 ( 
.A1(n_383),
.A2(n_25),
.B(n_30),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_413),
.B(n_34),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g458 ( 
.A1(n_402),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_458)
);

OAI21x1_ASAP7_75t_L g459 ( 
.A1(n_392),
.A2(n_39),
.B(n_40),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_389),
.B(n_41),
.Y(n_460)
);

AOI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_432),
.A2(n_43),
.B(n_46),
.Y(n_461)
);

AOI21xp5_ASAP7_75t_L g462 ( 
.A1(n_409),
.A2(n_47),
.B(n_49),
.Y(n_462)
);

AOI21x1_ASAP7_75t_L g463 ( 
.A1(n_401),
.A2(n_50),
.B(n_51),
.Y(n_463)
);

NAND3xp33_ASAP7_75t_L g464 ( 
.A(n_406),
.B(n_387),
.C(n_385),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_417),
.A2(n_53),
.B(n_55),
.Y(n_465)
);

INVx4_ASAP7_75t_L g466 ( 
.A(n_427),
.Y(n_466)
);

OAI21x1_ASAP7_75t_L g467 ( 
.A1(n_393),
.A2(n_56),
.B(n_57),
.Y(n_467)
);

OAI21x1_ASAP7_75t_L g468 ( 
.A1(n_400),
.A2(n_58),
.B(n_61),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_426),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_404),
.A2(n_405),
.B(n_399),
.Y(n_470)
);

OAI21x1_ASAP7_75t_L g471 ( 
.A1(n_423),
.A2(n_63),
.B(n_64),
.Y(n_471)
);

HB1xp67_ASAP7_75t_L g472 ( 
.A(n_446),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_419),
.A2(n_65),
.B(n_67),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_388),
.B(n_68),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_416),
.A2(n_69),
.B(n_70),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g476 ( 
.A1(n_440),
.A2(n_73),
.B(n_74),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_407),
.B(n_75),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g478 ( 
.A1(n_445),
.A2(n_77),
.B(n_78),
.Y(n_478)
);

OAI21x1_ASAP7_75t_SL g479 ( 
.A1(n_449),
.A2(n_79),
.B(n_80),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_450),
.B(n_82),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_408),
.Y(n_481)
);

AND2x4_ASAP7_75t_L g482 ( 
.A(n_425),
.B(n_83),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_451),
.A2(n_88),
.B(n_89),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_431),
.B(n_90),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_390),
.B(n_91),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_436),
.B(n_92),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_415),
.A2(n_94),
.B(n_95),
.Y(n_487)
);

OAI21x1_ASAP7_75t_L g488 ( 
.A1(n_391),
.A2(n_97),
.B(n_98),
.Y(n_488)
);

A2O1A1Ixp33_ASAP7_75t_L g489 ( 
.A1(n_443),
.A2(n_99),
.B(n_100),
.C(n_105),
.Y(n_489)
);

A2O1A1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_444),
.A2(n_106),
.B(n_107),
.C(n_108),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_428),
.A2(n_109),
.B(n_110),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_436),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.Y(n_492)
);

AO31x2_ASAP7_75t_L g493 ( 
.A1(n_386),
.A2(n_117),
.A3(n_118),
.B(n_119),
.Y(n_493)
);

A2O1A1Ixp33_ASAP7_75t_L g494 ( 
.A1(n_384),
.A2(n_125),
.B(n_126),
.C(n_128),
.Y(n_494)
);

OAI21x1_ASAP7_75t_L g495 ( 
.A1(n_435),
.A2(n_129),
.B(n_132),
.Y(n_495)
);

AND2x2_ASAP7_75t_SL g496 ( 
.A(n_427),
.B(n_439),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_441),
.B(n_442),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_424),
.Y(n_498)
);

OAI21x1_ASAP7_75t_L g499 ( 
.A1(n_437),
.A2(n_136),
.B(n_137),
.Y(n_499)
);

O2A1O1Ixp33_ASAP7_75t_L g500 ( 
.A1(n_420),
.A2(n_138),
.B(n_139),
.C(n_143),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_410),
.Y(n_501)
);

OAI21x1_ASAP7_75t_L g502 ( 
.A1(n_433),
.A2(n_144),
.B(n_145),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_396),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g504 ( 
.A1(n_394),
.A2(n_147),
.B(n_149),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

OAI21x1_ASAP7_75t_L g506 ( 
.A1(n_455),
.A2(n_447),
.B(n_421),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_395),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_486),
.Y(n_508)
);

AO21x2_ASAP7_75t_L g509 ( 
.A1(n_491),
.A2(n_411),
.B(n_438),
.Y(n_509)
);

BUFx6f_ASAP7_75t_L g510 ( 
.A(n_496),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_498),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_464),
.A2(n_414),
.B(n_397),
.Y(n_512)
);

OAI21x1_ASAP7_75t_L g513 ( 
.A1(n_487),
.A2(n_438),
.B(n_418),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_481),
.B(n_434),
.Y(n_514)
);

INVx8_ASAP7_75t_L g515 ( 
.A(n_482),
.Y(n_515)
);

CKINVDCx6p67_ASAP7_75t_R g516 ( 
.A(n_482),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_505),
.Y(n_517)
);

OAI21x1_ASAP7_75t_L g518 ( 
.A1(n_467),
.A2(n_430),
.B(n_442),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_468),
.A2(n_441),
.B(n_412),
.Y(n_519)
);

INVx1_ASAP7_75t_SL g520 ( 
.A(n_469),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

OAI21x1_ASAP7_75t_L g522 ( 
.A1(n_459),
.A2(n_448),
.B(n_427),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_452),
.Y(n_523)
);

OA21x2_ASAP7_75t_L g524 ( 
.A1(n_470),
.A2(n_439),
.B(n_156),
.Y(n_524)
);

A2O1A1Ixp33_ASAP7_75t_L g525 ( 
.A1(n_504),
.A2(n_439),
.B(n_155),
.C(n_160),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_471),
.A2(n_499),
.B(n_488),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_486),
.Y(n_527)
);

BUFx12f_ASAP7_75t_L g528 ( 
.A(n_466),
.Y(n_528)
);

BUFx3_ASAP7_75t_L g529 ( 
.A(n_466),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_452),
.Y(n_530)
);

NOR2xp67_ASAP7_75t_L g531 ( 
.A(n_453),
.B(n_484),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_503),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_502),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_497),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_453),
.B(n_485),
.Y(n_535)
);

INVx2_ASAP7_75t_SL g536 ( 
.A(n_497),
.Y(n_536)
);

OAI21x1_ASAP7_75t_SL g537 ( 
.A1(n_477),
.A2(n_454),
.B(n_479),
.Y(n_537)
);

OAI21x1_ASAP7_75t_L g538 ( 
.A1(n_456),
.A2(n_478),
.B(n_462),
.Y(n_538)
);

INVx3_ASAP7_75t_L g539 ( 
.A(n_463),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_457),
.Y(n_540)
);

NOR4xp25_ASAP7_75t_L g541 ( 
.A(n_500),
.B(n_464),
.C(n_490),
.D(n_494),
.Y(n_541)
);

INVx6_ASAP7_75t_L g542 ( 
.A(n_461),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_480),
.Y(n_543)
);

A2O1A1Ixp33_ASAP7_75t_L g544 ( 
.A1(n_489),
.A2(n_483),
.B(n_460),
.C(n_474),
.Y(n_544)
);

NAND2x1p5_ASAP7_75t_L g545 ( 
.A(n_495),
.B(n_465),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_475),
.A2(n_476),
.B(n_473),
.Y(n_546)
);

OA21x2_ASAP7_75t_L g547 ( 
.A1(n_452),
.A2(n_458),
.B(n_492),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_493),
.Y(n_548)
);

AOI21xp33_ASAP7_75t_L g549 ( 
.A1(n_493),
.A2(n_318),
.B(n_265),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_528),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_521),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_517),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_514),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_514),
.Y(n_554)
);

BUFx2_ASAP7_75t_L g555 ( 
.A(n_508),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_516),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_527),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_526),
.A2(n_493),
.B(n_519),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_517),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_523),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_532),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_523),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_530),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_515),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_534),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_515),
.Y(n_566)
);

OAI21x1_ASAP7_75t_L g567 ( 
.A1(n_526),
.A2(n_519),
.B(n_522),
.Y(n_567)
);

NAND2x1p5_ASAP7_75t_L g568 ( 
.A(n_508),
.B(n_510),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_516),
.Y(n_569)
);

OAI21x1_ASAP7_75t_L g570 ( 
.A1(n_522),
.A2(n_506),
.B(n_513),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_530),
.Y(n_571)
);

INVx2_ASAP7_75t_SL g572 ( 
.A(n_515),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g573 ( 
.A(n_511),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_507),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_538),
.A2(n_531),
.B(n_506),
.Y(n_575)
);

AO21x1_ASAP7_75t_SL g576 ( 
.A1(n_540),
.A2(n_512),
.B(n_549),
.Y(n_576)
);

AOI22xp33_ASAP7_75t_SL g577 ( 
.A1(n_535),
.A2(n_515),
.B1(n_508),
.B2(n_510),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_510),
.Y(n_578)
);

OAI22xp33_ASAP7_75t_L g579 ( 
.A1(n_535),
.A2(n_520),
.B1(n_510),
.B2(n_528),
.Y(n_579)
);

AND2x4_ASAP7_75t_L g580 ( 
.A(n_511),
.B(n_529),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_536),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_536),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_529),
.Y(n_583)
);

OA21x2_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_538),
.B(n_513),
.Y(n_584)
);

HB1xp67_ASAP7_75t_L g585 ( 
.A(n_524),
.Y(n_585)
);

OAI221xp5_ASAP7_75t_L g586 ( 
.A1(n_525),
.A2(n_541),
.B1(n_544),
.B2(n_543),
.C(n_547),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_524),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_542),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_524),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_518),
.Y(n_590)
);

OAI221xp5_ASAP7_75t_L g591 ( 
.A1(n_525),
.A2(n_544),
.B1(n_543),
.B2(n_547),
.C(n_542),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_574),
.B(n_547),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_588),
.Y(n_593)
);

BUFx2_ASAP7_75t_SL g594 ( 
.A(n_556),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_551),
.Y(n_595)
);

OAI21xp33_ASAP7_75t_SL g596 ( 
.A1(n_591),
.A2(n_546),
.B(n_518),
.Y(n_596)
);

BUFx12f_ASAP7_75t_L g597 ( 
.A(n_550),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_571),
.Y(n_598)
);

AND2x2_ASAP7_75t_L g599 ( 
.A(n_553),
.B(n_548),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_571),
.Y(n_600)
);

BUFx6f_ASAP7_75t_L g601 ( 
.A(n_588),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g602 ( 
.A(n_556),
.Y(n_602)
);

INVxp67_ASAP7_75t_L g603 ( 
.A(n_557),
.Y(n_603)
);

AOI22xp33_ASAP7_75t_L g604 ( 
.A1(n_579),
.A2(n_509),
.B1(n_542),
.B2(n_537),
.Y(n_604)
);

AOI22xp33_ASAP7_75t_L g605 ( 
.A1(n_554),
.A2(n_509),
.B1(n_542),
.B2(n_539),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g606 ( 
.A(n_560),
.B(n_509),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_561),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_SL g608 ( 
.A1(n_586),
.A2(n_533),
.B1(n_545),
.B2(n_539),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_559),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_552),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_555),
.B(n_533),
.Y(n_613)
);

AND2x4_ASAP7_75t_L g614 ( 
.A(n_578),
.B(n_539),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g615 ( 
.A(n_562),
.B(n_563),
.Y(n_615)
);

BUFx2_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

AND2x2_ASAP7_75t_L g617 ( 
.A(n_577),
.B(n_533),
.Y(n_617)
);

AND2x2_ASAP7_75t_L g618 ( 
.A(n_576),
.B(n_533),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_576),
.B(n_533),
.Y(n_619)
);

OR2x2_ASAP7_75t_L g620 ( 
.A(n_563),
.B(n_581),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_568),
.B(n_545),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_587),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_568),
.B(n_546),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_583),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_568),
.B(n_582),
.Y(n_625)
);

BUFx6f_ASAP7_75t_L g626 ( 
.A(n_564),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_569),
.A2(n_580),
.B1(n_573),
.B2(n_564),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_580),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_589),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_580),
.Y(n_630)
);

AND2x4_ASAP7_75t_L g631 ( 
.A(n_566),
.B(n_572),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_585),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_558),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_566),
.Y(n_634)
);

INVx2_ASAP7_75t_SL g635 ( 
.A(n_550),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_572),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_575),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_584),
.B(n_575),
.Y(n_638)
);

BUFx2_ASAP7_75t_L g639 ( 
.A(n_584),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_592),
.B(n_584),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_598),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_594),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_612),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_595),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_607),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_598),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_609),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_624),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_599),
.A2(n_590),
.B1(n_558),
.B2(n_567),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_600),
.Y(n_651)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_632),
.B(n_590),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_622),
.Y(n_653)
);

BUFx3_ASAP7_75t_L g654 ( 
.A(n_597),
.Y(n_654)
);

OR2x2_ASAP7_75t_L g655 ( 
.A(n_592),
.B(n_616),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_622),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_613),
.B(n_570),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_603),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_613),
.B(n_617),
.Y(n_659)
);

OAI22xp5_ASAP7_75t_L g660 ( 
.A1(n_602),
.A2(n_567),
.B1(n_570),
.B2(n_608),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_597),
.Y(n_661)
);

AOI22xp33_ASAP7_75t_L g662 ( 
.A1(n_599),
.A2(n_617),
.B1(n_605),
.B2(n_593),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_616),
.B(n_639),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_593),
.A2(n_601),
.B1(n_628),
.B2(n_630),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g665 ( 
.A1(n_602),
.A2(n_627),
.B1(n_604),
.B2(n_635),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_620),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_620),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_625),
.B(n_593),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_618),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_593),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_625),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_629),
.B(n_639),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_629),
.Y(n_673)
);

INVx5_ASAP7_75t_L g674 ( 
.A(n_618),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_610),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_623),
.B(n_619),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_606),
.B(n_615),
.Y(n_677)
);

HB1xp67_ASAP7_75t_L g678 ( 
.A(n_614),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_659),
.B(n_623),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_643),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_659),
.B(n_619),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_653),
.Y(n_682)
);

AND2x2_ASAP7_75t_L g683 ( 
.A(n_676),
.B(n_633),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_644),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_658),
.B(n_635),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_670),
.B(n_601),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_653),
.Y(n_688)
);

AND2x2_ASAP7_75t_L g689 ( 
.A(n_676),
.B(n_633),
.Y(n_689)
);

NAND2x1p5_ASAP7_75t_SL g690 ( 
.A(n_663),
.B(n_621),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_641),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_648),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_649),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_673),
.Y(n_694)
);

NAND2x1p5_ASAP7_75t_L g695 ( 
.A(n_670),
.B(n_621),
.Y(n_695)
);

INVx3_ASAP7_75t_L g696 ( 
.A(n_674),
.Y(n_696)
);

NAND2x1p5_ASAP7_75t_L g697 ( 
.A(n_670),
.B(n_593),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_674),
.B(n_669),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_641),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_655),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_669),
.B(n_637),
.Y(n_701)
);

HB1xp67_ASAP7_75t_L g702 ( 
.A(n_655),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_646),
.Y(n_703)
);

INVx3_ASAP7_75t_L g704 ( 
.A(n_674),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_657),
.B(n_637),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_663),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_646),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_674),
.B(n_614),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_680),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_685),
.A2(n_665),
.B1(n_664),
.B2(n_662),
.C(n_660),
.Y(n_710)
);

OAI33xp33_ASAP7_75t_L g711 ( 
.A1(n_684),
.A2(n_667),
.A3(n_666),
.B1(n_672),
.B2(n_668),
.B3(n_675),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_686),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_692),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_693),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_706),
.B(n_642),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_682),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_700),
.B(n_640),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_702),
.B(n_640),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_682),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_688),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_681),
.B(n_674),
.Y(n_723)
);

INVxp67_ASAP7_75t_SL g724 ( 
.A(n_688),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_679),
.B(n_678),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_681),
.B(n_657),
.Y(n_726)
);

OR2x2_ASAP7_75t_L g727 ( 
.A(n_690),
.B(n_672),
.Y(n_727)
);

OAI21xp33_ASAP7_75t_L g728 ( 
.A1(n_727),
.A2(n_705),
.B(n_679),
.Y(n_728)
);

OAI21xp33_ASAP7_75t_L g729 ( 
.A1(n_722),
.A2(n_705),
.B(n_683),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_716),
.Y(n_730)
);

AOI21xp33_ASAP7_75t_L g731 ( 
.A1(n_710),
.A2(n_694),
.B(n_671),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_719),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_722),
.B(n_698),
.Y(n_733)
);

OAI21xp33_ASAP7_75t_L g734 ( 
.A1(n_724),
.A2(n_689),
.B(n_683),
.Y(n_734)
);

NOR2xp67_ASAP7_75t_L g735 ( 
.A(n_717),
.B(n_704),
.Y(n_735)
);

NOR2x1p5_ASAP7_75t_L g736 ( 
.A(n_725),
.B(n_661),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_715),
.A2(n_698),
.B1(n_704),
.B2(n_696),
.Y(n_737)
);

NAND2x1_ASAP7_75t_L g738 ( 
.A(n_723),
.B(n_698),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_731),
.A2(n_711),
.B1(n_601),
.B2(n_671),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_734),
.B(n_724),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_736),
.A2(n_711),
.B1(n_715),
.B2(n_689),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_738),
.B(n_726),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_728),
.A2(n_713),
.B1(n_709),
.B2(n_712),
.C(n_714),
.Y(n_743)
);

AOI21xp5_ASAP7_75t_L g744 ( 
.A1(n_733),
.A2(n_687),
.B(n_718),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_742),
.B(n_735),
.Y(n_745)
);

NOR4xp25_ASAP7_75t_SL g746 ( 
.A(n_743),
.B(n_729),
.C(n_732),
.D(n_730),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_741),
.B(n_739),
.Y(n_747)
);

OAI221xp5_ASAP7_75t_L g748 ( 
.A1(n_740),
.A2(n_737),
.B1(n_720),
.B2(n_661),
.C(n_654),
.Y(n_748)
);

O2A1O1Ixp5_ASAP7_75t_L g749 ( 
.A1(n_744),
.A2(n_704),
.B(n_696),
.C(n_701),
.Y(n_749)
);

AOI221xp5_ASAP7_75t_L g750 ( 
.A1(n_739),
.A2(n_690),
.B1(n_694),
.B2(n_596),
.C(n_654),
.Y(n_750)
);

NAND4xp25_ASAP7_75t_SL g751 ( 
.A(n_750),
.B(n_701),
.C(n_650),
.D(n_634),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_747),
.B(n_636),
.Y(n_752)
);

OR2x2_ASAP7_75t_L g753 ( 
.A(n_748),
.B(n_652),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_745),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_746),
.B(n_670),
.C(n_626),
.Y(n_755)
);

NAND3xp33_ASAP7_75t_L g756 ( 
.A(n_752),
.B(n_755),
.C(n_749),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_754),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_753),
.Y(n_758)
);

NAND4xp75_ASAP7_75t_L g759 ( 
.A(n_757),
.B(n_751),
.C(n_673),
.D(n_651),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_758),
.Y(n_760)
);

OAI22xp5_ASAP7_75t_L g761 ( 
.A1(n_756),
.A2(n_696),
.B1(n_708),
.B2(n_697),
.Y(n_761)
);

AND2x4_ASAP7_75t_L g762 ( 
.A(n_760),
.B(n_708),
.Y(n_762)
);

NAND4xp75_ASAP7_75t_L g763 ( 
.A(n_759),
.B(n_651),
.C(n_721),
.D(n_638),
.Y(n_763)
);

NOR2x1p5_ASAP7_75t_L g764 ( 
.A(n_761),
.B(n_626),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_760),
.Y(n_765)
);

OR2x2_ASAP7_75t_L g766 ( 
.A(n_760),
.B(n_652),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_763),
.A2(n_670),
.B1(n_614),
.B2(n_631),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_765),
.Y(n_768)
);

XOR2x1_ASAP7_75t_L g769 ( 
.A(n_762),
.B(n_697),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_766),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_764),
.Y(n_771)
);

AO22x2_ASAP7_75t_L g772 ( 
.A1(n_765),
.A2(n_631),
.B1(n_708),
.B2(n_703),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_768),
.B(n_697),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_770),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_771),
.B(n_631),
.Y(n_775)
);

OR3x2_ASAP7_75t_L g776 ( 
.A(n_769),
.B(n_677),
.C(n_626),
.Y(n_776)
);

AO22x2_ASAP7_75t_L g777 ( 
.A1(n_772),
.A2(n_707),
.B1(n_703),
.B2(n_699),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_775),
.A2(n_767),
.B1(n_601),
.B2(n_626),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_774),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_773),
.B(n_695),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_776),
.Y(n_781)
);

INVx1_ASAP7_75t_SL g782 ( 
.A(n_777),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_779),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_781),
.A2(n_777),
.B1(n_626),
.B2(n_699),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_778),
.A2(n_695),
.B1(n_707),
.B2(n_691),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_783),
.A2(n_782),
.B1(n_780),
.B2(n_695),
.Y(n_786)
);

HB1xp67_ASAP7_75t_L g787 ( 
.A(n_786),
.Y(n_787)
);

XNOR2x1_ASAP7_75t_L g788 ( 
.A(n_787),
.B(n_785),
.Y(n_788)
);

AOI221xp5_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_784),
.B1(n_637),
.B2(n_611),
.C(n_656),
.Y(n_789)
);

AOI211xp5_ASAP7_75t_L g790 ( 
.A1(n_789),
.A2(n_656),
.B(n_647),
.C(n_606),
.Y(n_790)
);


endmodule