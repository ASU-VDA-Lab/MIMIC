module fake_netlist_1_7235_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_15, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_15;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_16;
wire n_33;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
INVx6_ASAP7_75t_L g16 ( .A(n_11), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_9), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_0), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_7), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_5), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_7), .Y(n_21) );
INVx2_ASAP7_75t_L g22 ( .A(n_6), .Y(n_22) );
INVxp67_ASAP7_75t_L g23 ( .A(n_8), .Y(n_23) );
AOI21xp5_ASAP7_75t_L g24 ( .A1(n_23), .A2(n_15), .B(n_14), .Y(n_24) );
NAND2xp5_ASAP7_75t_L g25 ( .A(n_17), .B(n_22), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_21), .B(n_0), .Y(n_26) );
NAND2xp5_ASAP7_75t_SL g27 ( .A(n_20), .B(n_1), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_19), .B1(n_18), .B2(n_20), .Y(n_28) );
AOI21x1_ASAP7_75t_L g29 ( .A1(n_24), .A2(n_19), .B(n_18), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_25), .Y(n_30) );
INVx2_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
AND2x2_ASAP7_75t_L g32 ( .A(n_30), .B(n_20), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_28), .Y(n_33) );
INVx1_ASAP7_75t_L g34 ( .A(n_31), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_33), .Y(n_35) );
OR2x2_ASAP7_75t_L g36 ( .A(n_33), .B(n_27), .Y(n_36) );
INVx2_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AOI31xp67_ASAP7_75t_SL g38 ( .A1(n_35), .A2(n_1), .A3(n_2), .B(n_3), .Y(n_38) );
AND2x2_ASAP7_75t_SL g39 ( .A(n_37), .B(n_34), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_36), .A2(n_16), .B1(n_29), .B2(n_4), .Y(n_40) );
NOR4xp75_ASAP7_75t_L g41 ( .A(n_38), .B(n_2), .C(n_3), .D(n_4), .Y(n_41) );
INVx1_ASAP7_75t_L g42 ( .A(n_39), .Y(n_42) );
INVx1_ASAP7_75t_L g43 ( .A(n_40), .Y(n_43) );
XNOR2xp5_ASAP7_75t_L g44 ( .A(n_41), .B(n_40), .Y(n_44) );
AOI21x1_ASAP7_75t_L g45 ( .A1(n_43), .A2(n_37), .B(n_16), .Y(n_45) );
OAI22x1_ASAP7_75t_L g46 ( .A1(n_44), .A2(n_42), .B1(n_6), .B2(n_5), .Y(n_46) );
OA331x2_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_44), .A3(n_45), .B1(n_42), .B2(n_13), .B3(n_10), .C1(n_12), .Y(n_47) );
endmodule