module fake_jpeg_3514_n_722 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_722);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_722;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_716;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_717;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_718;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_713;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_704;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_715;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_720;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_710;
wire n_610;
wire n_174;
wire n_714;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_709;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_708;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_650;
wire n_344;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_398;
wire n_240;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_719;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_707;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_705;
wire n_665;
wire n_706;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_721;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_712;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_711;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx12_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_7),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_15),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_4),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_9),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_9),
.Y(n_61)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_62),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_63),
.Y(n_136)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_21),
.Y(n_64)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_64),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx4f_ASAP7_75t_SL g176 ( 
.A(n_65),
.Y(n_176)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g196 ( 
.A(n_66),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_35),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_67),
.Y(n_147)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_68),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_69),
.Y(n_148)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_70),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_71),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_29),
.B(n_19),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_72),
.B(n_75),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_28),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_37),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_76),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_77),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_37),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_78),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_28),
.B(n_19),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_79),
.B(n_85),
.Y(n_153)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_37),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_81),
.Y(n_212)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_21),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g171 ( 
.A(n_84),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_18),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_86),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_48),
.B(n_18),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_87),
.B(n_101),
.Y(n_182)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_88),
.Y(n_155)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_89),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_42),
.Y(n_90)
);

INVx5_ASAP7_75t_L g163 ( 
.A(n_90),
.Y(n_163)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_91),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_61),
.B(n_18),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_92),
.B(n_100),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_93),
.Y(n_219)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_94),
.Y(n_140)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_21),
.Y(n_95)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_95),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_96),
.Y(n_228)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_24),
.Y(n_97)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_97),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_40),
.Y(n_98)
);

INVx5_ASAP7_75t_L g209 ( 
.A(n_98),
.Y(n_209)
);

BUFx12_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_22),
.B(n_18),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_53),
.B(n_17),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_21),
.Y(n_102)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_102),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_23),
.B(n_17),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_103),
.B(n_109),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_104),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_55),
.Y(n_106)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_106),
.Y(n_206)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_31),
.Y(n_107)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_107),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_58),
.Y(n_108)
);

INVx6_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_17),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_23),
.B(n_17),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_110),
.B(n_126),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_58),
.Y(n_111)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_111),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_58),
.Y(n_112)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_58),
.Y(n_113)
);

INVx3_ASAP7_75t_SL g154 ( 
.A(n_113),
.Y(n_154)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_114),
.Y(n_188)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_31),
.Y(n_115)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_115),
.Y(n_158)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_31),
.Y(n_116)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_116),
.Y(n_177)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_117),
.Y(n_218)
);

BUFx5_ASAP7_75t_L g118 ( 
.A(n_24),
.Y(n_118)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_119),
.Y(n_204)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_50),
.Y(n_120)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_120),
.Y(n_226)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

INVx4_ASAP7_75t_L g221 ( 
.A(n_121),
.Y(n_221)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_50),
.Y(n_122)
);

INVx8_ASAP7_75t_L g168 ( 
.A(n_122),
.Y(n_168)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_50),
.Y(n_123)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_123),
.Y(n_185)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_23),
.Y(n_124)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_124),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_125),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_16),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_38),
.Y(n_127)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_127),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_23),
.Y(n_128)
);

CKINVDCx14_ASAP7_75t_R g205 ( 
.A(n_128),
.Y(n_205)
);

BUFx12f_ASAP7_75t_L g129 ( 
.A(n_40),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_129),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_56),
.Y(n_130)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_130),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_131),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_38),
.Y(n_132)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_132),
.Y(n_229)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_38),
.Y(n_133)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_133),
.Y(n_159)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_23),
.Y(n_134)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_134),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_128),
.A2(n_32),
.B1(n_51),
.B2(n_54),
.Y(n_141)
);

OA22x2_ASAP7_75t_L g299 ( 
.A1(n_141),
.A2(n_156),
.B1(n_180),
.B2(n_1),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_103),
.A2(n_36),
.B1(n_49),
.B2(n_54),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_144),
.A2(n_160),
.B1(n_170),
.B2(n_181),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_32),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_145),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_86),
.A2(n_36),
.B1(n_49),
.B2(n_52),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g257 ( 
.A(n_146),
.B(n_150),
.Y(n_257)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_99),
.B(n_43),
.CON(n_150),
.SN(n_150)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_152),
.B(n_157),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_97),
.A2(n_64),
.B1(n_62),
.B2(n_117),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_130),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_96),
.A2(n_61),
.B1(n_30),
.B2(n_52),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_68),
.B(n_132),
.C(n_83),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_162),
.B(n_175),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_105),
.A2(n_22),
.B1(n_39),
.B2(n_34),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_71),
.Y(n_173)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_173),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_131),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_107),
.A2(n_51),
.B1(n_32),
.B2(n_34),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_89),
.A2(n_91),
.B1(n_69),
.B2(n_67),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_106),
.A2(n_39),
.B1(n_30),
.B2(n_60),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_187),
.A2(n_200),
.B1(n_211),
.B2(n_160),
.Y(n_276)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_63),
.A2(n_60),
.B1(n_20),
.B2(n_44),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_129),
.B(n_98),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_215),
.Y(n_288)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_112),
.Y(n_207)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_108),
.A2(n_113),
.B1(n_73),
.B2(n_76),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_208),
.A2(n_225),
.B1(n_41),
.B2(n_47),
.Y(n_239)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_84),
.Y(n_210)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_210),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g211 ( 
.A1(n_77),
.A2(n_20),
.B1(n_46),
.B2(n_45),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_65),
.B(n_46),
.Y(n_215)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_90),
.B(n_45),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_216),
.B(n_217),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_129),
.B(n_44),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_L g225 ( 
.A1(n_78),
.A2(n_43),
.B1(n_47),
.B2(n_41),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_136),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_231),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_220),
.A2(n_32),
.B1(n_51),
.B2(n_41),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_232),
.A2(n_242),
.B1(n_244),
.B2(n_248),
.Y(n_312)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_203),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g321 ( 
.A(n_233),
.Y(n_321)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_234),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_202),
.B(n_47),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_246),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_176),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_236),
.B(n_280),
.Y(n_329)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_168),
.Y(n_237)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_237),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_205),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_238),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_239),
.A2(n_277),
.B1(n_281),
.B2(n_292),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_184),
.A2(n_192),
.B1(n_153),
.B2(n_182),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g342 ( 
.A(n_241),
.Y(n_342)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_143),
.A2(n_32),
.B1(n_51),
.B2(n_122),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_243),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_196),
.A2(n_51),
.B1(n_123),
.B2(n_120),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_222),
.Y(n_245)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_245),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_145),
.B(n_65),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_216),
.A2(n_99),
.B(n_98),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g369 ( 
.A(n_247),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_196),
.A2(n_119),
.B1(n_95),
.B2(n_124),
.Y(n_248)
);

INVx3_ASAP7_75t_L g249 ( 
.A(n_169),
.Y(n_249)
);

BUFx4f_ASAP7_75t_SL g336 ( 
.A(n_249),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_140),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_250),
.B(n_256),
.Y(n_347)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_186),
.Y(n_251)
);

INVx4_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

INVx11_ASAP7_75t_L g253 ( 
.A(n_161),
.Y(n_253)
);

INVx11_ASAP7_75t_L g360 ( 
.A(n_253),
.Y(n_360)
);

INVx4_ASAP7_75t_SL g254 ( 
.A(n_161),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_255),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_141),
.A2(n_205),
.B(n_180),
.Y(n_256)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_168),
.Y(n_260)
);

BUFx12f_ASAP7_75t_L g334 ( 
.A(n_260),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_135),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_262),
.B(n_271),
.Y(n_317)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_159),
.Y(n_263)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_263),
.Y(n_367)
);

INVx5_ASAP7_75t_L g266 ( 
.A(n_186),
.Y(n_266)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_266),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_158),
.B(n_0),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_267),
.B(n_272),
.Y(n_351)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_154),
.Y(n_268)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_268),
.Y(n_372)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_161),
.Y(n_269)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_269),
.Y(n_349)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_154),
.Y(n_270)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_270),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_135),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_177),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_183),
.B(n_1),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_274),
.B(n_275),
.Y(n_352)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_150),
.A2(n_24),
.B(n_27),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_276),
.A2(n_283),
.B1(n_284),
.B2(n_299),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_170),
.A2(n_93),
.B1(n_81),
.B2(n_43),
.Y(n_277)
);

BUFx3_ASAP7_75t_L g278 ( 
.A(n_189),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g344 ( 
.A(n_278),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_189),
.Y(n_279)
);

INVx6_ASAP7_75t_L g314 ( 
.A(n_279),
.Y(n_314)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_137),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_187),
.A2(n_43),
.B1(n_27),
.B2(n_40),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_222),
.Y(n_282)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_282),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_SL g283 ( 
.A1(n_174),
.A2(n_43),
.B1(n_27),
.B2(n_40),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_188),
.A2(n_16),
.B1(n_15),
.B2(n_13),
.Y(n_284)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_136),
.Y(n_285)
);

INVx8_ASAP7_75t_L g346 ( 
.A(n_285),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_208),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_286),
.A2(n_290),
.B1(n_224),
.B2(n_206),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_138),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_287),
.B(n_291),
.Y(n_322)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_185),
.Y(n_289)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_289),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_225),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_142),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_211),
.A2(n_12),
.B1(n_11),
.B2(n_3),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_147),
.Y(n_293)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_293),
.Y(n_359)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_139),
.Y(n_294)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_294),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_147),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_295),
.Y(n_361)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_229),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_296),
.B(n_297),
.Y(n_325)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_190),
.Y(n_297)
);

BUFx12_ASAP7_75t_L g298 ( 
.A(n_176),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_298),
.Y(n_362)
);

INVx8_ASAP7_75t_L g300 ( 
.A(n_228),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_SL g327 ( 
.A1(n_300),
.A2(n_308),
.B1(n_309),
.B2(n_191),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_151),
.B(n_2),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_301),
.B(n_303),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_155),
.B(n_2),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_209),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_304),
.B(n_305),
.Y(n_331)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_213),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_172),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_306),
.B(n_307),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_171),
.Y(n_307)
);

INVx5_ASAP7_75t_L g308 ( 
.A(n_163),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g309 ( 
.A1(n_178),
.A2(n_11),
.B1(n_4),
.B2(n_5),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_213),
.B(n_214),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_310),
.B(n_286),
.Y(n_375)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_166),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_148),
.B1(n_219),
.B2(n_198),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_252),
.A2(n_228),
.B1(n_179),
.B2(n_167),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_313),
.A2(n_316),
.B1(n_343),
.B2(n_247),
.Y(n_376)
);

AOI22xp33_ASAP7_75t_L g316 ( 
.A1(n_256),
.A2(n_179),
.B1(n_167),
.B2(n_219),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_323),
.A2(n_345),
.B1(n_356),
.B2(n_363),
.Y(n_377)
);

AO22x1_ASAP7_75t_L g324 ( 
.A1(n_277),
.A2(n_171),
.B1(n_197),
.B2(n_193),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_324),
.B(n_245),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_274),
.B(n_235),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_326),
.B(n_272),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_327),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_250),
.B(n_221),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_328),
.B(n_375),
.Y(n_379)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_261),
.A2(n_226),
.B1(n_204),
.B2(n_164),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_333),
.A2(n_335),
.B1(n_350),
.B2(n_357),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g335 ( 
.A1(n_299),
.A2(n_164),
.B1(n_218),
.B2(n_165),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_L g343 ( 
.A1(n_239),
.A2(n_149),
.B1(n_148),
.B2(n_212),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_257),
.A2(n_214),
.B1(n_224),
.B2(n_206),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_299),
.A2(n_156),
.B1(n_212),
.B2(n_198),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_299),
.A2(n_149),
.B1(n_166),
.B2(n_6),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_302),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_358)
);

OAI211xp5_ASAP7_75t_L g403 ( 
.A1(n_358),
.A2(n_373),
.B(n_245),
.C(n_270),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_257),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_363)
);

OR2x2_ASAP7_75t_SL g368 ( 
.A(n_241),
.B(n_7),
.Y(n_368)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_368),
.Y(n_386)
);

AOI22xp33_ASAP7_75t_SL g371 ( 
.A1(n_288),
.A2(n_9),
.B1(n_7),
.B2(n_8),
.Y(n_371)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_371),
.Y(n_413)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_264),
.A2(n_9),
.B1(n_246),
.B2(n_275),
.Y(n_373)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_260),
.A2(n_249),
.B1(n_258),
.B2(n_237),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_374),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_376),
.A2(n_387),
.B1(n_401),
.B2(n_402),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_321),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_378),
.B(n_396),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_347),
.A2(n_290),
.B(n_291),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_380),
.A2(n_392),
.B(n_404),
.Y(n_432)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_381),
.Y(n_427)
);

A2O1A1Ixp33_ASAP7_75t_SL g383 ( 
.A1(n_347),
.A2(n_309),
.B(n_310),
.C(n_253),
.Y(n_383)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_383),
.Y(n_468)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_338),
.Y(n_384)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_384),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_385),
.B(n_399),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_375),
.A2(n_303),
.B1(n_301),
.B2(n_267),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_338),
.Y(n_388)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_388),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_351),
.B(n_255),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_389),
.B(n_393),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g390 ( 
.A(n_340),
.Y(n_390)
);

INVx6_ASAP7_75t_L g435 ( 
.A(n_390),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_320),
.A2(n_305),
.B1(n_234),
.B2(n_243),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g434 ( 
.A1(n_391),
.A2(n_409),
.B1(n_412),
.B2(n_353),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_352),
.A2(n_287),
.B(n_289),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_351),
.B(n_233),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_325),
.Y(n_394)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_394),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_263),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_395),
.B(n_415),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_340),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_319),
.B(n_265),
.C(n_259),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_397),
.B(n_416),
.Y(n_469)
);

BUFx12f_ASAP7_75t_L g398 ( 
.A(n_349),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_398),
.B(n_407),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_230),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_320),
.A2(n_318),
.B1(n_352),
.B2(n_356),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_373),
.A2(n_285),
.B1(n_300),
.B2(n_293),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_403),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_369),
.A2(n_273),
.B(n_240),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_336),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_405),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_L g406 ( 
.A1(n_369),
.A2(n_231),
.B1(n_295),
.B2(n_268),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g452 ( 
.A1(n_406),
.A2(n_410),
.B1(n_423),
.B2(n_372),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_321),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_336),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_408),
.Y(n_451)
);

AOI22xp33_ASAP7_75t_L g409 ( 
.A1(n_369),
.A2(n_297),
.B1(n_308),
.B2(n_296),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_364),
.A2(n_307),
.B1(n_282),
.B2(n_266),
.Y(n_410)
);

AND2x2_ASAP7_75t_L g411 ( 
.A(n_345),
.B(n_269),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_411),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_328),
.A2(n_251),
.B1(n_304),
.B2(n_254),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_321),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_422),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_326),
.B(n_278),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_319),
.B(n_298),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g418 ( 
.A(n_342),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_418),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_342),
.B(n_279),
.C(n_298),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_419),
.B(n_366),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_312),
.A2(n_363),
.B(n_317),
.Y(n_420)
);

AOI21xp5_ASAP7_75t_L g442 ( 
.A1(n_420),
.A2(n_330),
.B(n_341),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_355),
.B(n_337),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_367),
.Y(n_462)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_323),
.A2(n_324),
.B1(n_358),
.B2(n_361),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_322),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_424),
.B(n_425),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_331),
.Y(n_425)
);

AOI32xp33_ASAP7_75t_L g426 ( 
.A1(n_368),
.A2(n_329),
.A3(n_330),
.B1(n_332),
.B2(n_353),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_334),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_399),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_428),
.B(n_443),
.Y(n_474)
);

MAJx2_ASAP7_75t_L g430 ( 
.A(n_416),
.B(n_370),
.C(n_362),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_433),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_SL g433 ( 
.A(n_379),
.B(n_329),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_434),
.B(n_452),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_425),
.C(n_419),
.Y(n_475)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_442),
.A2(n_465),
.B(n_403),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_421),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_380),
.A2(n_324),
.B1(n_361),
.B2(n_346),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_445),
.A2(n_454),
.B1(n_459),
.B2(n_463),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_410),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_448),
.B(n_411),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g453 ( 
.A1(n_392),
.A2(n_362),
.B(n_349),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_453),
.A2(n_426),
.B(n_381),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_SL g454 ( 
.A1(n_377),
.A2(n_346),
.B1(n_348),
.B2(n_359),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_387),
.B(n_366),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_455),
.B(n_462),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_404),
.B(n_332),
.Y(n_457)
);

CKINVDCx16_ASAP7_75t_R g471 ( 
.A(n_457),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_401),
.A2(n_346),
.B1(n_336),
.B2(n_359),
.Y(n_458)
);

OAI22xp5_ASAP7_75t_L g476 ( 
.A1(n_458),
.A2(n_461),
.B1(n_464),
.B2(n_466),
.Y(n_476)
);

OAI22xp5_ASAP7_75t_SL g459 ( 
.A1(n_377),
.A2(n_348),
.B1(n_359),
.B2(n_341),
.Y(n_459)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_423),
.A2(n_336),
.B1(n_348),
.B2(n_372),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_379),
.A2(n_367),
.B1(n_315),
.B2(n_339),
.Y(n_463)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_376),
.A2(n_315),
.B1(n_339),
.B2(n_354),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_L g466 ( 
.A1(n_391),
.A2(n_334),
.B1(n_354),
.B2(n_365),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_470),
.A2(n_480),
.B(n_505),
.Y(n_537)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_472),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_438),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_473),
.B(n_479),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_475),
.B(n_478),
.C(n_486),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_446),
.A2(n_382),
.B1(n_420),
.B2(n_383),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g518 ( 
.A1(n_477),
.A2(n_497),
.B1(n_456),
.B2(n_445),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_469),
.B(n_393),
.C(n_395),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_438),
.Y(n_479)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_481),
.Y(n_525)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_465),
.A2(n_417),
.B(n_400),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g520 ( 
.A1(n_482),
.A2(n_491),
.B(n_503),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_444),
.B(n_389),
.Y(n_483)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_483),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_467),
.B(n_415),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_484),
.B(n_485),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_467),
.B(n_385),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_469),
.B(n_397),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_394),
.Y(n_487)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_487),
.Y(n_533)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_429),
.Y(n_490)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_490),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_436),
.A2(n_383),
.B(n_381),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_428),
.B(n_424),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_493),
.B(n_443),
.Y(n_513)
);

CKINVDCx20_ASAP7_75t_R g494 ( 
.A(n_431),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g524 ( 
.A(n_494),
.B(n_502),
.Y(n_524)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_495),
.Y(n_544)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_441),
.Y(n_496)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_496),
.Y(n_548)
);

OAI22x1_ASAP7_75t_SL g497 ( 
.A1(n_468),
.A2(n_383),
.B1(n_412),
.B2(n_411),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_446),
.A2(n_402),
.B1(n_411),
.B2(n_383),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_498),
.A2(n_500),
.B1(n_468),
.B2(n_458),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_446),
.A2(n_383),
.B1(n_406),
.B2(n_413),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_463),
.Y(n_501)
);

INVx1_ASAP7_75t_SL g538 ( 
.A(n_501),
.Y(n_538)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_449),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_432),
.A2(n_386),
.B(n_405),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_469),
.B(n_440),
.C(n_430),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_504),
.B(n_506),
.C(n_508),
.Y(n_531)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_432),
.A2(n_408),
.B(n_388),
.Y(n_505)
);

XOR2xp5_ASAP7_75t_L g506 ( 
.A(n_433),
.B(n_422),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_453),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_507),
.B(n_509),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_433),
.B(n_384),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_439),
.B(n_414),
.Y(n_509)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_511),
.A2(n_514),
.B1(n_516),
.B2(n_534),
.Y(n_565)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_513),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g514 ( 
.A1(n_498),
.A2(n_468),
.B1(n_452),
.B2(n_458),
.Y(n_514)
);

CKINVDCx20_ASAP7_75t_R g515 ( 
.A(n_509),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_515),
.B(n_523),
.Y(n_557)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_499),
.A2(n_452),
.B1(n_448),
.B2(n_461),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_470),
.B(n_457),
.Y(n_517)
);

INVx1_ASAP7_75t_SL g563 ( 
.A(n_517),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_518),
.A2(n_471),
.B1(n_507),
.B2(n_505),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_L g521 ( 
.A1(n_499),
.A2(n_500),
.B1(n_492),
.B2(n_487),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_L g577 ( 
.A1(n_521),
.A2(n_526),
.B1(n_528),
.B2(n_542),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_474),
.Y(n_523)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_497),
.A2(n_454),
.B1(n_459),
.B2(n_457),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_477),
.A2(n_439),
.B1(n_461),
.B2(n_427),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_473),
.B(n_449),
.Y(n_529)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_529),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_479),
.B(n_462),
.Y(n_530)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_530),
.Y(n_561)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_474),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_532),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_SL g534 ( 
.A1(n_499),
.A2(n_455),
.B1(n_464),
.B2(n_442),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_493),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_535),
.B(n_545),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_494),
.B(n_483),
.Y(n_539)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_539),
.Y(n_567)
);

CKINVDCx16_ASAP7_75t_R g540 ( 
.A(n_481),
.Y(n_540)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_540),
.Y(n_570)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_476),
.A2(n_427),
.B1(n_434),
.B2(n_464),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_504),
.B(n_440),
.C(n_430),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_543),
.B(n_486),
.C(n_508),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_484),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_489),
.B(n_450),
.Y(n_546)
);

INVxp33_ASAP7_75t_L g574 ( 
.A(n_546),
.Y(n_574)
);

XNOR2xp5_ASAP7_75t_SL g547 ( 
.A(n_488),
.B(n_450),
.Y(n_547)
);

XOR2xp5_ASAP7_75t_L g578 ( 
.A(n_547),
.B(n_472),
.Y(n_578)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_536),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_549),
.B(n_575),
.Y(n_593)
);

A2O1A1O1Ixp25_ASAP7_75t_L g550 ( 
.A1(n_545),
.A2(n_478),
.B(n_485),
.C(n_488),
.D(n_475),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_550),
.A2(n_576),
.B(n_530),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_551),
.A2(n_555),
.B1(n_562),
.B2(n_571),
.Y(n_585)
);

INVxp67_ASAP7_75t_L g552 ( 
.A(n_524),
.Y(n_552)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_552),
.Y(n_603)
);

OAI22xp5_ASAP7_75t_SL g555 ( 
.A1(n_518),
.A2(n_471),
.B1(n_507),
.B2(n_492),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_536),
.B(n_460),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_559),
.B(n_564),
.Y(n_587)
);

XNOR2xp5_ASAP7_75t_L g588 ( 
.A(n_560),
.B(n_531),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_526),
.A2(n_501),
.B1(n_491),
.B2(n_480),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_512),
.B(n_502),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_512),
.B(n_506),
.C(n_503),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g591 ( 
.A(n_566),
.B(n_543),
.C(n_531),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_535),
.B(n_396),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g605 ( 
.A(n_568),
.Y(n_605)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_513),
.Y(n_569)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_569),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_528),
.A2(n_491),
.B1(n_476),
.B2(n_489),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_524),
.Y(n_572)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_572),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_515),
.A2(n_496),
.B1(n_495),
.B2(n_490),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g586 ( 
.A1(n_573),
.A2(n_581),
.B1(n_540),
.B2(n_525),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_546),
.B(n_390),
.Y(n_575)
);

OAI21xp5_ASAP7_75t_L g576 ( 
.A1(n_537),
.A2(n_482),
.B(n_431),
.Y(n_576)
);

XOR2xp5_ASAP7_75t_L g594 ( 
.A(n_578),
.B(n_510),
.Y(n_594)
);

CKINVDCx20_ASAP7_75t_R g579 ( 
.A(n_529),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_579),
.A2(n_580),
.B1(n_583),
.B2(n_542),
.Y(n_600)
);

AOI22x1_ASAP7_75t_L g580 ( 
.A1(n_511),
.A2(n_466),
.B1(n_451),
.B2(n_447),
.Y(n_580)
);

OAI22xp5_ASAP7_75t_SL g581 ( 
.A1(n_525),
.A2(n_437),
.B1(n_386),
.B2(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_539),
.Y(n_582)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_582),
.Y(n_595)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_521),
.A2(n_437),
.B1(n_407),
.B2(n_378),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_510),
.Y(n_584)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_584),
.Y(n_604)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_586),
.Y(n_615)
);

XNOR2xp5_ASAP7_75t_L g627 ( 
.A(n_588),
.B(n_591),
.Y(n_627)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_590),
.Y(n_616)
);

XNOR2x1_ASAP7_75t_L g634 ( 
.A(n_594),
.B(n_609),
.Y(n_634)
);

MAJIxp5_ASAP7_75t_L g596 ( 
.A(n_560),
.B(n_547),
.C(n_532),
.Y(n_596)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_597),
.C(n_606),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_566),
.B(n_523),
.C(n_538),
.Y(n_597)
);

AOI22xp5_ASAP7_75t_L g598 ( 
.A1(n_577),
.A2(n_514),
.B1(n_538),
.B2(n_533),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g628 ( 
.A1(n_598),
.A2(n_583),
.B1(n_554),
.B2(n_553),
.Y(n_628)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_584),
.Y(n_599)
);

CKINVDCx14_ASAP7_75t_R g630 ( 
.A(n_599),
.Y(n_630)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_600),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g601 ( 
.A(n_556),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_601),
.B(n_572),
.Y(n_618)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_578),
.B(n_520),
.Y(n_602)
);

XOR2xp5_ASAP7_75t_L g637 ( 
.A(n_602),
.B(n_581),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_563),
.B(n_520),
.C(n_537),
.Y(n_606)
);

OAI22x1_ASAP7_75t_L g607 ( 
.A1(n_565),
.A2(n_517),
.B1(n_522),
.B2(n_533),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_607),
.A2(n_571),
.B1(n_555),
.B2(n_551),
.Y(n_620)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_608),
.Y(n_633)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_563),
.A2(n_522),
.B(n_517),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_576),
.B(n_527),
.C(n_534),
.Y(n_610)
);

MAJIxp5_ASAP7_75t_L g621 ( 
.A(n_610),
.B(n_614),
.C(n_552),
.Y(n_621)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_558),
.Y(n_611)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_611),
.Y(n_624)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_557),
.Y(n_612)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_612),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_556),
.B(n_527),
.Y(n_613)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_613),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g614 ( 
.A(n_570),
.B(n_516),
.C(n_519),
.Y(n_614)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_618),
.B(n_586),
.Y(n_645)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_620),
.B(n_637),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_621),
.B(n_622),
.Y(n_660)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_597),
.B(n_570),
.C(n_565),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_599),
.Y(n_623)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_623),
.Y(n_646)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_628),
.A2(n_636),
.B1(n_640),
.B2(n_592),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_596),
.B(n_562),
.C(n_574),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_629),
.B(n_631),
.Y(n_662)
);

MAJIxp5_ASAP7_75t_L g631 ( 
.A(n_588),
.B(n_554),
.C(n_580),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_613),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_632),
.B(n_635),
.Y(n_650)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_604),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_590),
.A2(n_553),
.B1(n_582),
.B2(n_567),
.Y(n_636)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_591),
.B(n_580),
.C(n_567),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g647 ( 
.A(n_638),
.B(n_639),
.C(n_589),
.Y(n_647)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_594),
.B(n_561),
.C(n_573),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_593),
.Y(n_640)
);

CKINVDCx16_ASAP7_75t_R g641 ( 
.A(n_618),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_641),
.B(n_642),
.Y(n_666)
);

OAI21xp5_ASAP7_75t_L g642 ( 
.A1(n_633),
.A2(n_608),
.B(n_550),
.Y(n_642)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_643),
.Y(n_674)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_633),
.A2(n_587),
.B(n_610),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_L g673 ( 
.A1(n_644),
.A2(n_548),
.B1(n_544),
.B2(n_541),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g678 ( 
.A1(n_645),
.A2(n_544),
.B(n_541),
.Y(n_678)
);

XNOR2xp5_ASAP7_75t_L g675 ( 
.A(n_647),
.B(n_649),
.Y(n_675)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_634),
.B(n_602),
.Y(n_649)
);

XOR2xp5_ASAP7_75t_L g651 ( 
.A(n_634),
.B(n_598),
.Y(n_651)
);

XOR2xp5_ASAP7_75t_L g667 ( 
.A(n_651),
.B(n_657),
.Y(n_667)
);

MAJIxp5_ASAP7_75t_L g652 ( 
.A(n_627),
.B(n_619),
.C(n_622),
.Y(n_652)
);

MAJIxp5_ASAP7_75t_L g663 ( 
.A(n_652),
.B(n_653),
.C(n_654),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g653 ( 
.A(n_627),
.B(n_614),
.C(n_585),
.Y(n_653)
);

MAJIxp5_ASAP7_75t_L g654 ( 
.A(n_619),
.B(n_585),
.C(n_607),
.Y(n_654)
);

XNOR2xp5_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_629),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_655),
.B(n_656),
.Y(n_677)
);

XNOR2xp5_ASAP7_75t_L g656 ( 
.A(n_637),
.B(n_639),
.Y(n_656)
);

XOR2xp5_ASAP7_75t_L g657 ( 
.A(n_638),
.B(n_606),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g658 ( 
.A(n_631),
.B(n_603),
.C(n_609),
.Y(n_658)
);

MAJIxp5_ASAP7_75t_L g665 ( 
.A(n_658),
.B(n_659),
.C(n_623),
.Y(n_665)
);

MAJIxp5_ASAP7_75t_L g659 ( 
.A(n_615),
.B(n_603),
.C(n_595),
.Y(n_659)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_620),
.B(n_561),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g671 ( 
.A(n_661),
.B(n_601),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g664 ( 
.A1(n_645),
.A2(n_617),
.B1(n_626),
.B2(n_615),
.Y(n_664)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_664),
.A2(n_668),
.B1(n_670),
.B2(n_651),
.Y(n_693)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_665),
.Y(n_682)
);

AOI21x1_ASAP7_75t_L g668 ( 
.A1(n_650),
.A2(n_625),
.B(n_624),
.Y(n_668)
);

AOI21xp5_ASAP7_75t_L g669 ( 
.A1(n_659),
.A2(n_616),
.B(n_636),
.Y(n_669)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_669),
.A2(n_666),
.B(n_678),
.Y(n_694)
);

AOI22xp5_ASAP7_75t_L g670 ( 
.A1(n_661),
.A2(n_628),
.B1(n_630),
.B2(n_654),
.Y(n_670)
);

XNOR2xp5_ASAP7_75t_L g684 ( 
.A(n_671),
.B(n_658),
.Y(n_684)
);

MAJIxp5_ASAP7_75t_L g672 ( 
.A(n_652),
.B(n_605),
.C(n_548),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_672),
.B(n_679),
.Y(n_686)
);

AOI22xp5_ASAP7_75t_L g688 ( 
.A1(n_673),
.A2(n_676),
.B1(n_678),
.B2(n_671),
.Y(n_688)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_646),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g679 ( 
.A(n_653),
.B(n_519),
.C(n_390),
.Y(n_679)
);

MAJIxp5_ASAP7_75t_L g680 ( 
.A(n_655),
.B(n_396),
.C(n_435),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_680),
.B(n_649),
.Y(n_691)
);

XOR2xp5_ASAP7_75t_L g681 ( 
.A(n_679),
.B(n_656),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_681),
.B(n_683),
.Y(n_697)
);

XOR2xp5_ASAP7_75t_L g683 ( 
.A(n_665),
.B(n_657),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g695 ( 
.A(n_684),
.B(n_691),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_663),
.B(n_660),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_685),
.B(n_687),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_663),
.B(n_672),
.Y(n_687)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_688),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_677),
.B(n_647),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_SL g701 ( 
.A(n_689),
.B(n_680),
.Y(n_701)
);

MAJIxp5_ASAP7_75t_L g690 ( 
.A(n_675),
.B(n_667),
.C(n_662),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_690),
.B(n_693),
.Y(n_696)
);

XOR2xp5_ASAP7_75t_L g692 ( 
.A(n_667),
.B(n_648),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_692),
.B(n_648),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g699 ( 
.A1(n_694),
.A2(n_669),
.B(n_664),
.Y(n_699)
);

NOR2x1_ASAP7_75t_L g698 ( 
.A(n_684),
.B(n_675),
.Y(n_698)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_698),
.A2(n_702),
.B(n_696),
.Y(n_705)
);

MAJx2_ASAP7_75t_L g708 ( 
.A(n_699),
.B(n_690),
.C(n_692),
.Y(n_708)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_701),
.Y(n_710)
);

OAI21xp5_ASAP7_75t_SL g702 ( 
.A1(n_682),
.A2(n_670),
.B(n_674),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_704),
.B(n_398),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_705),
.B(n_706),
.Y(n_712)
);

XNOR2xp5_ASAP7_75t_L g706 ( 
.A(n_695),
.B(n_681),
.Y(n_706)
);

OAI22xp5_ASAP7_75t_SL g707 ( 
.A1(n_700),
.A2(n_694),
.B1(n_686),
.B2(n_683),
.Y(n_707)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_707),
.B(n_696),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_708),
.B(n_709),
.Y(n_714)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_703),
.A2(n_435),
.B(n_314),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_SL g715 ( 
.A(n_711),
.B(n_697),
.Y(n_715)
);

OAI21xp5_ASAP7_75t_L g716 ( 
.A1(n_713),
.A2(n_715),
.B(n_695),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g718 ( 
.A1(n_716),
.A2(n_717),
.B(n_712),
.Y(n_718)
);

MAJIxp5_ASAP7_75t_L g717 ( 
.A(n_714),
.B(n_710),
.C(n_708),
.Y(n_717)
);

MAJIxp5_ASAP7_75t_L g719 ( 
.A(n_718),
.B(n_365),
.C(n_344),
.Y(n_719)
);

OAI321xp33_ASAP7_75t_L g720 ( 
.A1(n_719),
.A2(n_398),
.A3(n_360),
.B1(n_334),
.B2(n_314),
.C(n_344),
.Y(n_720)
);

MAJIxp5_ASAP7_75t_L g721 ( 
.A(n_720),
.B(n_360),
.C(n_398),
.Y(n_721)
);

AOI21xp5_ASAP7_75t_L g722 ( 
.A1(n_721),
.A2(n_398),
.B(n_334),
.Y(n_722)
);


endmodule