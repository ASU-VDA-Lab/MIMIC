module real_jpeg_19210_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_243;
wire n_197;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_188;
wire n_139;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_262;
wire n_148;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_70;
wire n_80;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_277;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_52;
wire n_58;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_0),
.A2(n_46),
.B1(n_47),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_0),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_27),
.B1(n_30),
.B2(n_54),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_1),
.A2(n_46),
.B1(n_47),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_1),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_1),
.A2(n_27),
.B1(n_30),
.B2(n_52),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_52),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_2),
.A2(n_73),
.B1(n_79),
.B2(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_2),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_97),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_97),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_2),
.A2(n_27),
.B1(n_30),
.B2(n_97),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_3),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_4),
.A2(n_27),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_4),
.A2(n_38),
.B1(n_73),
.B2(n_79),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_38),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_4),
.A2(n_38),
.B1(n_46),
.B2(n_47),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_5),
.A2(n_73),
.B1(n_79),
.B2(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_5),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_5),
.A2(n_46),
.B1(n_47),
.B2(n_152),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_5),
.A2(n_27),
.B1(n_30),
.B2(n_152),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_5),
.A2(n_33),
.B1(n_34),
.B2(n_152),
.Y(n_204)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_6),
.Y(n_61)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_6),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_88),
.B(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_6),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_29),
.B2(n_30),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_7),
.A2(n_29),
.B1(n_33),
.B2(n_34),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_7),
.A2(n_29),
.B1(n_73),
.B2(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_7),
.A2(n_29),
.B1(n_46),
.B2(n_47),
.Y(n_125)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_9),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_9),
.A2(n_14),
.B(n_34),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_9),
.A2(n_27),
.B1(n_30),
.B2(n_150),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_9),
.A2(n_60),
.B1(n_204),
.B2(n_208),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_9),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_9),
.B(n_46),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_9),
.A2(n_46),
.B(n_231),
.Y(n_235)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_11),
.A2(n_73),
.B1(n_79),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_11),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_11),
.A2(n_46),
.B1(n_47),
.B2(n_130),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_11),
.A2(n_33),
.B1(n_34),
.B2(n_130),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_11),
.A2(n_27),
.B1(n_30),
.B2(n_130),
.Y(n_222)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx13_ASAP7_75t_L g72 ( 
.A(n_13),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_13),
.A2(n_46),
.B1(n_47),
.B2(n_72),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_14),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_32)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

A2O1A1Ixp33_ASAP7_75t_L g40 ( 
.A1(n_14),
.A2(n_30),
.B(n_32),
.C(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_14),
.B(n_30),
.Y(n_41)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_15),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_133),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_132),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_106),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_20),
.B(n_106),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_84),
.B2(n_105),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_56),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_42),
.B(n_55),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_24),
.B(n_42),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_36),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_25),
.A2(n_40),
.B(n_238),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_31),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_26),
.Y(n_143)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_27),
.A2(n_30),
.B1(n_44),
.B2(n_50),
.Y(n_49)
);

A2O1A1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_27),
.A2(n_35),
.B(n_150),
.C(n_196),
.Y(n_195)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_27),
.B(n_44),
.Y(n_232)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_30),
.A2(n_47),
.A3(n_50),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_31),
.B(n_37),
.Y(n_66)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_32),
.A2(n_40),
.B1(n_65),
.B2(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_32),
.A2(n_36),
.B(n_93),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_32),
.A2(n_40),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_32),
.B(n_150),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_32),
.A2(n_40),
.B1(n_200),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_32),
.A2(n_40),
.B1(n_222),
.B2(n_238),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_33),
.B(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_39),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_65),
.B(n_66),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_40),
.A2(n_66),
.B(n_143),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_53),
.Y(n_42)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_43),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_43),
.A2(n_49),
.B1(n_146),
.B2(n_147),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_43),
.A2(n_49),
.B1(n_146),
.B2(n_176),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_43),
.A2(n_49),
.B1(n_176),
.B2(n_235),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B(n_48),
.C(n_49),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_46),
.Y(n_48)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_44),
.Y(n_50)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_46),
.B(n_72),
.Y(n_156)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_47),
.A2(n_75),
.B1(n_149),
.B2(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_51),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_49),
.B(n_104),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_49),
.B(n_125),
.Y(n_167)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_49),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_67),
.B2(n_68),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_59),
.A2(n_69),
.B1(n_82),
.B2(n_83),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_59),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_64),
.B1(n_83),
.B2(n_111),
.Y(n_110)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_61),
.B(n_62),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_60),
.A2(n_119),
.B1(n_122),
.B2(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_60),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_60),
.A2(n_122),
.B1(n_190),
.B2(n_204),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_60),
.A2(n_90),
.B(n_192),
.Y(n_223)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_61),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_61),
.B(n_150),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_63),
.B(n_91),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_121),
.B(n_188),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_64),
.Y(n_111)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_69),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_77),
.B(n_80),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_70),
.A2(n_96),
.B(n_98),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_96),
.B1(n_129),
.B2(n_131),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_70),
.A2(n_129),
.B1(n_131),
.B2(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_71),
.A2(n_76),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_75),
.C(n_76),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_73),
.Y(n_75)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

HAxp5_ASAP7_75t_SL g149 ( 
.A(n_73),
.B(n_150),
.CON(n_149),
.SN(n_149)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_76),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_76),
.B(n_78),
.Y(n_98)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_84),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_94),
.C(n_99),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_92),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_86),
.B(n_92),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_90),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_89),
.B(n_122),
.Y(n_121)
);

INVx4_ASAP7_75t_L g208 ( 
.A(n_91),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_94),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_102),
.A2(n_124),
.B(n_126),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_102),
.A2(n_166),
.B(n_167),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.C(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_107),
.A2(n_108),
.B1(n_110),
.B2(n_281),
.Y(n_280)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_110),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_112),
.B(n_280),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_123),
.C(n_127),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_113),
.A2(n_114),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_115),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_123),
.A2(n_127),
.B1(n_128),
.B2(n_273),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_123),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_125),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_131),
.B(n_150),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_277),
.B(n_282),
.Y(n_133)
);

O2A1O1Ixp33_ASAP7_75t_SL g134 ( 
.A1(n_135),
.A2(n_180),
.B(n_262),
.C(n_276),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_169),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_136),
.B(n_169),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_138),
.B1(n_153),
.B2(n_168),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_139),
.B(n_140),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_139),
.B(n_140),
.C(n_168),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_144),
.C(n_148),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_141),
.A2(n_142),
.B1(n_144),
.B2(n_145),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_SL g170 ( 
.A(n_148),
.B(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_151),
.Y(n_163)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_153),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_160),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_154),
.B(n_161),
.C(n_165),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_157),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_164),
.B2(n_165),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.C(n_174),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_170),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_172),
.A2(n_173),
.B1(n_174),
.B2(n_259),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_174),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.C(n_178),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_175),
.B(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_177),
.A2(n_178),
.B1(n_179),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_177),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_261),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_255),
.B(n_260),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_183),
.A2(n_243),
.B(n_254),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_225),
.B(n_242),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_213),
.B(n_224),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_201),
.B(n_212),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_193),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_187),
.B(n_193),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_197),
.B2(n_198),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_195),
.B(n_197),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_206),
.B(n_211),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_205),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_203),
.B(n_205),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_209),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_214),
.B(n_215),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_223),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_217),
.A2(n_218),
.B1(n_220),
.B2(n_221),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_217),
.B(n_221),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_240),
.B2(n_241),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_229),
.B(n_230),
.Y(n_252)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_252),
.C(n_253),
.Y(n_256)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_256),
.B(n_257),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_263),
.B(n_264),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_274),
.B2(n_275),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_270),
.C(n_275),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);


endmodule