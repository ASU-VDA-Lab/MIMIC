module fake_jpeg_29179_n_216 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_216);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_216;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_122;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_12),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_1),
.B(n_5),
.Y(n_35)
);

INVx11_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_37),
.Y(n_84)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_38),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_2),
.B(n_4),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_40),
.B(n_26),
.Y(n_70)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_41),
.Y(n_81)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_42),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_30),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_48),
.Y(n_69)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_2),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

AND2x2_ASAP7_75t_SL g51 ( 
.A(n_27),
.B(n_5),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_53),
.Y(n_87)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_52),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_13),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_14),
.B(n_5),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_60),
.Y(n_88)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_17),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_58),
.A2(n_64),
.B1(n_20),
.B2(n_28),
.Y(n_71)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_61),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_15),
.B(n_8),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_62),
.B(n_65),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_19),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_64)
);

CKINVDCx12_ASAP7_75t_R g65 ( 
.A(n_22),
.Y(n_65)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_18),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_67),
.B(n_20),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_78),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_71),
.A2(n_102),
.B1(n_105),
.B2(n_98),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_74),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_62),
.B(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_31),
.B1(n_22),
.B2(n_28),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_79),
.A2(n_97),
.B1(n_99),
.B2(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_56),
.B(n_26),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_80),
.B(n_85),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_55),
.B(n_23),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_82),
.B(n_92),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_15),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_32),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_86),
.B(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_21),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_81),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_49),
.A2(n_21),
.B1(n_24),
.B2(n_31),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_95),
.A2(n_103),
.B1(n_72),
.B2(n_68),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_42),
.A2(n_22),
.B1(n_31),
.B2(n_24),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_46),
.A2(n_31),
.B1(n_10),
.B2(n_12),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_9),
.B1(n_12),
.B2(n_64),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_37),
.A2(n_9),
.B1(n_61),
.B2(n_52),
.Y(n_104)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_107),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_54),
.C(n_63),
.Y(n_109)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_109),
.B(n_130),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_110),
.A2(n_111),
.B1(n_123),
.B2(n_128),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_102),
.A2(n_104),
.B1(n_79),
.B2(n_97),
.Y(n_111)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_83),
.Y(n_112)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_112),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_93),
.A2(n_39),
.B1(n_47),
.B2(n_41),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g114 ( 
.A(n_77),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_124),
.Y(n_136)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_84),
.Y(n_118)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_118),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g153 ( 
.A(n_119),
.B(n_122),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_127),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_73),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_90),
.A2(n_106),
.B1(n_99),
.B2(n_91),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_69),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_125),
.B(n_126),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_75),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_93),
.A2(n_91),
.B1(n_77),
.B2(n_103),
.Y(n_128)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g130 ( 
.A(n_75),
.B(n_100),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_72),
.A2(n_68),
.B1(n_83),
.B2(n_98),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_134),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_105),
.B(n_81),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_96),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_96),
.B(n_70),
.Y(n_134)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_130),
.B(n_115),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_140),
.B(n_142),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_119),
.B(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_132),
.B1(n_120),
.B2(n_107),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_109),
.B(n_120),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_146),
.B(n_117),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_133),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_122),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_116),
.B(n_125),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_160),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_140),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_159),
.B(n_166),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_152),
.A2(n_111),
.B1(n_122),
.B2(n_131),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_171),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_138),
.Y(n_162)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_162),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_148),
.B(n_133),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_137),
.B(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_167),
.B(n_168),
.Y(n_173)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_138),
.Y(n_169)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_169),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_144),
.A2(n_152),
.B1(n_151),
.B2(n_156),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_170),
.A2(n_139),
.B(n_141),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_137),
.B(n_124),
.Y(n_171)
);

NAND3xp33_ASAP7_75t_L g172 ( 
.A(n_142),
.B(n_155),
.C(n_150),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_172),
.B(n_153),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_162),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_180),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_SL g187 ( 
.A(n_178),
.B(n_164),
.C(n_163),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_164),
.B(n_146),
.Y(n_180)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_169),
.Y(n_182)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_182),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_170),
.A2(n_154),
.B(n_156),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_183),
.A2(n_184),
.B(n_168),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_175),
.A2(n_143),
.B1(n_160),
.B2(n_157),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_185),
.A2(n_145),
.B1(n_190),
.B2(n_182),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_181),
.B(n_159),
.C(n_166),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_186),
.B(n_187),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_SL g199 ( 
.A(n_188),
.B(n_189),
.C(n_136),
.Y(n_199)
);

MAJx2_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_163),
.C(n_153),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_181),
.B(n_136),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_192),
.B(n_193),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_176),
.B(n_165),
.C(n_147),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_194),
.A2(n_179),
.B1(n_147),
.B2(n_143),
.Y(n_205)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_197),
.B(n_200),
.Y(n_203)
);

AOI321xp33_ASAP7_75t_L g198 ( 
.A1(n_187),
.A2(n_173),
.A3(n_183),
.B1(n_184),
.B2(n_174),
.C(n_176),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_198),
.A2(n_199),
.B(n_186),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_193),
.B(n_179),
.Y(n_200)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_201),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_196),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_202),
.A2(n_204),
.B(n_205),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_199),
.A2(n_188),
.B1(n_192),
.B2(n_175),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_202),
.A2(n_198),
.B(n_197),
.Y(n_208)
);

AO21x1_ASAP7_75t_L g210 ( 
.A1(n_208),
.A2(n_189),
.B(n_157),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_204),
.B(n_195),
.C(n_203),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_209),
.B(n_149),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_210),
.B(n_211),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_207),
.A2(n_149),
.B(n_126),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_212),
.B(n_206),
.C(n_118),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_214),
.B(n_112),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_215),
.A2(n_213),
.B(n_114),
.Y(n_216)
);


endmodule