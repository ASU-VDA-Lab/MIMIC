module fake_jpeg_24334_n_318 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_318);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_318;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx2_ASAP7_75t_SL g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx11_ASAP7_75t_SL g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_5),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_38),
.B(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_19),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_43),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_0),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_0),
.Y(n_52)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_44),
.B(n_45),
.Y(n_47)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_39),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_48),
.B(n_59),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_27),
.B1(n_20),
.B2(n_33),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_50),
.A2(n_55),
.B1(n_57),
.B2(n_61),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_18),
.C(n_17),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_51),
.B(n_66),
.C(n_69),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_52),
.B(n_64),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_39),
.A2(n_21),
.B1(n_20),
.B2(n_34),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_44),
.A2(n_21),
.B1(n_30),
.B2(n_19),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_21),
.B1(n_33),
.B2(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_45),
.B1(n_40),
.B2(n_37),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_62),
.B(n_63),
.Y(n_90)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_33),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_65),
.B(n_43),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_45),
.A2(n_29),
.B1(n_35),
.B2(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_40),
.A2(n_29),
.B1(n_35),
.B2(n_25),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

INVx5_ASAP7_75t_L g94 ( 
.A(n_70),
.Y(n_94)
);

AO22x2_ASAP7_75t_L g71 ( 
.A1(n_50),
.A2(n_43),
.B1(n_36),
.B2(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_71),
.A2(n_92),
.B1(n_39),
.B2(n_60),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx8_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_70),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

NAND2x1_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_22),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_SL g111 ( 
.A(n_77),
.B(n_84),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_52),
.B(n_38),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_79),
.B(n_82),
.Y(n_110)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_80),
.B(n_81),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_38),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

OR2x2_ASAP7_75t_SL g84 ( 
.A(n_51),
.B(n_23),
.Y(n_84)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_86),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_47),
.B(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_87),
.B(n_98),
.Y(n_137)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_89),
.Y(n_126)
);

AOI21xp33_ASAP7_75t_L g91 ( 
.A1(n_68),
.A2(n_18),
.B(n_23),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_91),
.B(n_22),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_40),
.B1(n_25),
.B2(n_37),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_96),
.A2(n_36),
.B1(n_30),
.B2(n_24),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_66),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_54),
.B(n_26),
.Y(n_101)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_101),
.B(n_103),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_61),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_56),
.B(n_1),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_105),
.B(n_23),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_54),
.B(n_26),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_39),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_69),
.B(n_31),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_107),
.B(n_28),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_60),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_118),
.Y(n_141)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_108),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_115),
.B(n_119),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_123),
.B1(n_71),
.B2(n_74),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_39),
.Y(n_118)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_78),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_121),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_65),
.B1(n_37),
.B2(n_41),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_104),
.B(n_41),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_127),
.Y(n_146)
);

CKINVDCx12_ASAP7_75t_R g129 ( 
.A(n_72),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_129),
.Y(n_143)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_132),
.B(n_86),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_100),
.A2(n_28),
.B1(n_32),
.B2(n_31),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_133),
.B(n_22),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_136),
.B(n_105),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_139),
.A2(n_125),
.B1(n_90),
.B2(n_96),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_124),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_150),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_118),
.B(n_85),
.C(n_71),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_157),
.C(n_120),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_122),
.B(n_109),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_153),
.Y(n_171)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_145),
.B(n_147),
.Y(n_189)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_123),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_117),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_127),
.B(n_88),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_151),
.B(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_117),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g153 ( 
.A(n_136),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_116),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_111),
.A2(n_102),
.B(n_100),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_156),
.A2(n_161),
.B(n_163),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_88),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_110),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_158),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_126),
.Y(n_159)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_160),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_131),
.A2(n_102),
.B(n_77),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_115),
.B(n_75),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_164),
.B(n_165),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_131),
.A2(n_84),
.B(n_98),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_32),
.B(n_22),
.Y(n_190)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_126),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_168),
.Y(n_194)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_112),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_169),
.B(n_26),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g170 ( 
.A1(n_139),
.A2(n_71),
.B1(n_113),
.B2(n_125),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_170),
.A2(n_179),
.B1(n_188),
.B2(n_197),
.Y(n_204)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_138),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_176),
.B(n_183),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_113),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_177),
.B(n_180),
.C(n_186),
.Y(n_214)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_150),
.Y(n_181)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_181),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_97),
.Y(n_182)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_182),
.Y(n_220)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_154),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_159),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_184),
.B(n_187),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_80),
.B(n_132),
.Y(n_185)
);

A2O1A1Ixp33_ASAP7_75t_SL g227 ( 
.A1(n_185),
.A2(n_141),
.B(n_30),
.C(n_24),
.Y(n_227)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_147),
.A2(n_119),
.B1(n_83),
.B2(n_93),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_190),
.B(n_195),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_120),
.C(n_135),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_199),
.Y(n_226)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_166),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_196),
.B(n_163),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_155),
.A2(n_89),
.B1(n_94),
.B2(n_130),
.Y(n_197)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_141),
.B(n_30),
.C(n_24),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_152),
.B(n_128),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_144),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_191),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_202),
.B(n_221),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_200),
.B(n_143),
.Y(n_205)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_170),
.A2(n_162),
.B1(n_165),
.B2(n_151),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_216),
.B1(n_185),
.B2(n_193),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_207),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_200),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_209),
.Y(n_238)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_210),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_183),
.B(n_143),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_211),
.B(n_212),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_195),
.B1(n_162),
.B2(n_175),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_217),
.B(n_218),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_184),
.B(n_94),
.Y(n_218)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_189),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_222),
.B(n_225),
.Y(n_236)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_188),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_223),
.A2(n_224),
.B1(n_227),
.B2(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_198),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_171),
.B(n_157),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_186),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_228),
.B(n_235),
.Y(n_250)
);

BUFx24_ASAP7_75t_SL g229 ( 
.A(n_221),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_229),
.B(n_10),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_192),
.C(n_180),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_230),
.B(n_231),
.C(n_232),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_174),
.C(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_174),
.C(n_182),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_207),
.B(n_172),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_242),
.B1(n_224),
.B2(n_215),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_197),
.B1(n_187),
.B2(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_172),
.C(n_199),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_245),
.C(n_248),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_204),
.A2(n_198),
.B1(n_190),
.B2(n_173),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_173),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_244),
.B(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_130),
.C(n_36),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_247),
.B(n_213),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_73),
.C(n_24),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_251),
.B(n_7),
.C(n_15),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_253),
.B(n_261),
.Y(n_269)
);

OAI22x1_ASAP7_75t_SL g254 ( 
.A1(n_234),
.A2(n_216),
.B1(n_227),
.B2(n_204),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_254),
.A2(n_245),
.B1(n_244),
.B2(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_238),
.B(n_209),
.Y(n_255)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_255),
.Y(n_271)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_208),
.Y(n_257)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_257),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_239),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_246),
.A2(n_212),
.B(n_222),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_259),
.A2(n_267),
.B(n_10),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_230),
.B(n_206),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_262),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_241),
.A2(n_227),
.B1(n_219),
.B2(n_203),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_228),
.B(n_227),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_240),
.A2(n_227),
.B1(n_243),
.B2(n_249),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_263),
.B(n_264),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_202),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_270),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_254),
.A2(n_231),
.B1(n_236),
.B2(n_203),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_272),
.A2(n_279),
.B1(n_269),
.B2(n_268),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_26),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_275),
.B(n_278),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_8),
.B(n_15),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g291 ( 
.A1(n_276),
.A2(n_11),
.B1(n_3),
.B2(n_4),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_272),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_1),
.C(n_2),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_280),
.B(n_266),
.C(n_265),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_282),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_271),
.B(n_263),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_283),
.B(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_266),
.C(n_250),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_287),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_281),
.B(n_251),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_273),
.Y(n_299)
);

BUFx4f_ASAP7_75t_SL g290 ( 
.A(n_274),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_290),
.A2(n_292),
.B(n_278),
.Y(n_294)
);

OAI321xp33_ASAP7_75t_L g297 ( 
.A1(n_291),
.A2(n_12),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_7),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_250),
.C(n_3),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_11),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_293),
.A2(n_276),
.B(n_275),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_294),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_296),
.B(n_302),
.Y(n_305)
);

AOI222xp33_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_291),
.B1(n_6),
.B2(n_7),
.C1(n_13),
.C2(n_14),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_301),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_290),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_289),
.A2(n_4),
.B(n_6),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_295),
.Y(n_304)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_304),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_290),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_307),
.A2(n_308),
.B(n_293),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_SL g308 ( 
.A(n_298),
.B(n_289),
.Y(n_308)
);

OAI221xp5_ASAP7_75t_L g312 ( 
.A1(n_309),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.C(n_1),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_312),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g313 ( 
.A1(n_306),
.A2(n_1),
.A3(n_13),
.B1(n_14),
.B2(n_16),
.C1(n_285),
.C2(n_307),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_313),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_310),
.C(n_303),
.Y(n_316)
);

OAI21xp5_ASAP7_75t_SL g317 ( 
.A1(n_316),
.A2(n_314),
.B(n_305),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_317),
.B(n_285),
.Y(n_318)
);


endmodule