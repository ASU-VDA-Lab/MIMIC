module fake_ariane_2453_n_1558 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_49, n_20, n_283, n_50, n_187, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_251, n_116, n_39, n_155, n_127, n_1558);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1558;

wire n_913;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_1495;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_1548;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_1253;
wire n_762;
wire n_1468;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_1506;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1467;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1489;
wire n_1218;
wire n_321;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_845;
wire n_888;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_1552;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1482;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_318;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_1067;
wire n_968;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1551;
wire n_1285;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1003;
wire n_701;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_323;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_1477;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_1479;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1474;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_201),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_96),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_15),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_142),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_162),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_50),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_184),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_166),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_109),
.Y(n_324)
);

CKINVDCx14_ASAP7_75t_R g325 ( 
.A(n_227),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_250),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_83),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_246),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_173),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_77),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_31),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_50),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_218),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_8),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_145),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_87),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_72),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_304),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_186),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_279),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_16),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_110),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_197),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_161),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_222),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_232),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_298),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_262),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_309),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_285),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_71),
.Y(n_351)
);

CKINVDCx14_ASAP7_75t_R g352 ( 
.A(n_170),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_18),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_245),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_56),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_69),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_263),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_177),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g359 ( 
.A(n_265),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_293),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_43),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_176),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_93),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_206),
.Y(n_364)
);

BUFx3_ASAP7_75t_L g365 ( 
.A(n_284),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_69),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_155),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_137),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_103),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_178),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_39),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_175),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_0),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_68),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_299),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_13),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_169),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_138),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_18),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_124),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_241),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_278),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_151),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_216),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_168),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_300),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_115),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_182),
.Y(n_388)
);

BUFx6f_ASAP7_75t_L g389 ( 
.A(n_266),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_223),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_140),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_65),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g393 ( 
.A(n_226),
.Y(n_393)
);

INVx1_ASAP7_75t_SL g394 ( 
.A(n_205),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_204),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_267),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g397 ( 
.A(n_89),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_153),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_131),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_272),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_43),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_234),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_106),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_9),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_58),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_314),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_82),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_66),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_217),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_47),
.Y(n_410)
);

INVx2_ASAP7_75t_SL g411 ( 
.A(n_125),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_230),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_59),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_294),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_31),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_53),
.Y(n_416)
);

CKINVDCx16_ASAP7_75t_R g417 ( 
.A(n_315),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_133),
.Y(n_418)
);

BUFx5_ASAP7_75t_L g419 ( 
.A(n_286),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g420 ( 
.A(n_191),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_307),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_62),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_296),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_104),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_192),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_52),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_199),
.Y(n_427)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_248),
.Y(n_428)
);

CKINVDCx20_ASAP7_75t_R g429 ( 
.A(n_220),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_67),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_188),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_268),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_114),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_256),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_221),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_158),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g437 ( 
.A(n_303),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_1),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_163),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_144),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_88),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_187),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_123),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_264),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_258),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_75),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_34),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_73),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_134),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_49),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_16),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_277),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_71),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_14),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_135),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_126),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_282),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_85),
.Y(n_458)
);

BUFx10_ASAP7_75t_L g459 ( 
.A(n_160),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_39),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_25),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_308),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_310),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_48),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_107),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_274),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_157),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_261),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_49),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_291),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_76),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_128),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_129),
.Y(n_473)
);

INVx2_ASAP7_75t_SL g474 ( 
.A(n_154),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_23),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_276),
.Y(n_476)
);

INVx1_ASAP7_75t_SL g477 ( 
.A(n_228),
.Y(n_477)
);

BUFx10_ASAP7_75t_L g478 ( 
.A(n_214),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_180),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_254),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_78),
.Y(n_481)
);

INVx2_ASAP7_75t_SL g482 ( 
.A(n_312),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_219),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_57),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_260),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_301),
.Y(n_486)
);

BUFx10_ASAP7_75t_L g487 ( 
.A(n_95),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_313),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_33),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_14),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_64),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_311),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_46),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_55),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_9),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_122),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_30),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_302),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_167),
.Y(n_499)
);

INVx1_ASAP7_75t_SL g500 ( 
.A(n_239),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_1),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_136),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_100),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_224),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_141),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_146),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_297),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_229),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_288),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_21),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_159),
.Y(n_511)
);

BUFx10_ASAP7_75t_L g512 ( 
.A(n_77),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_209),
.Y(n_513)
);

BUFx10_ASAP7_75t_L g514 ( 
.A(n_99),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_47),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g516 ( 
.A(n_98),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_195),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_171),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_30),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_76),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_61),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_152),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_198),
.Y(n_523)
);

BUFx2_ASAP7_75t_L g524 ( 
.A(n_189),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_305),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_275),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_287),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_94),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_174),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_225),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_28),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_91),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_295),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_306),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_165),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_25),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_82),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_231),
.Y(n_538)
);

BUFx3_ASAP7_75t_L g539 ( 
.A(n_280),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_28),
.Y(n_540)
);

CKINVDCx16_ASAP7_75t_R g541 ( 
.A(n_194),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_271),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_139),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_283),
.Y(n_544)
);

CKINVDCx16_ASAP7_75t_R g545 ( 
.A(n_270),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_90),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_38),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_92),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_149),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_46),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_86),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_45),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g553 ( 
.A(n_381),
.B(n_0),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_318),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_332),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_512),
.B(n_2),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g557 ( 
.A(n_462),
.B(n_2),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_470),
.B(n_3),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_398),
.Y(n_559)
);

AND2x4_ASAP7_75t_L g560 ( 
.A(n_392),
.B(n_3),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g561 ( 
.A(n_321),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_524),
.Y(n_562)
);

AND2x4_ASAP7_75t_L g563 ( 
.A(n_392),
.B(n_494),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_332),
.Y(n_564)
);

BUFx3_ASAP7_75t_L g565 ( 
.A(n_398),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_494),
.B(n_4),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_399),
.B(n_4),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_521),
.B(n_5),
.Y(n_568)
);

BUFx8_ASAP7_75t_SL g569 ( 
.A(n_408),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_332),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_332),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_430),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_430),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_508),
.B(n_5),
.Y(n_574)
);

BUFx6f_ASAP7_75t_L g575 ( 
.A(n_326),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_398),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_393),
.B(n_6),
.Y(n_577)
);

AND2x6_ASAP7_75t_L g578 ( 
.A(n_372),
.B(n_97),
.Y(n_578)
);

INVx5_ASAP7_75t_L g579 ( 
.A(n_459),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_430),
.Y(n_580)
);

INVx5_ASAP7_75t_L g581 ( 
.A(n_459),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g582 ( 
.A(n_512),
.B(n_6),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_326),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_521),
.B(n_7),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_430),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_365),
.B(n_539),
.Y(n_586)
);

BUFx3_ASAP7_75t_L g587 ( 
.A(n_459),
.Y(n_587)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_326),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_478),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_327),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_326),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_478),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_317),
.B(n_7),
.Y(n_593)
);

INVx5_ASAP7_75t_L g594 ( 
.A(n_478),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_324),
.B(n_8),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_342),
.B(n_10),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_365),
.Y(n_597)
);

INVx5_ASAP7_75t_L g598 ( 
.A(n_487),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_343),
.B(n_348),
.Y(n_599)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_340),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_512),
.B(n_10),
.Y(n_601)
);

INVx4_ASAP7_75t_L g602 ( 
.A(n_340),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_323),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_325),
.B(n_11),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_323),
.Y(n_605)
);

BUFx6f_ASAP7_75t_L g606 ( 
.A(n_340),
.Y(n_606)
);

HB1xp67_ASAP7_75t_L g607 ( 
.A(n_330),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_349),
.B(n_11),
.Y(n_608)
);

CKINVDCx6p67_ASAP7_75t_R g609 ( 
.A(n_487),
.Y(n_609)
);

INVx5_ASAP7_75t_L g610 ( 
.A(n_487),
.Y(n_610)
);

BUFx3_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

INVx5_ASAP7_75t_L g612 ( 
.A(n_514),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_350),
.B(n_12),
.Y(n_613)
);

INVx5_ASAP7_75t_L g614 ( 
.A(n_514),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_363),
.B(n_12),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_539),
.B(n_13),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_546),
.B(n_15),
.Y(n_617)
);

AND2x4_ASAP7_75t_L g618 ( 
.A(n_546),
.B(n_17),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_364),
.B(n_17),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_368),
.B(n_19),
.Y(n_620)
);

BUFx12f_ASAP7_75t_L g621 ( 
.A(n_331),
.Y(n_621)
);

HB1xp67_ASAP7_75t_L g622 ( 
.A(n_337),
.Y(n_622)
);

INVx4_ASAP7_75t_L g623 ( 
.A(n_340),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_370),
.B(n_19),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_341),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_328),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_334),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_389),
.Y(n_628)
);

AND2x4_ASAP7_75t_L g629 ( 
.A(n_336),
.B(n_361),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_328),
.Y(n_630)
);

INVx5_ASAP7_75t_L g631 ( 
.A(n_389),
.Y(n_631)
);

BUFx6f_ASAP7_75t_L g632 ( 
.A(n_389),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_380),
.B(n_20),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_374),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_386),
.B(n_20),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_435),
.Y(n_636)
);

BUFx6f_ASAP7_75t_L g637 ( 
.A(n_389),
.Y(n_637)
);

BUFx6f_ASAP7_75t_L g638 ( 
.A(n_372),
.Y(n_638)
);

BUFx6f_ASAP7_75t_L g639 ( 
.A(n_435),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_388),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_325),
.B(n_21),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_465),
.Y(n_642)
);

INVx2_ASAP7_75t_L g643 ( 
.A(n_410),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_465),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_499),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_400),
.B(n_22),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_402),
.B(n_22),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_417),
.Y(n_648)
);

INVx4_ASAP7_75t_L g649 ( 
.A(n_319),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_422),
.Y(n_650)
);

HB1xp67_ASAP7_75t_L g651 ( 
.A(n_351),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_418),
.B(n_23),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_425),
.B(n_24),
.Y(n_653)
);

BUFx6f_ASAP7_75t_L g654 ( 
.A(n_499),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_447),
.B(n_24),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_431),
.B(n_26),
.Y(n_656)
);

INVxp67_ASAP7_75t_L g657 ( 
.A(n_469),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_479),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_L g659 ( 
.A(n_433),
.B(n_26),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_439),
.B(n_27),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_509),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_352),
.B(n_27),
.Y(n_662)
);

XNOR2x2_ASAP7_75t_L g663 ( 
.A(n_371),
.B(n_29),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_352),
.B(n_29),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_353),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_509),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_355),
.Y(n_667)
);

INVx3_ASAP7_75t_L g668 ( 
.A(n_471),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_SL g669 ( 
.A(n_541),
.B(n_32),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_484),
.B(n_32),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_356),
.Y(n_671)
);

INVx6_ASAP7_75t_L g672 ( 
.A(n_545),
.Y(n_672)
);

BUFx6f_ASAP7_75t_L g673 ( 
.A(n_528),
.Y(n_673)
);

BUFx12f_ASAP7_75t_L g674 ( 
.A(n_366),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_528),
.Y(n_675)
);

INVx4_ASAP7_75t_L g676 ( 
.A(n_320),
.Y(n_676)
);

AND2x4_ASAP7_75t_L g677 ( 
.A(n_489),
.B(n_33),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_440),
.Y(n_678)
);

BUFx8_ASAP7_75t_L g679 ( 
.A(n_329),
.Y(n_679)
);

BUFx8_ASAP7_75t_SL g680 ( 
.A(n_408),
.Y(n_680)
);

BUFx12f_ASAP7_75t_L g681 ( 
.A(n_373),
.Y(n_681)
);

HB1xp67_ASAP7_75t_L g682 ( 
.A(n_376),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_449),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_490),
.B(n_34),
.Y(n_684)
);

INVx5_ASAP7_75t_L g685 ( 
.A(n_411),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_452),
.B(n_35),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_322),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_493),
.B(n_35),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_501),
.Y(n_689)
);

INVx5_ASAP7_75t_L g690 ( 
.A(n_474),
.Y(n_690)
);

BUFx12f_ASAP7_75t_L g691 ( 
.A(n_379),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_515),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_467),
.B(n_472),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_476),
.B(n_36),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_485),
.B(n_36),
.Y(n_695)
);

INVx5_ASAP7_75t_L g696 ( 
.A(n_482),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_492),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_531),
.B(n_37),
.Y(n_698)
);

AND2x4_ASAP7_75t_L g699 ( 
.A(n_551),
.B(n_38),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_401),
.Y(n_700)
);

INVx5_ASAP7_75t_L g701 ( 
.A(n_516),
.Y(n_701)
);

INVx4_ASAP7_75t_L g702 ( 
.A(n_333),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_502),
.Y(n_703)
);

AND2x4_ASAP7_75t_L g704 ( 
.A(n_532),
.B(n_40),
.Y(n_704)
);

INVx5_ASAP7_75t_L g705 ( 
.A(n_428),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_503),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_506),
.Y(n_707)
);

BUFx6f_ASAP7_75t_L g708 ( 
.A(n_507),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_404),
.Y(n_709)
);

BUFx12f_ASAP7_75t_L g710 ( 
.A(n_405),
.Y(n_710)
);

INVx5_ASAP7_75t_L g711 ( 
.A(n_428),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_517),
.Y(n_712)
);

AND2x2_ASAP7_75t_L g713 ( 
.A(n_648),
.B(n_658),
.Y(n_713)
);

AO22x2_ASAP7_75t_L g714 ( 
.A1(n_604),
.A2(n_394),
.B1(n_477),
.B2(n_397),
.Y(n_714)
);

AND2x2_ASAP7_75t_L g715 ( 
.A(n_648),
.B(n_407),
.Y(n_715)
);

OAI22xp33_ASAP7_75t_L g716 ( 
.A1(n_577),
.A2(n_669),
.B1(n_574),
.B2(n_609),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_648),
.B(n_500),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_570),
.Y(n_718)
);

OAI22xp33_ASAP7_75t_SL g719 ( 
.A1(n_577),
.A2(n_415),
.B1(n_416),
.B2(n_413),
.Y(n_719)
);

OAI22xp33_ASAP7_75t_L g720 ( 
.A1(n_669),
.A2(n_574),
.B1(n_562),
.B2(n_672),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_658),
.B(n_565),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_658),
.B(n_426),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_556),
.A2(n_495),
.B1(n_460),
.B2(n_409),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_587),
.B(n_438),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_641),
.A2(n_518),
.B1(n_523),
.B2(n_522),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_589),
.B(n_441),
.Y(n_726)
);

OAI22xp33_ASAP7_75t_L g727 ( 
.A1(n_672),
.A2(n_409),
.B1(n_429),
.B2(n_316),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_L g728 ( 
.A1(n_558),
.A2(n_429),
.B1(n_463),
.B2(n_316),
.Y(n_728)
);

OA22x2_ASAP7_75t_L g729 ( 
.A1(n_629),
.A2(n_448),
.B1(n_450),
.B2(n_446),
.Y(n_729)
);

AO22x2_ASAP7_75t_L g730 ( 
.A1(n_662),
.A2(n_535),
.B1(n_538),
.B2(n_533),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_570),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_L g732 ( 
.A1(n_582),
.A2(n_463),
.B1(n_347),
.B2(n_359),
.Y(n_732)
);

OAI22xp33_ASAP7_75t_SL g733 ( 
.A1(n_553),
.A2(n_552),
.B1(n_453),
.B2(n_454),
.Y(n_733)
);

OAI22xp5_ASAP7_75t_L g734 ( 
.A1(n_664),
.A2(n_458),
.B1(n_461),
.B2(n_451),
.Y(n_734)
);

AOI22xp5_ASAP7_75t_L g735 ( 
.A1(n_557),
.A2(n_387),
.B1(n_486),
.B2(n_344),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_L g736 ( 
.A(n_649),
.B(n_420),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_611),
.B(n_464),
.Y(n_737)
);

AOI22x1_ASAP7_75t_SL g738 ( 
.A1(n_569),
.A2(n_475),
.B1(n_491),
.B2(n_481),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_573),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_559),
.B(n_497),
.Y(n_740)
);

OAI22xp5_ASAP7_75t_SL g741 ( 
.A1(n_663),
.A2(n_519),
.B1(n_520),
.B2(n_510),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_567),
.A2(n_536),
.B1(n_540),
.B2(n_537),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_573),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_601),
.A2(n_547),
.B1(n_550),
.B2(n_432),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_616),
.A2(n_544),
.B1(n_548),
.B2(n_543),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_560),
.A2(n_549),
.B1(n_468),
.B2(n_436),
.Y(n_746)
);

OAI22xp33_ASAP7_75t_L g747 ( 
.A1(n_559),
.A2(n_338),
.B1(n_339),
.B2(n_335),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_559),
.B(n_345),
.Y(n_748)
);

INVx2_ASAP7_75t_L g749 ( 
.A(n_555),
.Y(n_749)
);

OR2x2_ASAP7_75t_L g750 ( 
.A(n_657),
.B(n_40),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_576),
.B(n_346),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_576),
.B(n_354),
.Y(n_752)
);

AOI22xp5_ASAP7_75t_L g753 ( 
.A1(n_560),
.A2(n_358),
.B1(n_360),
.B2(n_357),
.Y(n_753)
);

AND2x2_ASAP7_75t_L g754 ( 
.A(n_579),
.B(n_362),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_639),
.Y(n_755)
);

OAI22xp33_ASAP7_75t_SL g756 ( 
.A1(n_693),
.A2(n_369),
.B1(n_375),
.B2(n_367),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_564),
.Y(n_757)
);

AOI22xp5_ASAP7_75t_L g758 ( 
.A1(n_566),
.A2(n_378),
.B1(n_382),
.B2(n_377),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_579),
.B(n_383),
.Y(n_759)
);

AOI22xp5_ASAP7_75t_L g760 ( 
.A1(n_566),
.A2(n_385),
.B1(n_390),
.B2(n_384),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_649),
.B(n_391),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_579),
.A2(n_542),
.B1(n_534),
.B2(n_530),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_581),
.B(n_395),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_572),
.Y(n_764)
);

BUFx10_ASAP7_75t_L g765 ( 
.A(n_616),
.Y(n_765)
);

OAI22xp5_ASAP7_75t_SL g766 ( 
.A1(n_592),
.A2(n_529),
.B1(n_527),
.B2(n_526),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_639),
.Y(n_767)
);

AO22x2_ASAP7_75t_L g768 ( 
.A1(n_617),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_575),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_581),
.B(n_396),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_403),
.Y(n_771)
);

AOI22xp5_ASAP7_75t_L g772 ( 
.A1(n_568),
.A2(n_525),
.B1(n_513),
.B2(n_511),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_676),
.B(n_406),
.Y(n_773)
);

OAI22xp33_ASAP7_75t_SL g774 ( 
.A1(n_693),
.A2(n_505),
.B1(n_504),
.B2(n_498),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_594),
.B(n_412),
.Y(n_775)
);

OAI22xp33_ASAP7_75t_L g776 ( 
.A1(n_594),
.A2(n_496),
.B1(n_488),
.B2(n_483),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_598),
.B(n_414),
.Y(n_777)
);

OAI22xp33_ASAP7_75t_L g778 ( 
.A1(n_598),
.A2(n_612),
.B1(n_614),
.B2(n_610),
.Y(n_778)
);

INVx2_ASAP7_75t_L g779 ( 
.A(n_575),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_598),
.B(n_610),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

AOI22xp5_ASAP7_75t_L g782 ( 
.A1(n_568),
.A2(n_480),
.B1(n_473),
.B2(n_466),
.Y(n_782)
);

INVx1_ASAP7_75t_SL g783 ( 
.A(n_680),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_642),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_610),
.B(n_421),
.Y(n_785)
);

AO22x2_ASAP7_75t_L g786 ( 
.A1(n_617),
.A2(n_41),
.B1(n_42),
.B2(n_44),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_575),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_SL g788 ( 
.A(n_618),
.B(n_423),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_642),
.Y(n_789)
);

OA22x2_ASAP7_75t_L g790 ( 
.A1(n_629),
.A2(n_457),
.B1(n_456),
.B2(n_455),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_612),
.B(n_424),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_642),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_584),
.A2(n_445),
.B1(n_444),
.B2(n_443),
.Y(n_793)
);

OAI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_595),
.A2(n_442),
.B1(n_434),
.B2(n_427),
.Y(n_794)
);

AOI22xp5_ASAP7_75t_L g795 ( 
.A1(n_584),
.A2(n_437),
.B1(n_419),
.B2(n_51),
.Y(n_795)
);

OR2x2_ASAP7_75t_L g796 ( 
.A(n_561),
.B(n_45),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_614),
.B(n_419),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_644),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_704),
.A2(n_618),
.B1(n_599),
.B2(n_593),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_586),
.B(n_419),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_676),
.B(n_419),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_583),
.Y(n_802)
);

AO22x2_ASAP7_75t_L g803 ( 
.A1(n_586),
.A2(n_48),
.B1(n_51),
.B2(n_52),
.Y(n_803)
);

AOI22xp5_ASAP7_75t_L g804 ( 
.A1(n_704),
.A2(n_437),
.B1(n_419),
.B2(n_55),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_687),
.B(n_702),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_638),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_583),
.Y(n_807)
);

OAI22xp33_ASAP7_75t_L g808 ( 
.A1(n_595),
.A2(n_53),
.B1(n_54),
.B2(n_56),
.Y(n_808)
);

OAI22xp33_ASAP7_75t_SL g809 ( 
.A1(n_608),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_655),
.A2(n_59),
.B1(n_60),
.B2(n_61),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_644),
.Y(n_811)
);

NOR2xp33_ASAP7_75t_L g812 ( 
.A(n_687),
.B(n_419),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

OAI22xp33_ASAP7_75t_L g814 ( 
.A1(n_608),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_596),
.A2(n_437),
.B1(n_419),
.B2(n_65),
.Y(n_815)
);

OR2x6_ASAP7_75t_L g816 ( 
.A(n_621),
.B(n_674),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_619),
.A2(n_437),
.B1(n_64),
.B2(n_66),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_806),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_718),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_806),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_805),
.B(n_702),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_765),
.Y(n_822)
);

XOR2xp5_ASAP7_75t_L g823 ( 
.A(n_735),
.B(n_590),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_731),
.Y(n_824)
);

CKINVDCx20_ASAP7_75t_R g825 ( 
.A(n_766),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_739),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_554),
.Y(n_827)
);

OAI21xp5_ASAP7_75t_L g828 ( 
.A1(n_800),
.A2(n_578),
.B(n_613),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_801),
.A2(n_615),
.B(n_613),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_723),
.Y(n_830)
);

INVx2_ASAP7_75t_L g831 ( 
.A(n_743),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_812),
.A2(n_620),
.B(n_615),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_749),
.Y(n_833)
);

NAND2x1p5_ASAP7_75t_L g834 ( 
.A(n_795),
.B(n_655),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_755),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_767),
.Y(n_836)
);

NOR2xp33_ASAP7_75t_L g837 ( 
.A(n_736),
.B(n_705),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_726),
.B(n_625),
.Y(n_838)
);

OR2x6_ASAP7_75t_L g839 ( 
.A(n_816),
.B(n_681),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_781),
.Y(n_840)
);

BUFx6f_ASAP7_75t_L g841 ( 
.A(n_769),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_784),
.Y(n_842)
);

HB1xp67_ASAP7_75t_L g843 ( 
.A(n_737),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_789),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_779),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_792),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_798),
.Y(n_847)
);

NOR2xp33_ASAP7_75t_L g848 ( 
.A(n_753),
.B(n_705),
.Y(n_848)
);

OR2x2_ASAP7_75t_L g849 ( 
.A(n_723),
.B(n_607),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_811),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_764),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_783),
.Y(n_853)
);

OR2x2_ASAP7_75t_L g854 ( 
.A(n_732),
.B(n_622),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_797),
.B(n_799),
.Y(n_855)
);

XNOR2x2_ASAP7_75t_L g856 ( 
.A(n_714),
.B(n_695),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_787),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_753),
.B(n_705),
.Y(n_858)
);

INVxp67_ASAP7_75t_SL g859 ( 
.A(n_795),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_758),
.B(n_711),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_802),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_721),
.B(n_640),
.Y(n_862)
);

XOR2xp5_ASAP7_75t_L g863 ( 
.A(n_727),
.B(n_651),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_715),
.B(n_711),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_807),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_765),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_740),
.B(n_665),
.Y(n_867)
);

INVx1_ASAP7_75t_SL g868 ( 
.A(n_722),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_813),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_761),
.B(n_711),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_744),
.B(n_667),
.Y(n_871)
);

NOR2xp67_ASAP7_75t_L g872 ( 
.A(n_804),
.B(n_691),
.Y(n_872)
);

XOR2x2_ASAP7_75t_L g873 ( 
.A(n_744),
.B(n_682),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_780),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_759),
.A2(n_633),
.B(n_620),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_799),
.B(n_578),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_750),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_804),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_758),
.B(n_671),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_796),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_713),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_748),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_751),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_752),
.Y(n_884)
);

CKINVDCx14_ASAP7_75t_R g885 ( 
.A(n_816),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_754),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_763),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_760),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_770),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_771),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_775),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_746),
.B(n_683),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_777),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_785),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_773),
.B(n_700),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_791),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_734),
.B(n_709),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_746),
.B(n_578),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_760),
.B(n_697),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_772),
.B(n_679),
.Y(n_900)
);

INVxp67_ASAP7_75t_SL g901 ( 
.A(n_720),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_729),
.Y(n_902)
);

INVxp67_ASAP7_75t_SL g903 ( 
.A(n_815),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_772),
.B(n_685),
.Y(n_904)
);

NOR2xp33_ASAP7_75t_L g905 ( 
.A(n_782),
.B(n_679),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_815),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_725),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_738),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_725),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_821),
.B(n_782),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_843),
.Y(n_911)
);

INVx2_ASAP7_75t_L g912 ( 
.A(n_833),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_827),
.Y(n_913)
);

OAI21xp5_ASAP7_75t_L g914 ( 
.A1(n_829),
.A2(n_793),
.B(n_578),
.Y(n_914)
);

AND2x2_ASAP7_75t_L g915 ( 
.A(n_901),
.B(n_745),
.Y(n_915)
);

BUFx6f_ASAP7_75t_L g916 ( 
.A(n_841),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_838),
.Y(n_917)
);

AND2x2_ASAP7_75t_L g918 ( 
.A(n_901),
.B(n_745),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_851),
.Y(n_919)
);

INVxp67_ASAP7_75t_SL g920 ( 
.A(n_834),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_SL g921 ( 
.A(n_829),
.B(n_716),
.Y(n_921)
);

AND2x6_ASAP7_75t_L g922 ( 
.A(n_876),
.B(n_817),
.Y(n_922)
);

INVx4_ASAP7_75t_L g923 ( 
.A(n_841),
.Y(n_923)
);

BUFx3_ASAP7_75t_L g924 ( 
.A(n_841),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_859),
.B(n_872),
.Y(n_925)
);

INVx1_ASAP7_75t_SL g926 ( 
.A(n_853),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_821),
.B(n_793),
.Y(n_927)
);

OAI21xp5_ASAP7_75t_L g928 ( 
.A1(n_832),
.A2(n_742),
.B(n_635),
.Y(n_928)
);

AND2x4_ASAP7_75t_L g929 ( 
.A(n_859),
.B(n_670),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_852),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_845),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_899),
.B(n_730),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_819),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_895),
.B(n_756),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_824),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_845),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_831),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_826),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_855),
.B(n_730),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_SL g940 ( 
.A(n_900),
.B(n_728),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_869),
.Y(n_941)
);

AND2x2_ASAP7_75t_L g942 ( 
.A(n_855),
.B(n_768),
.Y(n_942)
);

HB1xp67_ASAP7_75t_L g943 ( 
.A(n_843),
.Y(n_943)
);

AND2x2_ASAP7_75t_L g944 ( 
.A(n_906),
.B(n_768),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_835),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_878),
.B(n_786),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_836),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_840),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_875),
.B(n_670),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_903),
.B(n_677),
.Y(n_950)
);

OR2x2_ASAP7_75t_L g951 ( 
.A(n_849),
.B(n_741),
.Y(n_951)
);

AND2x2_ASAP7_75t_L g952 ( 
.A(n_892),
.B(n_786),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_892),
.B(n_803),
.Y(n_953)
);

AND2x2_ASAP7_75t_SL g954 ( 
.A(n_876),
.B(n_817),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_842),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_834),
.B(n_803),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_903),
.B(n_714),
.Y(n_957)
);

INVx1_ASAP7_75t_SL g958 ( 
.A(n_862),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_844),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_868),
.B(n_774),
.Y(n_960)
);

BUFx6f_ASAP7_75t_L g961 ( 
.A(n_845),
.Y(n_961)
);

AND2x4_ASAP7_75t_L g962 ( 
.A(n_907),
.B(n_677),
.Y(n_962)
);

AND2x2_ASAP7_75t_L g963 ( 
.A(n_867),
.B(n_684),
.Y(n_963)
);

AND2x2_ASAP7_75t_L g964 ( 
.A(n_879),
.B(n_684),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_879),
.B(n_688),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_862),
.Y(n_966)
);

INVx3_ASAP7_75t_L g967 ( 
.A(n_891),
.Y(n_967)
);

AND2x4_ASAP7_75t_L g968 ( 
.A(n_909),
.B(n_688),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_894),
.B(n_698),
.Y(n_969)
);

OAI21xp5_ASAP7_75t_L g970 ( 
.A1(n_832),
.A2(n_646),
.B(n_624),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_877),
.B(n_698),
.Y(n_971)
);

AND2x2_ASAP7_75t_L g972 ( 
.A(n_896),
.B(n_699),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_880),
.B(n_699),
.Y(n_973)
);

INVx2_ASAP7_75t_L g974 ( 
.A(n_846),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_847),
.Y(n_975)
);

INVx2_ASAP7_75t_SL g976 ( 
.A(n_822),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_850),
.Y(n_977)
);

HB1xp67_ASAP7_75t_L g978 ( 
.A(n_866),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_818),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_820),
.Y(n_980)
);

NOR2xp67_ASAP7_75t_R g981 ( 
.A(n_902),
.B(n_710),
.Y(n_981)
);

AND2x2_ASAP7_75t_L g982 ( 
.A(n_848),
.B(n_790),
.Y(n_982)
);

OR2x2_ASAP7_75t_SL g983 ( 
.A(n_871),
.B(n_719),
.Y(n_983)
);

INVx2_ASAP7_75t_SL g984 ( 
.A(n_874),
.Y(n_984)
);

BUFx3_ASAP7_75t_L g985 ( 
.A(n_839),
.Y(n_985)
);

AND2x4_ASAP7_75t_L g986 ( 
.A(n_882),
.B(n_717),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_857),
.Y(n_987)
);

AND2x4_ASAP7_75t_L g988 ( 
.A(n_883),
.B(n_884),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_861),
.Y(n_989)
);

NAND2xp5_ASAP7_75t_L g990 ( 
.A(n_875),
.B(n_788),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_865),
.Y(n_991)
);

INVx2_ASAP7_75t_SL g992 ( 
.A(n_881),
.Y(n_992)
);

INVxp67_ASAP7_75t_L g993 ( 
.A(n_863),
.Y(n_993)
);

OAI21xp5_ASAP7_75t_L g994 ( 
.A1(n_828),
.A2(n_656),
.B(n_647),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_886),
.Y(n_995)
);

AND2x6_ASAP7_75t_L g996 ( 
.A(n_898),
.B(n_638),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_887),
.Y(n_997)
);

INVx4_ASAP7_75t_L g998 ( 
.A(n_839),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_889),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_848),
.B(n_706),
.Y(n_1000)
);

HB1xp67_ASAP7_75t_L g1001 ( 
.A(n_854),
.Y(n_1001)
);

BUFx6f_ASAP7_75t_L g1002 ( 
.A(n_890),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_858),
.B(n_707),
.Y(n_1003)
);

INVx2_ASAP7_75t_L g1004 ( 
.A(n_893),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_823),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_905),
.B(n_712),
.Y(n_1006)
);

INVxp67_ASAP7_75t_SL g1007 ( 
.A(n_920),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_937),
.Y(n_1008)
);

OR2x6_ASAP7_75t_L g1009 ( 
.A(n_925),
.B(n_839),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_913),
.B(n_873),
.Y(n_1010)
);

INVx5_ASAP7_75t_L g1011 ( 
.A(n_925),
.Y(n_1011)
);

AND2x4_ASAP7_75t_L g1012 ( 
.A(n_925),
.B(n_888),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_917),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_910),
.B(n_858),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_927),
.B(n_860),
.Y(n_1015)
);

AND2x2_ASAP7_75t_L g1016 ( 
.A(n_964),
.B(n_897),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_SL g1017 ( 
.A(n_940),
.B(n_860),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_937),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_954),
.B(n_904),
.Y(n_1019)
);

BUFx4f_ASAP7_75t_L g1020 ( 
.A(n_950),
.Y(n_1020)
);

OR2x2_ASAP7_75t_L g1021 ( 
.A(n_951),
.B(n_911),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_954),
.B(n_904),
.Y(n_1022)
);

BUFx6f_ASAP7_75t_L g1023 ( 
.A(n_916),
.Y(n_1023)
);

BUFx3_ASAP7_75t_L g1024 ( 
.A(n_926),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_967),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_943),
.Y(n_1026)
);

OR2x6_ASAP7_75t_L g1027 ( 
.A(n_998),
.B(n_885),
.Y(n_1027)
);

AND2x4_ASAP7_75t_L g1028 ( 
.A(n_950),
.B(n_825),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_1004),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_916),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_985),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_934),
.B(n_830),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_923),
.Y(n_1033)
);

OR2x6_ASAP7_75t_L g1034 ( 
.A(n_998),
.B(n_810),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_958),
.Y(n_1035)
);

NOR2xp33_ASAP7_75t_L g1036 ( 
.A(n_951),
.B(n_794),
.Y(n_1036)
);

OR2x6_ASAP7_75t_L g1037 ( 
.A(n_998),
.B(n_563),
.Y(n_1037)
);

NAND2xp33_ASAP7_75t_L g1038 ( 
.A(n_990),
.B(n_828),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_912),
.Y(n_1039)
);

OR2x6_ASAP7_75t_L g1040 ( 
.A(n_985),
.B(n_563),
.Y(n_1040)
);

INVx3_ASAP7_75t_L g1041 ( 
.A(n_923),
.Y(n_1041)
);

OR2x2_ASAP7_75t_L g1042 ( 
.A(n_1001),
.B(n_856),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_933),
.Y(n_1043)
);

INVx5_ASAP7_75t_L g1044 ( 
.A(n_996),
.Y(n_1044)
);

AO21x2_ASAP7_75t_L g1045 ( 
.A1(n_994),
.A2(n_605),
.B(n_603),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1003),
.B(n_837),
.Y(n_1046)
);

OR2x2_ASAP7_75t_L g1047 ( 
.A(n_1005),
.B(n_597),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_923),
.Y(n_1048)
);

NOR2xp33_ASAP7_75t_SL g1049 ( 
.A(n_914),
.B(n_908),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_L g1050 ( 
.A(n_1003),
.B(n_864),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_912),
.Y(n_1051)
);

OR2x6_ASAP7_75t_L g1052 ( 
.A(n_956),
.B(n_634),
.Y(n_1052)
);

INVxp67_ASAP7_75t_SL g1053 ( 
.A(n_916),
.Y(n_1053)
);

INVx2_ASAP7_75t_L g1054 ( 
.A(n_941),
.Y(n_1054)
);

NOR2xp33_ASAP7_75t_SL g1055 ( 
.A(n_922),
.B(n_809),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_941),
.Y(n_1056)
);

OR2x6_ASAP7_75t_L g1057 ( 
.A(n_956),
.B(n_643),
.Y(n_1057)
);

INVxp67_ASAP7_75t_L g1058 ( 
.A(n_963),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_966),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_933),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_950),
.B(n_689),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_964),
.B(n_778),
.Y(n_1062)
);

BUFx4f_ASAP7_75t_L g1063 ( 
.A(n_929),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1000),
.B(n_733),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_916),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_929),
.B(n_689),
.Y(n_1066)
);

OR2x2_ASAP7_75t_L g1067 ( 
.A(n_965),
.B(n_692),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_965),
.B(n_627),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_921),
.B(n_870),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_999),
.Y(n_1070)
);

AND2x4_ASAP7_75t_L g1071 ( 
.A(n_929),
.B(n_692),
.Y(n_1071)
);

INVxp67_ASAP7_75t_L g1072 ( 
.A(n_963),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_999),
.Y(n_1073)
);

OR2x6_ASAP7_75t_L g1074 ( 
.A(n_966),
.B(n_650),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_916),
.Y(n_1075)
);

HB1xp67_ASAP7_75t_L g1076 ( 
.A(n_952),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_936),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_SL g1078 ( 
.A(n_997),
.B(n_747),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_947),
.Y(n_1079)
);

BUFx8_ASAP7_75t_SL g1080 ( 
.A(n_988),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_947),
.Y(n_1081)
);

NAND2x1p5_ASAP7_75t_L g1082 ( 
.A(n_924),
.B(n_644),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_935),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_948),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_SL g1085 ( 
.A(n_922),
.B(n_808),
.Y(n_1085)
);

BUFx6f_ASAP7_75t_L g1086 ( 
.A(n_936),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_936),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_936),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_1008),
.Y(n_1089)
);

BUFx3_ASAP7_75t_L g1090 ( 
.A(n_1024),
.Y(n_1090)
);

NOR2xp67_ASAP7_75t_L g1091 ( 
.A(n_1011),
.B(n_976),
.Y(n_1091)
);

CKINVDCx16_ASAP7_75t_R g1092 ( 
.A(n_1027),
.Y(n_1092)
);

NAND2x1p5_ASAP7_75t_L g1093 ( 
.A(n_1011),
.B(n_1020),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_1007),
.Y(n_1094)
);

BUFx4_ASAP7_75t_SL g1095 ( 
.A(n_1009),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_1018),
.Y(n_1096)
);

INVxp67_ASAP7_75t_SL g1097 ( 
.A(n_1014),
.Y(n_1097)
);

INVx2_ASAP7_75t_L g1098 ( 
.A(n_1039),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1043),
.Y(n_1099)
);

NAND2x1p5_ASAP7_75t_L g1100 ( 
.A(n_1011),
.B(n_924),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1060),
.Y(n_1101)
);

NAND2x1p5_ASAP7_75t_L g1102 ( 
.A(n_1020),
.B(n_931),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1036),
.A2(n_922),
.B1(n_957),
.B2(n_942),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1026),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_1063),
.B(n_931),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_1023),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_1063),
.Y(n_1107)
);

BUFx3_ASAP7_75t_L g1108 ( 
.A(n_1080),
.Y(n_1108)
);

BUFx6f_ASAP7_75t_L g1109 ( 
.A(n_1023),
.Y(n_1109)
);

BUFx3_ASAP7_75t_L g1110 ( 
.A(n_1027),
.Y(n_1110)
);

INVx5_ASAP7_75t_L g1111 ( 
.A(n_1044),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_1013),
.Y(n_1112)
);

INVx1_ASAP7_75t_L g1113 ( 
.A(n_1070),
.Y(n_1113)
);

BUFx2_ASAP7_75t_L g1114 ( 
.A(n_1009),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_1009),
.B(n_915),
.Y(n_1115)
);

INVx6_ASAP7_75t_L g1116 ( 
.A(n_1012),
.Y(n_1116)
);

NAND2x1p5_ASAP7_75t_L g1117 ( 
.A(n_1044),
.B(n_1033),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1016),
.B(n_915),
.Y(n_1118)
);

BUFx6f_ASAP7_75t_L g1119 ( 
.A(n_1023),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1051),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_1031),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_1030),
.Y(n_1122)
);

BUFx12f_ASAP7_75t_L g1123 ( 
.A(n_1028),
.Y(n_1123)
);

BUFx6f_ASAP7_75t_L g1124 ( 
.A(n_1030),
.Y(n_1124)
);

CKINVDCx16_ASAP7_75t_R g1125 ( 
.A(n_1040),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_1061),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1073),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1044),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1032),
.A2(n_922),
.B1(n_957),
.B2(n_942),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_1028),
.Y(n_1130)
);

BUFx6f_ASAP7_75t_L g1131 ( 
.A(n_1030),
.Y(n_1131)
);

INVx3_ASAP7_75t_L g1132 ( 
.A(n_1075),
.Y(n_1132)
);

INVx5_ASAP7_75t_L g1133 ( 
.A(n_1075),
.Y(n_1133)
);

BUFx6f_ASAP7_75t_L g1134 ( 
.A(n_1075),
.Y(n_1134)
);

INVx5_ASAP7_75t_SL g1135 ( 
.A(n_1040),
.Y(n_1135)
);

INVx2_ASAP7_75t_SL g1136 ( 
.A(n_1012),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_1083),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1021),
.B(n_918),
.Y(n_1138)
);

INVx4_ASAP7_75t_L g1139 ( 
.A(n_1077),
.Y(n_1139)
);

INVxp67_ASAP7_75t_SL g1140 ( 
.A(n_1014),
.Y(n_1140)
);

INVx3_ASAP7_75t_L g1141 ( 
.A(n_1077),
.Y(n_1141)
);

BUFx3_ASAP7_75t_L g1142 ( 
.A(n_1059),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1035),
.Y(n_1143)
);

INVx4_ASAP7_75t_L g1144 ( 
.A(n_1077),
.Y(n_1144)
);

BUFx6f_ASAP7_75t_L g1145 ( 
.A(n_1086),
.Y(n_1145)
);

INVx2_ASAP7_75t_SL g1146 ( 
.A(n_1047),
.Y(n_1146)
);

BUFx6f_ASAP7_75t_L g1147 ( 
.A(n_1086),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_L g1148 ( 
.A(n_1086),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_1040),
.Y(n_1149)
);

INVx8_ASAP7_75t_L g1150 ( 
.A(n_1074),
.Y(n_1150)
);

BUFx2_ASAP7_75t_L g1151 ( 
.A(n_1034),
.Y(n_1151)
);

INVx3_ASAP7_75t_SL g1152 ( 
.A(n_1034),
.Y(n_1152)
);

BUFx4_ASAP7_75t_SL g1153 ( 
.A(n_1034),
.Y(n_1153)
);

INVx1_ASAP7_75t_SL g1154 ( 
.A(n_1010),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1087),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_1087),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1087),
.Y(n_1157)
);

INVx3_ASAP7_75t_L g1158 ( 
.A(n_1088),
.Y(n_1158)
);

INVxp67_ASAP7_75t_SL g1159 ( 
.A(n_1015),
.Y(n_1159)
);

BUFx3_ASAP7_75t_L g1160 ( 
.A(n_1088),
.Y(n_1160)
);

NAND2x1p5_ASAP7_75t_L g1161 ( 
.A(n_1033),
.B(n_936),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_1137),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1154),
.A2(n_1017),
.B1(n_1049),
.B2(n_922),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1099),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1101),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1104),
.Y(n_1166)
);

BUFx12f_ASAP7_75t_L g1167 ( 
.A(n_1108),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1113),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1127),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1089),
.Y(n_1170)
);

AOI22xp33_ASAP7_75t_L g1171 ( 
.A1(n_1129),
.A2(n_1017),
.B1(n_1015),
.B2(n_1049),
.Y(n_1171)
);

BUFx6f_ASAP7_75t_L g1172 ( 
.A(n_1111),
.Y(n_1172)
);

CKINVDCx11_ASAP7_75t_R g1173 ( 
.A(n_1108),
.Y(n_1173)
);

CKINVDCx6p67_ASAP7_75t_R g1174 ( 
.A(n_1090),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_1138),
.B(n_1076),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_1121),
.Y(n_1176)
);

CKINVDCx11_ASAP7_75t_R g1177 ( 
.A(n_1090),
.Y(n_1177)
);

AO22x1_ASAP7_75t_L g1178 ( 
.A1(n_1097),
.A2(n_922),
.B1(n_1006),
.B2(n_1061),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_1097),
.A2(n_1022),
.B1(n_1019),
.B2(n_921),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1129),
.A2(n_1022),
.B1(n_1019),
.B2(n_1042),
.Y(n_1180)
);

OAI22xp5_ASAP7_75t_L g1181 ( 
.A1(n_1140),
.A2(n_1067),
.B1(n_1072),
.B2(n_1046),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_SL g1182 ( 
.A1(n_1140),
.A2(n_928),
.B(n_970),
.Y(n_1182)
);

INVx6_ASAP7_75t_SL g1183 ( 
.A(n_1115),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1159),
.A2(n_1103),
.B1(n_1118),
.B2(n_1064),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1159),
.A2(n_1072),
.B1(n_1046),
.B2(n_949),
.Y(n_1185)
);

INVx2_ASAP7_75t_L g1186 ( 
.A(n_1089),
.Y(n_1186)
);

BUFx6f_ASAP7_75t_L g1187 ( 
.A(n_1111),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1096),
.Y(n_1188)
);

BUFx4f_ASAP7_75t_SL g1189 ( 
.A(n_1142),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_L g1190 ( 
.A1(n_1123),
.A2(n_1055),
.B1(n_960),
.B2(n_1006),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1096),
.Y(n_1191)
);

INVx5_ASAP7_75t_L g1192 ( 
.A(n_1111),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1103),
.B(n_1050),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1098),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1098),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1126),
.B(n_952),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1123),
.A2(n_1055),
.B1(n_1006),
.B2(n_932),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1111),
.Y(n_1198)
);

BUFx12f_ASAP7_75t_L g1199 ( 
.A(n_1130),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1120),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1120),
.Y(n_1201)
);

CKINVDCx6p67_ASAP7_75t_R g1202 ( 
.A(n_1092),
.Y(n_1202)
);

INVx2_ASAP7_75t_SL g1203 ( 
.A(n_1095),
.Y(n_1203)
);

INVx6_ASAP7_75t_L g1204 ( 
.A(n_1133),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_SL g1205 ( 
.A1(n_1151),
.A2(n_814),
.B(n_982),
.Y(n_1205)
);

BUFx8_ASAP7_75t_L g1206 ( 
.A(n_1130),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1094),
.Y(n_1207)
);

AOI22xp33_ASAP7_75t_SL g1208 ( 
.A1(n_1116),
.A2(n_1085),
.B1(n_939),
.B2(n_982),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1112),
.Y(n_1209)
);

OAI22x1_ASAP7_75t_L g1210 ( 
.A1(n_1152),
.A2(n_1066),
.B1(n_1071),
.B2(n_944),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1136),
.A2(n_1085),
.B1(n_939),
.B2(n_932),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_1093),
.Y(n_1212)
);

BUFx12f_ASAP7_75t_L g1213 ( 
.A(n_1143),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1116),
.A2(n_918),
.B1(n_944),
.B2(n_946),
.Y(n_1214)
);

INVx8_ASAP7_75t_L g1215 ( 
.A(n_1150),
.Y(n_1215)
);

BUFx3_ASAP7_75t_L g1216 ( 
.A(n_1142),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1094),
.Y(n_1217)
);

BUFx12f_ASAP7_75t_L g1218 ( 
.A(n_1146),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1126),
.A2(n_1050),
.B1(n_1058),
.B2(n_983),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1116),
.A2(n_946),
.B1(n_1081),
.B2(n_1079),
.Y(n_1220)
);

BUFx2_ASAP7_75t_L g1221 ( 
.A(n_1152),
.Y(n_1221)
);

INVx6_ASAP7_75t_L g1222 ( 
.A(n_1133),
.Y(n_1222)
);

BUFx12f_ASAP7_75t_L g1223 ( 
.A(n_1110),
.Y(n_1223)
);

INVx2_ASAP7_75t_L g1224 ( 
.A(n_1115),
.Y(n_1224)
);

BUFx4_ASAP7_75t_R g1225 ( 
.A(n_1110),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_L g1226 ( 
.A1(n_1115),
.A2(n_1084),
.B1(n_1066),
.B2(n_1071),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1155),
.Y(n_1227)
);

AOI22xp33_ASAP7_75t_L g1228 ( 
.A1(n_1150),
.A2(n_1029),
.B1(n_997),
.B2(n_1002),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1114),
.Y(n_1229)
);

INVx3_ASAP7_75t_L g1230 ( 
.A(n_1128),
.Y(n_1230)
);

CKINVDCx6p67_ASAP7_75t_R g1231 ( 
.A(n_1133),
.Y(n_1231)
);

CKINVDCx11_ASAP7_75t_R g1232 ( 
.A(n_1125),
.Y(n_1232)
);

INVx2_ASAP7_75t_L g1233 ( 
.A(n_1155),
.Y(n_1233)
);

AOI22xp33_ASAP7_75t_SL g1234 ( 
.A1(n_1219),
.A2(n_1150),
.B1(n_1135),
.B2(n_953),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1162),
.Y(n_1235)
);

BUFx3_ASAP7_75t_L g1236 ( 
.A(n_1177),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1171),
.A2(n_1057),
.B1(n_1052),
.B2(n_993),
.Y(n_1237)
);

AOI21xp33_ASAP7_75t_L g1238 ( 
.A1(n_1171),
.A2(n_1069),
.B(n_1078),
.Y(n_1238)
);

OAI21xp33_ASAP7_75t_SL g1239 ( 
.A1(n_1193),
.A2(n_1069),
.B(n_1139),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1184),
.A2(n_976),
.B1(n_983),
.B2(n_992),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1164),
.Y(n_1241)
);

BUFx4f_ASAP7_75t_SL g1242 ( 
.A(n_1167),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1184),
.A2(n_1163),
.B1(n_1181),
.B2(n_1193),
.Y(n_1243)
);

BUFx4f_ASAP7_75t_SL g1244 ( 
.A(n_1206),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1165),
.Y(n_1245)
);

OAI222xp33_ASAP7_75t_L g1246 ( 
.A1(n_1208),
.A2(n_1057),
.B1(n_1052),
.B2(n_1074),
.C1(n_953),
.C2(n_1037),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1168),
.Y(n_1247)
);

OAI21xp5_ASAP7_75t_SL g1248 ( 
.A1(n_1219),
.A2(n_1153),
.B(n_652),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1175),
.B(n_1135),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1208),
.A2(n_1057),
.B1(n_1052),
.B2(n_997),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1180),
.A2(n_997),
.B1(n_1002),
.B2(n_992),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_SL g1252 ( 
.A1(n_1181),
.A2(n_1135),
.B1(n_1149),
.B2(n_1153),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_L g1253 ( 
.A1(n_1180),
.A2(n_1002),
.B1(n_997),
.B2(n_988),
.Y(n_1253)
);

NOR2xp33_ASAP7_75t_L g1254 ( 
.A(n_1209),
.B(n_978),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1196),
.B(n_1037),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_1189),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1166),
.B(n_1068),
.Y(n_1257)
);

BUFx2_ASAP7_75t_L g1258 ( 
.A(n_1221),
.Y(n_1258)
);

AOI22xp33_ASAP7_75t_SL g1259 ( 
.A1(n_1179),
.A2(n_1002),
.B1(n_996),
.B2(n_1107),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1190),
.A2(n_1002),
.B1(n_988),
.B2(n_995),
.Y(n_1260)
);

BUFx2_ASAP7_75t_L g1261 ( 
.A(n_1216),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1179),
.A2(n_996),
.B1(n_1107),
.B2(n_1093),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1169),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1166),
.B(n_1209),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_L g1265 ( 
.A1(n_1197),
.A2(n_1210),
.B1(n_1211),
.B2(n_1226),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1173),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1185),
.A2(n_948),
.B1(n_974),
.B2(n_959),
.Y(n_1267)
);

OAI21xp33_ASAP7_75t_L g1268 ( 
.A1(n_1182),
.A2(n_652),
.B(n_633),
.Y(n_1268)
);

OAI22xp5_ASAP7_75t_L g1269 ( 
.A1(n_1185),
.A2(n_1091),
.B1(n_1074),
.B2(n_938),
.Y(n_1269)
);

OR2x2_ASAP7_75t_L g1270 ( 
.A(n_1207),
.B(n_1037),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1226),
.A2(n_919),
.B1(n_974),
.B2(n_959),
.Y(n_1271)
);

BUFx4f_ASAP7_75t_SL g1272 ( 
.A(n_1206),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1203),
.B(n_984),
.Y(n_1273)
);

INVx2_ASAP7_75t_L g1274 ( 
.A(n_1170),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1214),
.A2(n_919),
.B1(n_975),
.B2(n_1054),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1214),
.A2(n_975),
.B1(n_1056),
.B2(n_991),
.Y(n_1276)
);

OAI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_1205),
.A2(n_659),
.B(n_653),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1220),
.A2(n_989),
.B1(n_991),
.B2(n_930),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1186),
.Y(n_1279)
);

AOI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1218),
.A2(n_989),
.B1(n_930),
.B2(n_986),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1217),
.Y(n_1281)
);

INVxp67_ASAP7_75t_L g1282 ( 
.A(n_1229),
.Y(n_1282)
);

BUFx4f_ASAP7_75t_SL g1283 ( 
.A(n_1174),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1189),
.Y(n_1284)
);

BUFx5_ASAP7_75t_L g1285 ( 
.A(n_1188),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1220),
.A2(n_986),
.B1(n_955),
.B2(n_977),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1191),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1228),
.A2(n_984),
.B1(n_1062),
.B2(n_1102),
.Y(n_1288)
);

AOI22xp33_ASAP7_75t_L g1289 ( 
.A1(n_1224),
.A2(n_986),
.B1(n_945),
.B2(n_987),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1195),
.Y(n_1290)
);

AOI22xp33_ASAP7_75t_L g1291 ( 
.A1(n_1199),
.A2(n_969),
.B1(n_996),
.B2(n_1025),
.Y(n_1291)
);

AOI22xp33_ASAP7_75t_SL g1292 ( 
.A1(n_1223),
.A2(n_996),
.B1(n_1038),
.B2(n_969),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1232),
.A2(n_969),
.B1(n_703),
.B2(n_708),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1213),
.A2(n_703),
.B1(n_708),
.B2(n_678),
.Y(n_1294)
);

AND2x2_ASAP7_75t_L g1295 ( 
.A(n_1202),
.B(n_973),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1228),
.A2(n_1105),
.B1(n_1102),
.B2(n_653),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1201),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_SL g1298 ( 
.A1(n_1215),
.A2(n_996),
.B1(n_972),
.B2(n_686),
.Y(n_1298)
);

BUFx8_ASAP7_75t_L g1299 ( 
.A(n_1227),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1194),
.A2(n_972),
.B1(n_980),
.B2(n_979),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_1172),
.Y(n_1301)
);

NAND3xp33_ASAP7_75t_L g1302 ( 
.A(n_1277),
.B(n_694),
.C(n_660),
.Y(n_1302)
);

NAND3xp33_ASAP7_75t_L g1303 ( 
.A(n_1248),
.B(n_694),
.C(n_660),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1243),
.A2(n_1237),
.B1(n_1265),
.B2(n_1238),
.Y(n_1304)
);

OAI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1268),
.A2(n_707),
.B(n_1082),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1250),
.A2(n_1200),
.B1(n_1183),
.B2(n_1233),
.Y(n_1306)
);

HB1xp67_ASAP7_75t_L g1307 ( 
.A(n_1282),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1281),
.Y(n_1308)
);

AOI22xp33_ASAP7_75t_L g1309 ( 
.A1(n_1240),
.A2(n_1183),
.B1(n_979),
.B2(n_703),
.Y(n_1309)
);

AOI22xp33_ASAP7_75t_L g1310 ( 
.A1(n_1234),
.A2(n_979),
.B1(n_708),
.B2(n_678),
.Y(n_1310)
);

AOI22xp33_ASAP7_75t_L g1311 ( 
.A1(n_1260),
.A2(n_979),
.B1(n_678),
.B2(n_654),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1235),
.B(n_1045),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_SL g1313 ( 
.A1(n_1266),
.A2(n_1225),
.B1(n_1178),
.B2(n_1095),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_L g1314 ( 
.A1(n_1252),
.A2(n_979),
.B1(n_654),
.B2(n_661),
.Y(n_1314)
);

OAI22xp5_ASAP7_75t_L g1315 ( 
.A1(n_1293),
.A2(n_1105),
.B1(n_1230),
.B2(n_1192),
.Y(n_1315)
);

AOI22xp33_ASAP7_75t_L g1316 ( 
.A1(n_1293),
.A2(n_654),
.B1(n_661),
.B2(n_645),
.Y(n_1316)
);

AOI222xp33_ASAP7_75t_L g1317 ( 
.A1(n_1246),
.A2(n_973),
.B1(n_971),
.B2(n_603),
.C1(n_636),
.C2(n_675),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1241),
.B(n_1045),
.Y(n_1318)
);

AOI22xp33_ASAP7_75t_L g1319 ( 
.A1(n_1269),
.A2(n_666),
.B1(n_673),
.B2(n_645),
.Y(n_1319)
);

OAI221xp5_ASAP7_75t_L g1320 ( 
.A1(n_1280),
.A2(n_668),
.B1(n_627),
.B2(n_971),
.C(n_605),
.Y(n_1320)
);

OAI222xp33_ASAP7_75t_L g1321 ( 
.A1(n_1288),
.A2(n_630),
.B1(n_636),
.B2(n_675),
.C1(n_626),
.C2(n_1082),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_SL g1322 ( 
.A1(n_1296),
.A2(n_1215),
.B1(n_1192),
.B2(n_1212),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1286),
.A2(n_673),
.B1(n_666),
.B2(n_630),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1253),
.A2(n_673),
.B1(n_626),
.B2(n_1212),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1255),
.A2(n_1212),
.B1(n_1215),
.B2(n_961),
.Y(n_1325)
);

OAI21xp5_ASAP7_75t_SL g1326 ( 
.A1(n_1256),
.A2(n_668),
.B(n_1230),
.Y(n_1326)
);

AOI22xp33_ASAP7_75t_SL g1327 ( 
.A1(n_1239),
.A2(n_1192),
.B1(n_1222),
.B2(n_1204),
.Y(n_1327)
);

OAI22xp33_ASAP7_75t_L g1328 ( 
.A1(n_1257),
.A2(n_1192),
.B1(n_1231),
.B2(n_1198),
.Y(n_1328)
);

NAND3xp33_ASAP7_75t_L g1329 ( 
.A(n_1282),
.B(n_638),
.C(n_580),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1275),
.A2(n_961),
.B1(n_1048),
.B2(n_1041),
.Y(n_1330)
);

AOI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1276),
.A2(n_961),
.B1(n_1048),
.B2(n_1041),
.Y(n_1331)
);

AOI22xp33_ASAP7_75t_L g1332 ( 
.A1(n_1295),
.A2(n_961),
.B1(n_1100),
.B2(n_1160),
.Y(n_1332)
);

AOI22xp33_ASAP7_75t_L g1333 ( 
.A1(n_1267),
.A2(n_961),
.B1(n_1100),
.B2(n_1160),
.Y(n_1333)
);

NAND3xp33_ASAP7_75t_L g1334 ( 
.A(n_1254),
.B(n_580),
.C(n_571),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1267),
.A2(n_571),
.B1(n_585),
.B2(n_968),
.Y(n_1335)
);

OAI22xp33_ASAP7_75t_L g1336 ( 
.A1(n_1249),
.A2(n_1198),
.B1(n_1187),
.B2(n_1172),
.Y(n_1336)
);

OAI22x1_ASAP7_75t_L g1337 ( 
.A1(n_1245),
.A2(n_962),
.B1(n_968),
.B2(n_1128),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1298),
.A2(n_1161),
.B1(n_1204),
.B2(n_1222),
.Y(n_1338)
);

AOI22x1_ASAP7_75t_L g1339 ( 
.A1(n_1258),
.A2(n_1144),
.B1(n_1139),
.B2(n_1161),
.Y(n_1339)
);

AOI222xp33_ASAP7_75t_L g1340 ( 
.A1(n_1247),
.A2(n_962),
.B1(n_981),
.B2(n_776),
.C1(n_762),
.C2(n_685),
.Y(n_1340)
);

AOI22xp33_ASAP7_75t_SL g1341 ( 
.A1(n_1299),
.A2(n_1222),
.B1(n_1204),
.B2(n_1198),
.Y(n_1341)
);

OAI221xp5_ASAP7_75t_SL g1342 ( 
.A1(n_1294),
.A2(n_1106),
.B1(n_1132),
.B2(n_1141),
.C(n_1158),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1264),
.B(n_1106),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1263),
.B(n_1132),
.Y(n_1344)
);

AOI22xp33_ASAP7_75t_L g1345 ( 
.A1(n_1278),
.A2(n_1053),
.B1(n_1176),
.B2(n_1141),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1251),
.A2(n_1158),
.B1(n_1139),
.B2(n_1144),
.Y(n_1346)
);

OAI222xp33_ASAP7_75t_L g1347 ( 
.A1(n_1294),
.A2(n_701),
.B1(n_685),
.B2(n_690),
.C1(n_696),
.C2(n_1128),
.Y(n_1347)
);

OAI222xp33_ASAP7_75t_L g1348 ( 
.A1(n_1259),
.A2(n_701),
.B1(n_696),
.B2(n_690),
.C1(n_1144),
.C2(n_1117),
.Y(n_1348)
);

AOI22xp33_ASAP7_75t_L g1349 ( 
.A1(n_1271),
.A2(n_1176),
.B1(n_1187),
.B2(n_1172),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1274),
.A2(n_1187),
.B1(n_1065),
.B2(n_1088),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1285),
.Y(n_1351)
);

AOI22xp33_ASAP7_75t_L g1352 ( 
.A1(n_1279),
.A2(n_1065),
.B1(n_701),
.B2(n_696),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1287),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1262),
.A2(n_1133),
.B1(n_1117),
.B2(n_1148),
.Y(n_1354)
);

OAI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1283),
.A2(n_1157),
.B1(n_1156),
.B2(n_1148),
.Y(n_1355)
);

OAI22xp5_ASAP7_75t_L g1356 ( 
.A1(n_1283),
.A2(n_1157),
.B1(n_1156),
.B2(n_1148),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1289),
.A2(n_690),
.B1(n_1156),
.B2(n_1148),
.Y(n_1357)
);

OAI21xp33_ASAP7_75t_L g1358 ( 
.A1(n_1292),
.A2(n_63),
.B(n_67),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1290),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1285),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1261),
.B(n_1109),
.Y(n_1361)
);

INVx1_ASAP7_75t_SL g1362 ( 
.A(n_1284),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1300),
.A2(n_1157),
.B1(n_1156),
.B2(n_1147),
.Y(n_1363)
);

OAI22xp5_ASAP7_75t_L g1364 ( 
.A1(n_1291),
.A2(n_1157),
.B1(n_1147),
.B2(n_1145),
.Y(n_1364)
);

OAI22xp5_ASAP7_75t_L g1365 ( 
.A1(n_1244),
.A2(n_1147),
.B1(n_1145),
.B2(n_1134),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1297),
.A2(n_1147),
.B1(n_1145),
.B2(n_1134),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1285),
.Y(n_1367)
);

OAI22xp5_ASAP7_75t_L g1368 ( 
.A1(n_1244),
.A2(n_1145),
.B1(n_1134),
.B2(n_1131),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1307),
.B(n_1285),
.Y(n_1369)
);

NAND2xp5_ASAP7_75t_L g1370 ( 
.A(n_1343),
.B(n_1285),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1308),
.B(n_1285),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1308),
.B(n_1299),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1353),
.B(n_1273),
.Y(n_1373)
);

AND2x2_ASAP7_75t_L g1374 ( 
.A(n_1362),
.B(n_1236),
.Y(n_1374)
);

NAND2xp5_ASAP7_75t_L g1375 ( 
.A(n_1353),
.B(n_1270),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1359),
.B(n_1301),
.Y(n_1376)
);

AND2x2_ASAP7_75t_L g1377 ( 
.A(n_1359),
.B(n_1301),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1351),
.B(n_1301),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1361),
.B(n_1301),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1312),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_SL g1381 ( 
.A1(n_1313),
.A2(n_1272),
.B1(n_1242),
.B2(n_437),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1344),
.B(n_70),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_L g1383 ( 
.A(n_1312),
.B(n_70),
.Y(n_1383)
);

NOR2xp33_ASAP7_75t_L g1384 ( 
.A(n_1326),
.B(n_1272),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1318),
.B(n_1109),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1360),
.B(n_1109),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_L g1387 ( 
.A(n_1304),
.B(n_1328),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1327),
.B(n_1336),
.Y(n_1388)
);

OAI21xp5_ASAP7_75t_SL g1389 ( 
.A1(n_1303),
.A2(n_1242),
.B(n_73),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1351),
.B(n_74),
.Y(n_1390)
);

AND2x2_ASAP7_75t_L g1391 ( 
.A(n_1360),
.B(n_1119),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1360),
.B(n_1119),
.Y(n_1392)
);

AOI221xp5_ASAP7_75t_L g1393 ( 
.A1(n_1302),
.A2(n_623),
.B1(n_602),
.B2(n_600),
.C(n_591),
.Y(n_1393)
);

NOR2xp33_ASAP7_75t_R g1394 ( 
.A(n_1332),
.B(n_1119),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_SL g1395 ( 
.A(n_1322),
.B(n_1122),
.Y(n_1395)
);

OAI21xp5_ASAP7_75t_SL g1396 ( 
.A1(n_1358),
.A2(n_74),
.B(n_75),
.Y(n_1396)
);

AOI221xp5_ASAP7_75t_L g1397 ( 
.A1(n_1358),
.A2(n_602),
.B1(n_623),
.B2(n_591),
.C(n_600),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1366),
.B(n_78),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1340),
.A2(n_1134),
.B1(n_1131),
.B2(n_1124),
.C(n_1122),
.Y(n_1399)
);

NOR3xp33_ASAP7_75t_L g1400 ( 
.A(n_1342),
.B(n_79),
.C(n_80),
.Y(n_1400)
);

OAI221xp5_ASAP7_75t_L g1401 ( 
.A1(n_1320),
.A2(n_1131),
.B1(n_1124),
.B2(n_1122),
.C(n_83),
.Y(n_1401)
);

OAI221xp5_ASAP7_75t_L g1402 ( 
.A1(n_1349),
.A2(n_1131),
.B1(n_1124),
.B2(n_81),
.C(n_84),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1317),
.A2(n_437),
.B1(n_1124),
.B2(n_632),
.Y(n_1403)
);

NOR2xp33_ASAP7_75t_L g1404 ( 
.A(n_1365),
.B(n_79),
.Y(n_1404)
);

OAI221xp5_ASAP7_75t_SL g1405 ( 
.A1(n_1309),
.A2(n_80),
.B1(n_81),
.B2(n_84),
.C(n_85),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1367),
.B(n_86),
.Y(n_1406)
);

OAI21xp5_ASAP7_75t_SL g1407 ( 
.A1(n_1341),
.A2(n_1305),
.B(n_1347),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1345),
.A2(n_1310),
.B1(n_1333),
.B2(n_1306),
.Y(n_1408)
);

NAND3xp33_ASAP7_75t_L g1409 ( 
.A(n_1329),
.B(n_1334),
.C(n_1367),
.Y(n_1409)
);

NOR3xp33_ASAP7_75t_L g1410 ( 
.A(n_1368),
.B(n_87),
.C(n_88),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1354),
.B(n_437),
.Y(n_1411)
);

OAI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1314),
.A2(n_606),
.B1(n_632),
.B2(n_591),
.Y(n_1412)
);

AOI221xp5_ASAP7_75t_L g1413 ( 
.A1(n_1337),
.A2(n_637),
.B1(n_632),
.B2(n_628),
.C(n_606),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1315),
.B(n_588),
.Y(n_1414)
);

NOR3xp33_ASAP7_75t_L g1415 ( 
.A(n_1396),
.B(n_1356),
.C(n_1355),
.Y(n_1415)
);

NAND3xp33_ASAP7_75t_L g1416 ( 
.A(n_1400),
.B(n_1339),
.C(n_1319),
.Y(n_1416)
);

BUFx2_ASAP7_75t_L g1417 ( 
.A(n_1378),
.Y(n_1417)
);

NAND3xp33_ASAP7_75t_L g1418 ( 
.A(n_1410),
.B(n_1339),
.C(n_1363),
.Y(n_1418)
);

AO21x2_ASAP7_75t_L g1419 ( 
.A1(n_1414),
.A2(n_1364),
.B(n_1348),
.Y(n_1419)
);

AND2x4_ASAP7_75t_L g1420 ( 
.A(n_1377),
.B(n_1325),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1373),
.B(n_1338),
.Y(n_1421)
);

NAND4xp75_ASAP7_75t_L g1422 ( 
.A(n_1387),
.B(n_1337),
.C(n_1321),
.D(n_1357),
.Y(n_1422)
);

AOI221xp5_ASAP7_75t_L g1423 ( 
.A1(n_1389),
.A2(n_1335),
.B1(n_1323),
.B2(n_1346),
.C(n_1316),
.Y(n_1423)
);

BUFx2_ASAP7_75t_SL g1424 ( 
.A(n_1377),
.Y(n_1424)
);

OAI211xp5_ASAP7_75t_SL g1425 ( 
.A1(n_1372),
.A2(n_1352),
.B(n_1330),
.C(n_1331),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1380),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1378),
.B(n_1350),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1380),
.B(n_1324),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1385),
.B(n_1311),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1369),
.B(n_637),
.Y(n_1430)
);

NOR3xp33_ASAP7_75t_L g1431 ( 
.A(n_1405),
.B(n_101),
.C(n_102),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1390),
.B(n_588),
.Y(n_1432)
);

NAND4xp75_ASAP7_75t_L g1433 ( 
.A(n_1411),
.B(n_105),
.C(n_108),
.D(n_111),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1375),
.Y(n_1434)
);

AOI221xp5_ASAP7_75t_L g1435 ( 
.A1(n_1383),
.A2(n_637),
.B1(n_628),
.B2(n_606),
.C(n_600),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1371),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1370),
.B(n_112),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1376),
.Y(n_1438)
);

NAND3xp33_ASAP7_75t_L g1439 ( 
.A(n_1382),
.B(n_1406),
.C(n_1404),
.Y(n_1439)
);

NOR2x1_ASAP7_75t_L g1440 ( 
.A(n_1409),
.B(n_113),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1379),
.B(n_116),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1386),
.B(n_117),
.Y(n_1442)
);

AOI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1422),
.A2(n_1407),
.B1(n_1388),
.B2(n_1411),
.Y(n_1443)
);

XOR2x2_ASAP7_75t_L g1444 ( 
.A(n_1422),
.B(n_1374),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1417),
.B(n_1391),
.Y(n_1445)
);

XOR2x2_ASAP7_75t_L g1446 ( 
.A(n_1439),
.B(n_1399),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1436),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1434),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1417),
.B(n_1392),
.Y(n_1449)
);

NAND4xp75_ASAP7_75t_L g1450 ( 
.A(n_1440),
.B(n_1395),
.C(n_1384),
.D(n_1404),
.Y(n_1450)
);

NAND4xp75_ASAP7_75t_L g1451 ( 
.A(n_1421),
.B(n_1395),
.C(n_1384),
.D(n_1397),
.Y(n_1451)
);

XOR2x2_ASAP7_75t_L g1452 ( 
.A(n_1431),
.B(n_1402),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1438),
.B(n_1398),
.Y(n_1453)
);

NAND4xp75_ASAP7_75t_SL g1454 ( 
.A(n_1430),
.B(n_1381),
.C(n_1401),
.D(n_1394),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1427),
.Y(n_1455)
);

HB1xp67_ASAP7_75t_L g1456 ( 
.A(n_1430),
.Y(n_1456)
);

XNOR2xp5_ASAP7_75t_L g1457 ( 
.A(n_1427),
.B(n_1408),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1420),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1413),
.B2(n_1393),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1438),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1424),
.B(n_1394),
.Y(n_1461)
);

XNOR2xp5_ASAP7_75t_L g1462 ( 
.A(n_1420),
.B(n_1403),
.Y(n_1462)
);

INVx2_ASAP7_75t_L g1463 ( 
.A(n_1426),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1447),
.Y(n_1464)
);

INVxp67_ASAP7_75t_L g1465 ( 
.A(n_1456),
.Y(n_1465)
);

INVxp67_ASAP7_75t_L g1466 ( 
.A(n_1456),
.Y(n_1466)
);

INVxp67_ASAP7_75t_L g1467 ( 
.A(n_1450),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1448),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1455),
.Y(n_1469)
);

OA22x2_ASAP7_75t_L g1470 ( 
.A1(n_1443),
.A2(n_1457),
.B1(n_1462),
.B2(n_1444),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1449),
.B(n_1424),
.Y(n_1471)
);

XOR2x2_ASAP7_75t_L g1472 ( 
.A(n_1444),
.B(n_1415),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1445),
.Y(n_1473)
);

XNOR2xp5_ASAP7_75t_L g1474 ( 
.A(n_1446),
.B(n_1420),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1455),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1449),
.B(n_1442),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1453),
.Y(n_1477)
);

INVx2_ASAP7_75t_L g1478 ( 
.A(n_1458),
.Y(n_1478)
);

AO22x2_ASAP7_75t_L g1479 ( 
.A1(n_1458),
.A2(n_1428),
.B1(n_1429),
.B2(n_1416),
.Y(n_1479)
);

XOR2x2_ASAP7_75t_L g1480 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1480)
);

XOR2x2_ASAP7_75t_L g1481 ( 
.A(n_1452),
.B(n_1433),
.Y(n_1481)
);

OAI22x1_ASAP7_75t_L g1482 ( 
.A1(n_1474),
.A2(n_1461),
.B1(n_1460),
.B2(n_1459),
.Y(n_1482)
);

AOI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1480),
.A2(n_1451),
.B1(n_1425),
.B2(n_1429),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1464),
.Y(n_1484)
);

BUFx3_ASAP7_75t_L g1485 ( 
.A(n_1469),
.Y(n_1485)
);

OAI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1467),
.A2(n_1479),
.B1(n_1470),
.B2(n_1469),
.Y(n_1486)
);

NOR2xp33_ASAP7_75t_L g1487 ( 
.A(n_1467),
.B(n_1437),
.Y(n_1487)
);

OA22x2_ASAP7_75t_L g1488 ( 
.A1(n_1475),
.A2(n_1441),
.B1(n_1463),
.B2(n_1454),
.Y(n_1488)
);

OA22x2_ASAP7_75t_L g1489 ( 
.A1(n_1475),
.A2(n_1441),
.B1(n_1463),
.B2(n_1432),
.Y(n_1489)
);

AOI22x1_ASAP7_75t_L g1490 ( 
.A1(n_1479),
.A2(n_1428),
.B1(n_1423),
.B2(n_1419),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1480),
.Y(n_1491)
);

OA22x2_ASAP7_75t_L g1492 ( 
.A1(n_1472),
.A2(n_1419),
.B1(n_1412),
.B2(n_1435),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1465),
.B(n_118),
.Y(n_1493)
);

AOI22x1_ASAP7_75t_L g1494 ( 
.A1(n_1479),
.A2(n_1465),
.B1(n_1466),
.B2(n_1481),
.Y(n_1494)
);

OA22x2_ASAP7_75t_L g1495 ( 
.A1(n_1478),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_1495)
);

AOI22x1_ASAP7_75t_SL g1496 ( 
.A1(n_1481),
.A2(n_127),
.B1(n_130),
.B2(n_132),
.Y(n_1496)
);

CKINVDCx16_ASAP7_75t_R g1497 ( 
.A(n_1476),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1491),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1484),
.Y(n_1499)
);

XNOR2xp5_ASAP7_75t_L g1500 ( 
.A(n_1496),
.B(n_1470),
.Y(n_1500)
);

BUFx2_ASAP7_75t_L g1501 ( 
.A(n_1485),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1493),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1489),
.Y(n_1503)
);

OAI322xp33_ASAP7_75t_L g1504 ( 
.A1(n_1494),
.A2(n_1466),
.A3(n_1468),
.B1(n_1477),
.B2(n_1473),
.C1(n_1471),
.C2(n_143),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1486),
.Y(n_1505)
);

INVxp33_ASAP7_75t_SL g1506 ( 
.A(n_1496),
.Y(n_1506)
);

AOI211x1_ASAP7_75t_SL g1507 ( 
.A1(n_1504),
.A2(n_1490),
.B(n_1482),
.C(n_1488),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1499),
.Y(n_1508)
);

OAI322xp33_ASAP7_75t_L g1509 ( 
.A1(n_1505),
.A2(n_1490),
.A3(n_1483),
.B1(n_1492),
.B2(n_1487),
.C1(n_1497),
.C2(n_1495),
.Y(n_1509)
);

AOI22xp5_ASAP7_75t_L g1510 ( 
.A1(n_1506),
.A2(n_631),
.B1(n_147),
.B2(n_148),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1501),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1498),
.Y(n_1512)
);

AOI221xp5_ASAP7_75t_L g1513 ( 
.A1(n_1509),
.A2(n_1500),
.B1(n_1498),
.B2(n_1503),
.C(n_1502),
.Y(n_1513)
);

NAND4xp25_ASAP7_75t_SL g1514 ( 
.A(n_1512),
.B(n_1511),
.C(n_1507),
.D(n_1508),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1510),
.B(n_150),
.Y(n_1515)
);

NOR3xp33_ASAP7_75t_L g1516 ( 
.A(n_1515),
.B(n_156),
.C(n_164),
.Y(n_1516)
);

NOR4xp25_ASAP7_75t_L g1517 ( 
.A(n_1514),
.B(n_172),
.C(n_179),
.D(n_181),
.Y(n_1517)
);

NOR2x1_ASAP7_75t_L g1518 ( 
.A(n_1514),
.B(n_183),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_SL g1519 ( 
.A(n_1513),
.B(n_185),
.Y(n_1519)
);

NOR2x2_ASAP7_75t_L g1520 ( 
.A(n_1517),
.B(n_190),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1518),
.Y(n_1521)
);

INVxp67_ASAP7_75t_L g1522 ( 
.A(n_1519),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1516),
.Y(n_1523)
);

INVxp67_ASAP7_75t_SL g1524 ( 
.A(n_1521),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1523),
.Y(n_1525)
);

CKINVDCx20_ASAP7_75t_R g1526 ( 
.A(n_1522),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1520),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1524),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1526),
.Y(n_1529)
);

INVx3_ASAP7_75t_L g1530 ( 
.A(n_1527),
.Y(n_1530)
);

HB1xp67_ASAP7_75t_L g1531 ( 
.A(n_1525),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1527),
.Y(n_1532)
);

OAI22x1_ASAP7_75t_L g1533 ( 
.A1(n_1529),
.A2(n_193),
.B1(n_196),
.B2(n_200),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1530),
.A2(n_202),
.B1(n_203),
.B2(n_207),
.Y(n_1534)
);

INVx1_ASAP7_75t_SL g1535 ( 
.A(n_1531),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1530),
.A2(n_208),
.B1(n_210),
.B2(n_211),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1532),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1528),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1530),
.A2(n_233),
.B1(n_235),
.B2(n_236),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1529),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1535),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1540),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1538),
.Y(n_1543)
);

INVx2_ASAP7_75t_L g1544 ( 
.A(n_1533),
.Y(n_1544)
);

AO22x2_ASAP7_75t_L g1545 ( 
.A1(n_1541),
.A2(n_1539),
.B1(n_1536),
.B2(n_1537),
.Y(n_1545)
);

AOI31xp33_ASAP7_75t_L g1546 ( 
.A1(n_1543),
.A2(n_1534),
.A3(n_238),
.B(n_240),
.Y(n_1546)
);

NAND4xp25_ASAP7_75t_L g1547 ( 
.A(n_1542),
.B(n_237),
.C(n_242),
.D(n_243),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1544),
.A2(n_244),
.B1(n_247),
.B2(n_249),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1545),
.Y(n_1549)
);

BUFx2_ASAP7_75t_L g1550 ( 
.A(n_1547),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1546),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1548),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_SL g1553 ( 
.A1(n_1549),
.A2(n_1550),
.B1(n_1552),
.B2(n_253),
.Y(n_1553)
);

AOI22xp5_ASAP7_75t_L g1554 ( 
.A1(n_1551),
.A2(n_251),
.B1(n_252),
.B2(n_255),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1549),
.A2(n_257),
.B1(n_259),
.B2(n_269),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1553),
.Y(n_1556)
);

AOI221xp5_ASAP7_75t_L g1557 ( 
.A1(n_1556),
.A2(n_1555),
.B1(n_1554),
.B2(n_273),
.C(n_281),
.Y(n_1557)
);

AOI211xp5_ASAP7_75t_L g1558 ( 
.A1(n_1557),
.A2(n_289),
.B(n_290),
.C(n_292),
.Y(n_1558)
);


endmodule