module fake_jpeg_13556_n_289 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_289);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_289;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_19;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_127;
wire n_154;
wire n_76;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_266;
wire n_218;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_100;
wire n_128;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx5_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx10_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx6_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_1),
.Y(n_42)
);

OR2x2_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_44),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_27),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_1),
.B(n_2),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_45),
.B(n_7),
.C(n_8),
.Y(n_108)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_1),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_48),
.B(n_49),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_2),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_3),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_51),
.B(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_55),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_19),
.B(n_17),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_56),
.B(n_58),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_57),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_19),
.B(n_17),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_18),
.Y(n_59)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_41),
.B(n_5),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_61),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_23),
.Y(n_62)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_29),
.B(n_5),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_63),
.B(n_66),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_30),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_33),
.Y(n_88)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_25),
.Y(n_65)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_29),
.B(n_6),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g68 ( 
.A(n_31),
.Y(n_68)
);

INVx6_ASAP7_75t_SL g80 ( 
.A(n_68),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_54),
.A2(n_26),
.B1(n_31),
.B2(n_37),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_41),
.B1(n_28),
.B2(n_33),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_71),
.A2(n_81),
.B1(n_90),
.B2(n_105),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_26),
.B1(n_30),
.B2(n_37),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_74),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_50),
.A2(n_37),
.B1(n_30),
.B2(n_27),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g125 ( 
.A(n_75),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g81 ( 
.A1(n_47),
.A2(n_33),
.B1(n_28),
.B2(n_27),
.Y(n_81)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_89),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_88),
.B(n_108),
.Y(n_137)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_52),
.B(n_27),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_53),
.A2(n_42),
.B1(n_39),
.B2(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_65),
.Y(n_92)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_43),
.B(n_42),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_93),
.B(n_96),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_46),
.A2(n_35),
.B1(n_24),
.B2(n_36),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g136 ( 
.A(n_94),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_48),
.B(n_39),
.Y(n_96)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_57),
.Y(n_102)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_103),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_38),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_104),
.B(n_7),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_62),
.A2(n_36),
.B1(n_32),
.B2(n_25),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_64),
.A2(n_32),
.B1(n_20),
.B2(n_18),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_106),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_51),
.A2(n_20),
.B1(n_25),
.B2(n_9),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_107),
.B(n_109),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_59),
.B(n_25),
.Y(n_109)
);

INVx4_ASAP7_75t_SL g110 ( 
.A(n_67),
.Y(n_110)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_110),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_112),
.B(n_118),
.Y(n_174)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_113),
.Y(n_167)
);

A2O1A1Ixp33_ASAP7_75t_L g114 ( 
.A1(n_86),
.A2(n_7),
.B(n_8),
.C(n_9),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_114),
.B(n_139),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_99),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g172 ( 
.A(n_117),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_84),
.Y(n_118)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_95),
.B(n_9),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_126),
.Y(n_162)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_91),
.Y(n_127)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_127),
.Y(n_148)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_99),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_132),
.Y(n_170)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_80),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_135),
.B(n_140),
.Y(n_150)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_138),
.B(n_110),
.Y(n_155)
);

A2O1A1Ixp33_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_84),
.B(n_89),
.C(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_91),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_80),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_141),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_88),
.A2(n_10),
.B(n_12),
.C(n_13),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_143),
.B(n_73),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_69),
.C(n_14),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_144),
.B(n_137),
.C(n_142),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_82),
.B(n_12),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_72),
.Y(n_161)
);

INVx3_ASAP7_75t_SL g146 ( 
.A(n_101),
.Y(n_146)
);

INVxp33_ASAP7_75t_L g153 ( 
.A(n_146),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_121),
.Y(n_198)
);

XNOR2x1_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_139),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_149),
.B(n_158),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_142),
.A2(n_98),
.B1(n_77),
.B2(n_85),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_154),
.A2(n_165),
.B(n_123),
.Y(n_185)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_155),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_124),
.A2(n_100),
.B1(n_101),
.B2(n_111),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_96),
.B1(n_103),
.B2(n_76),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_164),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_129),
.A2(n_98),
.B1(n_85),
.B2(n_97),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_160),
.A2(n_131),
.B(n_123),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_161),
.B(n_119),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_129),
.A2(n_76),
.B1(n_79),
.B2(n_72),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_115),
.A2(n_79),
.B(n_87),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_137),
.B(n_111),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_166),
.B(n_168),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_144),
.B(n_87),
.C(n_15),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_14),
.C(n_16),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_169),
.B(n_176),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_134),
.A2(n_14),
.B1(n_120),
.B2(n_124),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_169),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_120),
.A2(n_143),
.B1(n_114),
.B2(n_116),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_164),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_163),
.B(n_117),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_180),
.B(n_182),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_184),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_198),
.B(n_199),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_128),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_190),
.Y(n_207)
);

A2O1A1Ixp33_ASAP7_75t_L g188 ( 
.A1(n_173),
.A2(n_138),
.B(n_113),
.C(n_146),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_188),
.B(n_165),
.Y(n_211)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_189),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_155),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_170),
.Y(n_192)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_192),
.Y(n_218)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_175),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_194),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_156),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_155),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_200),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_196),
.B(n_197),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_166),
.A2(n_133),
.B(n_122),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_151),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_201),
.B(n_202),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_151),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_167),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_179),
.A2(n_158),
.B1(n_173),
.B2(n_171),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_205),
.A2(n_212),
.B1(n_217),
.B2(n_190),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_209),
.A2(n_211),
.B(n_172),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_149),
.C(n_186),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_224),
.C(n_194),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_160),
.B1(n_168),
.B2(n_159),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_185),
.A2(n_147),
.B(n_153),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_213),
.A2(n_215),
.B(n_222),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_198),
.A2(n_153),
.B(n_162),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_183),
.A2(n_174),
.B1(n_122),
.B2(n_130),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_219),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g221 ( 
.A1(n_191),
.A2(n_119),
.A3(n_132),
.B1(n_172),
.B2(n_186),
.C1(n_177),
.C2(n_196),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_221),
.B(n_197),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_199),
.B(n_191),
.C(n_181),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_211),
.A2(n_183),
.B1(n_181),
.B2(n_188),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_225),
.A2(n_212),
.B1(n_224),
.B2(n_209),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_226),
.B(n_228),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_213),
.Y(n_227)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_205),
.A2(n_195),
.B1(n_200),
.B2(n_184),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_216),
.B1(n_204),
.B2(n_206),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_231),
.B(n_233),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_209),
.B(n_178),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_207),
.B(n_202),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_232),
.B(n_239),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_214),
.A2(n_189),
.B(n_192),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_203),
.B1(n_193),
.B2(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_235),
.B(n_240),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_236),
.B(n_238),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_201),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_201),
.B(n_215),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_207),
.Y(n_241)
);

INVxp33_ASAP7_75t_L g247 ( 
.A(n_241),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_246),
.A2(n_252),
.B1(n_228),
.B2(n_233),
.Y(n_258)
);

XNOR2x1_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_214),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_249),
.B(n_253),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_240),
.A2(n_217),
.B1(n_220),
.B2(n_204),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_253),
.B(n_232),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_254),
.B(n_257),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_236),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_255),
.B(n_256),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_230),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_229),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_258),
.A2(n_250),
.B1(n_231),
.B2(n_244),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_252),
.A2(n_237),
.B1(n_227),
.B2(n_223),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_259),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_235),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_260),
.B(n_262),
.Y(n_269)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_225),
.CI(n_231),
.CON(n_261),
.SN(n_261)
);

AOI21xp5_ASAP7_75t_L g271 ( 
.A1(n_261),
.A2(n_250),
.B(n_247),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_243),
.C(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_262),
.Y(n_265)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_265),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_267),
.B(n_270),
.Y(n_273)
);

AOI21x1_ASAP7_75t_SL g276 ( 
.A1(n_271),
.A2(n_263),
.B(n_223),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_267),
.A2(n_247),
.B(n_261),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_275),
.Y(n_278)
);

NAND4xp25_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_237),
.C(n_256),
.D(n_260),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_276),
.B(n_269),
.Y(n_281)
);

OAI221xp5_ASAP7_75t_L g277 ( 
.A1(n_264),
.A2(n_255),
.B1(n_218),
.B2(n_206),
.C(n_208),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_277),
.B(n_270),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_280),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_268),
.C(n_269),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_281),
.B(n_276),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_282),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_278),
.C(n_272),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_284),
.B(n_268),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_286),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_287),
.A2(n_283),
.B(n_208),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_288),
.B(n_218),
.Y(n_289)
);


endmodule