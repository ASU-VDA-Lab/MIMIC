module real_jpeg_909_n_13 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_13);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_13;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_126;
wire n_113;
wire n_120;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_135;
wire n_134;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_1),
.A2(n_23),
.B1(n_24),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_26),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_4),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_54),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g30 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_5),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_5),
.A2(n_31),
.B1(n_37),
.B2(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_7),
.A2(n_33),
.B(n_34),
.C(n_40),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_7),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_7),
.B(n_59),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_7),
.B(n_24),
.C(n_48),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_7),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_7),
.B(n_21),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_7),
.B(n_69),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_52),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_52),
.Y(n_126)
);

BUFx10_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_11),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_91),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_90),
.Y(n_14)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_16),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_63),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_17),
.B(n_63),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_44),
.C(n_55),
.Y(n_17)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_18),
.B(n_104),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_32),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_32),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B(n_27),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_24),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_20),
.A2(n_22),
.B1(n_29),
.B2(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_20),
.B(n_30),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_20),
.A2(n_29),
.B1(n_100),
.B2(n_131),
.Y(n_130)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_21),
.A2(n_28),
.B(n_126),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g50 ( 
.A1(n_23),
.A2(n_24),
.B1(n_48),
.B2(n_49),
.Y(n_50)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_24),
.B(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_30),
.Y(n_28)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_29),
.A2(n_100),
.B(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_29),
.Y(n_123)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

O2A1O1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_40),
.B(n_58),
.C(n_59),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_33),
.B(n_40),
.Y(n_58)
);

AO22x1_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_36),
.B(n_37),
.Y(n_34)
);

AOI21xp5_ASAP7_75t_L g122 ( 
.A1(n_36),
.A2(n_102),
.B(n_123),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_38),
.B1(n_48),
.B2(n_49),
.Y(n_47)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_38),
.B(n_110),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OA22x2_ASAP7_75t_L g82 ( 
.A1(n_40),
.A2(n_41),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_44),
.B(n_55),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_50),
.B1(n_51),
.B2(n_53),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_45),
.A2(n_68),
.B(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_46),
.A2(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_46),
.B(n_70),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

INVx13_ASAP7_75t_L g49 ( 
.A(n_48),
.Y(n_49)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_51),
.B(n_96),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_61),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_57),
.B(n_62),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_59),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_72),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_71),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_78),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_77),
.Y(n_73)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_86),
.B2(n_87),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g85 ( 
.A(n_83),
.Y(n_85)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_105),
.B(n_136),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_103),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_97),
.C(n_98),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_95),
.B1(n_97),
.B2(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_98),
.A2(n_99),
.B1(n_114),
.B2(n_116),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_117),
.B(n_135),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_113),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_113),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_111),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_108),
.A2(n_109),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_129),
.B(n_134),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g118 ( 
.A1(n_119),
.A2(n_124),
.B(n_128),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_120),
.B(n_122),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_127),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_126),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_132),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_132),
.Y(n_134)
);


endmodule