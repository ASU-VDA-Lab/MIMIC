module fake_jpeg_30400_n_339 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_339);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_8),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_14),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_11),
.Y(n_37)
);

BUFx8_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_3),
.B(n_9),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_49),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_52),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_53),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g82 ( 
.A(n_56),
.Y(n_82)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g112 ( 
.A(n_57),
.Y(n_112)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_58),
.Y(n_91)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx3_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_62),
.B(n_64),
.Y(n_94)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_7),
.Y(n_64)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_67),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_23),
.Y(n_68)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_69),
.Y(n_105)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_25),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_73),
.Y(n_98)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_79),
.Y(n_90)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_75),
.B(n_77),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_38),
.Y(n_77)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_37),
.B(n_7),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_62),
.A2(n_24),
.B1(n_26),
.B2(n_40),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_100),
.B(n_106),
.Y(n_119)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_0),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_64),
.B(n_45),
.C(n_43),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_116),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_80),
.A2(n_21),
.B1(n_31),
.B2(n_30),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g117 ( 
.A(n_111),
.B(n_21),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_66),
.B(n_31),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_117),
.B(n_120),
.Y(n_149)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_85),
.Y(n_118)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_81),
.Y(n_120)
);

CKINVDCx5p33_ASAP7_75t_R g121 ( 
.A(n_89),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_121),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_122),
.Y(n_156)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_103),
.Y(n_123)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_123),
.Y(n_162)
);

INVx8_ASAP7_75t_L g124 ( 
.A(n_103),
.Y(n_124)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_124),
.Y(n_164)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_95),
.A2(n_53),
.B1(n_48),
.B2(n_49),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_125),
.A2(n_138),
.B1(n_144),
.B2(n_146),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_102),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_126),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_50),
.B1(n_71),
.B2(n_68),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_127),
.A2(n_145),
.B1(n_112),
.B2(n_89),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_131),
.Y(n_151)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_132),
.B(n_133),
.Y(n_153)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_92),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_134),
.Y(n_160)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_137),
.B1(n_141),
.B2(n_143),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_106),
.B(n_35),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_136),
.B(n_142),
.Y(n_161)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_98),
.Y(n_137)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_114),
.A2(n_115),
.B1(n_73),
.B2(n_54),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_106),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_139),
.B(n_140),
.Y(n_157)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_109),
.A2(n_70),
.B1(n_65),
.B2(n_60),
.Y(n_145)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_83),
.Y(n_146)
);

BUFx3_ASAP7_75t_L g147 ( 
.A(n_104),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_148),
.B1(n_84),
.B2(n_82),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_113),
.B(n_43),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_90),
.C(n_82),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_150),
.B(n_163),
.C(n_168),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_96),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_119),
.B(n_112),
.C(n_94),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_125),
.A2(n_114),
.B1(n_115),
.B2(n_108),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_167),
.A2(n_108),
.B1(n_122),
.B2(n_133),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_119),
.B(n_136),
.C(n_118),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_169),
.A2(n_132),
.B1(n_123),
.B2(n_147),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_117),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_179),
.Y(n_195)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_159),
.Y(n_171)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_171),
.Y(n_203)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_173),
.Y(n_188)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_174),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_142),
.C(n_129),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_175),
.B(n_161),
.C(n_157),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_176),
.A2(n_177),
.B1(n_183),
.B2(n_184),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_168),
.A2(n_134),
.B1(n_131),
.B2(n_83),
.Y(n_177)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_178),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_140),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_110),
.B1(n_143),
.B2(n_141),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_180),
.A2(n_185),
.B1(n_186),
.B2(n_154),
.Y(n_189)
);

INVx4_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_181),
.Y(n_192)
);

CKINVDCx14_ASAP7_75t_R g182 ( 
.A(n_158),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_182),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_163),
.A2(n_122),
.B1(n_135),
.B2(n_110),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_169),
.A2(n_137),
.B1(n_124),
.B2(n_40),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_163),
.B1(n_155),
.B2(n_167),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_187),
.A2(n_184),
.B1(n_178),
.B2(n_171),
.Y(n_210)
);

INVxp33_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_158),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_170),
.A2(n_175),
.B1(n_172),
.B2(n_180),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_200),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_172),
.B(n_150),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_198),
.B(n_183),
.Y(n_204)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_174),
.Y(n_199)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_185),
.A2(n_167),
.B1(n_161),
.B2(n_157),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_149),
.C(n_153),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_152),
.B1(n_151),
.B2(n_149),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_184),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_214),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_206),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_151),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_197),
.A2(n_154),
.B1(n_152),
.B2(n_177),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_209),
.A2(n_210),
.B1(n_215),
.B2(n_200),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_194),
.A2(n_184),
.B(n_164),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_211),
.A2(n_191),
.B(n_199),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_212),
.B(n_213),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_197),
.A2(n_176),
.B1(n_173),
.B2(n_153),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_195),
.B(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_217),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_203),
.Y(n_218)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_218),
.B(n_191),
.C(n_195),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_220),
.B(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_216),
.Y(n_223)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_223),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_209),
.A2(n_187),
.B1(n_196),
.B2(n_189),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_224),
.B(n_228),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_232),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_204),
.B(n_198),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_229),
.Y(n_237)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_216),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_230),
.Y(n_246)
);

NAND3xp33_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_202),
.C(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_201),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_217),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_228),
.B(n_204),
.C(n_214),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_235),
.B(n_238),
.C(n_239),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_236),
.B(n_192),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_219),
.B(n_205),
.C(n_210),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_205),
.C(n_213),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_227),
.B(n_215),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_240),
.B(n_242),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_225),
.A2(n_190),
.B(n_188),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g262 ( 
.A(n_241),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_211),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_232),
.B(n_211),
.C(n_212),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_162),
.C(n_192),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_221),
.A2(n_208),
.B1(n_218),
.B2(n_188),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_247),
.A2(n_222),
.B1(n_223),
.B2(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_243),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_244),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_250),
.B(n_253),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_237),
.A2(n_226),
.B1(n_222),
.B2(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_251),
.A2(n_166),
.B1(n_41),
.B2(n_28),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_239),
.B(n_164),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_265),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_260),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_246),
.B(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_257),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_245),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_259),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_235),
.B(n_162),
.Y(n_260)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_247),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_264),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_234),
.B(n_165),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_263),
.B(n_165),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_240),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_242),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_238),
.C(n_234),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_272),
.C(n_273),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_274),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_262),
.A2(n_181),
.B1(n_160),
.B2(n_26),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_270),
.A2(n_280),
.B1(n_91),
.B2(n_17),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_181),
.C(n_126),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_260),
.B(n_121),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_256),
.B(n_166),
.C(n_28),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_275),
.B(n_277),
.C(n_279),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_254),
.B(n_41),
.C(n_30),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_255),
.B(n_263),
.C(n_253),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_257),
.A2(n_24),
.B1(n_40),
.B2(n_35),
.Y(n_280)
);

OR2x2_ASAP7_75t_L g284 ( 
.A(n_282),
.B(n_251),
.Y(n_284)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_284),
.Y(n_299)
);

AOI22x1_ASAP7_75t_L g285 ( 
.A1(n_281),
.A2(n_261),
.B1(n_255),
.B2(n_96),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_285),
.A2(n_20),
.B1(n_6),
.B2(n_13),
.Y(n_306)
);

OAI21x1_ASAP7_75t_L g286 ( 
.A1(n_278),
.A2(n_14),
.B(n_13),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_279),
.B(n_110),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_290),
.C(n_55),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_288),
.B(n_289),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_276),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_266),
.B(n_89),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_294),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_272),
.A2(n_275),
.B(n_277),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_292),
.A2(n_296),
.B(n_284),
.Y(n_297)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_267),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_269),
.A2(n_91),
.B(n_12),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_297),
.B(n_300),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_293),
.A2(n_269),
.B(n_271),
.Y(n_298)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_298),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_283),
.A2(n_12),
.B1(n_19),
.B2(n_16),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_12),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_302),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_295),
.A2(n_6),
.B(n_19),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_307),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_295),
.A2(n_19),
.B(n_16),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_299),
.B(n_290),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_309),
.B(n_0),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_283),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_311),
.B(n_313),
.Y(n_319)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_285),
.B(n_287),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_312),
.A2(n_315),
.B(n_318),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_305),
.B(n_15),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_308),
.B(n_15),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_317),
.B(n_6),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_320),
.B(n_321),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_322),
.B(n_324),
.Y(n_330)
);

AOI21x1_ASAP7_75t_L g323 ( 
.A1(n_309),
.A2(n_0),
.B(n_1),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g328 ( 
.A1(n_323),
.A2(n_2),
.B(n_3),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_20),
.C(n_2),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_325),
.A2(n_4),
.B(n_5),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_20),
.B(n_2),
.Y(n_326)
);

O2A1O1Ixp33_ASAP7_75t_SL g327 ( 
.A1(n_326),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_319),
.Y(n_332)
);

O2A1O1Ixp33_ASAP7_75t_SL g333 ( 
.A1(n_328),
.A2(n_331),
.B(n_322),
.C(n_5),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_332),
.B(n_333),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_329),
.B(n_4),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_330),
.C(n_5),
.Y(n_335)
);

AOI21x1_ASAP7_75t_L g337 ( 
.A1(n_335),
.A2(n_4),
.B(n_5),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_336),
.B(n_4),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_20),
.Y(n_339)
);


endmodule