module real_jpeg_707_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_1),
.B(n_27),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_1),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_1),
.B(n_69),
.Y(n_139)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_2),
.B(n_35),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_2),
.B(n_42),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_2),
.B(n_27),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_67),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_2),
.B(n_32),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_4),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_4),
.B(n_39),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_4),
.B(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_4),
.B(n_45),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_4),
.B(n_42),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_4),
.B(n_67),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_4),
.B(n_27),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_4),
.B(n_32),
.Y(n_277)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_5),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_5),
.B(n_39),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_5),
.B(n_69),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_5),
.B(n_45),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_5),
.B(n_42),
.Y(n_271)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_6),
.Y(n_45)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_39),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_8),
.B(n_69),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_8),
.B(n_45),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_8),
.B(n_42),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_8),
.B(n_67),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_9),
.B(n_27),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_9),
.B(n_45),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_9),
.B(n_32),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_9),
.B(n_69),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_9),
.B(n_67),
.Y(n_103)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_9),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_10),
.B(n_27),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_10),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_10),
.B(n_32),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_10),
.B(n_42),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_10),
.B(n_45),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g67 ( 
.A(n_11),
.Y(n_67)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_12),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_13),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_14),
.B(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_45),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_14),
.B(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_14),
.B(n_42),
.Y(n_102)
);

AND2x2_ASAP7_75t_SL g117 ( 
.A(n_14),
.B(n_27),
.Y(n_117)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_14),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_14),
.B(n_67),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_14),
.B(n_35),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_168),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_166),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_19),
.B(n_132),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_80),
.C(n_113),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_20),
.A2(n_21),
.B1(n_113),
.B2(n_114),
.Y(n_172)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_57),
.B2(n_79),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_22),
.B(n_58),
.C(n_72),
.Y(n_133)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.C(n_46),
.Y(n_23)
);

FAx1_ASAP7_75t_SL g198 ( 
.A(n_24),
.B(n_37),
.CI(n_46),
.CON(n_198),
.SN(n_198)
);

XNOR2xp5_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_34),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_30),
.B1(n_31),
.B2(n_33),
.Y(n_25)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_26),
.B(n_31),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_26),
.A2(n_33),
.B1(n_184),
.B2(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_28),
.B(n_62),
.Y(n_275)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_30),
.A2(n_31),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

O2A1O1Ixp33_ASAP7_75t_L g124 ( 
.A1(n_30),
.A2(n_33),
.B(n_34),
.C(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_30),
.B(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_30),
.A2(n_31),
.B1(n_252),
.B2(n_253),
.Y(n_265)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_31),
.B(n_117),
.C(n_119),
.Y(n_161)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_32),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_33),
.B(n_184),
.Y(n_183)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_41),
.C(n_44),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_38),
.A2(n_44),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_38),
.Y(n_196)
);

INVx4_ASAP7_75t_SL g54 ( 
.A(n_39),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_41),
.A2(n_152),
.B1(n_153),
.B2(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_41),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_41),
.A2(n_153),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_42),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_44),
.Y(n_195)
);

INVx3_ASAP7_75t_SL g95 ( 
.A(n_45),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_50),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_52),
.C(n_55),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_105),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_49),
.B(n_185),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_54),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_95),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_53),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_54),
.B(n_120),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_54),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_55),
.Y(n_56)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

XNOR2xp5_ASAP7_75t_SL g57 ( 
.A(n_58),
.B(n_72),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_66),
.C(n_68),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_59),
.A2(n_60),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_65),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g83 ( 
.A(n_61),
.B(n_84),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_63),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_64),
.A2(n_65),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_64),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_65),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_65),
.A2(n_86),
.B1(n_117),
.B2(n_118),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_66),
.A2(n_68),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_66),
.Y(n_111)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

XOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_74),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_76),
.C(n_77),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_77),
.B2(n_78),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_76),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_76),
.A2(n_78),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_80),
.B(n_172),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_98),
.C(n_108),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_81),
.A2(n_82),
.B1(n_175),
.B2(n_176),
.Y(n_174)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_87),
.C(n_91),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_83),
.B(n_234),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_88),
.A2(n_89),
.B(n_90),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_91),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_96),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_92),
.A2(n_93),
.B1(n_96),
.B2(n_97),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g180 ( 
.A(n_94),
.B(n_181),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_98),
.B(n_108),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_104),
.C(n_106),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_99),
.B(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_102),
.C(n_103),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_100),
.B(n_212),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_101),
.B(n_185),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_101),
.B(n_105),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g212 ( 
.A1(n_102),
.A2(n_103),
.B1(n_127),
.B2(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_102),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_103),
.A2(n_127),
.B1(n_128),
.B2(n_131),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_103),
.B(n_129),
.C(n_130),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_104),
.B(n_106),
.Y(n_190)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_123),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_115),
.B(n_124),
.C(n_126),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_121),
.B2(n_122),
.Y(n_115)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_116),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_117),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_117),
.A2(n_118),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_126),
.Y(n_123)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_125),
.A2(n_207),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_128),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_130),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_156),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_137),
.B1(n_144),
.B2(n_155),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_142),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_142),
.B(n_187),
.C(n_188),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_142),
.A2(n_143),
.B1(n_187),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_145),
.B(n_146),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_152),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g326 ( 
.A(n_156),
.Y(n_326)
);

FAx1_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_158),
.CI(n_159),
.CON(n_156),
.SN(n_156)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_199),
.B(n_320),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_173),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_171),
.B(n_173),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.C(n_197),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_174),
.A2(n_197),
.B1(n_198),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_174),
.Y(n_315)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_177),
.B(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_189),
.C(n_191),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_178),
.B(n_230),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_182),
.C(n_186),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_179),
.A2(n_180),
.B1(n_215),
.B2(n_217),
.Y(n_214)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_182),
.A2(n_183),
.B1(n_186),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_184),
.Y(n_227)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_186),
.Y(n_216)
);

CKINVDCx14_ASAP7_75t_R g221 ( 
.A(n_187),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_220),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_191),
.B1(n_192),
.B2(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx24_ASAP7_75t_SL g324 ( 
.A(n_198),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_317),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_311),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_236),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_228),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_204),
.B(n_228),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_214),
.C(n_218),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_205),
.B(n_308),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g322 ( 
.A(n_205),
.Y(n_322)
);

FAx1_ASAP7_75t_SL g205 ( 
.A(n_206),
.B(n_210),
.CI(n_211),
.CON(n_205),
.SN(n_205)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_210),
.C(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.C(n_209),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_208),
.B(n_209),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_214),
.B(n_218),
.Y(n_308)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_215),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_222),
.C(n_226),
.Y(n_218)
);

FAx1_ASAP7_75t_SL g298 ( 
.A(n_219),
.B(n_222),
.CI(n_226),
.CON(n_298),
.SN(n_298)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.C(n_225),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_223),
.B(n_225),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_224),
.B(n_247),
.Y(n_246)
);

BUFx24_ASAP7_75t_SL g325 ( 
.A(n_228),
.Y(n_325)
);

FAx1_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_232),
.CI(n_233),
.CON(n_228),
.SN(n_228)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_229),
.B(n_232),
.C(n_233),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_306),
.B(n_310),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_294),
.B(n_305),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_266),
.B(n_293),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_257),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_240),
.B(n_257),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_250),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_242),
.A2(n_246),
.B1(n_248),
.B2(n_249),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_242),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.C(n_245),
.Y(n_242)
);

FAx1_ASAP7_75t_SL g258 ( 
.A(n_243),
.B(n_244),
.CI(n_245),
.CON(n_258),
.SN(n_258)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_246),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_246),
.B(n_248),
.C(n_250),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_254),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_251),
.B(n_255),
.C(n_256),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.C(n_265),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_258),
.B(n_290),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_258),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_259),
.A2(n_260),
.B1(n_265),
.B2(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_261),
.A2(n_262),
.B1(n_263),
.B2(n_264),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_262),
.Y(n_261)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_265),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_287),
.B(n_292),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_268),
.A2(n_278),
.B(n_286),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_274),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_269),
.B(n_274),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_272),
.C(n_273),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_280),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_275),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_281),
.B(n_285),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_283),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_288),
.B(n_289),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_301),
.C(n_302),
.Y(n_309)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_298),
.Y(n_328)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_307),
.B(n_309),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_316),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_313),
.B(n_316),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);


endmodule