module fake_jpeg_31001_n_35 (n_3, n_2, n_1, n_0, n_4, n_5, n_35);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_35;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g6 ( 
.A(n_4),
.Y(n_6)
);

INVx1_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx4_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NOR2xp33_ASAP7_75t_SL g13 ( 
.A(n_10),
.B(n_5),
.Y(n_13)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_11),
.B(n_0),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_14),
.B(n_17),
.Y(n_20)
);

INVx3_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_15),
.Y(n_21)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_16),
.B(n_18),
.C(n_6),
.Y(n_19)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g24 ( 
.A1(n_19),
.A2(n_16),
.B(n_14),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_21),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_23),
.B(n_25),
.C(n_18),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_14),
.C(n_20),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g25 ( 
.A1(n_19),
.A2(n_18),
.B(n_17),
.C(n_7),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_27),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_20),
.C(n_22),
.Y(n_27)
);

AOI21x1_ASAP7_75t_L g30 ( 
.A1(n_28),
.A2(n_13),
.B(n_17),
.Y(n_30)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_30),
.B(n_13),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_12),
.B2(n_15),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_29),
.A2(n_30),
.B(n_15),
.Y(n_32)
);

NOR2xp67_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_8),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_8),
.Y(n_35)
);


endmodule