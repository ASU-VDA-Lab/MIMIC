module real_jpeg_6441_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_1),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_1),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_1),
.Y(n_270)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_2),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_291),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_2),
.B(n_308),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_2),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_2),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_2),
.B(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_SL g27 ( 
.A(n_3),
.B(n_28),
.Y(n_27)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_3),
.B(n_48),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_3),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g139 ( 
.A(n_3),
.B(n_140),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_3),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_3),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_3),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_4),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_4),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_4),
.B(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_4),
.B(n_52),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_4),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_4),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_5),
.B(n_100),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_5),
.A2(n_30),
.B(n_283),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_5),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_5),
.B(n_354),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_5),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_5),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_5),
.B(n_431),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_5),
.B(n_414),
.Y(n_441)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_7),
.B(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_7),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_7),
.B(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_7),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g241 ( 
.A(n_7),
.B(n_242),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_7),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_7),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_7),
.B(n_351),
.Y(n_350)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_8),
.Y(n_153)
);

INVx8_ASAP7_75t_L g239 ( 
.A(n_8),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g351 ( 
.A(n_8),
.Y(n_351)
);

BUFx5_ASAP7_75t_L g414 ( 
.A(n_8),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_9),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_9),
.B(n_313),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_9),
.B(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_9),
.B(n_405),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_9),
.B(n_424),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_9),
.B(n_403),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_9),
.B(n_438),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_10),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g345 ( 
.A(n_10),
.Y(n_345)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_12),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_12),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_12),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_12),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_12),
.B(n_304),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_12),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_12),
.B(n_417),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_12),
.B(n_455),
.Y(n_454)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_13),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_13),
.Y(n_122)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_13),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_13),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_14),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_14),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_14),
.Y(n_403)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_14),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_15),
.B(n_22),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_15),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_15),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_15),
.B(n_122),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_15),
.B(n_124),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_15),
.B(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_111),
.B(n_127),
.C(n_499),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_39),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_19),
.B(n_103),
.CI(n_104),
.CON(n_102),
.SN(n_102)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_27),
.C(n_32),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_20),
.A2(n_21),
.B1(n_32),
.B2(n_79),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_20),
.A2(n_21),
.B1(n_107),
.B2(n_109),
.Y(n_106)
);

NOR3xp33_ASAP7_75t_L g499 ( 
.A(n_20),
.B(n_47),
.C(n_107),
.Y(n_499)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_21),
.B(n_185),
.C(n_186),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_21),
.B(n_231),
.Y(n_230)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_25),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_25),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_25),
.Y(n_265)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_26),
.Y(n_357)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_27),
.A2(n_89),
.B1(n_90),
.B2(n_91),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_27),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_27),
.A2(n_91),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_27),
.B(n_139),
.C(n_143),
.Y(n_168)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_31),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_32),
.A2(n_44),
.B1(n_79),
.B2(n_80),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_32),
.B(n_234),
.C(n_240),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_32),
.A2(n_79),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_34),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g405 ( 
.A(n_37),
.Y(n_405)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_38),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g275 ( 
.A(n_38),
.Y(n_275)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_38),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_40),
.B(n_102),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_86),
.C(n_87),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_41),
.B(n_497),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_64),
.C(n_76),
.Y(n_41)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_42),
.B(n_171),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_54),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_60),
.C(n_62),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_50),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_79),
.C(n_85),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_44),
.A2(n_80),
.B1(n_166),
.B2(n_167),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_44),
.A2(n_80),
.B1(n_261),
.B2(n_262),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx11_ASAP7_75t_L g133 ( 
.A(n_46),
.Y(n_133)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_46),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_46),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_47),
.A2(n_105),
.B1(n_106),
.B2(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_47),
.A2(n_50),
.B1(n_51),
.B2(n_110),
.Y(n_167)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_50),
.A2(n_51),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_50),
.B(n_121),
.C(n_128),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_50),
.A2(n_51),
.B1(n_307),
.B2(n_369),
.Y(n_368)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_51),
.B(n_303),
.C(n_307),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_60),
.B1(n_62),
.B2(n_63),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_55),
.Y(n_62)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_59),
.Y(n_246)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_59),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_64),
.B(n_76),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_69),
.C(n_74),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_65),
.A2(n_69),
.B1(n_70),
.B2(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_65),
.Y(n_147)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_69),
.A2(n_70),
.B1(n_217),
.B2(n_218),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_70),
.B(n_152),
.C(n_196),
.Y(n_195)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_73),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_81),
.B2(n_85),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_80),
.B(n_261),
.C(n_266),
.Y(n_260)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_81),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_81),
.B(n_128),
.C(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_81),
.A2(n_85),
.B1(n_130),
.B2(n_183),
.Y(n_182)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_86),
.B(n_87),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_87)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_96),
.C(n_101),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx4_ASAP7_75t_L g187 ( 
.A(n_99),
.Y(n_187)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx24_ASAP7_75t_SL g502 ( 
.A(n_102),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_107),
.Y(n_109)
);

MAJx2_ASAP7_75t_L g194 ( 
.A(n_107),
.B(n_195),
.C(n_199),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_107),
.A2(n_109),
.B1(n_160),
.B2(n_206),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_107),
.A2(n_109),
.B1(n_199),
.B2(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_150),
.C(n_160),
.Y(n_149)
);

AO21x1_ASAP7_75t_SL g111 ( 
.A1(n_112),
.A2(n_494),
.B(n_498),
.Y(n_111)
);

OAI21xp33_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_251),
.B(n_491),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_208),
.Y(n_113)
);

AOI21xp33_ASAP7_75t_SL g491 ( 
.A1(n_114),
.A2(n_492),
.B(n_493),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_115),
.B(n_172),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_115),
.B(n_172),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_163),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_116),
.B(n_164),
.C(n_170),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_145),
.C(n_148),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_117),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_129),
.C(n_134),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_118),
.B(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_123),
.B1(n_127),
.B2(n_128),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_121),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_123),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g180 ( 
.A1(n_123),
.A2(n_128),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g348 ( 
.A(n_123),
.B(n_235),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_123),
.A2(n_128),
.B1(n_234),
.B2(n_235),
.Y(n_459)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_126),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_134),
.Y(n_213)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_130),
.Y(n_183)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_132),
.Y(n_242)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_133),
.Y(n_376)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_139),
.B1(n_143),
.B2(n_144),
.Y(n_136)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_137),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g144 ( 
.A(n_139),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_139),
.B(n_222),
.Y(n_259)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_144),
.B(n_221),
.C(n_226),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_145),
.A2(n_148),
.B1(n_149),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_145),
.Y(n_175)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_150),
.A2(n_151),
.B1(n_205),
.B2(n_207),
.Y(n_204)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_152),
.A2(n_158),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_152),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_152),
.A2(n_190),
.B1(n_196),
.B2(n_219),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_152),
.A2(n_190),
.B1(n_416),
.B2(n_418),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_152),
.B(n_418),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_154),
.A2(n_189),
.B1(n_192),
.B2(n_193),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_154),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_154),
.B(n_273),
.C(n_276),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_154),
.A2(n_192),
.B1(n_273),
.B2(n_340),
.Y(n_339)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_156),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_170),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_169),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_176),
.C(n_178),
.Y(n_172)
);

FAx1_ASAP7_75t_SL g250 ( 
.A(n_173),
.B(n_176),
.CI(n_178),
.CON(n_250),
.SN(n_250)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_194),
.C(n_204),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_211),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_184),
.C(n_188),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_180),
.B(n_184),
.Y(n_324)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_186),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_188),
.B(n_324),
.Y(n_323)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_189),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_194),
.B(n_204),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_195),
.B(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_196),
.B(n_311),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_196),
.A2(n_219),
.B1(n_311),
.B2(n_312),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g410 ( 
.A(n_197),
.Y(n_410)
);

INVx8_ASAP7_75t_L g432 ( 
.A(n_197),
.Y(n_432)
);

BUFx8_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_198),
.Y(n_440)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_199),
.Y(n_249)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx8_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g308 ( 
.A(n_203),
.Y(n_308)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_205),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_250),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_209),
.B(n_250),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_212),
.C(n_214),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_210),
.B(n_212),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_214),
.B(n_331),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_232),
.C(n_247),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_215),
.B(n_326),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_220),
.C(n_230),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_216),
.Y(n_296)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_220),
.B(n_230),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_226),
.B(n_259),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_232),
.B(n_247),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_241),
.C(n_243),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_293),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_234),
.A2(n_235),
.B1(n_240),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_235),
.Y(n_234)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_239),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_240),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_241),
.Y(n_294)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx6_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx24_ASAP7_75t_SL g501 ( 
.A(n_250),
.Y(n_501)
);

AOI221xp5_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_389),
.B1(n_484),
.B2(n_489),
.C(n_490),
.Y(n_251)
);

NOR3xp33_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_328),
.C(n_332),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_253),
.A2(n_485),
.B(n_488),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_321),
.Y(n_253)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_254),
.B(n_321),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_295),
.C(n_298),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_255),
.B(n_295),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_256),
.B(n_280),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_256),
.B(n_281),
.C(n_292),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_271),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_258),
.B(n_272),
.Y(n_359)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_260),
.B(n_359),
.Y(n_358)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx5_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_266),
.B(n_301),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

INVx5_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

BUFx5_ASAP7_75t_L g417 ( 
.A(n_270),
.Y(n_417)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_273),
.Y(n_340)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_276),
.B(n_339),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_292),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_287),
.C(n_290),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_320),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_282),
.A2(n_283),
.B(n_342),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

INVx4_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_287),
.B(n_290),
.Y(n_320)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_289),
.B(n_343),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_298),
.B(n_361),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_315),
.C(n_319),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_299),
.B(n_336),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.C(n_309),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_300),
.B(n_385),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_302),
.A2(n_309),
.B1(n_310),
.B2(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_302),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g367 ( 
.A(n_303),
.B(n_368),
.Y(n_367)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx4_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_307),
.Y(n_369)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx6_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_315),
.B(n_319),
.Y(n_336)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_327),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_325),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_325),
.C(n_327),
.Y(n_329)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_328),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_329),
.B(n_330),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_329),
.B(n_330),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_333),
.B(n_362),
.Y(n_332)
);

AOI21xp5_ASAP7_75t_L g485 ( 
.A1(n_333),
.A2(n_486),
.B(n_487),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_360),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g487 ( 
.A(n_334),
.B(n_360),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.C(n_358),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_388),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_337),
.B(n_358),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_341),
.C(n_346),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_338),
.B(n_341),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_346),
.B(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.C(n_352),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_347),
.A2(n_348),
.B1(n_472),
.B2(n_473),
.Y(n_471)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_349),
.A2(n_350),
.B1(n_352),
.B2(n_353),
.Y(n_472)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_387),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_363),
.B(n_387),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.C(n_384),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_364),
.B(n_482),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_366),
.B(n_384),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.C(n_382),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_367),
.B(n_475),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_370),
.A2(n_382),
.B1(n_383),
.B2(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_370),
.Y(n_476)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_374),
.C(n_377),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g464 ( 
.A1(n_371),
.A2(n_372),
.B1(n_377),
.B2(n_378),
.Y(n_464)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g463 ( 
.A(n_374),
.B(n_464),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_L g374 ( 
.A(n_375),
.B(n_376),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_375),
.B(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx4_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_SL g389 ( 
.A1(n_390),
.A2(n_479),
.B(n_483),
.Y(n_389)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_466),
.B(n_478),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_392),
.A2(n_450),
.B(n_465),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_393),
.A2(n_426),
.B(n_449),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_419),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_394),
.B(n_419),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_406),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_395),
.B(n_407),
.C(n_415),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_401),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_396),
.B(n_402),
.C(n_404),
.Y(n_462)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_404),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_415),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_411),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_408),
.B(n_411),
.Y(n_420)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_413),
.Y(n_411)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_416),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_421),
.C(n_422),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_420),
.B(n_446),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g446 ( 
.A1(n_421),
.A2(n_422),
.B1(n_423),
.B2(n_447),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_421),
.Y(n_447)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_427),
.A2(n_443),
.B(n_448),
.Y(n_426)
);

AOI21xp5_ASAP7_75t_L g427 ( 
.A1(n_428),
.A2(n_436),
.B(n_442),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_429),
.B(n_435),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_435),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_433),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g444 ( 
.A(n_430),
.B(n_433),
.Y(n_444)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_441),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_439),
.Y(n_438)
);

INVx3_ASAP7_75t_L g439 ( 
.A(n_440),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_445),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_445),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_452),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_451),
.B(n_452),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_461),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g468 ( 
.A1(n_453),
.A2(n_469),
.B1(n_470),
.B2(n_471),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_453),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_462),
.C(n_463),
.Y(n_477)
);

FAx1_ASAP7_75t_SL g453 ( 
.A(n_454),
.B(n_459),
.CI(n_460),
.CON(n_453),
.SN(n_453)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_462),
.B(n_463),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_467),
.B(n_477),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_477),
.Y(n_478)
);

XOR2xp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_474),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_469),
.B(n_471),
.C(n_474),
.Y(n_480)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_472),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_481),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_480),
.B(n_481),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_495),
.B(n_496),
.Y(n_498)
);


endmodule