module fake_jpeg_25951_n_59 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

INVx3_ASAP7_75t_L g22 ( 
.A(n_19),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_9),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx5_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_22),
.Y(n_28)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_0),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_29),
.B(n_30),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_1),
.Y(n_31)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_31),
.A2(n_32),
.B(n_3),
.Y(n_41)
);

NAND2x1_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_1),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_26),
.B(n_2),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_22),
.B1(n_26),
.B2(n_31),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_20),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_36),
.B(n_38),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_34),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_41),
.A2(n_42),
.B(n_43),
.Y(n_47)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_15),
.B(n_5),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_SL g43 ( 
.A1(n_32),
.A2(n_24),
.B(n_25),
.C(n_4),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_8),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_44),
.B(n_47),
.C(n_48),
.Y(n_52)
);

OAI221xp5_ASAP7_75t_L g45 ( 
.A1(n_40),
.A2(n_4),
.B1(n_21),
.B2(n_11),
.C(n_12),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_46),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_13),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g51 ( 
.A(n_37),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_52),
.A2(n_49),
.B1(n_51),
.B2(n_50),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_49),
.B(n_16),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_14),
.B(n_17),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_55),
.Y(n_59)
);


endmodule