module fake_jpeg_21821_n_256 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_256);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_256;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx6_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_9),
.B(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_38),
.B(n_39),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_43),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_18),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_47),
.Y(n_54)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_26),
.B(n_0),
.Y(n_44)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_44),
.A2(n_36),
.B(n_27),
.Y(n_78)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_26),
.Y(n_46)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_46),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_29),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_46),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_60),
.Y(n_83)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_31),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_52),
.B(n_47),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_35),
.B1(n_33),
.B2(n_21),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_68),
.B1(n_73),
.B2(n_20),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_37),
.A2(n_19),
.B1(n_25),
.B2(n_36),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_55),
.A2(n_62),
.B(n_20),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_18),
.C(n_31),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_65),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_35),
.B1(n_33),
.B2(n_30),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_45),
.A2(n_19),
.B1(n_25),
.B2(n_33),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_69),
.A2(n_22),
.B1(n_27),
.B2(n_35),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_45),
.A2(n_19),
.B1(n_25),
.B2(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_75),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_39),
.B(n_23),
.Y(n_77)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_21),
.Y(n_108)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

CKINVDCx9p33_ASAP7_75t_R g80 ( 
.A(n_46),
.Y(n_80)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_62),
.A2(n_42),
.B1(n_40),
.B2(n_28),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_84),
.A2(n_104),
.B1(n_80),
.B2(n_72),
.Y(n_132)
);

AO22x1_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_44),
.B1(n_34),
.B2(n_42),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_85),
.A2(n_110),
.B1(n_24),
.B2(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_54),
.B(n_44),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_86),
.B(n_98),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_106),
.B1(n_24),
.B2(n_30),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_49),
.A2(n_36),
.B1(n_20),
.B2(n_22),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_29),
.Y(n_127)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_107),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_51),
.B(n_34),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_100),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_61),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_102),
.B(n_30),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_57),
.A2(n_28),
.B1(n_22),
.B2(n_27),
.Y(n_104)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_70),
.Y(n_107)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_108),
.A2(n_56),
.B(n_24),
.C(n_32),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_73),
.A2(n_47),
.B1(n_39),
.B2(n_21),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_52),
.B(n_23),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_111),
.B(n_58),
.Y(n_123)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_112),
.B(n_113),
.Y(n_143)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_83),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_98),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_114),
.B(n_118),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_116),
.B(n_121),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_117),
.A2(n_137),
.B1(n_91),
.B2(n_4),
.Y(n_166)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_119),
.A2(n_127),
.B1(n_131),
.B2(n_132),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_3),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_32),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_96),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_126),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g162 ( 
.A(n_123),
.B(n_125),
.Y(n_162)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_111),
.Y(n_126)
);

NAND3xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_75),
.C(n_16),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_130),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_87),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_85),
.A2(n_59),
.B1(n_72),
.B2(n_75),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_108),
.B(n_71),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_89),
.B(n_66),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_95),
.B(n_50),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_88),
.B(n_50),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_99),
.B(n_15),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_138),
.B(n_15),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_88),
.B(n_76),
.Y(n_139)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_139),
.Y(n_150)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_84),
.Y(n_140)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_140),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_119),
.A2(n_85),
.B1(n_101),
.B2(n_82),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_142),
.A2(n_149),
.B1(n_154),
.B2(n_156),
.Y(n_168)
);

OR2x4_ASAP7_75t_L g145 ( 
.A(n_133),
.B(n_97),
.Y(n_145)
);

A2O1A1Ixp33_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_165),
.B(n_5),
.C(n_7),
.Y(n_181)
);

AO22x2_ASAP7_75t_L g146 ( 
.A1(n_134),
.A2(n_82),
.B1(n_101),
.B2(n_81),
.Y(n_146)
);

AO22x1_ASAP7_75t_SL g173 ( 
.A1(n_146),
.A2(n_127),
.B1(n_136),
.B2(n_129),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_135),
.A2(n_97),
.B1(n_94),
.B2(n_105),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_147),
.A2(n_151),
.B1(n_166),
.B2(n_112),
.Y(n_177)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_155),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_140),
.A2(n_94),
.B1(n_105),
.B2(n_81),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_125),
.A2(n_109),
.B1(n_100),
.B2(n_103),
.Y(n_151)
);

AND2x6_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_3),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g174 ( 
.A1(n_153),
.A2(n_160),
.B(n_167),
.C(n_129),
.D(n_121),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_109),
.B1(n_103),
.B2(n_92),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_132),
.A2(n_92),
.B1(n_87),
.B2(n_107),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_123),
.A2(n_91),
.B(n_4),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_8),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_115),
.A2(n_3),
.B(n_5),
.Y(n_167)
);

NAND3xp33_ASAP7_75t_L g169 ( 
.A(n_145),
.B(n_126),
.C(n_115),
.Y(n_169)
);

OAI322xp33_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_165),
.A3(n_144),
.B1(n_146),
.B2(n_167),
.C1(n_160),
.C2(n_155),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g170 ( 
.A1(n_159),
.A2(n_120),
.B(n_118),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_146),
.B(n_152),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_139),
.Y(n_171)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_171),
.Y(n_190)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_172),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g201 ( 
.A1(n_173),
.A2(n_177),
.B1(n_185),
.B2(n_153),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_174),
.B(n_181),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_158),
.B(n_127),
.Y(n_176)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_176),
.Y(n_194)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_178),
.B(n_183),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_156),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g202 ( 
.A(n_179),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_142),
.A2(n_113),
.B1(n_124),
.B2(n_116),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_180),
.A2(n_186),
.B1(n_141),
.B2(n_154),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_149),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_146),
.B(n_8),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_184),
.B(n_11),
.Y(n_200)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_159),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_150),
.B(n_162),
.Y(n_187)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_187),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_150),
.B(n_11),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_189),
.B(n_181),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_173),
.B(n_183),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_171),
.B(n_141),
.C(n_152),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_193),
.B(n_198),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_196),
.B(n_200),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_176),
.B(n_147),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_187),
.B(n_163),
.Y(n_199)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_199),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_204),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_175),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_196),
.A2(n_168),
.B1(n_179),
.B2(n_173),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_218),
.B1(n_190),
.B2(n_188),
.Y(n_230)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_213),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_184),
.B(n_200),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_191),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_192),
.Y(n_217)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_217),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_193),
.A2(n_203),
.B1(n_195),
.B2(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_199),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_219),
.A2(n_220),
.B1(n_205),
.B2(n_203),
.Y(n_221)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_221),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_177),
.B1(n_170),
.B2(n_205),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_224),
.A2(n_230),
.B1(n_217),
.B2(n_186),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_210),
.B(n_198),
.C(n_194),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_226),
.B(n_227),
.C(n_228),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_210),
.B(n_218),
.C(n_194),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_190),
.C(n_195),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_229),
.A2(n_216),
.B1(n_211),
.B2(n_213),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_231),
.B(n_148),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_232),
.B(n_236),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_226),
.B(n_216),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_239),
.Y(n_242)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_161),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_235),
.A2(n_225),
.B1(n_229),
.B2(n_223),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_230),
.B(n_178),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_231),
.B(n_197),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_240),
.B(n_244),
.Y(n_247)
);

AOI322xp5_ASAP7_75t_L g241 ( 
.A1(n_237),
.A2(n_222),
.A3(n_233),
.B1(n_227),
.B2(n_232),
.C1(n_235),
.C2(n_228),
.Y(n_241)
);

AOI21xp33_ASAP7_75t_L g246 ( 
.A1(n_241),
.A2(n_238),
.B(n_12),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_237),
.A2(n_174),
.B(n_206),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_245),
.A2(n_11),
.B(n_14),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_246),
.B(n_248),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_238),
.C(n_13),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_249),
.B(n_244),
.Y(n_250)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_250),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_247),
.A2(n_243),
.B1(n_240),
.B2(n_14),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_251),
.B(n_14),
.C(n_252),
.Y(n_253)
);

BUFx24_ASAP7_75t_SL g255 ( 
.A(n_253),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_254),
.Y(n_256)
);


endmodule