module real_aes_5367_n_422 (n_76, n_113, n_187, n_90, n_257, n_390, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_386, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_421, n_329, n_132, n_1424, n_131, n_144, n_169, n_242, n_376, n_308, n_172, n_341, n_232, n_6, n_401, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_1425, n_379, n_374, n_26, n_235, n_399, n_378, n_245, n_161, n_189, n_271, n_2, n_145, n_415, n_227, n_92, n_330, n_388, n_395, n_332, n_292, n_400, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_408, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_384, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_409, n_298, n_49, n_43, n_297, n_383, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_381, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_398, n_89, n_277, n_331, n_93, n_182, n_363, n_417, n_323, n_199, n_350, n_142, n_223, n_67, n_405, n_368, n_250, n_85, n_406, n_45, n_5, n_244, n_118, n_139, n_402, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_416, n_410, n_120, n_261, n_238, n_391, n_360, n_58, n_165, n_361, n_246, n_176, n_412, n_163, n_29, n_52, n_1427, n_251, n_220, n_387, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_392, n_150, n_147, n_288, n_404, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_413, n_306, n_158, n_4, n_366, n_346, n_193, n_397, n_293, n_162, n_358, n_385, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_377, n_273, n_114, n_276, n_295, n_382, n_265, n_354, n_154, n_127, n_326, n_24, n_407, n_217, n_419, n_55, n_62, n_411, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_389, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_420, n_1426, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_418, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_1428, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_414, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_380, n_394, n_168, n_175, n_241, n_105, n_84, n_294, n_393, n_258, n_206, n_307, n_396, n_342, n_348, n_14, n_403, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_422);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_390;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_386;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_421;
input n_329;
input n_132;
input n_1424;
input n_131;
input n_144;
input n_169;
input n_242;
input n_376;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_401;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_1425;
input n_379;
input n_374;
input n_26;
input n_235;
input n_399;
input n_378;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_415;
input n_227;
input n_92;
input n_330;
input n_388;
input n_395;
input n_332;
input n_292;
input n_400;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_408;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_384;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_409;
input n_298;
input n_49;
input n_43;
input n_297;
input n_383;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_381;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_398;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_417;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_405;
input n_368;
input n_250;
input n_85;
input n_406;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_402;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_416;
input n_410;
input n_120;
input n_261;
input n_238;
input n_391;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_412;
input n_163;
input n_29;
input n_52;
input n_1427;
input n_251;
input n_220;
input n_387;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_392;
input n_150;
input n_147;
input n_288;
input n_404;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_413;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_397;
input n_293;
input n_162;
input n_358;
input n_385;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_377;
input n_273;
input n_114;
input n_276;
input n_295;
input n_382;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_407;
input n_217;
input n_419;
input n_55;
input n_62;
input n_411;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_389;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_420;
input n_1426;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_418;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_1428;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_414;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_380;
input n_394;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_393;
input n_258;
input n_206;
input n_307;
input n_396;
input n_342;
input n_348;
input n_14;
input n_403;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_422;
wire n_476;
wire n_887;
wire n_599;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_919;
wire n_1217;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_786;
wire n_512;
wire n_795;
wire n_1379;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_755;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1317;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_898;
wire n_562;
wire n_1022;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1209;
wire n_498;
wire n_765;
wire n_1397;
wire n_648;
wire n_939;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_591;
wire n_1366;
wire n_678;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_1368;
wire n_994;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_617;
wire n_602;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_895;
wire n_799;
wire n_490;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_1026;
wire n_492;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_526;
wire n_1194;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_721;
wire n_1133;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_943;
wire n_977;
wire n_905;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_816;
wire n_625;
wire n_953;
wire n_1373;
wire n_716;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_1207;
wire n_664;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_561;
wire n_437;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1060;
wire n_1154;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_563;
wire n_891;
wire n_568;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_1083;
wire n_727;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_1139;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1127;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1051;
wire n_1355;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1164;
wire n_433;
wire n_627;
wire n_771;
wire n_1378;
wire n_524;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1156;
wire n_988;
wire n_1396;
wire n_921;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1318;
wire n_1290;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_425;
wire n_879;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_542;
wire n_1256;
wire n_1077;
wire n_1111;
wire n_1249;
wire n_1416;
wire n_1239;
wire n_969;
wire n_1009;
wire n_1202;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_1183;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1345;
wire n_587;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_729;
wire n_1280;
wire n_1352;
wire n_1323;
wire n_1369;
wire n_703;
wire n_1097;
wire n_601;
wire n_463;
wire n_1236;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_0), .A2(n_373), .B1(n_590), .B2(n_951), .Y(n_1016) );
INVx1_ASAP7_75t_L g749 ( .A(n_1), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_2), .A2(n_349), .B1(n_558), .B2(n_559), .Y(n_1078) );
AOI22xp5_ASAP7_75t_L g762 ( .A1(n_3), .A2(n_314), .B1(n_618), .B2(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g1055 ( .A(n_4), .Y(n_1055) );
INVx1_ASAP7_75t_L g654 ( .A(n_5), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g1061 ( .A1(n_6), .A2(n_332), .B1(n_552), .B2(n_714), .Y(n_1061) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_7), .A2(n_353), .B1(n_505), .B2(n_538), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_8), .A2(n_260), .B1(n_687), .B2(n_718), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1412 ( .A1(n_9), .A2(n_193), .B1(n_526), .B2(n_714), .Y(n_1412) );
AOI22xp33_ASAP7_75t_SL g943 ( .A1(n_10), .A2(n_339), .B1(n_527), .B2(n_532), .Y(n_943) );
INVx1_ASAP7_75t_SL g1242 ( .A(n_11), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_12), .A2(n_164), .B1(n_491), .B2(n_634), .Y(n_665) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_13), .A2(n_242), .B1(n_618), .B2(n_619), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g648 ( .A1(n_14), .A2(n_327), .B1(n_649), .B2(n_650), .C(n_653), .Y(n_648) );
INVx1_ASAP7_75t_L g789 ( .A(n_15), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g1093 ( .A1(n_16), .A2(n_83), .B1(n_522), .B2(n_887), .Y(n_1093) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_17), .A2(n_269), .B1(n_600), .B2(n_601), .Y(n_599) );
INVx1_ASAP7_75t_L g752 ( .A(n_18), .Y(n_752) );
AOI22xp33_ASAP7_75t_L g929 ( .A1(n_19), .A2(n_345), .B1(n_522), .B2(n_772), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_20), .A2(n_22), .B1(n_772), .B2(n_774), .Y(n_868) );
AOI22xp5_ASAP7_75t_L g713 ( .A1(n_21), .A2(n_80), .B1(n_552), .B2(n_714), .Y(n_713) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_23), .B(n_438), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g877 ( .A1(n_24), .A2(n_813), .B(n_878), .Y(n_877) );
CKINVDCx20_ASAP7_75t_R g1152 ( .A(n_25), .Y(n_1152) );
AOI222xp33_ASAP7_75t_L g1368 ( .A1(n_25), .A2(n_1369), .B1(n_1375), .B2(n_1396), .C1(n_1399), .C2(n_1414), .Y(n_1368) );
INVx1_ASAP7_75t_L g746 ( .A(n_26), .Y(n_746) );
AOI221x1_ASAP7_75t_L g938 ( .A1(n_27), .A2(n_101), .B1(n_727), .B2(n_939), .C(n_940), .Y(n_938) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_28), .A2(n_402), .B1(n_555), .B2(n_556), .Y(n_716) );
AOI22xp33_ASAP7_75t_L g775 ( .A1(n_29), .A2(n_256), .B1(n_521), .B2(n_776), .Y(n_775) );
BUFx6f_ASAP7_75t_L g438 ( .A(n_30), .Y(n_438) );
AOI22xp33_ASAP7_75t_L g1110 ( .A1(n_31), .A2(n_39), .B1(n_621), .B2(n_774), .Y(n_1110) );
INVx1_ASAP7_75t_L g733 ( .A(n_32), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g1182 ( .A1(n_32), .A2(n_109), .B1(n_1140), .B2(n_1159), .Y(n_1182) );
AOI22xp5_ASAP7_75t_L g849 ( .A1(n_33), .A2(n_249), .B1(n_561), .B2(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g578 ( .A(n_34), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g551 ( .A1(n_35), .A2(n_317), .B1(n_552), .B2(n_553), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g1380 ( .A1(n_36), .A2(n_56), .B1(n_986), .B2(n_1087), .Y(n_1380) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_37), .A2(n_97), .B1(n_504), .B2(n_512), .Y(n_503) );
INVx1_ASAP7_75t_L g583 ( .A(n_38), .Y(n_583) );
AOI21xp33_ASAP7_75t_L g635 ( .A1(n_40), .A2(n_597), .B(n_636), .Y(n_635) );
AOI22xp33_ASAP7_75t_L g1075 ( .A1(n_41), .A2(n_233), .B1(n_470), .B2(n_663), .Y(n_1075) );
INVx1_ASAP7_75t_L g1021 ( .A(n_42), .Y(n_1021) );
AOI22xp33_ASAP7_75t_L g1046 ( .A1(n_43), .A2(n_142), .B1(n_570), .B2(n_663), .Y(n_1046) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_44), .A2(n_283), .B1(n_496), .B2(n_876), .Y(n_875) );
AOI22xp33_ASAP7_75t_SL g811 ( .A1(n_45), .A2(n_343), .B1(n_573), .B2(n_812), .Y(n_811) );
INVx1_ASAP7_75t_L g1054 ( .A(n_46), .Y(n_1054) );
CKINVDCx16_ASAP7_75t_R g701 ( .A(n_47), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g679 ( .A1(n_48), .A2(n_212), .B1(n_626), .B2(n_680), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g1244 ( .A1(n_49), .A2(n_277), .B1(n_1124), .B2(n_1179), .Y(n_1244) );
NAND2xp5_ASAP7_75t_L g1103 ( .A(n_50), .B(n_732), .Y(n_1103) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_51), .A2(n_354), .B1(n_505), .B2(n_870), .Y(n_885) );
INVx1_ASAP7_75t_L g786 ( .A(n_52), .Y(n_786) );
AOI22xp5_ASAP7_75t_L g620 ( .A1(n_53), .A2(n_65), .B1(n_621), .B2(n_623), .Y(n_620) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_54), .A2(n_261), .B1(n_556), .B2(n_618), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_55), .A2(n_346), .B1(n_500), .B2(n_992), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_57), .A2(n_157), .B1(n_609), .B2(n_610), .Y(n_1012) );
AOI22xp33_ASAP7_75t_L g822 ( .A1(n_58), .A2(n_390), .B1(n_512), .B2(n_823), .Y(n_822) );
INVx1_ASAP7_75t_L g1149 ( .A(n_59), .Y(n_1149) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_60), .A2(n_281), .B1(n_505), .B2(n_870), .Y(n_869) );
AOI22xp5_ASAP7_75t_L g1029 ( .A1(n_61), .A2(n_263), .B1(n_623), .B2(n_772), .Y(n_1029) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_62), .A2(n_413), .B1(n_634), .B2(n_693), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_63), .A2(n_421), .B1(n_485), .B2(n_491), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_64), .A2(n_405), .B1(n_588), .B2(n_754), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g999 ( .A1(n_66), .A2(n_125), .B1(n_555), .B2(n_556), .Y(n_999) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_67), .B(n_594), .Y(n_730) );
AOI21xp33_ASAP7_75t_L g814 ( .A1(n_68), .A2(n_815), .B(n_817), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g1385 ( .A1(n_69), .A2(n_163), .B1(n_846), .B2(n_1386), .Y(n_1385) );
AOI22xp5_ASAP7_75t_L g889 ( .A1(n_70), .A2(n_417), .B1(n_625), .B2(n_626), .Y(n_889) );
OA22x2_ASAP7_75t_L g443 ( .A1(n_71), .A2(n_186), .B1(n_438), .B2(n_442), .Y(n_443) );
INVx1_ASAP7_75t_L g483 ( .A(n_71), .Y(n_483) );
AOI22xp33_ASAP7_75t_L g1033 ( .A1(n_72), .A2(n_216), .B1(n_632), .B2(n_748), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1014 ( .A1(n_73), .A2(n_367), .B1(n_601), .B2(n_607), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g631 ( .A1(n_74), .A2(n_128), .B1(n_496), .B2(n_632), .Y(n_631) );
CKINVDCx5p33_ASAP7_75t_R g949 ( .A(n_75), .Y(n_949) );
NAND2xp33_ASAP7_75t_L g690 ( .A(n_76), .B(n_691), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g1088 ( .A1(n_77), .A2(n_175), .B1(n_630), .B2(n_1089), .Y(n_1088) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_78), .A2(n_411), .B1(n_606), .B2(n_618), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_79), .A2(n_252), .B1(n_505), .B2(n_538), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_81), .A2(n_359), .B1(n_505), .B2(n_513), .Y(n_924) );
INVx1_ASAP7_75t_L g441 ( .A(n_82), .Y(n_441) );
NOR2xp33_ASAP7_75t_L g477 ( .A(n_82), .B(n_205), .Y(n_477) );
OAI21xp33_ASAP7_75t_L g494 ( .A1(n_82), .A2(n_186), .B(n_468), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g928 ( .A1(n_84), .A2(n_386), .B1(n_625), .B2(n_626), .Y(n_928) );
AOI22xp5_ASAP7_75t_L g1027 ( .A1(n_85), .A2(n_293), .B1(n_513), .B2(n_522), .Y(n_1027) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_86), .A2(n_145), .B1(n_459), .B2(n_570), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g1393 ( .A1(n_87), .A2(n_290), .B1(n_1063), .B2(n_1394), .Y(n_1393) );
AOI22xp33_ASAP7_75t_L g865 ( .A1(n_88), .A2(n_300), .B1(n_625), .B2(n_626), .Y(n_865) );
AOI22xp33_ASAP7_75t_L g1094 ( .A1(n_89), .A2(n_251), .B1(n_625), .B2(n_830), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g720 ( .A1(n_90), .A2(n_206), .B1(n_649), .B2(n_721), .Y(n_720) );
AOI22xp33_ASAP7_75t_L g991 ( .A1(n_91), .A2(n_271), .B1(n_594), .B2(n_992), .Y(n_991) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_92), .A2(n_399), .B1(n_682), .B2(n_855), .Y(n_854) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_93), .A2(n_254), .B1(n_558), .B2(n_682), .Y(n_715) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_94), .A2(n_118), .B1(n_552), .B2(n_714), .Y(n_857) );
AOI21xp33_ASAP7_75t_L g896 ( .A1(n_95), .A2(n_649), .B(n_897), .Y(n_896) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_96), .B(n_313), .Y(n_1128) );
INVx1_ASAP7_75t_L g1142 ( .A(n_96), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1417 ( .A(n_96), .Y(n_1417) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_98), .A2(n_259), .B1(n_517), .B2(n_521), .Y(n_516) );
INVx1_ASAP7_75t_L g795 ( .A(n_99), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g1406 ( .A1(n_100), .A2(n_228), .B1(n_820), .B2(n_1407), .Y(n_1406) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_102), .A2(n_166), .B1(n_538), .B2(n_682), .Y(n_681) );
AOI22xp5_ASAP7_75t_L g1111 ( .A1(n_103), .A2(n_337), .B1(n_625), .B2(n_626), .Y(n_1111) );
INVx1_ASAP7_75t_L g979 ( .A(n_104), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g1032 ( .A1(n_105), .A2(n_181), .B1(n_630), .B2(n_992), .Y(n_1032) );
AOI22xp33_ASAP7_75t_SL g858 ( .A1(n_106), .A2(n_195), .B1(n_517), .B2(n_718), .Y(n_858) );
AOI22xp33_ASAP7_75t_L g995 ( .A1(n_107), .A2(n_404), .B1(n_552), .B2(n_626), .Y(n_995) );
AO22x1_ASAP7_75t_L g886 ( .A1(n_108), .A2(n_363), .B1(n_522), .B2(n_887), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_110), .A2(n_204), .B1(n_594), .B2(n_841), .Y(n_1090) );
AOI22xp33_ASAP7_75t_L g761 ( .A1(n_111), .A2(n_139), .B1(n_527), .B2(n_532), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_112), .A2(n_170), .B1(n_459), .B2(n_630), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g569 ( .A1(n_113), .A2(n_368), .B1(n_459), .B2(n_570), .Y(n_569) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_114), .A2(n_309), .B1(n_687), .B2(n_688), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_115), .A2(n_133), .B1(n_500), .B2(n_663), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_116), .A2(n_255), .B1(n_630), .B2(n_632), .Y(n_872) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_117), .B(n_816), .Y(n_914) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_119), .A2(n_162), .B1(n_540), .B2(n_621), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_120), .A2(n_344), .B1(n_517), .B2(n_1063), .Y(n_1062) );
INVx1_ASAP7_75t_L g1023 ( .A(n_121), .Y(n_1023) );
AOI22xp33_ASAP7_75t_SL g856 ( .A1(n_122), .A2(n_129), .B1(n_555), .B2(n_556), .Y(n_856) );
AOI22xp5_ASAP7_75t_L g1410 ( .A1(n_123), .A2(n_160), .B1(n_783), .B2(n_1411), .Y(n_1410) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_124), .A2(n_231), .B1(n_555), .B2(n_556), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g1030 ( .A1(n_126), .A2(n_148), .B1(n_559), .B2(n_870), .Y(n_1030) );
INVx1_ASAP7_75t_L g1127 ( .A(n_127), .Y(n_1127) );
INVx1_ASAP7_75t_SL g1143 ( .A(n_127), .Y(n_1143) );
AND2x4_ASAP7_75t_L g1146 ( .A(n_127), .B(n_1126), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_130), .A2(n_401), .B1(n_559), .B2(n_658), .Y(n_657) );
NAND2xp5_ASAP7_75t_SL g899 ( .A(n_131), .B(n_816), .Y(n_899) );
AOI21xp5_ASAP7_75t_L g839 ( .A1(n_132), .A2(n_840), .B(n_843), .Y(n_839) );
AOI22xp33_ASAP7_75t_SL g998 ( .A1(n_134), .A2(n_138), .B1(n_558), .B2(n_682), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_135), .A2(n_229), .B1(n_536), .B2(n_540), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_136), .B(n_593), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1409 ( .A1(n_137), .A2(n_322), .B1(n_1389), .B2(n_1390), .Y(n_1409) );
AO22x2_ASAP7_75t_L g778 ( .A1(n_140), .A2(n_173), .B1(n_680), .B2(n_779), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g915 ( .A1(n_141), .A2(n_916), .B(n_918), .Y(n_915) );
CKINVDCx16_ASAP7_75t_R g1173 ( .A(n_143), .Y(n_1173) );
XOR2x2_ASAP7_75t_L g767 ( .A(n_144), .B(n_768), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1203 ( .A1(n_144), .A2(n_169), .B1(n_1167), .B2(n_1204), .Y(n_1203) );
AOI33xp33_ASAP7_75t_R g1097 ( .A1(n_146), .A2(n_289), .A3(n_435), .B1(n_493), .B2(n_1098), .B3(n_1428), .Y(n_1097) );
AOI22xp33_ASAP7_75t_SL g1376 ( .A1(n_147), .A2(n_1377), .B1(n_1378), .B2(n_1395), .Y(n_1376) );
INVx1_ASAP7_75t_L g1395 ( .A(n_147), .Y(n_1395) );
INVx1_ASAP7_75t_L g862 ( .A(n_149), .Y(n_862) );
INVx1_ASAP7_75t_L g1144 ( .A(n_150), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_151), .A2(n_375), .B1(n_601), .B2(n_604), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_152), .A2(n_307), .B1(n_603), .B2(n_604), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1392 ( .A1(n_153), .A2(n_304), .B1(n_552), .B2(n_553), .Y(n_1392) );
AO22x1_ASAP7_75t_L g659 ( .A1(n_154), .A2(n_366), .B1(n_517), .B2(n_555), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_155), .A2(n_192), .B1(n_526), .B2(n_530), .Y(n_525) );
AOI22xp33_ASAP7_75t_L g808 ( .A1(n_156), .A2(n_276), .B1(n_809), .B2(n_810), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g549 ( .A1(n_158), .A2(n_258), .B1(n_517), .B2(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g1072 ( .A1(n_159), .A2(n_379), .B1(n_649), .B2(n_1073), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_161), .A2(n_221), .B1(n_693), .B2(n_732), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g1388 ( .A1(n_165), .A2(n_395), .B1(n_1389), .B2(n_1390), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g1059 ( .A1(n_167), .A2(n_171), .B1(n_555), .B2(n_556), .Y(n_1059) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_168), .A2(n_331), .B1(n_742), .B2(n_1087), .Y(n_1086) );
AOI22x1_ASAP7_75t_L g835 ( .A1(n_172), .A2(n_836), .B1(n_837), .B2(n_859), .Y(n_835) );
INVx1_ASAP7_75t_L g859 ( .A(n_172), .Y(n_859) );
INVx1_ASAP7_75t_L g844 ( .A(n_174), .Y(n_844) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_176), .B(n_816), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_177), .A2(n_318), .B1(n_558), .B2(n_559), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g1074 ( .A1(n_178), .A2(n_262), .B1(n_693), .B2(n_939), .Y(n_1074) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_179), .A2(n_352), .B1(n_625), .B2(n_626), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g1391 ( .A1(n_180), .A2(n_409), .B1(n_558), .B2(n_559), .Y(n_1391) );
AOI22xp5_ASAP7_75t_L g1108 ( .A1(n_182), .A2(n_198), .B1(n_522), .B2(n_556), .Y(n_1108) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_183), .A2(n_385), .B1(n_652), .B2(n_1106), .Y(n_1105) );
CKINVDCx6p67_ASAP7_75t_R g975 ( .A(n_184), .Y(n_975) );
INVx1_ASAP7_75t_L g455 ( .A(n_185), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_185), .B(n_245), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_185), .B(n_480), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_186), .B(n_326), .Y(n_476) );
XNOR2x1_ASAP7_75t_L g1008 ( .A(n_187), .B(n_1009), .Y(n_1008) );
INVx1_ASAP7_75t_L g614 ( .A(n_188), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_189), .A2(n_213), .B1(n_496), .B2(n_499), .Y(n_495) );
INVx1_ASAP7_75t_L g564 ( .A(n_190), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g1077 ( .A1(n_191), .A2(n_388), .B1(n_555), .B2(n_556), .Y(n_1077) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_194), .B(n_597), .Y(n_596) );
AOI22xp33_ASAP7_75t_L g1095 ( .A1(n_196), .A2(n_202), .B1(n_538), .B2(n_1096), .Y(n_1095) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_197), .A2(n_211), .B1(n_606), .B2(n_607), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_199), .A2(n_319), .B1(n_772), .B2(n_774), .Y(n_890) );
CKINVDCx5p33_ASAP7_75t_R g1040 ( .A(n_200), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g1160 ( .A1(n_201), .A2(n_381), .B1(n_1151), .B2(n_1154), .Y(n_1160) );
INVx1_ASAP7_75t_L g1048 ( .A(n_203), .Y(n_1048) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_205), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g1051 ( .A(n_207), .Y(n_1051) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_208), .A2(n_392), .B1(n_517), .B2(n_718), .Y(n_717) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_209), .A2(n_333), .B1(n_1151), .B2(n_1154), .Y(n_1183) );
AOI22xp33_ASAP7_75t_L g1381 ( .A1(n_210), .A2(n_374), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
INVx1_ASAP7_75t_L g699 ( .A(n_214), .Y(n_699) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_215), .A2(n_418), .B1(n_828), .B2(n_829), .Y(n_827) );
INVx1_ASAP7_75t_L g568 ( .A(n_217), .Y(n_568) );
INVx1_ASAP7_75t_L g1175 ( .A(n_218), .Y(n_1175) );
AOI22xp5_ASAP7_75t_L g996 ( .A1(n_219), .A2(n_351), .B1(n_517), .B2(n_718), .Y(n_996) );
INVx1_ASAP7_75t_L g637 ( .A(n_220), .Y(n_637) );
CKINVDCx5p33_ASAP7_75t_R g955 ( .A(n_222), .Y(n_955) );
AOI22xp33_ASAP7_75t_L g1026 ( .A1(n_223), .A2(n_267), .B1(n_625), .B2(n_626), .Y(n_1026) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_224), .B(n_634), .Y(n_633) );
AOI22xp33_ASAP7_75t_L g1011 ( .A1(n_225), .A2(n_410), .B1(n_600), .B2(n_606), .Y(n_1011) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_226), .A2(n_420), .B1(n_459), .B2(n_630), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_227), .A2(n_347), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
INVx1_ASAP7_75t_L g797 ( .A(n_230), .Y(n_797) );
INVx1_ASAP7_75t_L g740 ( .A(n_232), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_234), .A2(n_362), .B1(n_772), .B2(n_773), .Y(n_771) );
INVx1_ASAP7_75t_L g577 ( .A(n_235), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_236), .A2(n_397), .B1(n_1140), .B2(n_1159), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_237), .A2(n_364), .B1(n_540), .B2(n_558), .Y(n_667) );
AOI22xp33_ASAP7_75t_L g1202 ( .A1(n_238), .A2(n_324), .B1(n_1164), .B2(n_1179), .Y(n_1202) );
AOI22xp33_ASAP7_75t_L g831 ( .A1(n_239), .A2(n_286), .B1(n_783), .B2(n_832), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g946 ( .A1(n_240), .A2(n_321), .B1(n_603), .B2(n_607), .Y(n_946) );
XOR2x2_ASAP7_75t_L g1083 ( .A(n_241), .B(n_1084), .Y(n_1083) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_243), .B(n_820), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_244), .A2(n_403), .B1(n_609), .B2(n_610), .Y(n_608) );
INVx1_ASAP7_75t_L g439 ( .A(n_245), .Y(n_439) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_246), .B(n_1070), .Y(n_1384) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_247), .A2(n_383), .B1(n_630), .B2(n_696), .Y(n_921) );
INVx1_ASAP7_75t_L g646 ( .A(n_248), .Y(n_646) );
OAI222xp33_ASAP7_75t_L g660 ( .A1(n_248), .A2(n_661), .B1(n_666), .B2(n_667), .C1(n_1424), .C2(n_1425), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_248), .B(n_667), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g957 ( .A(n_250), .Y(n_957) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_253), .A2(n_400), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g1163 ( .A1(n_257), .A2(n_275), .B1(n_1164), .B2(n_1165), .Y(n_1163) );
XNOR2x1_ASAP7_75t_L g805 ( .A(n_264), .B(n_806), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1079 ( .A1(n_265), .A2(n_301), .B1(n_552), .B2(n_553), .Y(n_1079) );
INVx1_ASAP7_75t_L g729 ( .A(n_266), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g695 ( .A1(n_268), .A2(n_288), .B1(n_630), .B2(n_696), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g684 ( .A1(n_270), .A2(n_315), .B1(n_556), .B2(n_685), .Y(n_684) );
AOI22xp33_ASAP7_75t_SL g925 ( .A1(n_272), .A2(n_335), .B1(n_870), .B2(n_926), .Y(n_925) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_273), .A2(n_649), .B(n_698), .Y(n_697) );
AOI221xp5_ASAP7_75t_L g1034 ( .A1(n_274), .A2(n_296), .B1(n_649), .B2(n_727), .C(n_1035), .Y(n_1034) );
AOI21xp5_ASAP7_75t_L g429 ( .A1(n_278), .A2(n_430), .B(n_456), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g1413 ( .A1(n_279), .A2(n_341), .B1(n_517), .B2(n_774), .Y(n_1413) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_280), .A2(n_387), .B1(n_485), .B2(n_490), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g1018 ( .A1(n_282), .A2(n_407), .B1(n_591), .B2(n_597), .Y(n_1018) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_284), .A2(n_310), .B1(n_1167), .B2(n_1168), .Y(n_1188) );
OAI21x1_ASAP7_75t_L g881 ( .A1(n_285), .A2(n_882), .B(n_900), .Y(n_881) );
NAND2xp5_ASAP7_75t_L g903 ( .A(n_285), .B(n_885), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1404 ( .A1(n_287), .A2(n_365), .B1(n_649), .B2(n_721), .Y(n_1404) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_291), .A2(n_369), .B1(n_558), .B2(n_682), .Y(n_1060) );
NAND2xp5_ASAP7_75t_L g1069 ( .A(n_292), .B(n_1070), .Y(n_1069) );
INVx1_ASAP7_75t_L g457 ( .A(n_294), .Y(n_457) );
INVx1_ASAP7_75t_L g987 ( .A(n_295), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_297), .B(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g879 ( .A(n_298), .Y(n_879) );
INVx1_ASAP7_75t_L g818 ( .A(n_299), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g758 ( .A1(n_302), .A2(n_342), .B1(n_505), .B2(n_538), .Y(n_758) );
INVx1_ASAP7_75t_L g1044 ( .A(n_303), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g1403 ( .A1(n_305), .A2(n_414), .B1(n_490), .B2(n_1050), .Y(n_1403) );
INVx1_ASAP7_75t_L g794 ( .A(n_306), .Y(n_794) );
INVx1_ASAP7_75t_L g1036 ( .A(n_308), .Y(n_1036) );
INVx1_ASAP7_75t_L g911 ( .A(n_310), .Y(n_911) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_310), .B(n_927), .Y(n_931) );
AOI22xp33_ASAP7_75t_L g1187 ( .A1(n_311), .A2(n_334), .B1(n_1124), .B2(n_1165), .Y(n_1187) );
AOI21xp5_ASAP7_75t_L g724 ( .A1(n_312), .A2(n_725), .B(n_728), .Y(n_724) );
AND2x4_ASAP7_75t_L g1141 ( .A(n_313), .B(n_1142), .Y(n_1141) );
HB1xp67_ASAP7_75t_L g1374 ( .A(n_313), .Y(n_1374) );
CKINVDCx5p33_ASAP7_75t_R g952 ( .A(n_316), .Y(n_952) );
AOI211x1_ASAP7_75t_L g560 ( .A1(n_320), .A2(n_561), .B(n_563), .C(n_571), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g845 ( .A(n_323), .B(n_846), .Y(n_845) );
INVx1_ASAP7_75t_L g781 ( .A(n_325), .Y(n_781) );
INVx1_ASAP7_75t_L g453 ( .A(n_326), .Y(n_453) );
INVxp67_ASAP7_75t_L g467 ( .A(n_326), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_328), .A2(n_412), .B1(n_825), .B2(n_826), .Y(n_824) );
INVx1_ASAP7_75t_L g898 ( .A(n_329), .Y(n_898) );
INVx1_ASAP7_75t_L g980 ( .A(n_330), .Y(n_980) );
INVxp67_ASAP7_75t_R g1177 ( .A(n_336), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g666 ( .A1(n_338), .A2(n_380), .B1(n_552), .B2(n_553), .Y(n_666) );
INVx2_ASAP7_75t_L g1126 ( .A(n_340), .Y(n_1126) );
INVx1_ASAP7_75t_SL g937 ( .A(n_347), .Y(n_937) );
NOR3xp33_ASAP7_75t_L g963 ( .A(n_347), .B(n_964), .C(n_965), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_348), .A2(n_394), .B1(n_573), .B2(n_813), .Y(n_920) );
INVx1_ASAP7_75t_L g743 ( .A(n_350), .Y(n_743) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_355), .A2(n_357), .B1(n_590), .B2(n_591), .Y(n_589) );
XNOR2x2_ASAP7_75t_L g1066 ( .A(n_356), .B(n_1067), .Y(n_1066) );
AOI21xp33_ASAP7_75t_L g1019 ( .A1(n_358), .A2(n_587), .B(n_1020), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_360), .A2(n_378), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g1104 ( .A1(n_361), .A2(n_382), .B1(n_632), .B2(n_742), .Y(n_1104) );
INVx1_ASAP7_75t_L g919 ( .A(n_370), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g1091 ( .A(n_371), .B(n_634), .Y(n_1091) );
INVx1_ASAP7_75t_L g984 ( .A(n_372), .Y(n_984) );
INVx1_ASAP7_75t_L g791 ( .A(n_376), .Y(n_791) );
NAND2xp5_ASAP7_75t_L g1405 ( .A(n_377), .B(n_799), .Y(n_1405) );
INVx1_ASAP7_75t_L g1147 ( .A(n_384), .Y(n_1147) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_389), .A2(n_393), .B1(n_632), .B2(n_748), .Y(n_893) );
INVx1_ASAP7_75t_L g1112 ( .A(n_391), .Y(n_1112) );
AOI22xp33_ASAP7_75t_L g592 ( .A1(n_396), .A2(n_416), .B1(n_593), .B2(n_594), .Y(n_592) );
AO22x2_ASAP7_75t_L g734 ( .A1(n_397), .A2(n_735), .B1(n_736), .B2(n_737), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_397), .Y(n_735) );
AND2x2_ASAP7_75t_L g940 ( .A(n_398), .B(n_846), .Y(n_940) );
INVx1_ASAP7_75t_L g575 ( .A(n_406), .Y(n_575) );
INVx1_ASAP7_75t_L g1243 ( .A(n_408), .Y(n_1243) );
INVx1_ASAP7_75t_L g989 ( .A(n_415), .Y(n_989) );
XOR2x2_ASAP7_75t_L g426 ( .A(n_419), .B(n_427), .Y(n_426) );
OAI22xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_1118), .B1(n_1419), .B2(n_1422), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_704), .B(n_1117), .Y(n_423) );
INVxp67_ASAP7_75t_L g1119 ( .A(n_424), .Y(n_1119) );
OA21x2_ASAP7_75t_L g1419 ( .A1(n_424), .A2(n_704), .B(n_1420), .Y(n_1419) );
XNOR2xp5_ASAP7_75t_L g424 ( .A(n_425), .B(n_543), .Y(n_424) );
HB1xp67_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2x1_ASAP7_75t_L g427 ( .A(n_428), .B(n_502), .Y(n_427) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_484), .C(n_495), .Y(n_428) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g563 ( .A1(n_431), .A2(n_564), .B(n_565), .Y(n_563) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx3_ASAP7_75t_SL g691 ( .A(n_433), .Y(n_691) );
INVx2_ASAP7_75t_L g727 ( .A(n_433), .Y(n_727) );
INVx2_ASAP7_75t_L g816 ( .A(n_433), .Y(n_816) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
BUFx3_ASAP7_75t_L g652 ( .A(n_434), .Y(n_652) );
INVx2_ASAP7_75t_L g842 ( .A(n_434), .Y(n_842) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_444), .Y(n_434) );
AND2x2_ASAP7_75t_L g501 ( .A(n_435), .B(n_498), .Y(n_501) );
AND2x2_ASAP7_75t_L g518 ( .A(n_435), .B(n_519), .Y(n_518) );
AND2x4_ASAP7_75t_L g523 ( .A(n_435), .B(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g590 ( .A(n_435), .B(n_498), .Y(n_590) );
AND2x2_ASAP7_75t_L g597 ( .A(n_435), .B(n_444), .Y(n_597) );
AND2x4_ASAP7_75t_L g600 ( .A(n_435), .B(n_509), .Y(n_600) );
AND2x4_ASAP7_75t_L g606 ( .A(n_435), .B(n_519), .Y(n_606) );
AND2x2_ASAP7_75t_L g622 ( .A(n_435), .B(n_519), .Y(n_622) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_443), .Y(n_435) );
INVx1_ASAP7_75t_L g489 ( .A(n_436), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
NAND2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx2_ASAP7_75t_L g442 ( .A(n_438), .Y(n_442) );
INVx3_ASAP7_75t_L g448 ( .A(n_438), .Y(n_448) );
NAND2xp33_ASAP7_75t_L g454 ( .A(n_438), .B(n_455), .Y(n_454) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_438), .Y(n_463) );
INVx1_ASAP7_75t_L g468 ( .A(n_438), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_439), .B(n_483), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_441), .B(n_442), .Y(n_440) );
OAI21xp5_ASAP7_75t_L g466 ( .A1(n_441), .A2(n_467), .B(n_468), .Y(n_466) );
AND2x2_ASAP7_75t_L g465 ( .A(n_443), .B(n_466), .Y(n_465) );
AND2x2_ASAP7_75t_L g488 ( .A(n_443), .B(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g508 ( .A(n_443), .Y(n_508) );
AND2x4_ASAP7_75t_L g487 ( .A(n_444), .B(n_488), .Y(n_487) );
AND2x4_ASAP7_75t_L g492 ( .A(n_444), .B(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g534 ( .A(n_444), .B(n_507), .Y(n_534) );
AND2x4_ASAP7_75t_L g591 ( .A(n_444), .B(n_493), .Y(n_591) );
AND2x2_ASAP7_75t_L g593 ( .A(n_444), .B(n_488), .Y(n_593) );
AND2x4_ASAP7_75t_L g610 ( .A(n_444), .B(n_507), .Y(n_610) );
AND2x4_ASAP7_75t_L g444 ( .A(n_445), .B(n_450), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x2_ASAP7_75t_L g461 ( .A(n_446), .B(n_462), .Y(n_461) );
AND2x4_ASAP7_75t_L g498 ( .A(n_446), .B(n_450), .Y(n_498) );
OR2x2_ASAP7_75t_L g510 ( .A(n_446), .B(n_511), .Y(n_510) );
AND2x4_ASAP7_75t_L g519 ( .A(n_446), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g446 ( .A(n_447), .B(n_449), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_448), .B(n_453), .Y(n_452) );
INVxp67_ASAP7_75t_L g480 ( .A(n_448), .Y(n_480) );
NAND3xp33_ASAP7_75t_L g478 ( .A(n_449), .B(n_479), .C(n_481), .Y(n_478) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g511 ( .A(n_451), .Y(n_511) );
AND2x2_ASAP7_75t_L g451 ( .A(n_452), .B(n_454), .Y(n_451) );
OAI21xp33_ASAP7_75t_L g456 ( .A1(n_457), .A2(n_458), .B(n_469), .Y(n_456) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
BUFx4f_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx5_ASAP7_75t_L g664 ( .A(n_460), .Y(n_664) );
BUFx2_ASAP7_75t_L g992 ( .A(n_460), .Y(n_992) );
BUFx2_ASAP7_75t_L g1089 ( .A(n_460), .Y(n_1089) );
AND2x4_ASAP7_75t_L g460 ( .A(n_461), .B(n_465), .Y(n_460) );
AND2x2_ASAP7_75t_L g588 ( .A(n_461), .B(n_465), .Y(n_588) );
AND2x4_ASAP7_75t_L g951 ( .A(n_461), .B(n_465), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
INVx1_ASAP7_75t_L g474 ( .A(n_463), .Y(n_474) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx4_ASAP7_75t_L g570 ( .A(n_471), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_471), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g820 ( .A(n_471), .Y(n_820) );
NOR2xp33_ASAP7_75t_L g878 ( .A(n_471), .B(n_879), .Y(n_878) );
INVx4_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx3_ASAP7_75t_L g847 ( .A(n_472), .Y(n_847) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_473), .Y(n_595) );
AO21x2_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_478), .Y(n_473) );
HB1xp67_ASAP7_75t_L g1398 ( .A(n_475), .Y(n_1398) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_480), .B(n_482), .Y(n_481) );
AND2x2_ASAP7_75t_L g493 ( .A(n_481), .B(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx3_ASAP7_75t_L g732 ( .A(n_486), .Y(n_732) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g567 ( .A(n_487), .Y(n_567) );
BUFx3_ASAP7_75t_L g634 ( .A(n_487), .Y(n_634) );
BUFx6f_ASAP7_75t_L g748 ( .A(n_487), .Y(n_748) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_487), .Y(n_813) );
BUFx8_ASAP7_75t_SL g939 ( .A(n_487), .Y(n_939) );
AND2x4_ASAP7_75t_L g497 ( .A(n_488), .B(n_498), .Y(n_497) );
AND2x4_ASAP7_75t_L g587 ( .A(n_488), .B(n_498), .Y(n_587) );
AND2x4_ASAP7_75t_L g507 ( .A(n_489), .B(n_508), .Y(n_507) );
BUFx3_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx4_ASAP7_75t_L g1052 ( .A(n_491), .Y(n_1052) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
INVx3_ASAP7_75t_L g574 ( .A(n_492), .Y(n_574) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_492), .Y(n_632) );
AND2x4_ASAP7_75t_L g515 ( .A(n_493), .B(n_509), .Y(n_515) );
AND2x4_ASAP7_75t_L g542 ( .A(n_493), .B(n_519), .Y(n_542) );
AND2x4_ASAP7_75t_L g601 ( .A(n_493), .B(n_509), .Y(n_601) );
AND2x4_ASAP7_75t_L g607 ( .A(n_493), .B(n_519), .Y(n_607) );
INVx2_ASAP7_75t_L g562 ( .A(n_496), .Y(n_562) );
BUFx3_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_497), .Y(n_649) );
BUFx3_ASAP7_75t_L g742 ( .A(n_497), .Y(n_742) );
INVx1_ASAP7_75t_L g917 ( .A(n_497), .Y(n_917) );
AND2x4_ASAP7_75t_L g529 ( .A(n_498), .B(n_507), .Y(n_529) );
AND2x4_ASAP7_75t_L g609 ( .A(n_498), .B(n_507), .Y(n_609) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx2_ASAP7_75t_L g576 ( .A(n_500), .Y(n_576) );
BUFx3_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
BUFx6f_ASAP7_75t_L g630 ( .A(n_501), .Y(n_630) );
INVx2_ASAP7_75t_L g723 ( .A(n_501), .Y(n_723) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_503), .B(n_516), .C(n_525), .D(n_535), .Y(n_502) );
BUFx3_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
BUFx6f_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
BUFx6f_ASAP7_75t_L g559 ( .A(n_506), .Y(n_559) );
BUFx6f_ASAP7_75t_L g682 ( .A(n_506), .Y(n_682) );
BUFx6f_ASAP7_75t_L g1096 ( .A(n_506), .Y(n_1096) );
AND2x4_ASAP7_75t_L g506 ( .A(n_507), .B(n_509), .Y(n_506) );
AND2x4_ASAP7_75t_L g539 ( .A(n_507), .B(n_519), .Y(n_539) );
AND2x4_ASAP7_75t_L g603 ( .A(n_507), .B(n_519), .Y(n_603) );
AND2x4_ASAP7_75t_L g604 ( .A(n_507), .B(n_524), .Y(n_604) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g524 ( .A(n_510), .Y(n_524) );
INVx1_ASAP7_75t_L g520 ( .A(n_511), .Y(n_520) );
BUFx2_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx2_ASAP7_75t_L g619 ( .A(n_514), .Y(n_619) );
INVx1_ASAP7_75t_L g658 ( .A(n_514), .Y(n_658) );
INVx3_ASAP7_75t_L g763 ( .A(n_514), .Y(n_763) );
INVx5_ASAP7_75t_L g887 ( .A(n_514), .Y(n_887) );
INVx1_ASAP7_75t_L g1390 ( .A(n_514), .Y(n_1390) );
INVx6_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
BUFx12f_ASAP7_75t_L g556 ( .A(n_515), .Y(n_556) );
BUFx8_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
BUFx6f_ASAP7_75t_L g687 ( .A(n_518), .Y(n_687) );
HB1xp67_ASAP7_75t_L g1098 ( .A(n_519), .Y(n_1098) );
BUFx3_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx6f_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
BUFx6f_ASAP7_75t_L g555 ( .A(n_523), .Y(n_555) );
BUFx6f_ASAP7_75t_L g618 ( .A(n_523), .Y(n_618) );
BUFx12f_ASAP7_75t_L g685 ( .A(n_523), .Y(n_685) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_523), .Y(n_1389) );
BUFx4f_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g680 ( .A(n_528), .Y(n_680) );
INVx3_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_529), .Y(n_552) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_529), .Y(n_625) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_532), .Y(n_714) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
BUFx5_ASAP7_75t_L g553 ( .A(n_534), .Y(n_553) );
BUFx6f_ASAP7_75t_L g626 ( .A(n_534), .Y(n_626) );
BUFx3_ASAP7_75t_L g830 ( .A(n_534), .Y(n_830) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx6f_ASAP7_75t_L g783 ( .A(n_538), .Y(n_783) );
BUFx12f_ASAP7_75t_L g855 ( .A(n_538), .Y(n_855) );
BUFx12f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
BUFx6f_ASAP7_75t_L g558 ( .A(n_539), .Y(n_558) );
BUFx6f_ASAP7_75t_L g870 ( .A(n_539), .Y(n_870) );
INVx4_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g550 ( .A(n_541), .Y(n_550) );
INVx2_ASAP7_75t_SL g623 ( .A(n_541), .Y(n_623) );
INVx2_ASAP7_75t_L g688 ( .A(n_541), .Y(n_688) );
INVx4_ASAP7_75t_L g718 ( .A(n_541), .Y(n_718) );
INVx4_ASAP7_75t_L g774 ( .A(n_541), .Y(n_774) );
INVx1_ASAP7_75t_L g926 ( .A(n_541), .Y(n_926) );
INVx1_ASAP7_75t_L g1063 ( .A(n_541), .Y(n_1063) );
INVx8_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AOI22xp33_ASAP7_75t_SL g543 ( .A1(n_544), .A2(n_642), .B1(n_702), .B2(n_703), .Y(n_543) );
INVx2_ASAP7_75t_SL g702 ( .A(n_544), .Y(n_702) );
OA22x2_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_579), .B1(n_580), .B2(n_641), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g641 ( .A(n_546), .Y(n_641) );
XNOR2x1_ASAP7_75t_L g546 ( .A(n_547), .B(n_578), .Y(n_546) );
NAND2x1_ASAP7_75t_L g547 ( .A(n_548), .B(n_560), .Y(n_547) );
AND4x1_ASAP7_75t_L g548 ( .A(n_549), .B(n_551), .C(n_554), .D(n_557), .Y(n_548) );
BUFx2_ASAP7_75t_L g832 ( .A(n_550), .Y(n_832) );
BUFx3_ASAP7_75t_L g776 ( .A(n_556), .Y(n_776) );
BUFx3_ASAP7_75t_L g785 ( .A(n_559), .Y(n_785) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
OAI21xp5_ASAP7_75t_SL g566 ( .A1(n_567), .A2(n_568), .B(n_569), .Y(n_566) );
INVx2_ASAP7_75t_SL g986 ( .A(n_567), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g571 ( .A1(n_572), .A2(n_575), .B1(n_576), .B2(n_577), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx3_ASAP7_75t_L g693 ( .A(n_574), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_574), .A2(n_747), .B1(n_794), .B2(n_795), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g983 ( .A1(n_574), .A2(n_984), .B1(n_985), .B2(n_987), .Y(n_983) );
INVx2_ASAP7_75t_L g1087 ( .A(n_574), .Y(n_1087) );
INVx2_ASAP7_75t_L g810 ( .A(n_576), .Y(n_810) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AOI22x1_ASAP7_75t_L g580 ( .A1(n_581), .A2(n_611), .B1(n_639), .B2(n_640), .Y(n_580) );
INVx2_ASAP7_75t_L g640 ( .A(n_581), .Y(n_640) );
INVx3_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
XNOR2x1_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_598), .Y(n_584) );
NAND4xp25_ASAP7_75t_L g585 ( .A(n_586), .B(n_589), .C(n_592), .D(n_596), .Y(n_585) );
INVx2_ASAP7_75t_L g956 ( .A(n_587), .Y(n_956) );
INVx2_ASAP7_75t_L g958 ( .A(n_590), .Y(n_958) );
INVx2_ASAP7_75t_L g953 ( .A(n_591), .Y(n_953) );
INVx3_ASAP7_75t_L g700 ( .A(n_594), .Y(n_700) );
INVx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
BUFx6f_ASAP7_75t_L g638 ( .A(n_595), .Y(n_638) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_595), .Y(n_755) );
NOR2xp33_ASAP7_75t_L g1020 ( .A(n_595), .B(n_1021), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .C(n_605), .D(n_608), .Y(n_598) );
INVxp67_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
BUFx2_ASAP7_75t_L g639 ( .A(n_612), .Y(n_639) );
XOR2xp5_ASAP7_75t_L g675 ( .A(n_612), .B(n_676), .Y(n_675) );
XNOR2x1_ASAP7_75t_L g612 ( .A(n_613), .B(n_615), .Y(n_612) );
CKINVDCx5p33_ASAP7_75t_R g613 ( .A(n_614), .Y(n_613) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_628), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_617), .B(n_620), .C(n_624), .D(n_627), .Y(n_616) );
BUFx4f_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
BUFx6f_ASAP7_75t_L g772 ( .A(n_622), .Y(n_772) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_625), .Y(n_828) );
BUFx2_ASAP7_75t_SL g779 ( .A(n_626), .Y(n_779) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_629), .B(n_631), .C(n_633), .D(n_635), .Y(n_628) );
INVx3_ASAP7_75t_L g744 ( .A(n_630), .Y(n_744) );
INVx3_ASAP7_75t_L g750 ( .A(n_632), .Y(n_750) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_638), .Y(n_636) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_638), .B(n_898), .Y(n_897) );
NOR2xp33_ASAP7_75t_L g918 ( .A(n_638), .B(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g1106 ( .A(n_638), .Y(n_1106) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_643), .Y(n_703) );
XNOR2x1_ASAP7_75t_L g643 ( .A(n_644), .B(n_675), .Y(n_643) );
AND2x4_ASAP7_75t_L g644 ( .A(n_645), .B(n_668), .Y(n_644) );
AOI21x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B(n_660), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_648), .B(n_655), .Y(n_647) );
BUFx2_ASAP7_75t_L g669 ( .A(n_648), .Y(n_669) );
INVx4_ASAP7_75t_L g790 ( .A(n_649), .Y(n_790) );
INVx1_ASAP7_75t_L g1045 ( .A(n_650), .Y(n_1045) );
INVx2_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
OAI21xp33_ASAP7_75t_L g751 ( .A1(n_651), .A2(n_752), .B(n_753), .Y(n_751) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
INVx1_ASAP7_75t_L g800 ( .A(n_652), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_659), .Y(n_655) );
INVxp67_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
AND2x2_ASAP7_75t_L g673 ( .A(n_657), .B(n_666), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_659), .Y(n_674) );
INVx1_ASAP7_75t_L g672 ( .A(n_661), .Y(n_672) );
AND2x2_ASAP7_75t_L g661 ( .A(n_662), .B(n_665), .Y(n_661) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx2_ASAP7_75t_L g696 ( .A(n_664), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g728 ( .A1(n_664), .A2(n_729), .B(n_730), .Y(n_728) );
OAI21xp5_ASAP7_75t_L g817 ( .A1(n_664), .A2(n_818), .B(n_819), .Y(n_817) );
OAI21xp33_ASAP7_75t_L g843 ( .A1(n_664), .A2(n_844), .B(n_845), .Y(n_843) );
INVx4_ASAP7_75t_L g876 ( .A(n_664), .Y(n_876) );
INVx2_ASAP7_75t_L g1386 ( .A(n_664), .Y(n_1386) );
INVx3_ASAP7_75t_L g1407 ( .A(n_664), .Y(n_1407) );
NAND4xp75_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .C(n_673), .D(n_674), .Y(n_668) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
XNOR2x1_ASAP7_75t_L g676 ( .A(n_677), .B(n_701), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_678), .B(n_683), .C(n_689), .D(n_694), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_681), .Y(n_678) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_682), .Y(n_823) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_686), .Y(n_683) );
BUFx3_ASAP7_75t_L g826 ( .A(n_685), .Y(n_826) );
BUFx3_ASAP7_75t_L g825 ( .A(n_687), .Y(n_825) );
HB1xp67_ASAP7_75t_L g1394 ( .A(n_687), .Y(n_1394) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
AND2x2_ASAP7_75t_L g694 ( .A(n_695), .B(n_697), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_905), .Y(n_704) );
NOR2xp67_ASAP7_75t_L g1117 ( .A(n_705), .B(n_905), .Y(n_1117) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
XNOR2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_803), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_709), .A2(n_766), .B1(n_767), .B2(n_802), .Y(n_708) );
INVx1_ASAP7_75t_L g802 ( .A(n_709), .Y(n_802) );
AO22x2_ASAP7_75t_L g709 ( .A1(n_710), .A2(n_734), .B1(n_764), .B2(n_765), .Y(n_709) );
INVx1_ASAP7_75t_L g764 ( .A(n_710), .Y(n_764) );
XOR2x2_ASAP7_75t_L g710 ( .A(n_711), .B(n_733), .Y(n_710) );
NOR2x1_ASAP7_75t_L g711 ( .A(n_712), .B(n_719), .Y(n_711) );
NAND4xp25_ASAP7_75t_L g712 ( .A(n_713), .B(n_715), .C(n_716), .D(n_717), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_724), .C(n_731), .Y(n_719) );
INVx2_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_722), .Y(n_792) );
INVx1_ASAP7_75t_L g1057 ( .A(n_722), .Y(n_1057) );
INVx2_ASAP7_75t_L g1073 ( .A(n_722), .Y(n_1073) );
INVx2_ASAP7_75t_L g1383 ( .A(n_722), .Y(n_1383) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g852 ( .A(n_723), .Y(n_852) );
INVx1_ASAP7_75t_L g982 ( .A(n_723), .Y(n_982) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g990 ( .A(n_727), .Y(n_990) );
INVx2_ASAP7_75t_L g765 ( .A(n_734), .Y(n_765) );
INVx1_ASAP7_75t_L g966 ( .A(n_734), .Y(n_966) );
INVx1_ASAP7_75t_L g969 ( .A(n_734), .Y(n_969) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_756), .Y(n_737) );
NOR3xp33_ASAP7_75t_SL g738 ( .A(n_739), .B(n_745), .C(n_751), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_739) );
INVx1_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
BUFx2_ASAP7_75t_L g809 ( .A(n_742), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B1(n_749), .B2(n_750), .Y(n_745) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
BUFx3_ASAP7_75t_L g1050 ( .A(n_748), .Y(n_1050) );
INVx1_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
NOR2xp33_ASAP7_75t_L g1035 ( .A(n_755), .B(n_1036), .Y(n_1035) );
NOR2xp33_ASAP7_75t_L g756 ( .A(n_757), .B(n_760), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_761), .B(n_762), .Y(n_760) );
INVx1_ASAP7_75t_L g766 ( .A(n_767), .Y(n_766) );
NAND3xp33_ASAP7_75t_L g768 ( .A(n_769), .B(n_777), .C(n_787), .Y(n_768) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g770 ( .A(n_771), .B(n_775), .Y(n_770) );
BUFx2_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NOR2x1_ASAP7_75t_L g777 ( .A(n_778), .B(n_780), .Y(n_777) );
OAI22x1_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_782), .B1(n_784), .B2(n_786), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g784 ( .A(n_785), .Y(n_784) );
NOR3xp33_ASAP7_75t_SL g787 ( .A(n_788), .B(n_793), .C(n_796), .Y(n_787) );
OAI22xp5_ASAP7_75t_SL g788 ( .A1(n_789), .A2(n_790), .B1(n_791), .B2(n_792), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g978 ( .A1(n_790), .A2(n_979), .B1(n_980), .B2(n_981), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1053 ( .A1(n_790), .A2(n_1054), .B1(n_1055), .B2(n_1056), .Y(n_1053) );
OAI21xp33_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_798), .B(n_801), .Y(n_796) );
INVx1_ASAP7_75t_L g798 ( .A(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_805), .B1(n_833), .B2(n_834), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
OR2x2_ASAP7_75t_L g806 ( .A(n_807), .B(n_821), .Y(n_806) );
NAND3xp33_ASAP7_75t_L g807 ( .A(n_808), .B(n_811), .C(n_814), .Y(n_807) );
BUFx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
HB1xp67_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
NAND4xp25_ASAP7_75t_L g821 ( .A(n_822), .B(n_824), .C(n_827), .D(n_831), .Y(n_821) );
BUFx2_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
XNOR2xp5_ASAP7_75t_L g834 ( .A(n_835), .B(n_860), .Y(n_834) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_838), .B(n_853), .Y(n_837) );
NAND3xp33_ASAP7_75t_L g838 ( .A(n_839), .B(n_848), .C(n_849), .Y(n_838) );
BUFx3_ASAP7_75t_L g840 ( .A(n_841), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_842), .Y(n_841) );
BUFx6f_ASAP7_75t_L g1071 ( .A(n_842), .Y(n_1071) );
INVx4_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g850 ( .A(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_852), .Y(n_851) );
NAND4xp25_ASAP7_75t_SL g853 ( .A(n_854), .B(n_856), .C(n_857), .D(n_858), .Y(n_853) );
OAI22xp5_ASAP7_75t_L g860 ( .A1(n_861), .A2(n_880), .B1(n_881), .B2(n_904), .Y(n_860) );
INVx1_ASAP7_75t_L g904 ( .A(n_861), .Y(n_904) );
XNOR2xp5_ASAP7_75t_L g861 ( .A(n_862), .B(n_863), .Y(n_861) );
NOR4xp75_ASAP7_75t_L g863 ( .A(n_864), .B(n_867), .C(n_871), .D(n_874), .Y(n_863) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_865), .B(n_866), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_869), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_872), .B(n_873), .Y(n_871) );
NAND2xp5_ASAP7_75t_SL g874 ( .A(n_875), .B(n_877), .Y(n_874) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
AND2x2_ASAP7_75t_L g882 ( .A(n_883), .B(n_891), .Y(n_882) );
NOR3xp33_ASAP7_75t_L g883 ( .A(n_884), .B(n_886), .C(n_888), .Y(n_883) );
INVx1_ASAP7_75t_L g884 ( .A(n_885), .Y(n_884) );
NOR3xp33_ASAP7_75t_L g902 ( .A(n_886), .B(n_895), .C(n_903), .Y(n_902) );
NOR2xp33_ASAP7_75t_L g901 ( .A(n_888), .B(n_892), .Y(n_901) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_889), .B(n_890), .Y(n_888) );
NOR2xp33_ASAP7_75t_L g891 ( .A(n_892), .B(n_895), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g892 ( .A(n_893), .B(n_894), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g895 ( .A(n_896), .B(n_899), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g900 ( .A(n_901), .B(n_902), .Y(n_900) );
XNOR2x1_ASAP7_75t_L g905 ( .A(n_906), .B(n_1002), .Y(n_905) );
AO22x2_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_908), .B1(n_970), .B2(n_1001), .Y(n_906) );
INVx2_ASAP7_75t_SL g907 ( .A(n_908), .Y(n_907) );
AO22x2_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_908) );
INVx1_ASAP7_75t_L g967 ( .A(n_909), .Y(n_967) );
XNOR2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_933), .Y(n_909) );
OAI21x1_ASAP7_75t_L g910 ( .A1(n_911), .A2(n_912), .B(n_930), .Y(n_910) );
AND2x2_ASAP7_75t_L g912 ( .A(n_913), .B(n_922), .Y(n_912) );
NAND3xp33_ASAP7_75t_L g930 ( .A(n_913), .B(n_931), .C(n_932), .Y(n_930) );
AND4x1_ASAP7_75t_L g913 ( .A(n_914), .B(n_915), .C(n_920), .D(n_921), .Y(n_913) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx2_ASAP7_75t_L g1382 ( .A(n_917), .Y(n_1382) );
NOR2xp33_ASAP7_75t_L g922 ( .A(n_923), .B(n_927), .Y(n_922) );
INVxp67_ASAP7_75t_SL g932 ( .A(n_923), .Y(n_932) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_928), .B(n_929), .Y(n_927) );
INVx1_ASAP7_75t_L g973 ( .A(n_933), .Y(n_973) );
NAND2x1_ASAP7_75t_L g933 ( .A(n_934), .B(n_959), .Y(n_933) );
NOR3xp33_ASAP7_75t_L g934 ( .A(n_935), .B(n_941), .C(n_945), .Y(n_934) );
OAI22xp33_ASAP7_75t_L g935 ( .A1(n_936), .A2(n_937), .B1(n_938), .B2(n_1426), .Y(n_935) );
INVx1_ASAP7_75t_L g964 ( .A(n_936), .Y(n_964) );
NOR2xp67_ASAP7_75t_L g941 ( .A(n_937), .B(n_942), .Y(n_941) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_937), .A2(n_946), .B1(n_947), .B2(n_1427), .Y(n_945) );
INVx1_ASAP7_75t_L g961 ( .A(n_938), .Y(n_961) );
NAND3xp33_ASAP7_75t_L g959 ( .A(n_942), .B(n_960), .C(n_963), .Y(n_959) );
AND2x2_ASAP7_75t_L g942 ( .A(n_943), .B(n_944), .Y(n_942) );
INVx1_ASAP7_75t_L g965 ( .A(n_946), .Y(n_965) );
INVx1_ASAP7_75t_L g962 ( .A(n_947), .Y(n_962) );
NOR2x1_ASAP7_75t_L g947 ( .A(n_948), .B(n_954), .Y(n_947) );
OAI22xp5_ASAP7_75t_L g948 ( .A1(n_949), .A2(n_950), .B1(n_952), .B2(n_953), .Y(n_948) );
INVx4_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI22xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_956), .B1(n_957), .B2(n_958), .Y(n_954) );
NOR2xp33_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
INVx1_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
INVx2_ASAP7_75t_L g970 ( .A(n_971), .Y(n_970) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_971), .Y(n_1001) );
OAI22xp5_ASAP7_75t_SL g971 ( .A1(n_972), .A2(n_973), .B1(n_974), .B2(n_1000), .Y(n_971) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVxp67_ASAP7_75t_SL g1000 ( .A(n_974), .Y(n_1000) );
XNOR2x1_ASAP7_75t_L g974 ( .A(n_975), .B(n_976), .Y(n_974) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_975), .A2(n_1145), .B1(n_1172), .B2(n_1173), .Y(n_1171) );
NAND2x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_993), .Y(n_976) );
NOR3xp33_ASAP7_75t_SL g977 ( .A(n_978), .B(n_983), .C(n_988), .Y(n_977) );
INVx2_ASAP7_75t_L g981 ( .A(n_982), .Y(n_981) );
INVx2_ASAP7_75t_L g985 ( .A(n_986), .Y(n_985) );
OAI21xp5_ASAP7_75t_L g988 ( .A1(n_989), .A2(n_990), .B(n_991), .Y(n_988) );
NOR2x1_ASAP7_75t_L g993 ( .A(n_994), .B(n_997), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_995), .B(n_996), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g997 ( .A(n_998), .B(n_999), .Y(n_997) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_1003), .A2(n_1065), .B1(n_1115), .B2(n_1116), .Y(n_1002) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1003), .Y(n_1115) );
OAI22xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B1(n_1038), .B2(n_1064), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1005), .Y(n_1004) );
INVx3_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
AO22x2_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1008), .B1(n_1022), .B2(n_1037), .Y(n_1006) );
INVx1_ASAP7_75t_L g1007 ( .A(n_1008), .Y(n_1007) );
OR2x2_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1015), .Y(n_1009) );
NAND4xp25_ASAP7_75t_L g1010 ( .A(n_1011), .B(n_1012), .C(n_1013), .D(n_1014), .Y(n_1010) );
NAND4xp25_ASAP7_75t_L g1015 ( .A(n_1016), .B(n_1017), .C(n_1018), .D(n_1019), .Y(n_1015) );
INVx1_ASAP7_75t_L g1037 ( .A(n_1022), .Y(n_1037) );
XNOR2x1_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1024), .Y(n_1022) );
NAND4xp75_ASAP7_75t_L g1024 ( .A(n_1025), .B(n_1028), .C(n_1031), .D(n_1034), .Y(n_1024) );
AND2x2_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1027), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1028 ( .A(n_1029), .B(n_1030), .Y(n_1028) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_1032), .B(n_1033), .Y(n_1031) );
BUFx3_ASAP7_75t_L g1038 ( .A(n_1039), .Y(n_1038) );
INVx4_ASAP7_75t_R g1064 ( .A(n_1039), .Y(n_1064) );
XNOR2x1_ASAP7_75t_L g1039 ( .A(n_1040), .B(n_1041), .Y(n_1039) );
AND2x4_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1058), .Y(n_1041) );
NOR3xp33_ASAP7_75t_L g1042 ( .A(n_1043), .B(n_1047), .C(n_1053), .Y(n_1042) );
OAI21xp5_ASAP7_75t_L g1043 ( .A1(n_1044), .A2(n_1045), .B(n_1046), .Y(n_1043) );
OAI22xp33_ASAP7_75t_L g1047 ( .A1(n_1048), .A2(n_1049), .B1(n_1051), .B2(n_1052), .Y(n_1047) );
INVx1_ASAP7_75t_L g1049 ( .A(n_1050), .Y(n_1049) );
INVxp67_ASAP7_75t_L g1056 ( .A(n_1057), .Y(n_1056) );
AND4x1_ASAP7_75t_L g1058 ( .A(n_1059), .B(n_1060), .C(n_1061), .D(n_1062), .Y(n_1058) );
OA21x2_ASAP7_75t_L g1065 ( .A1(n_1066), .A2(n_1081), .B(n_1113), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1113 ( .A(n_1066), .B(n_1114), .Y(n_1113) );
OAI21xp5_ASAP7_75t_L g1116 ( .A1(n_1066), .A2(n_1081), .B(n_1113), .Y(n_1116) );
OR2x2_ASAP7_75t_L g1067 ( .A(n_1068), .B(n_1076), .Y(n_1067) );
NAND4xp25_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1072), .C(n_1074), .D(n_1075), .Y(n_1068) );
INVx2_ASAP7_75t_L g1070 ( .A(n_1071), .Y(n_1070) );
NAND4xp25_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1078), .C(n_1079), .D(n_1080), .Y(n_1076) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1114 ( .A(n_1082), .Y(n_1114) );
XNOR2xp5_ASAP7_75t_L g1082 ( .A(n_1083), .B(n_1099), .Y(n_1082) );
NOR2x1_ASAP7_75t_L g1084 ( .A(n_1085), .B(n_1092), .Y(n_1084) );
NAND4xp25_ASAP7_75t_L g1085 ( .A(n_1086), .B(n_1088), .C(n_1090), .D(n_1091), .Y(n_1085) );
NAND4xp25_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1094), .C(n_1095), .D(n_1097), .Y(n_1092) );
BUFx3_ASAP7_75t_L g1411 ( .A(n_1096), .Y(n_1411) );
XOR2x2_ASAP7_75t_L g1099 ( .A(n_1100), .B(n_1112), .Y(n_1099) );
NOR2x1_ASAP7_75t_L g1100 ( .A(n_1101), .B(n_1107), .Y(n_1100) );
NAND4xp25_ASAP7_75t_L g1101 ( .A(n_1102), .B(n_1103), .C(n_1104), .D(n_1105), .Y(n_1101) );
NAND4xp25_ASAP7_75t_L g1107 ( .A(n_1108), .B(n_1109), .C(n_1110), .D(n_1111), .Y(n_1107) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1117), .Y(n_1120) );
OAI21xp5_ASAP7_75t_L g1118 ( .A1(n_1119), .A2(n_1120), .B(n_1121), .Y(n_1118) );
INVxp67_ASAP7_75t_L g1422 ( .A(n_1121), .Y(n_1422) );
OA21x2_ASAP7_75t_L g1121 ( .A1(n_1122), .A2(n_1129), .B(n_1368), .Y(n_1121) );
CKINVDCx5p33_ASAP7_75t_R g1122 ( .A(n_1123), .Y(n_1122) );
BUFx2_ASAP7_75t_L g1123 ( .A(n_1124), .Y(n_1123) );
INVx3_ASAP7_75t_L g1176 ( .A(n_1124), .Y(n_1176) );
AND2x4_ASAP7_75t_L g1124 ( .A(n_1125), .B(n_1128), .Y(n_1124) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1125), .B(n_1128), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1125), .B(n_1128), .Y(n_1164) );
AND2x4_ASAP7_75t_L g1167 ( .A(n_1125), .B(n_1141), .Y(n_1167) );
AND2x2_ASAP7_75t_L g1125 ( .A(n_1126), .B(n_1127), .Y(n_1125) );
AND3x4_ASAP7_75t_L g1140 ( .A(n_1126), .B(n_1141), .C(n_1143), .Y(n_1140) );
HB1xp67_ASAP7_75t_L g1372 ( .A(n_1126), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1128), .B(n_1146), .Y(n_1151) );
AND2x2_ASAP7_75t_L g1165 ( .A(n_1128), .B(n_1146), .Y(n_1165) );
AND2x4_ASAP7_75t_L g1179 ( .A(n_1128), .B(n_1146), .Y(n_1179) );
AOI21x1_ASAP7_75t_L g1129 ( .A1(n_1130), .A2(n_1283), .B(n_1332), .Y(n_1129) );
NAND5xp2_ASAP7_75t_L g1130 ( .A(n_1131), .B(n_1216), .C(n_1246), .D(n_1258), .E(n_1270), .Y(n_1130) );
AOI221xp5_ASAP7_75t_SL g1131 ( .A1(n_1132), .A2(n_1196), .B1(n_1206), .B2(n_1210), .C(n_1211), .Y(n_1131) );
A2O1A1Ixp33_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1180), .B(n_1184), .C(n_1189), .Y(n_1132) );
INVxp67_ASAP7_75t_SL g1366 ( .A(n_1133), .Y(n_1366) );
NAND2xp5_ASAP7_75t_L g1133 ( .A(n_1134), .B(n_1169), .Y(n_1133) );
INVx1_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
AOI211xp5_ASAP7_75t_L g1254 ( .A1(n_1135), .A2(n_1247), .B(n_1255), .C(n_1257), .Y(n_1254) );
OAI21xp33_ASAP7_75t_L g1273 ( .A1(n_1135), .A2(n_1274), .B(n_1276), .Y(n_1273) );
NAND2xp5_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1155), .Y(n_1135) );
INVx1_ASAP7_75t_L g1227 ( .A(n_1136), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1234 ( .A(n_1136), .B(n_1208), .Y(n_1234) );
AND2x2_ASAP7_75t_L g1251 ( .A(n_1136), .B(n_1223), .Y(n_1251) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1136), .B(n_1261), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1264 ( .A(n_1136), .B(n_1231), .Y(n_1264) );
NAND2xp5_ASAP7_75t_L g1293 ( .A(n_1136), .B(n_1195), .Y(n_1293) );
NAND2xp5_ASAP7_75t_L g1297 ( .A(n_1136), .B(n_1233), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1136), .B(n_1184), .Y(n_1345) );
CKINVDCx6p67_ASAP7_75t_R g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1194 ( .A(n_1137), .Y(n_1194) );
AND2x2_ASAP7_75t_L g1209 ( .A(n_1137), .B(n_1155), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1213 ( .A(n_1137), .B(n_1169), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1271 ( .A(n_1137), .B(n_1233), .Y(n_1271) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1137), .B(n_1286), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1137), .B(n_1208), .Y(n_1289) );
NOR2xp33_ASAP7_75t_L g1311 ( .A(n_1137), .B(n_1169), .Y(n_1311) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1137), .B(n_1170), .Y(n_1317) );
NAND2xp5_ASAP7_75t_L g1323 ( .A(n_1137), .B(n_1324), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1329 ( .A(n_1137), .B(n_1309), .Y(n_1329) );
OR2x6_ASAP7_75t_SL g1137 ( .A(n_1138), .B(n_1148), .Y(n_1137) );
OAI22xp5_ASAP7_75t_L g1138 ( .A1(n_1139), .A2(n_1144), .B1(n_1145), .B2(n_1147), .Y(n_1138) );
INVx1_ASAP7_75t_L g1139 ( .A(n_1140), .Y(n_1139) );
NAND2xp5_ASAP7_75t_L g1145 ( .A(n_1141), .B(n_1146), .Y(n_1145) );
AND2x4_ASAP7_75t_L g1159 ( .A(n_1141), .B(n_1146), .Y(n_1159) );
AND2x4_ASAP7_75t_L g1168 ( .A(n_1141), .B(n_1146), .Y(n_1168) );
AOI21xp5_ASAP7_75t_L g1418 ( .A1(n_1143), .A2(n_1371), .B(n_1374), .Y(n_1418) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_1145), .A2(n_1172), .B1(n_1242), .B2(n_1243), .C(n_1244), .Y(n_1241) );
OAI22xp5_ASAP7_75t_L g1148 ( .A1(n_1149), .A2(n_1150), .B1(n_1152), .B2(n_1153), .Y(n_1148) );
INVx1_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
XOR2x2_ASAP7_75t_L g1400 ( .A(n_1152), .B(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1153 ( .A(n_1154), .Y(n_1153) );
NAND2xp5_ASAP7_75t_L g1180 ( .A(n_1155), .B(n_1181), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1220 ( .A(n_1155), .B(n_1208), .Y(n_1220) );
AND2x2_ASAP7_75t_L g1250 ( .A(n_1155), .B(n_1251), .Y(n_1250) );
NAND2xp5_ASAP7_75t_L g1342 ( .A(n_1155), .B(n_1234), .Y(n_1342) );
AND2x2_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1161), .Y(n_1155) );
NOR2xp33_ASAP7_75t_L g1190 ( .A(n_1156), .B(n_1181), .Y(n_1190) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1156), .B(n_1162), .Y(n_1215) );
CKINVDCx5p33_ASAP7_75t_R g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1233 ( .A(n_1157), .B(n_1162), .Y(n_1233) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1157), .B(n_1161), .Y(n_1262) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1157), .B(n_1181), .Y(n_1300) );
OR2x2_ASAP7_75t_L g1340 ( .A(n_1157), .B(n_1181), .Y(n_1340) );
AND2x4_ASAP7_75t_SL g1157 ( .A(n_1158), .B(n_1160), .Y(n_1157) );
INVx2_ASAP7_75t_SL g1205 ( .A(n_1159), .Y(n_1205) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1161), .Y(n_1222) );
AND2x2_ASAP7_75t_L g1267 ( .A(n_1161), .B(n_1223), .Y(n_1267) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1161), .B(n_1223), .Y(n_1324) );
INVx1_ASAP7_75t_L g1161 ( .A(n_1162), .Y(n_1161) );
NAND2xp5_ASAP7_75t_L g1162 ( .A(n_1163), .B(n_1166), .Y(n_1162) );
INVx3_ASAP7_75t_L g1172 ( .A(n_1167), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1169), .B(n_1186), .Y(n_1210) );
NOR2xp33_ASAP7_75t_L g1269 ( .A(n_1169), .B(n_1225), .Y(n_1269) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1169), .B(n_1200), .Y(n_1272) );
NAND2xp5_ASAP7_75t_L g1291 ( .A(n_1169), .B(n_1199), .Y(n_1291) );
INVx3_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
AND2x2_ASAP7_75t_L g1195 ( .A(n_1170), .B(n_1185), .Y(n_1195) );
OR2x2_ASAP7_75t_L g1231 ( .A(n_1170), .B(n_1186), .Y(n_1231) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1170), .Y(n_1249) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1170), .B(n_1186), .Y(n_1305) );
OR2x2_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1174), .Y(n_1170) );
OAI22xp5_ASAP7_75t_L g1174 ( .A1(n_1175), .A2(n_1176), .B1(n_1177), .B2(n_1178), .Y(n_1174) );
INVx2_ASAP7_75t_L g1178 ( .A(n_1179), .Y(n_1178) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1180), .Y(n_1362) );
CKINVDCx6p67_ASAP7_75t_R g1208 ( .A(n_1181), .Y(n_1208) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1181), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1282 ( .A(n_1181), .B(n_1262), .Y(n_1282) );
AND2x2_ASAP7_75t_L g1286 ( .A(n_1181), .B(n_1215), .Y(n_1286) );
OAI322xp33_ASAP7_75t_L g1292 ( .A1(n_1181), .A2(n_1198), .A3(n_1293), .B1(n_1294), .B2(n_1297), .C1(n_1298), .C2(n_1300), .Y(n_1292) );
AND2x2_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1183), .Y(n_1181) );
AOI221xp5_ASAP7_75t_L g1270 ( .A1(n_1184), .A2(n_1271), .B1(n_1272), .B2(n_1273), .C(n_1277), .Y(n_1270) );
INVx3_ASAP7_75t_L g1312 ( .A(n_1184), .Y(n_1312) );
OAI21xp5_ASAP7_75t_L g1313 ( .A1(n_1184), .A2(n_1314), .B(n_1315), .Y(n_1313) );
INVx3_ASAP7_75t_L g1184 ( .A(n_1185), .Y(n_1184) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1185), .B(n_1201), .Y(n_1225) );
NAND2xp5_ASAP7_75t_L g1236 ( .A(n_1185), .B(n_1201), .Y(n_1236) );
INVx2_ASAP7_75t_L g1185 ( .A(n_1186), .Y(n_1185) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1186), .B(n_1201), .Y(n_1279) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1187), .B(n_1188), .Y(n_1186) );
NAND2xp5_ASAP7_75t_L g1189 ( .A(n_1190), .B(n_1191), .Y(n_1189) );
NAND2xp5_ASAP7_75t_L g1316 ( .A(n_1190), .B(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1192), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1245 ( .A(n_1192), .B(n_1221), .Y(n_1245) );
NOR2xp33_ASAP7_75t_L g1252 ( .A(n_1192), .B(n_1253), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1195), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1193), .B(n_1215), .Y(n_1237) );
NOR2xp33_ASAP7_75t_L g1328 ( .A(n_1193), .B(n_1201), .Y(n_1328) );
NOR2xp33_ASAP7_75t_L g1357 ( .A(n_1193), .B(n_1358), .Y(n_1357) );
O2A1O1Ixp33_ASAP7_75t_L g1367 ( .A1(n_1193), .A2(n_1228), .B(n_1237), .C(n_1281), .Y(n_1367) );
INVx3_ASAP7_75t_L g1193 ( .A(n_1194), .Y(n_1193) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1195), .B(n_1198), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1364 ( .A(n_1195), .B(n_1267), .C(n_1328), .Y(n_1364) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1196), .Y(n_1350) );
INVx3_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
INVx3_ASAP7_75t_L g1197 ( .A(n_1198), .Y(n_1197) );
NOR2xp33_ASAP7_75t_L g1211 ( .A(n_1198), .B(n_1212), .Y(n_1211) );
INVx3_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1238 ( .A(n_1200), .B(n_1239), .Y(n_1238) );
A2O1A1Ixp33_ASAP7_75t_L g1361 ( .A1(n_1200), .A2(n_1230), .B(n_1362), .C(n_1363), .Y(n_1361) );
INVx3_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1201), .B(n_1230), .Y(n_1229) );
INVx1_ASAP7_75t_L g1296 ( .A(n_1201), .Y(n_1296) );
NAND2xp5_ASAP7_75t_L g1337 ( .A(n_1201), .B(n_1305), .Y(n_1337) );
AND2x4_ASAP7_75t_L g1201 ( .A(n_1202), .B(n_1203), .Y(n_1201) );
INVx2_ASAP7_75t_L g1204 ( .A(n_1205), .Y(n_1204) );
INVx1_ASAP7_75t_L g1206 ( .A(n_1207), .Y(n_1206) );
NAND2xp5_ASAP7_75t_L g1207 ( .A(n_1208), .B(n_1209), .Y(n_1207) );
AND2x2_ASAP7_75t_SL g1214 ( .A(n_1208), .B(n_1215), .Y(n_1214) );
NOR2xp33_ASAP7_75t_L g1256 ( .A(n_1208), .B(n_1253), .Y(n_1256) );
AND2x2_ASAP7_75t_L g1261 ( .A(n_1208), .B(n_1262), .Y(n_1261) );
NAND2xp5_ASAP7_75t_L g1353 ( .A(n_1208), .B(n_1233), .Y(n_1353) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1209), .B(n_1223), .Y(n_1314) );
INVx1_ASAP7_75t_L g1339 ( .A(n_1209), .Y(n_1339) );
AOI322xp5_ASAP7_75t_L g1335 ( .A1(n_1210), .A2(n_1259), .A3(n_1299), .B1(n_1336), .B2(n_1338), .C1(n_1340), .C2(n_1341), .Y(n_1335) );
INVxp67_ASAP7_75t_SL g1302 ( .A(n_1212), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1212 ( .A(n_1213), .B(n_1214), .Y(n_1212) );
INVxp67_ASAP7_75t_L g1280 ( .A(n_1213), .Y(n_1280) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1214), .Y(n_1268) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1215), .B(n_1234), .Y(n_1239) );
AOI222xp33_ASAP7_75t_L g1258 ( .A1(n_1215), .A2(n_1259), .B1(n_1263), .B2(n_1264), .C1(n_1265), .C2(n_1269), .Y(n_1258) );
OR2x2_ASAP7_75t_L g1327 ( .A(n_1215), .B(n_1262), .Y(n_1327) );
INVxp33_ASAP7_75t_L g1358 ( .A(n_1215), .Y(n_1358) );
NOR3xp33_ASAP7_75t_L g1216 ( .A(n_1217), .B(n_1235), .C(n_1245), .Y(n_1216) );
OAI32xp33_ASAP7_75t_L g1217 ( .A1(n_1218), .A2(n_1225), .A3(n_1226), .B1(n_1228), .B2(n_1232), .Y(n_1217) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
NAND2xp5_ASAP7_75t_L g1219 ( .A(n_1220), .B(n_1221), .Y(n_1219) );
INVx1_ASAP7_75t_L g1319 ( .A(n_1220), .Y(n_1319) );
INVx1_ASAP7_75t_L g1346 ( .A(n_1221), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1223), .Y(n_1221) );
AOI321xp33_ASAP7_75t_L g1326 ( .A1(n_1223), .A2(n_1272), .A3(n_1327), .B1(n_1328), .B2(n_1329), .C(n_1330), .Y(n_1326) );
INVx1_ASAP7_75t_L g1223 ( .A(n_1224), .Y(n_1223) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1225), .Y(n_1263) );
OAI211xp5_ASAP7_75t_L g1360 ( .A1(n_1225), .A2(n_1316), .B(n_1361), .C(n_1364), .Y(n_1360) );
CKINVDCx14_ASAP7_75t_R g1226 ( .A(n_1227), .Y(n_1226) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1231), .Y(n_1230) );
OAI221xp5_ASAP7_75t_L g1303 ( .A1(n_1231), .A2(n_1304), .B1(n_1306), .B2(n_1307), .C(n_1310), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1232 ( .A(n_1233), .B(n_1234), .Y(n_1232) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1233), .Y(n_1253) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1233), .B(n_1288), .Y(n_1287) );
NAND3xp33_ASAP7_75t_L g1310 ( .A(n_1233), .B(n_1311), .C(n_1312), .Y(n_1310) );
AND2x2_ASAP7_75t_L g1349 ( .A(n_1233), .B(n_1251), .Y(n_1349) );
OAI211xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1237), .B(n_1238), .C(n_1240), .Y(n_1235) );
INVx1_ASAP7_75t_L g1257 ( .A(n_1236), .Y(n_1257) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1238), .Y(n_1363) );
INVx2_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
BUFx3_ASAP7_75t_L g1331 ( .A(n_1241), .Y(n_1331) );
AOI211xp5_ASAP7_75t_L g1246 ( .A1(n_1247), .A2(n_1250), .B(n_1252), .C(n_1254), .Y(n_1246) );
INVx2_ASAP7_75t_L g1247 ( .A(n_1248), .Y(n_1247) );
BUFx2_ASAP7_75t_L g1248 ( .A(n_1249), .Y(n_1248) );
INVx1_ASAP7_75t_L g1275 ( .A(n_1249), .Y(n_1275) );
NOR2xp33_ASAP7_75t_L g1295 ( .A(n_1249), .B(n_1296), .Y(n_1295) );
INVx1_ASAP7_75t_L g1276 ( .A(n_1250), .Y(n_1276) );
NOR2xp33_ASAP7_75t_L g1325 ( .A(n_1255), .B(n_1294), .Y(n_1325) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1257), .B(n_1275), .Y(n_1299) );
AOI221xp5_ASAP7_75t_L g1318 ( .A1(n_1257), .A2(n_1319), .B1(n_1320), .B2(n_1322), .C(n_1325), .Y(n_1318) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1262), .Y(n_1309) );
AOI21xp5_ASAP7_75t_L g1301 ( .A1(n_1263), .A2(n_1302), .B(n_1303), .Y(n_1301) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1268), .Y(n_1265) );
INVx1_ASAP7_75t_L g1266 ( .A(n_1267), .Y(n_1266) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1269), .Y(n_1359) );
INVx1_ASAP7_75t_L g1274 ( .A(n_1275), .Y(n_1274) );
NAND2xp5_ASAP7_75t_L g1348 ( .A(n_1275), .B(n_1349), .Y(n_1348) );
AOI21xp5_ASAP7_75t_L g1277 ( .A1(n_1278), .A2(n_1280), .B(n_1281), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
O2A1O1Ixp33_ASAP7_75t_L g1365 ( .A1(n_1279), .A2(n_1287), .B(n_1366), .C(n_1367), .Y(n_1365) );
INVx1_ASAP7_75t_L g1281 ( .A(n_1282), .Y(n_1281) );
NAND5xp2_ASAP7_75t_L g1283 ( .A(n_1284), .B(n_1301), .C(n_1313), .D(n_1318), .E(n_1326), .Y(n_1283) );
O2A1O1Ixp33_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1287), .B(n_1290), .C(n_1292), .Y(n_1284) );
INVx1_ASAP7_75t_L g1355 ( .A(n_1286), .Y(n_1355) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1287), .Y(n_1306) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1289), .Y(n_1288) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1289), .B(n_1309), .Y(n_1308) );
NAND2xp5_ASAP7_75t_SL g1338 ( .A(n_1289), .B(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1294 ( .A(n_1295), .Y(n_1294) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1304 ( .A(n_1305), .Y(n_1304) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
INVxp67_ASAP7_75t_SL g1315 ( .A(n_1316), .Y(n_1315) );
AOI21xp33_ASAP7_75t_L g1351 ( .A1(n_1320), .A2(n_1352), .B(n_1354), .Y(n_1351) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1323), .Y(n_1322) );
INVx1_ASAP7_75t_L g1330 ( .A(n_1331), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1332 ( .A(n_1333), .B(n_1365), .Y(n_1332) );
NOR2xp33_ASAP7_75t_L g1333 ( .A(n_1334), .B(n_1360), .Y(n_1333) );
NAND3xp33_ASAP7_75t_L g1334 ( .A(n_1335), .B(n_1343), .C(n_1351), .Y(n_1334) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1337), .Y(n_1336) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
A2O1A1Ixp33_ASAP7_75t_L g1343 ( .A1(n_1344), .A2(n_1346), .B(n_1347), .C(n_1350), .Y(n_1343) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1347 ( .A(n_1348), .Y(n_1347) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1353), .Y(n_1352) );
AOI21xp33_ASAP7_75t_L g1354 ( .A1(n_1355), .A2(n_1356), .B(n_1359), .Y(n_1354) );
INVxp33_ASAP7_75t_L g1356 ( .A(n_1357), .Y(n_1356) );
BUFx2_ASAP7_75t_SL g1369 ( .A(n_1370), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1371), .B(n_1373), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1396 ( .A(n_1371), .B(n_1397), .Y(n_1396) );
NAND3xp33_ASAP7_75t_L g1421 ( .A(n_1371), .B(n_1374), .C(n_1398), .Y(n_1421) );
INVx1_ASAP7_75t_L g1371 ( .A(n_1372), .Y(n_1371) );
AO21x1_ASAP7_75t_L g1415 ( .A1(n_1372), .A2(n_1416), .B(n_1418), .Y(n_1415) );
NOR2xp33_ASAP7_75t_L g1397 ( .A(n_1373), .B(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVxp67_ASAP7_75t_SL g1377 ( .A(n_1378), .Y(n_1377) );
OR2x2_ASAP7_75t_L g1378 ( .A(n_1379), .B(n_1387), .Y(n_1378) );
NAND4xp25_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1381), .C(n_1384), .D(n_1385), .Y(n_1379) );
NAND4xp25_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1391), .C(n_1392), .D(n_1393), .Y(n_1387) );
BUFx2_ASAP7_75t_L g1399 ( .A(n_1400), .Y(n_1399) );
NOR2x1_ASAP7_75t_L g1401 ( .A(n_1402), .B(n_1408), .Y(n_1401) );
NAND4xp25_ASAP7_75t_L g1402 ( .A(n_1403), .B(n_1404), .C(n_1405), .D(n_1406), .Y(n_1402) );
NAND4xp25_ASAP7_75t_L g1408 ( .A(n_1409), .B(n_1410), .C(n_1412), .D(n_1413), .Y(n_1408) );
BUFx2_ASAP7_75t_L g1414 ( .A(n_1415), .Y(n_1414) );
CKINVDCx5p33_ASAP7_75t_R g1416 ( .A(n_1417), .Y(n_1416) );
INVx2_ASAP7_75t_SL g1420 ( .A(n_1421), .Y(n_1420) );
endmodule