module fake_jpeg_2144_n_625 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_625);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_625;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_384;
wire n_296;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

BUFx4f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_18),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

BUFx12_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_8),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

BUFx12_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g49 ( 
.A(n_8),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_2),
.B(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_0),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_6),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx4f_ASAP7_75t_SL g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_5),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_62),
.Y(n_131)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_63),
.Y(n_166)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_65),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_31),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_66),
.B(n_71),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_67),
.Y(n_153)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_69),
.Y(n_173)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_49),
.Y(n_70)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_70),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_50),
.B(n_17),
.Y(n_71)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

INVx3_ASAP7_75t_SL g142 ( 
.A(n_72),
.Y(n_142)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_75),
.Y(n_163)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g159 ( 
.A(n_76),
.Y(n_159)
);

AOI21xp33_ASAP7_75t_L g77 ( 
.A1(n_23),
.A2(n_9),
.B(n_15),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_77),
.B(n_102),
.Y(n_136)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_78),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_79),
.Y(n_195)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx3_ASAP7_75t_SL g148 ( 
.A(n_81),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx6_ASAP7_75t_L g138 ( 
.A(n_82),
.Y(n_138)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_32),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_84),
.B(n_88),
.Y(n_188)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_85),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_86),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx6_ASAP7_75t_L g187 ( 
.A(n_87),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_32),
.B(n_16),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_31),
.B(n_8),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_90),
.B(n_106),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_91),
.Y(n_160)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_40),
.Y(n_92)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_92),
.Y(n_167)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_93),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_40),
.Y(n_94)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_94),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_97),
.Y(n_189)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_29),
.Y(n_98)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_98),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_53),
.Y(n_99)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_57),
.Y(n_100)
);

INVx8_ASAP7_75t_L g198 ( 
.A(n_100),
.Y(n_198)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_41),
.Y(n_101)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_52),
.B(n_10),
.Y(n_102)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_61),
.Y(n_103)
);

INVx4_ASAP7_75t_L g180 ( 
.A(n_103),
.Y(n_180)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_104),
.Y(n_171)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_29),
.Y(n_105)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_105),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_34),
.B(n_10),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_107),
.Y(n_156)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_43),
.Y(n_108)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_10),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_110),
.B(n_120),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_59),
.Y(n_111)
);

BUFx4f_ASAP7_75t_SL g144 ( 
.A(n_111),
.Y(n_144)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_48),
.Y(n_112)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_112),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx4_ASAP7_75t_L g206 ( 
.A(n_113),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_59),
.Y(n_114)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_114),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_60),
.Y(n_115)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_115),
.Y(n_176)
);

INVx11_ASAP7_75t_L g116 ( 
.A(n_48),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_34),
.Y(n_117)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_117),
.Y(n_179)
);

INVx11_ASAP7_75t_L g118 ( 
.A(n_58),
.Y(n_118)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_118),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_27),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_119),
.A2(n_51),
.B1(n_38),
.B2(n_54),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_25),
.B(n_7),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_27),
.Y(n_121)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_121),
.Y(n_183)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_43),
.Y(n_122)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_22),
.Y(n_123)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_123),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_60),
.Y(n_124)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_125),
.Y(n_207)
);

BUFx5_ASAP7_75t_L g126 ( 
.A(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_45),
.Y(n_127)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_27),
.Y(n_128)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_128),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g134 ( 
.A1(n_127),
.A2(n_20),
.B1(n_45),
.B2(n_44),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g275 ( 
.A1(n_134),
.A2(n_135),
.B1(n_149),
.B2(n_36),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_74),
.A2(n_20),
.B1(n_45),
.B2(n_44),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_64),
.B(n_33),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_146),
.B(n_152),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_79),
.A2(n_94),
.B1(n_124),
.B2(n_87),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_70),
.B(n_47),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_76),
.A2(n_20),
.B1(n_25),
.B2(n_33),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_154),
.A2(n_186),
.B1(n_114),
.B2(n_100),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_65),
.B(n_54),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_157),
.B(n_165),
.Y(n_216)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_85),
.B(n_20),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_162),
.B(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_80),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_67),
.B(n_39),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_112),
.B(n_22),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_0),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_72),
.B(n_39),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_170),
.B(n_178),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_116),
.A2(n_44),
.B1(n_38),
.B2(n_51),
.Y(n_175)
);

OA22x2_ASAP7_75t_L g229 ( 
.A1(n_175),
.A2(n_37),
.B1(n_56),
.B2(n_113),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_81),
.B(n_47),
.Y(n_178)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_92),
.Y(n_184)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_184),
.Y(n_217)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_122),
.Y(n_190)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_190),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_96),
.B(n_58),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_91),
.Y(n_202)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_202),
.Y(n_254)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_203),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_82),
.B(n_58),
.Y(n_209)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g344 ( 
.A(n_213),
.Y(n_344)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_174),
.Y(n_214)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_214),
.Y(n_287)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_136),
.A2(n_37),
.B(n_55),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_218),
.B(n_240),
.Y(n_291)
);

BUFx3_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g321 ( 
.A(n_219),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g220 ( 
.A(n_151),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_179),
.Y(n_221)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_221),
.Y(n_296)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_131),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g294 ( 
.A(n_222),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_169),
.A2(n_56),
.B(n_55),
.Y(n_223)
);

OA21x2_ASAP7_75t_L g332 ( 
.A1(n_223),
.A2(n_229),
.B(n_260),
.Y(n_332)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

INVx3_ASAP7_75t_L g225 ( 
.A(n_155),
.Y(n_225)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_225),
.Y(n_331)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_131),
.Y(n_226)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_226),
.Y(n_302)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_160),
.Y(n_227)
);

INVx3_ASAP7_75t_L g345 ( 
.A(n_227),
.Y(n_345)
);

INVx3_ASAP7_75t_L g228 ( 
.A(n_153),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_228),
.Y(n_320)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_230),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_133),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_231),
.B(n_234),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g233 ( 
.A(n_201),
.Y(n_233)
);

INVx5_ASAP7_75t_L g312 ( 
.A(n_233),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_188),
.B(n_115),
.Y(n_234)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_143),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g343 ( 
.A(n_236),
.Y(n_343)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_237),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_193),
.A2(n_103),
.B1(n_111),
.B2(n_107),
.Y(n_239)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_239),
.A2(n_248),
.B1(n_251),
.B2(n_275),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_241),
.A2(n_156),
.B1(n_144),
.B2(n_195),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_201),
.Y(n_243)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_243),
.Y(n_315)
);

INVx2_ASAP7_75t_SL g244 ( 
.A(n_147),
.Y(n_244)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_244),
.Y(n_289)
);

AOI22xp33_ASAP7_75t_L g245 ( 
.A1(n_134),
.A2(n_99),
.B1(n_97),
.B2(n_95),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_245),
.A2(n_239),
.B1(n_187),
.B2(n_212),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_145),
.A2(n_86),
.B1(n_26),
.B2(n_30),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g299 ( 
.A(n_246),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_133),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_208),
.A2(n_211),
.B1(n_204),
.B2(n_143),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_177),
.B(n_12),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_249),
.B(n_255),
.Y(n_305)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_250),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_204),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_129),
.Y(n_252)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_252),
.Y(n_335)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_199),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_253),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_142),
.Y(n_255)
);

INVx8_ASAP7_75t_L g256 ( 
.A(n_132),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

BUFx8_ASAP7_75t_L g257 ( 
.A(n_142),
.Y(n_257)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_257),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_166),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_258),
.Y(n_334)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_199),
.Y(n_259)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_259),
.Y(n_304)
);

NAND2xp33_ASAP7_75t_SL g260 ( 
.A(n_162),
.B(n_0),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_159),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_262),
.B(n_267),
.Y(n_311)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_130),
.Y(n_263)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_137),
.Y(n_266)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_266),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_140),
.B(n_13),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

OAI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_135),
.A2(n_26),
.B1(n_30),
.B2(n_36),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_144),
.B1(n_156),
.B2(n_148),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_163),
.B(n_13),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_270),
.B(n_273),
.Y(n_317)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_176),
.Y(n_271)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_271),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_132),
.Y(n_272)
);

INVx8_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_161),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_139),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_277),
.Y(n_322)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_175),
.A2(n_30),
.B1(n_24),
.B2(n_36),
.Y(n_276)
);

AOI22xp33_ASAP7_75t_SL g313 ( 
.A1(n_276),
.A2(n_284),
.B1(n_286),
.B2(n_180),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_168),
.B(n_7),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_159),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_278),
.B(n_279),
.Y(n_326)
);

INVx5_ASAP7_75t_L g279 ( 
.A(n_181),
.Y(n_279)
);

INVx5_ASAP7_75t_L g280 ( 
.A(n_181),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_280),
.B(n_281),
.Y(n_338)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_200),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_282),
.B(n_283),
.Y(n_339)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_148),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_141),
.Y(n_284)
);

HB1xp67_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_285),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_342)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_192),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_265),
.B(n_205),
.C(n_191),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_292),
.B(n_300),
.C(n_255),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_297),
.A2(n_303),
.B1(n_319),
.B2(n_325),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_216),
.B(n_191),
.C(n_206),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_218),
.B(n_210),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_301),
.B(n_341),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g303 ( 
.A1(n_241),
.A2(n_158),
.B1(n_187),
.B2(n_212),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_313),
.Y(n_362)
);

AOI22xp33_ASAP7_75t_L g376 ( 
.A1(n_314),
.A2(n_222),
.B1(n_283),
.B2(n_257),
.Y(n_376)
);

AOI32xp33_ASAP7_75t_L g318 ( 
.A1(n_261),
.A2(n_206),
.A3(n_180),
.B1(n_194),
.B2(n_24),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_318),
.B(n_219),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_246),
.A2(n_138),
.B1(n_158),
.B2(n_210),
.Y(n_319)
);

AOI22xp33_ASAP7_75t_L g323 ( 
.A1(n_223),
.A2(n_195),
.B1(n_196),
.B2(n_198),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_323),
.A2(n_330),
.B1(n_336),
.B2(n_337),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_238),
.A2(n_138),
.B1(n_167),
.B2(n_189),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_229),
.A2(n_167),
.B1(n_196),
.B2(n_189),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_229),
.A2(n_198),
.B1(n_24),
.B2(n_11),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_L g337 ( 
.A1(n_215),
.A2(n_24),
.B1(n_2),
.B2(n_3),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_260),
.B(n_1),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g368 ( 
.A(n_342),
.Y(n_368)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_343),
.Y(n_346)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_346),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_298),
.B(n_264),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_347),
.B(n_357),
.C(n_302),
.Y(n_419)
);

OAI32xp33_ASAP7_75t_L g348 ( 
.A1(n_301),
.A2(n_317),
.A3(n_311),
.B1(n_291),
.B2(n_322),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_348),
.B(n_359),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_299),
.A2(n_248),
.B1(n_251),
.B2(n_276),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_349),
.A2(n_371),
.B1(n_303),
.B2(n_328),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g350 ( 
.A1(n_314),
.A2(n_236),
.B1(n_259),
.B2(n_253),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g422 ( 
.A1(n_350),
.A2(n_312),
.B1(n_331),
.B2(n_295),
.Y(n_422)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_289),
.Y(n_352)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_299),
.A2(n_276),
.B1(n_280),
.B2(n_279),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_354),
.A2(n_360),
.B(n_369),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_387),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_292),
.B(n_254),
.C(n_242),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_289),
.Y(n_358)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_358),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_300),
.B(n_213),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_305),
.B(n_235),
.Y(n_361)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_361),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g364 ( 
.A(n_344),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_364),
.B(n_365),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g365 ( 
.A(n_339),
.Y(n_365)
);

INVx4_ASAP7_75t_L g366 ( 
.A(n_343),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_366),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_332),
.A2(n_232),
.B1(n_217),
.B2(n_281),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_367),
.A2(n_376),
.B1(n_383),
.B2(n_297),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_291),
.A2(n_224),
.B1(n_225),
.B2(n_228),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g423 ( 
.A(n_370),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_330),
.A2(n_237),
.B1(n_250),
.B2(n_272),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_294),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_372),
.B(n_381),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_341),
.B(n_244),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_373),
.B(n_375),
.Y(n_402)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_374),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_326),
.B(n_332),
.Y(n_375)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_327),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_377),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_332),
.B(n_282),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_378),
.B(n_379),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_338),
.B(n_227),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_291),
.B(n_220),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_380),
.B(n_385),
.Y(n_401)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_294),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_329),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_382),
.B(n_388),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_319),
.A2(n_256),
.B1(n_257),
.B2(n_243),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_325),
.A2(n_318),
.B1(n_293),
.B2(n_343),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_384),
.A2(n_389),
.B(n_320),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_316),
.B(n_233),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_336),
.A2(n_11),
.B(n_15),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g404 ( 
.A1(n_386),
.A2(n_320),
.B(n_290),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_329),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_328),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_304),
.A2(n_5),
.B1(n_14),
.B2(n_15),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g390 ( 
.A(n_344),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_390),
.Y(n_424)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_344),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_391),
.B(n_315),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_362),
.A2(n_324),
.B1(n_290),
.B2(n_304),
.Y(n_392)
);

OAI21xp5_ASAP7_75t_L g458 ( 
.A1(n_392),
.A2(n_393),
.B(n_397),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g393 ( 
.A1(n_375),
.A2(n_310),
.B(n_309),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_378),
.A2(n_309),
.B(n_324),
.Y(n_397)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_400),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_355),
.B(n_306),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_403),
.B(n_429),
.C(n_308),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_404),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_406),
.B(n_413),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_SL g408 ( 
.A1(n_384),
.A2(n_345),
.B(n_312),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_408),
.A2(n_410),
.B(n_368),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_SL g409 ( 
.A(n_347),
.B(n_306),
.Y(n_409)
);

XNOR2x1_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_419),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g410 ( 
.A1(n_353),
.A2(n_334),
.B(n_327),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_387),
.B(n_359),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_373),
.B(n_340),
.Y(n_415)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_415),
.Y(n_433)
);

OAI22xp33_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_422),
.B1(n_426),
.B2(n_356),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_351),
.A2(n_340),
.B1(n_331),
.B2(n_295),
.Y(n_418)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_418),
.A2(n_371),
.B1(n_363),
.B2(n_352),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_353),
.B(n_357),
.Y(n_420)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_420),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_SL g426 ( 
.A1(n_362),
.A2(n_321),
.B1(n_345),
.B2(n_315),
.Y(n_426)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_351),
.A2(n_363),
.B1(n_367),
.B2(n_354),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_428),
.A2(n_383),
.B1(n_369),
.B2(n_386),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_380),
.B(n_287),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_430),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_434),
.A2(n_441),
.B(n_404),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_SL g435 ( 
.A(n_395),
.B(n_349),
.C(n_348),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g489 ( 
.A(n_435),
.B(n_437),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_398),
.B(n_395),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_425),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_438),
.B(n_439),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g439 ( 
.A(n_425),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_408),
.A2(n_368),
.B(n_379),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_442),
.B(n_445),
.Y(n_474)
);

OAI32xp33_ASAP7_75t_L g443 ( 
.A1(n_402),
.A2(n_358),
.A3(n_356),
.B1(n_382),
.B2(n_346),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_443),
.B(n_451),
.Y(n_475)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_444),
.A2(n_460),
.B1(n_461),
.B2(n_401),
.Y(n_469)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_399),
.Y(n_446)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_446),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_428),
.A2(n_381),
.B1(n_372),
.B2(n_364),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_447),
.A2(n_392),
.B1(n_421),
.B2(n_396),
.Y(n_480)
);

MAJx2_ASAP7_75t_L g449 ( 
.A(n_416),
.B(n_388),
.C(n_391),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g481 ( 
.A(n_449),
.B(n_450),
.Y(n_481)
);

MAJx2_ASAP7_75t_L g450 ( 
.A(n_416),
.B(n_403),
.C(n_409),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g451 ( 
.A(n_407),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_399),
.Y(n_452)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_452),
.Y(n_492)
);

OAI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_411),
.A2(n_389),
.B1(n_370),
.B2(n_366),
.Y(n_453)
);

AOI22xp5_ASAP7_75t_SL g488 ( 
.A1(n_453),
.A2(n_444),
.B1(n_463),
.B2(n_451),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_454),
.B(n_403),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_407),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_455),
.B(n_462),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_420),
.B(n_302),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_424),
.Y(n_470)
);

OAI22xp5_ASAP7_75t_L g457 ( 
.A1(n_411),
.A2(n_417),
.B1(n_402),
.B2(n_415),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_457),
.A2(n_463),
.B1(n_424),
.B2(n_412),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_413),
.A2(n_374),
.B1(n_377),
.B2(n_370),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_393),
.A2(n_397),
.B1(n_410),
.B2(n_394),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_430),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_400),
.A2(n_321),
.B1(n_308),
.B2(n_296),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_427),
.Y(n_464)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_464),
.Y(n_494)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_427),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_465),
.B(n_307),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_466),
.B(n_476),
.C(n_468),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_SL g506 ( 
.A1(n_467),
.A2(n_471),
.B(n_488),
.Y(n_506)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_440),
.B(n_409),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g505 ( 
.A(n_468),
.B(n_487),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_469),
.A2(n_478),
.B1(n_479),
.B2(n_482),
.Y(n_515)
);

CKINVDCx14_ASAP7_75t_R g503 ( 
.A(n_470),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g471 ( 
.A1(n_434),
.A2(n_394),
.B(n_406),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_460),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_472),
.B(n_483),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_440),
.B(n_419),
.C(n_429),
.Y(n_476)
);

AOI21xp33_ASAP7_75t_L g477 ( 
.A1(n_459),
.A2(n_401),
.B(n_421),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_477),
.B(n_432),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g478 ( 
.A1(n_431),
.A2(n_418),
.B1(n_412),
.B2(n_396),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_480),
.A2(n_484),
.B1(n_490),
.B2(n_448),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g482 ( 
.A1(n_431),
.A2(n_419),
.B1(n_421),
.B2(n_405),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_438),
.B(n_421),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_447),
.A2(n_426),
.B1(n_422),
.B2(n_405),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_457),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_485),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g487 ( 
.A(n_450),
.B(n_414),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_433),
.A2(n_423),
.B1(n_405),
.B2(n_414),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_461),
.A2(n_423),
.B1(n_296),
.B2(n_307),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_491),
.A2(n_442),
.B1(n_439),
.B2(n_465),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g493 ( 
.A1(n_458),
.A2(n_287),
.B(n_335),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_493),
.A2(n_465),
.B(n_452),
.Y(n_523)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_496),
.Y(n_501)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_454),
.B(n_335),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_497),
.B(n_446),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_521),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_436),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_499),
.B(n_494),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_500),
.A2(n_509),
.B1(n_480),
.B2(n_483),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_436),
.Y(n_502)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_502),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_466),
.B(n_449),
.C(n_435),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_504),
.B(n_513),
.C(n_514),
.Y(n_535)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_507),
.A2(n_474),
.B1(n_482),
.B2(n_472),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_SL g509 ( 
.A1(n_469),
.A2(n_485),
.B1(n_488),
.B2(n_475),
.Y(n_509)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_473),
.Y(n_511)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_511),
.Y(n_542)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_473),
.Y(n_512)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_512),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_459),
.C(n_433),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_497),
.B(n_455),
.C(n_458),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_474),
.A2(n_448),
.B1(n_462),
.B2(n_432),
.Y(n_516)
);

OAI22xp5_ASAP7_75t_L g530 ( 
.A1(n_516),
.A2(n_517),
.B1(n_519),
.B2(n_520),
.Y(n_530)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_486),
.Y(n_518)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_518),
.Y(n_533)
);

AOI21xp5_ASAP7_75t_L g519 ( 
.A1(n_475),
.A2(n_441),
.B(n_443),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_495),
.Y(n_520)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_520),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_487),
.B(n_464),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_495),
.Y(n_522)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_522),
.Y(n_550)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_523),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_524),
.B(n_493),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_481),
.B(n_2),
.C(n_3),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_525),
.B(n_526),
.C(n_494),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_481),
.B(n_4),
.C(n_5),
.Y(n_526)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_527),
.A2(n_531),
.B1(n_515),
.B2(n_509),
.Y(n_556)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_528),
.Y(n_563)
);

OR2x2_ASAP7_75t_L g553 ( 
.A(n_530),
.B(n_544),
.Y(n_553)
);

OAI22xp5_ASAP7_75t_SL g531 ( 
.A1(n_507),
.A2(n_474),
.B1(n_478),
.B2(n_491),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g568 ( 
.A(n_536),
.B(n_539),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g537 ( 
.A(n_503),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_537),
.B(n_543),
.Y(n_559)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_518),
.Y(n_538)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_538),
.Y(n_552)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_505),
.B(n_467),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_SL g540 ( 
.A(n_505),
.B(n_471),
.Y(n_540)
);

XNOR2xp5_ASAP7_75t_SL g551 ( 
.A(n_540),
.B(n_541),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_498),
.B(n_479),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_522),
.B(n_490),
.Y(n_547)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_547),
.Y(n_555)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_513),
.B(n_486),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_548),
.B(n_549),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_514),
.B(n_492),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_541),
.B(n_532),
.C(n_548),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_554),
.B(n_566),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g576 ( 
.A1(n_556),
.A2(n_550),
.B1(n_546),
.B2(n_545),
.Y(n_576)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_533),
.Y(n_557)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_557),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_529),
.B(n_519),
.Y(n_558)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_558),
.B(n_564),
.Y(n_577)
);

OA21x2_ASAP7_75t_L g560 ( 
.A1(n_528),
.A2(n_511),
.B(n_512),
.Y(n_560)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_560),
.Y(n_583)
);

XNOR2xp5_ASAP7_75t_SL g561 ( 
.A(n_540),
.B(n_504),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_506),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_SL g562 ( 
.A1(n_527),
.A2(n_510),
.B1(n_508),
.B2(n_484),
.Y(n_562)
);

OR2x2_ASAP7_75t_L g575 ( 
.A(n_562),
.B(n_565),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_532),
.B(n_510),
.Y(n_564)
);

AO21x1_ASAP7_75t_L g565 ( 
.A1(n_534),
.A2(n_516),
.B(n_508),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_535),
.B(n_524),
.C(n_521),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_535),
.B(n_539),
.C(n_536),
.Y(n_567)
);

HB1xp67_ASAP7_75t_L g572 ( 
.A(n_567),
.Y(n_572)
);

OAI21x1_ASAP7_75t_L g569 ( 
.A1(n_542),
.A2(n_523),
.B(n_501),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_569),
.B(n_565),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_570),
.B(n_538),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_571),
.B(n_578),
.Y(n_592)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_574),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_576),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_559),
.B(n_533),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_568),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_SL g580 ( 
.A1(n_555),
.A2(n_534),
.B(n_547),
.Y(n_580)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_580),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g582 ( 
.A(n_553),
.B(n_500),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_584),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_SL g584 ( 
.A(n_566),
.B(n_543),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g585 ( 
.A1(n_563),
.A2(n_553),
.B1(n_560),
.B2(n_556),
.Y(n_585)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_585),
.A2(n_501),
.B1(n_560),
.B2(n_531),
.Y(n_589)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_586),
.Y(n_597)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_577),
.Y(n_587)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_587),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_574),
.B(n_562),
.Y(n_588)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_588),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g603 ( 
.A(n_589),
.B(n_598),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_572),
.B(n_554),
.C(n_567),
.Y(n_593)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_593),
.B(n_551),
.C(n_580),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_SL g596 ( 
.A(n_581),
.B(n_568),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_SL g601 ( 
.A(n_596),
.B(n_599),
.Y(n_601)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_576),
.Y(n_599)
);

NOR2xp67_ASAP7_75t_L g600 ( 
.A(n_594),
.B(n_561),
.Y(n_600)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_600),
.A2(n_604),
.B(n_605),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_602),
.B(n_607),
.Y(n_612)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_587),
.A2(n_575),
.B(n_579),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g605 ( 
.A1(n_590),
.A2(n_575),
.B(n_583),
.Y(n_605)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_593),
.B(n_586),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_SL g608 ( 
.A1(n_595),
.A2(n_585),
.B(n_583),
.Y(n_608)
);

AOI21xp5_ASAP7_75t_SL g615 ( 
.A1(n_608),
.A2(n_588),
.B(n_597),
.Y(n_615)
);

AND2x2_ASAP7_75t_L g610 ( 
.A(n_606),
.B(n_592),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_610),
.A2(n_611),
.B(n_605),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_601),
.B(n_591),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g613 ( 
.A(n_602),
.B(n_588),
.C(n_598),
.Y(n_613)
);

XNOR2xp5_ASAP7_75t_L g619 ( 
.A(n_613),
.B(n_603),
.Y(n_619)
);

OAI21xp5_ASAP7_75t_L g618 ( 
.A1(n_615),
.A2(n_609),
.B(n_573),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g616 ( 
.A(n_612),
.Y(n_616)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_616),
.Y(n_621)
);

AOI21x1_ASAP7_75t_L g620 ( 
.A1(n_617),
.A2(n_618),
.B(n_619),
.Y(n_620)
);

MAJIxp5_ASAP7_75t_L g622 ( 
.A(n_621),
.B(n_614),
.C(n_603),
.Y(n_622)
);

AOI321xp33_ASAP7_75t_SL g623 ( 
.A1(n_622),
.A2(n_620),
.A3(n_589),
.B1(n_551),
.B2(n_573),
.C(n_506),
.Y(n_623)
);

AOI21xp5_ASAP7_75t_SL g624 ( 
.A1(n_623),
.A2(n_526),
.B(n_525),
.Y(n_624)
);

AOI311xp33_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_492),
.A3(n_496),
.B(n_5),
.C(n_16),
.Y(n_625)
);


endmodule