module fake_jpeg_28116_n_136 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx4f_ASAP7_75t_SL g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_17),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_29),
.Y(n_35)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_17),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_21),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_29),
.B(n_12),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_33),
.B(n_41),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_26),
.A2(n_21),
.B1(n_11),
.B2(n_20),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_20),
.B1(n_11),
.B2(n_31),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_30),
.B(n_23),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_23),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_42),
.B(n_15),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_35),
.B(n_19),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_46),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_38),
.A2(n_26),
.B1(n_32),
.B2(n_24),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_50),
.Y(n_58)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_32),
.B1(n_24),
.B2(n_25),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_22),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_37),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_34),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_52),
.A2(n_56),
.B1(n_43),
.B2(n_34),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_42),
.C(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_30),
.B1(n_11),
.B2(n_20),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_35),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_57),
.B(n_59),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_51),
.A2(n_27),
.B1(n_31),
.B2(n_44),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_60),
.A2(n_63),
.B1(n_67),
.B2(n_56),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_68),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_33),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_65),
.B(n_45),
.Y(n_71)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_SL g69 ( 
.A(n_65),
.B(n_55),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_73),
.C(n_66),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_75),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_72),
.A2(n_79),
.B(n_71),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_40),
.C(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_58),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_77),
.B(n_78),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_61),
.B(n_48),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_68),
.A2(n_19),
.B1(n_14),
.B2(n_53),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_80),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_81),
.B(n_83),
.Y(n_99)
);

A2O1A1O1Ixp25_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_67),
.B(n_66),
.C(n_28),
.D(n_13),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_82),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_49),
.B1(n_36),
.B2(n_39),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_85),
.A2(n_74),
.B1(n_48),
.B2(n_39),
.Y(n_93)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

MAJx2_ASAP7_75t_L g92 ( 
.A(n_73),
.B(n_13),
.C(n_43),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_22),
.C(n_18),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_93),
.A2(n_94),
.B1(n_96),
.B2(n_88),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_83),
.A2(n_34),
.B1(n_27),
.B2(n_62),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_84),
.A2(n_62),
.B1(n_22),
.B2(n_18),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_93),
.C(n_95),
.Y(n_110)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_91),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_102),
.B(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

FAx1_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_89),
.CI(n_82),
.CON(n_104),
.SN(n_104)
);

AOI31xp67_ASAP7_75t_L g113 ( 
.A1(n_104),
.A2(n_111),
.A3(n_94),
.B(n_112),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_100),
.A2(n_86),
.B1(n_92),
.B2(n_87),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_105),
.B(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_88),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_107),
.B(n_108),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_97),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_109),
.A2(n_0),
.B(n_1),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_96),
.C(n_22),
.Y(n_114)
);

NOR3xp33_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_90),
.C(n_10),
.Y(n_111)
);

OAI31xp33_ASAP7_75t_L g125 ( 
.A1(n_113),
.A2(n_5),
.A3(n_7),
.B(n_8),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_114),
.B(n_2),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_115),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_18),
.C(n_10),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_118),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_0),
.C(n_2),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_119),
.A2(n_108),
.B(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_124),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_116),
.C(n_7),
.Y(n_128)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_123),
.B(n_125),
.Y(n_126)
);

OA21x2_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_3),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_128),
.B(n_129),
.Y(n_132)
);

NOR2xp67_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_9),
.Y(n_129)
);

NOR2xp67_ASAP7_75t_SL g130 ( 
.A(n_127),
.B(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_130),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_126),
.A2(n_121),
.B(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_9),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_134),
.B(n_132),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule