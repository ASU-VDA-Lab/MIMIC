module fake_jpeg_28787_n_412 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_412);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_412;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_19),
.Y(n_22)
);

BUFx6f_ASAP7_75t_SL g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_19),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx11_ASAP7_75t_SL g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_21),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_51),
.B(n_54),
.Y(n_92)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_52),
.Y(n_134)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx11_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_55),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_57),
.Y(n_112)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

CKINVDCx6p67_ASAP7_75t_R g131 ( 
.A(n_59),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_31),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_61),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_62),
.Y(n_129)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_63),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_31),
.Y(n_64)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_64),
.Y(n_115)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g98 ( 
.A(n_65),
.Y(n_98)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_31),
.Y(n_67)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_67),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_28),
.B(n_0),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_85),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_69),
.Y(n_104)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_36),
.Y(n_72)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_72),
.Y(n_95)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_74),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

INVx11_ASAP7_75t_L g76 ( 
.A(n_23),
.Y(n_76)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_76),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_34),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g123 ( 
.A(n_77),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_34),
.Y(n_78)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_38),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_82),
.Y(n_102)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_47),
.Y(n_80)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_81),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_22),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_83),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_84),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_28),
.B(n_0),
.Y(n_85)
);

BUFx4f_ASAP7_75t_L g86 ( 
.A(n_40),
.Y(n_86)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_42),
.Y(n_87)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_88),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_59),
.B(n_43),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g151 ( 
.A(n_99),
.B(n_106),
.Y(n_151)
);

HAxp5_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_29),
.CON(n_105),
.SN(n_105)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_117),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_88),
.A2(n_24),
.B1(n_78),
.B2(n_77),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_108),
.A2(n_113),
.B1(n_120),
.B2(n_57),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_65),
.B(n_43),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_29),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_84),
.A2(n_50),
.B1(n_40),
.B2(n_37),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g117 ( 
.A1(n_74),
.A2(n_42),
.B1(n_47),
.B2(n_52),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_55),
.A2(n_24),
.B1(n_37),
.B2(n_26),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_56),
.B(n_48),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_45),
.Y(n_156)
);

NAND2xp33_ASAP7_75t_SL g126 ( 
.A(n_58),
.B(n_42),
.Y(n_126)
);

NAND2xp33_ASAP7_75t_SL g143 ( 
.A(n_126),
.B(n_83),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_63),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_96),
.B(n_48),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_136),
.B(n_147),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_137),
.A2(n_139),
.B1(n_154),
.B2(n_93),
.Y(n_181)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g186 ( 
.A(n_138),
.Y(n_186)
);

OAI22xp33_ASAP7_75t_L g139 ( 
.A1(n_107),
.A2(n_60),
.B1(n_69),
.B2(n_67),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_132),
.Y(n_140)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_90),
.Y(n_142)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_142),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_163),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_146),
.B(n_148),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_27),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_92),
.B(n_32),
.Y(n_148)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_32),
.B(n_49),
.C(n_45),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_149),
.B(n_156),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_150),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_89),
.B(n_49),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_152),
.B(n_165),
.Y(n_183)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_131),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_153),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_117),
.A2(n_62),
.B1(n_61),
.B2(n_64),
.Y(n_154)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_90),
.Y(n_155)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

CKINVDCx12_ASAP7_75t_R g157 ( 
.A(n_119),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_157),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx8_ASAP7_75t_L g192 ( 
.A(n_158),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g159 ( 
.A(n_98),
.Y(n_159)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_159),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_102),
.B(n_33),
.Y(n_160)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_100),
.Y(n_161)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_161),
.Y(n_177)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_95),
.Y(n_164)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_164),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_98),
.B(n_33),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g166 ( 
.A(n_119),
.Y(n_166)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_166),
.Y(n_193)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_125),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_128),
.Y(n_179)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_118),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_179),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_181),
.A2(n_187),
.B1(n_123),
.B2(n_115),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_152),
.B(n_117),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_184),
.B(n_139),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_162),
.A2(n_115),
.B1(n_107),
.B2(n_113),
.Y(n_187)
);

AO22x1_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_93),
.B1(n_129),
.B2(n_112),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_191),
.B(n_128),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_184),
.A2(n_181),
.B1(n_162),
.B2(n_191),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_195),
.A2(n_213),
.B1(n_207),
.B2(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_175),
.B(n_151),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_197),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_136),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_188),
.B(n_147),
.C(n_164),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_140),
.C(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_199),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_200),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_183),
.B(n_145),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_202),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_138),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_203),
.B(n_169),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_163),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_204),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_205),
.A2(n_208),
.B1(n_213),
.B2(n_186),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_211),
.Y(n_219)
);

OAI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_191),
.A2(n_149),
.B1(n_123),
.B2(n_168),
.Y(n_208)
);

INVx8_ASAP7_75t_L g209 ( 
.A(n_192),
.Y(n_209)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_209),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g210 ( 
.A(n_193),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_185),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_172),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

AND2x6_ASAP7_75t_L g214 ( 
.A(n_173),
.B(n_166),
.Y(n_214)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_214),
.A2(n_171),
.B(n_194),
.C(n_166),
.D(n_98),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_216),
.A2(n_217),
.B1(n_223),
.B2(n_199),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_173),
.B1(n_190),
.B2(n_141),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_210),
.Y(n_218)
);

OR2x2_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_222),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_203),
.A2(n_206),
.B(n_214),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_229),
.B(n_198),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_210),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_195),
.A2(n_97),
.B1(n_112),
.B2(n_114),
.Y(n_223)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_228),
.B(n_182),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_208),
.A2(n_194),
.B(n_185),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_212),
.B1(n_186),
.B2(n_200),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_203),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_159),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_SL g252 ( 
.A(n_235),
.B(n_177),
.Y(n_252)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_236),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_214),
.A3(n_204),
.B1(n_205),
.B2(n_201),
.Y(n_237)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_237),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_238),
.A2(n_239),
.B(n_218),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_221),
.A2(n_211),
.B(n_198),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_196),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_215),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_241),
.A2(n_176),
.B1(n_158),
.B2(n_104),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_242),
.A2(n_233),
.B1(n_223),
.B2(n_220),
.Y(n_263)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_232),
.A2(n_209),
.B1(n_193),
.B2(n_166),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_182),
.B1(n_118),
.B2(n_170),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_235),
.B(n_197),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_252),
.C(n_230),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_225),
.B(n_174),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_246),
.B(n_254),
.Y(n_262)
);

NOR2x1_ASAP7_75t_L g248 ( 
.A(n_228),
.B(n_144),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_251),
.Y(n_264)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_225),
.B(n_35),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_250),
.B(n_1),
.Y(n_279)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_231),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_255),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_35),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_226),
.B(n_177),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_258),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_228),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_219),
.B(n_170),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_219),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_260),
.B(n_261),
.Y(n_298)
);

A2O1A1O1Ixp25_ASAP7_75t_L g261 ( 
.A1(n_247),
.A2(n_217),
.B(n_224),
.C(n_216),
.D(n_229),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_266),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_242),
.A2(n_230),
.B1(n_220),
.B2(n_222),
.Y(n_266)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_268),
.B(n_269),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_247),
.A2(n_215),
.B1(n_209),
.B2(n_192),
.Y(n_271)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_272),
.B(n_20),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_274),
.A2(n_275),
.B1(n_189),
.B2(n_257),
.Y(n_284)
);

OA22x2_ASAP7_75t_L g276 ( 
.A1(n_236),
.A2(n_161),
.B1(n_104),
.B2(n_155),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_276),
.B(n_116),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_243),
.B(n_167),
.Y(n_277)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_277),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_243),
.B(n_176),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_280),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g281 ( 
.A1(n_238),
.A2(n_189),
.B(n_153),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_281),
.A2(n_248),
.B(n_249),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_239),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_283),
.B(n_292),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g314 ( 
.A1(n_284),
.A2(n_274),
.B1(n_276),
.B2(n_278),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_269),
.A2(n_236),
.B(n_241),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_285),
.A2(n_287),
.B(n_273),
.Y(n_316)
);

INVx3_ASAP7_75t_L g286 ( 
.A(n_270),
.Y(n_286)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_286),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_281),
.A2(n_250),
.B(n_253),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_288),
.B(n_290),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g290 ( 
.A(n_270),
.Y(n_290)
);

HB1xp67_ASAP7_75t_L g291 ( 
.A(n_280),
.Y(n_291)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_291),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_260),
.B(n_245),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_237),
.B1(n_240),
.B2(n_255),
.Y(n_293)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_259),
.A2(n_127),
.B(n_134),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_294),
.B(n_299),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_267),
.B(n_264),
.C(n_259),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_297),
.B(n_301),
.C(n_306),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_264),
.B(n_142),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_266),
.B(n_94),
.C(n_135),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_277),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_303),
.B(n_278),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_304),
.Y(n_319)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_271),
.B(n_129),
.C(n_97),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_261),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_309),
.B(n_315),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_307),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_311),
.B(n_3),
.Y(n_341)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_286),
.A2(n_296),
.B1(n_302),
.B2(n_295),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_313),
.B(n_317),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_314),
.A2(n_300),
.B1(n_306),
.B2(n_294),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_282),
.Y(n_315)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_316),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_282),
.B(n_276),
.C(n_265),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_322),
.B(n_330),
.C(n_121),
.Y(n_340)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_298),
.B(n_263),
.CI(n_276),
.CON(n_323),
.SN(n_323)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_323),
.B(n_329),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_265),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_325),
.B(n_326),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_299),
.B(n_262),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_301),
.B(n_279),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_288),
.B(n_127),
.Y(n_330)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_289),
.B(n_304),
.Y(n_331)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_333),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_336),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_323),
.B(n_24),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_327),
.A2(n_24),
.B1(n_37),
.B2(n_26),
.Y(n_336)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_SL g339 ( 
.A1(n_308),
.A2(n_121),
.B1(n_114),
.B2(n_101),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_339),
.B(n_341),
.Y(n_356)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_340),
.B(n_324),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_319),
.A2(n_322),
.B1(n_311),
.B2(n_328),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_345),
.Y(n_362)
);

BUFx12_ASAP7_75t_L g345 ( 
.A(n_330),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_47),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_348),
.Y(n_358)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_324),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g375 ( 
.A(n_349),
.B(n_50),
.Y(n_375)
);

NOR2xp67_ASAP7_75t_R g350 ( 
.A(n_335),
.B(n_326),
.Y(n_350)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_350),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_343),
.B(n_310),
.C(n_320),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_353),
.B(n_357),
.Y(n_374)
);

NOR2x1p5_ASAP7_75t_L g355 ( 
.A(n_331),
.B(n_309),
.Y(n_355)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_334),
.A2(n_337),
.B1(n_340),
.B2(n_310),
.Y(n_357)
);

BUFx24_ASAP7_75t_SL g359 ( 
.A(n_346),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_SL g365 ( 
.A(n_359),
.B(n_339),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_346),
.B(n_342),
.C(n_320),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_360),
.B(n_20),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g361 ( 
.A1(n_347),
.A2(n_325),
.B1(n_315),
.B2(n_26),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_361),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_362),
.B(n_342),
.C(n_333),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_364),
.B(n_369),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_370),
.Y(n_384)
);

NOR2xp67_ASAP7_75t_L g367 ( 
.A(n_355),
.B(n_345),
.Y(n_367)
);

NOR3xp33_ASAP7_75t_L g385 ( 
.A(n_367),
.B(n_373),
.C(n_364),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_345),
.Y(n_368)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_368),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_50),
.C(n_40),
.Y(n_369)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_358),
.B(n_3),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_371),
.B(n_4),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_351),
.B(n_4),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_372),
.B(n_375),
.C(n_356),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_376),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_378),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_366),
.A2(n_354),
.B1(n_352),
.B2(n_50),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_368),
.B(n_5),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g390 ( 
.A1(n_379),
.A2(n_386),
.B(n_41),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_374),
.B(n_53),
.C(n_8),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_7),
.C(n_8),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_383),
.B(n_12),
.C(n_13),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_385),
.A2(n_41),
.B1(n_15),
.B2(n_16),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_369),
.A2(n_59),
.B(n_41),
.Y(n_386)
);

AND2x4_ASAP7_75t_L g387 ( 
.A(n_375),
.B(n_7),
.Y(n_387)
);

OAI221xp5_ASAP7_75t_L g388 ( 
.A1(n_387),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_388),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_390),
.B(n_391),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_381),
.B(n_10),
.Y(n_391)
);

INVx6_ASAP7_75t_L g400 ( 
.A(n_393),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_379),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_394),
.A2(n_384),
.B(n_387),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_376),
.B(n_395),
.Y(n_397)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_397),
.Y(n_403)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_392),
.B(n_380),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_399),
.B(n_13),
.Y(n_405)
);

AOI322xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_13),
.A3(n_15),
.B1(n_16),
.B2(n_17),
.C1(n_18),
.C2(n_63),
.Y(n_406)
);

NOR3xp33_ASAP7_75t_L g404 ( 
.A(n_398),
.B(n_394),
.C(n_389),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_404),
.A2(n_405),
.B(n_406),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g408 ( 
.A1(n_403),
.A2(n_401),
.B(n_400),
.Y(n_408)
);

AOI322xp5_ASAP7_75t_L g409 ( 
.A1(n_408),
.A2(n_16),
.A3(n_17),
.B1(n_18),
.B2(n_39),
.C1(n_76),
.C2(n_407),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_409),
.Y(n_410)
);

AOI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_410),
.A2(n_17),
.B(n_39),
.Y(n_411)
);

O2A1O1Ixp33_ASAP7_75t_SL g412 ( 
.A1(n_411),
.A2(n_39),
.B(n_341),
.C(n_280),
.Y(n_412)
);


endmodule