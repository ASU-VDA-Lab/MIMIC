module fake_jpeg_27412_n_224 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_224);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_224;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVxp33_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_13),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_SL g31 ( 
.A(n_12),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_28),
.Y(n_34)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_29),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_0),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_36),
.B(n_39),
.Y(n_45)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_16),
.B(n_1),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_40),
.B(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

OR2x2_ASAP7_75t_L g44 ( 
.A(n_40),
.B(n_16),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_44),
.B(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_46),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_37),
.A2(n_30),
.B1(n_19),
.B2(n_20),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_49),
.A2(n_30),
.B1(n_31),
.B2(n_17),
.Y(n_62)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_38),
.A2(n_30),
.B1(n_19),
.B2(n_20),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_L g70 ( 
.A1(n_53),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_27),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_58),
.Y(n_86)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_39),
.B(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_60),
.B(n_27),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_70),
.B1(n_52),
.B2(n_22),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_60),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_63),
.B(n_66),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g64 ( 
.A1(n_55),
.A2(n_39),
.B1(n_43),
.B2(n_42),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_64),
.A2(n_71),
.B1(n_47),
.B2(n_51),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_69),
.Y(n_87)
);

NAND3xp33_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_22),
.C(n_32),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_55),
.A2(n_17),
.B1(n_22),
.B2(n_26),
.Y(n_71)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_82),
.Y(n_101)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_77),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_44),
.B(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_48),
.Y(n_79)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_52),
.A2(n_22),
.B1(n_26),
.B2(n_25),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_81),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_54),
.B(n_21),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_56),
.C(n_25),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_48),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_84),
.B(n_33),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_66),
.B(n_44),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_89),
.B(n_90),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_71),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_34),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_97),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_56),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_93),
.B(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_18),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_64),
.B(n_34),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_64),
.B(n_41),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_102),
.A2(n_62),
.B1(n_47),
.B2(n_77),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_58),
.B(n_26),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g112 ( 
.A1(n_103),
.A2(n_84),
.B(n_65),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_43),
.C(n_42),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_104),
.B(n_95),
.Y(n_129)
);

AOI32xp33_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_33),
.A3(n_50),
.B1(n_47),
.B2(n_29),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_91),
.B1(n_102),
.B2(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

FAx1_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_33),
.CI(n_25),
.CON(n_107),
.SN(n_107)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_108),
.Y(n_118)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_112),
.A2(n_123),
.B(n_92),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_117),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_116),
.A2(n_120),
.B1(n_124),
.B2(n_128),
.Y(n_139)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_103),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_121),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_111),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_75),
.B(n_79),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_90),
.A2(n_61),
.B1(n_74),
.B2(n_73),
.Y(n_124)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_110),
.Y(n_125)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_93),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_126),
.B(n_130),
.Y(n_147)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_104),
.Y(n_127)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_100),
.A2(n_92),
.B1(n_97),
.B2(n_89),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_129),
.B(n_87),
.Y(n_145)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_107),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_100),
.A2(n_61),
.B1(n_74),
.B2(n_73),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_132),
.A2(n_98),
.B1(n_108),
.B2(n_96),
.Y(n_142)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_133),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g134 ( 
.A(n_98),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_134),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_SL g136 ( 
.A(n_117),
.B(n_107),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_138),
.B(n_146),
.Y(n_168)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_124),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_143),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_142),
.A2(n_127),
.B1(n_134),
.B2(n_119),
.Y(n_158)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_145),
.B(n_153),
.C(n_113),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g146 ( 
.A1(n_118),
.A2(n_88),
.B(n_18),
.Y(n_146)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_112),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_149),
.B(n_152),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_125),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_150),
.Y(n_171)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_120),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_99),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

NOR3xp33_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_29),
.C(n_50),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_131),
.A2(n_18),
.B(n_99),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_155),
.A2(n_109),
.B(n_29),
.Y(n_165)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_113),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_4),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_158),
.A2(n_162),
.B1(n_170),
.B2(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_151),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_159),
.B(n_172),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_161),
.B(n_174),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_139),
.A2(n_128),
.B1(n_115),
.B2(n_116),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_153),
.B(n_131),
.C(n_123),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_166),
.C(n_140),
.Y(n_176)
);

OA21x2_ASAP7_75t_L g164 ( 
.A1(n_149),
.A2(n_122),
.B(n_109),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_167),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_173),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_140),
.B(n_96),
.C(n_85),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_136),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_169),
.A2(n_170),
.B1(n_174),
.B2(n_165),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_152),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_170)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_5),
.B(n_8),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_175),
.B(n_177),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_178),
.Y(n_192)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_160),
.Y(n_177)
);

AOI321xp33_ASAP7_75t_L g178 ( 
.A1(n_168),
.A2(n_145),
.A3(n_148),
.B1(n_156),
.B2(n_147),
.C(n_143),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_179),
.B(n_188),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_141),
.C(n_137),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_184),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_161),
.B(n_135),
.C(n_144),
.Y(n_184)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_187),
.A2(n_157),
.B1(n_166),
.B2(n_10),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_162),
.B(n_8),
.C(n_9),
.Y(n_188)
);

AOI321xp33_ASAP7_75t_L g189 ( 
.A1(n_186),
.A2(n_168),
.A3(n_164),
.B1(n_158),
.B2(n_157),
.C(n_171),
.Y(n_189)
);

NAND4xp25_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_10),
.C(n_11),
.D(n_12),
.Y(n_205)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_191),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_188),
.A2(n_171),
.B1(n_164),
.B2(n_173),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_193),
.A2(n_198),
.B(n_9),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_197),
.A2(n_186),
.B1(n_184),
.B2(n_11),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_8),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_194),
.A2(n_182),
.B1(n_180),
.B2(n_176),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_200),
.A2(n_193),
.B1(n_192),
.B2(n_196),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_201),
.B(n_202),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_9),
.C(n_10),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_203),
.B(n_204),
.Y(n_207)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_190),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_13),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_198),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_202),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_212),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_209),
.B(n_211),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_204),
.B(n_191),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_212),
.B(n_199),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_213),
.B(n_215),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_200),
.C(n_201),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_216),
.A2(n_210),
.B(n_207),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_217),
.B(n_219),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_214),
.A2(n_199),
.B(n_205),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_218),
.A2(n_203),
.B1(n_14),
.B2(n_15),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_221),
.B(n_13),
.C(n_14),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_222),
.B(n_220),
.C(n_15),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_15),
.Y(n_224)
);


endmodule