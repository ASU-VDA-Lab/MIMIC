module fake_jpeg_4846_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx2_ASAP7_75t_SL g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx16f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

INVx8_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx13_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

INVx4_ASAP7_75t_SL g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_43),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_7),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_25),
.B(n_0),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_45),
.B(n_61),
.Y(n_79)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_48),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_49),
.Y(n_91)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_53),
.A2(n_57),
.B1(n_64),
.B2(n_37),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_26),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_26),
.Y(n_56)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx9p33_ASAP7_75t_R g59 ( 
.A(n_29),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_60),
.Y(n_82)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

OR2x2_ASAP7_75t_SL g61 ( 
.A(n_18),
.B(n_16),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_62),
.B(n_32),
.Y(n_68)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_63),
.Y(n_72)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g65 ( 
.A1(n_58),
.A2(n_29),
.B1(n_32),
.B2(n_24),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_65),
.A2(n_32),
.B1(n_24),
.B2(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_85),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_68),
.B(n_90),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_20),
.Y(n_69)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_62),
.B(n_40),
.C(n_20),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_71),
.B(n_32),
.C(n_8),
.Y(n_119)
);

NOR2x1_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_21),
.Y(n_73)
);

NAND3xp33_ASAP7_75t_L g137 ( 
.A(n_73),
.B(n_7),
.C(n_13),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_78),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_64),
.A2(n_37),
.B1(n_22),
.B2(n_39),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_80),
.A2(n_83),
.B1(n_84),
.B2(n_101),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_37),
.B1(n_39),
.B2(n_28),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_60),
.A2(n_28),
.B1(n_30),
.B2(n_27),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_33),
.Y(n_86)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_86),
.Y(n_132)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_87),
.B(n_94),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_59),
.B(n_21),
.Y(n_90)
);

AOI211xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_33),
.B(n_27),
.C(n_30),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_92),
.A2(n_105),
.B1(n_108),
.B2(n_6),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_29),
.Y(n_93)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_93),
.Y(n_135)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_63),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_96),
.Y(n_129)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_43),
.B(n_25),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_97),
.B(n_6),
.Y(n_141)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_99),
.Y(n_133)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_51),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_53),
.B(n_29),
.Y(n_100)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_100),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_57),
.A2(n_28),
.B1(n_40),
.B2(n_38),
.Y(n_101)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_104),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_43),
.A2(n_38),
.B1(n_36),
.B2(n_23),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_45),
.B(n_36),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_45),
.B(n_31),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_107),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_56),
.A2(n_23),
.B1(n_31),
.B2(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_109),
.B(n_85),
.Y(n_114)
);

OAI21xp33_ASAP7_75t_L g110 ( 
.A1(n_73),
.A2(n_41),
.B(n_8),
.Y(n_110)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_110),
.A2(n_9),
.B(n_15),
.C(n_10),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_114),
.B(n_119),
.Y(n_157)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_115),
.B(n_118),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_117),
.A2(n_124),
.B1(n_90),
.B2(n_99),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_74),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_120),
.B(n_121),
.Y(n_164)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_79),
.B(n_0),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_131),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_79),
.B(n_24),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_70),
.C(n_96),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_79),
.B(n_68),
.Y(n_131)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_136),
.B(n_139),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g167 ( 
.A(n_137),
.B(n_141),
.Y(n_167)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_65),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_92),
.A2(n_7),
.B1(n_13),
.B2(n_11),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_140),
.A2(n_15),
.B1(n_11),
.B2(n_10),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_69),
.B(n_0),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_90),
.Y(n_150)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_65),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_143),
.B(n_144),
.Y(n_176)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_146),
.A2(n_4),
.B(n_5),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_129),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_148),
.B(n_152),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_149),
.A2(n_155),
.B1(n_156),
.B2(n_171),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_150),
.B(n_172),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g151 ( 
.A(n_144),
.Y(n_151)
);

BUFx2_ASAP7_75t_L g196 ( 
.A(n_151),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_112),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_139),
.A2(n_87),
.B1(n_76),
.B2(n_94),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_153),
.A2(n_174),
.B1(n_178),
.B2(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_71),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_154),
.B(n_158),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_136),
.A2(n_104),
.B1(n_81),
.B2(n_82),
.Y(n_155)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_117),
.A2(n_77),
.B1(n_66),
.B2(n_103),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_114),
.B(n_89),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_127),
.C(n_135),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_161),
.B(n_165),
.Y(n_189)
);

AOI32xp33_ASAP7_75t_L g163 ( 
.A1(n_134),
.A2(n_76),
.A3(n_98),
.B1(n_75),
.B2(n_88),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_163),
.B(n_178),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_131),
.B(n_89),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_170),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_168),
.B(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_126),
.B(n_95),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_75),
.B1(n_77),
.B2(n_88),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_143),
.A2(n_103),
.B1(n_91),
.B2(n_72),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_126),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_175),
.B(n_179),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_126),
.B(n_72),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_177),
.B(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_134),
.A2(n_91),
.B1(n_2),
.B2(n_3),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_116),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_125),
.B(n_0),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_142),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_179),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_182),
.A2(n_145),
.B(n_172),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g183 ( 
.A(n_166),
.B(n_154),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_183),
.A2(n_210),
.B(n_192),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_149),
.B1(n_169),
.B2(n_171),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_187),
.B1(n_188),
.B2(n_195),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_175),
.A2(n_130),
.B1(n_119),
.B2(n_138),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_156),
.A2(n_130),
.B1(n_138),
.B2(n_116),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_159),
.C(n_177),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_158),
.B(n_141),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_193),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_147),
.B(n_141),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_156),
.A2(n_135),
.B1(n_113),
.B2(n_132),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_147),
.B(n_132),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_197),
.B(n_206),
.Y(n_221)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_164),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_201),
.Y(n_217)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_176),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_176),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_202),
.B(n_211),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_181),
.B(n_115),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_203),
.B(n_201),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_156),
.A2(n_113),
.B1(n_121),
.B2(n_3),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_170),
.B(n_122),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_152),
.B(n_8),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_209),
.Y(n_231)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_208),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_180),
.B(n_122),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_162),
.Y(n_211)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_212),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_184),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_182),
.B1(n_156),
.B2(n_155),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_215),
.A2(n_230),
.B1(n_194),
.B2(n_186),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_218),
.B(n_191),
.C(n_187),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_163),
.B1(n_168),
.B2(n_148),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_219),
.B(n_227),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_185),
.A2(n_150),
.B(n_157),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_222),
.A2(n_226),
.B(n_232),
.Y(n_252)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_185),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_228),
.B(n_235),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_194),
.A2(n_157),
.B1(n_153),
.B2(n_174),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_184),
.A2(n_167),
.B(n_160),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_151),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g254 ( 
.A(n_233),
.Y(n_254)
);

NOR4xp25_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_167),
.C(n_151),
.D(n_160),
.Y(n_234)
);

NAND3xp33_ASAP7_75t_L g243 ( 
.A(n_234),
.B(n_198),
.C(n_188),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_214),
.B(n_199),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_193),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_214),
.B(n_203),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_238),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_190),
.B(n_197),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_183),
.B(n_190),
.Y(n_239)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_239),
.Y(n_242)
);

OA21x2_ASAP7_75t_SL g240 ( 
.A1(n_226),
.A2(n_183),
.B(n_198),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_240),
.B(n_251),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_241),
.A2(n_257),
.B1(n_229),
.B2(n_216),
.Y(n_270)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_243),
.B(n_232),
.CI(n_222),
.CON(n_261),
.SN(n_261)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_244),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_220),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g247 ( 
.A(n_217),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_247),
.A2(n_253),
.B1(n_259),
.B2(n_237),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_255),
.C(n_260),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_238),
.Y(n_250)
);

INVxp33_ASAP7_75t_SL g273 ( 
.A(n_250),
.Y(n_273)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_221),
.A2(n_202),
.B(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_221),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_195),
.C(n_200),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_196),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_256),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g257 ( 
.A1(n_239),
.A2(n_204),
.B(n_208),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_217),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_236),
.B(n_205),
.C(n_189),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_261),
.B(n_274),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_269),
.Y(n_286)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_263),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_258),
.B(n_218),
.C(n_220),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_266),
.B(n_272),
.C(n_248),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_260),
.A2(n_224),
.B1(n_230),
.B2(n_216),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_268),
.A2(n_246),
.B1(n_231),
.B2(n_259),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_219),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_270),
.A2(n_226),
.B1(n_257),
.B2(n_242),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_245),
.B(n_215),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g274 ( 
.A(n_241),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_257),
.A2(n_229),
.B1(n_234),
.B2(n_226),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_257),
.Y(n_277)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_277),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_274),
.A2(n_242),
.B1(n_252),
.B2(n_240),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_279),
.A2(n_288),
.B1(n_267),
.B2(n_261),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_255),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_285),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_273),
.A2(n_253),
.B1(n_250),
.B2(n_254),
.Y(n_282)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_282),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_252),
.B(n_249),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_284),
.B(n_262),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_265),
.A2(n_244),
.B(n_249),
.Y(n_287)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_287),
.A2(n_228),
.B1(n_267),
.B2(n_235),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_288),
.B(n_225),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_291),
.A2(n_294),
.B(n_296),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_293),
.A2(n_295),
.B1(n_278),
.B2(n_284),
.Y(n_297)
);

OAI31xp33_ASAP7_75t_L g296 ( 
.A1(n_279),
.A2(n_283),
.A3(n_280),
.B(n_261),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_297),
.A2(n_299),
.B1(n_301),
.B2(n_294),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_289),
.B(n_281),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_298),
.B(n_289),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_290),
.A2(n_278),
.B1(n_287),
.B2(n_264),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_292),
.A2(n_264),
.B1(n_285),
.B2(n_282),
.Y(n_301)
);

NAND3xp33_ASAP7_75t_L g302 ( 
.A(n_296),
.B(n_269),
.C(n_266),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_286),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_271),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_304),
.B(n_305),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_307),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_205),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_310),
.B(n_305),
.C(n_301),
.Y(n_311)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_311),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_309),
.B(n_223),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_308),
.C(n_223),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_SL g315 ( 
.A1(n_314),
.A2(n_231),
.B(n_312),
.Y(n_315)
);


endmodule