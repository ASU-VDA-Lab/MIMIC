module real_jpeg_20194_n_16 (n_5, n_4, n_8, n_0, n_12, n_339, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_339;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_1),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_1),
.A2(n_23),
.B1(n_40),
.B2(n_41),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g66 ( 
.A1(n_1),
.A2(n_23),
.B1(n_26),
.B2(n_28),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_1),
.A2(n_23),
.B1(n_46),
.B2(n_47),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_2),
.A2(n_22),
.B1(n_24),
.B2(n_123),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_2),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_2),
.A2(n_26),
.B1(n_28),
.B2(n_123),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_2),
.A2(n_40),
.B1(n_41),
.B2(n_123),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_2),
.A2(n_46),
.B1(n_47),
.B2(n_123),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_3),
.A2(n_26),
.B1(n_28),
.B2(n_116),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_3),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_22),
.B1(n_24),
.B2(n_116),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_46),
.B1(n_47),
.B2(n_116),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_116),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_4),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_4),
.B(n_25),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g171 ( 
.A1(n_4),
.A2(n_14),
.B(n_47),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_4),
.A2(n_40),
.B1(n_41),
.B2(n_121),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_4),
.A2(n_95),
.B1(n_100),
.B2(n_180),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_4),
.B(n_75),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_4),
.B(n_28),
.Y(n_207)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_28),
.B(n_207),
.Y(n_211)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_6),
.A2(n_22),
.B1(n_24),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_6),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_46),
.B1(n_47),
.B2(n_57),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g247 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_57),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g293 ( 
.A1(n_6),
.A2(n_26),
.B1(n_28),
.B2(n_57),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_7),
.A2(n_22),
.B1(n_24),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_7),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_55),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_46),
.B1(n_47),
.B2(n_55),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g272 ( 
.A1(n_7),
.A2(n_26),
.B1(n_28),
.B2(n_55),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_8),
.B(n_46),
.Y(n_96)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_8),
.Y(n_100)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_8),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_8),
.B(n_199),
.Y(n_198)
);

BUFx8_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_10),
.A2(n_26),
.B1(n_28),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_10),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_10),
.A2(n_46),
.B1(n_47),
.B2(n_118),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_118),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_10),
.A2(n_22),
.B1(n_24),
.B2(n_118),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_12),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_25)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g30 ( 
.A1(n_13),
.A2(n_22),
.B1(n_24),
.B2(n_31),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_13),
.A2(n_26),
.B1(n_28),
.B2(n_31),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_31),
.B1(n_46),
.B2(n_47),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_13),
.A2(n_31),
.B1(n_40),
.B2(n_41),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_L g39 ( 
.A1(n_14),
.A2(n_40),
.B(n_44),
.C(n_45),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_14),
.B(n_40),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_14),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g48 ( 
.A(n_14),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_15),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_83),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_81),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_34),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_19),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_29),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g274 ( 
.A1(n_20),
.A2(n_53),
.B(n_255),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_25),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_22),
.Y(n_24)
);

O2A1O1Ixp33_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_25),
.B(n_27),
.C(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_27),
.Y(n_33)
);

HAxp5_ASAP7_75t_SL g120 ( 
.A(n_22),
.B(n_121),
.CON(n_120),
.SN(n_120)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_25),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_25),
.B(n_30),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_32),
.B1(n_120),
.B2(n_122),
.Y(n_119)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_26),
.A2(n_33),
.B1(n_120),
.B2(n_127),
.Y(n_126)
);

AOI32xp33_ASAP7_75t_L g206 ( 
.A1(n_26),
.A2(n_40),
.A3(n_65),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_27),
.B(n_28),
.Y(n_127)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_28),
.A2(n_63),
.B(n_64),
.C(n_70),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_64),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_29),
.A2(n_54),
.B(n_58),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_32),
.Y(n_29)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_32),
.A2(n_78),
.B(n_79),
.Y(n_77)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_35),
.B(n_82),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_73),
.C(n_77),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_36),
.A2(n_37),
.B1(n_333),
.B2(n_335),
.Y(n_332)
);

CKINVDCx16_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_51),
.C(n_59),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_38),
.A2(n_313),
.B1(n_314),
.B2(n_315),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_38),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_38),
.A2(n_59),
.B1(n_60),
.B2(n_313),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_45),
.B(n_49),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_39),
.A2(n_49),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_39),
.A2(n_45),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_39),
.A2(n_45),
.B1(n_175),
.B2(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_39),
.A2(n_45),
.B1(n_196),
.B2(n_214),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_39),
.A2(n_214),
.B(n_229),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_39),
.A2(n_45),
.B1(n_103),
.B2(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g281 ( 
.A1(n_39),
.A2(n_111),
.B(n_247),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_41),
.B1(n_64),
.B2(n_65),
.Y(n_63)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_41),
.A2(n_48),
.B(n_121),
.C(n_171),
.Y(n_170)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_41),
.B(n_64),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g102 ( 
.A1(n_45),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_45),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_45),
.B(n_121),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_46),
.B(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_50),
.B(n_112),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_51),
.A2(n_52),
.B1(n_321),
.B2(n_322),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_56),
.B2(n_58),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_53),
.A2(n_58),
.B1(n_133),
.B2(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_53),
.A2(n_58),
.B1(n_134),
.B2(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_53),
.A2(n_80),
.B(n_301),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_67),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_62),
.A2(n_68),
.B(n_137),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_66),
.Y(n_62)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_63),
.A2(n_69),
.B1(n_115),
.B2(n_117),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_63),
.A2(n_69),
.B1(n_153),
.B2(n_211),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_63),
.B(n_72),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_63),
.A2(n_67),
.B(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_63),
.A2(n_69),
.B1(n_272),
.B2(n_293),
.Y(n_292)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_71),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_68),
.A2(n_75),
.B(n_76),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_68),
.A2(n_75),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_68),
.A2(n_76),
.B(n_258),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_68),
.A2(n_258),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_73),
.A2(n_74),
.B1(n_77),
.B2(n_334),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_77),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g79 ( 
.A(n_80),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_330),
.B(n_336),
.Y(n_83)
);

OAI321xp33_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_306),
.A3(n_325),
.B1(n_328),
.B2(n_329),
.C(n_339),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_285),
.B(n_305),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_87),
.A2(n_263),
.B(n_284),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_155),
.B(n_238),
.C(n_262),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_139),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_89),
.B(n_139),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B1(n_124),
.B2(n_138),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_108),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_92),
.B(n_108),
.C(n_138),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B1(n_102),
.B2(n_107),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_93),
.B(n_107),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_95),
.A2(n_97),
.B(n_98),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_97),
.B1(n_100),
.B2(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_95),
.A2(n_164),
.B1(n_180),
.B2(n_181),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_95),
.A2(n_167),
.B(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_95),
.A2(n_181),
.B(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_96),
.B(n_149),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_96),
.A2(n_163),
.B1(n_165),
.B2(n_166),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g205 ( 
.A1(n_96),
.A2(n_99),
.B(n_199),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_101),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_100),
.A2(n_129),
.B(n_148),
.Y(n_147)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_100),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_100),
.B(n_121),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_102),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_104),
.B(n_229),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_106),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_105),
.B(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_113),
.C(n_119),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_109),
.A2(n_110),
.B1(n_113),
.B2(n_114),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_117),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_119),
.B(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_122),
.Y(n_133)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_125),
.B(n_131),
.C(n_136),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_128),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_128),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_130)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_142),
.C(n_144),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_140),
.B(n_235),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_150),
.C(n_151),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_146),
.A2(n_147),
.B1(n_150),
.B2(n_225),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_148),
.B(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_150),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_151),
.B(n_224),
.Y(n_223)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_156),
.B(n_237),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_157),
.A2(n_232),
.B(n_236),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_219),
.B(n_231),
.Y(n_157)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_201),
.B(n_218),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_160),
.A2(n_188),
.B(n_200),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_176),
.B(n_187),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_168),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_162),
.B(n_168),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_170),
.B1(n_172),
.B2(n_173),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_170),
.B(n_172),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_182),
.B(n_186),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_178),
.B(n_179),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_190),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_189),
.B(n_190),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_197),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_192),
.A2(n_193),
.B1(n_194),
.B2(n_195),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_192),
.B(n_195),
.C(n_197),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_199),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_203),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_203),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_209),
.B1(n_216),
.B2(n_217),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_204),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_206),
.Y(n_230)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_212),
.B1(n_213),
.B2(n_215),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_210),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_212),
.B(n_215),
.C(n_216),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_220),
.B(n_221),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_226),
.B2(n_227),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_228),
.C(n_230),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_223),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_230),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_233),
.B(n_234),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_239),
.B(n_240),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_241),
.A2(n_242),
.B1(n_260),
.B2(n_261),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_249),
.C(n_261),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_245),
.B(n_246),
.Y(n_269)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_251),
.B1(n_252),
.B2(n_259),
.Y(n_249)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_250),
.Y(n_259)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_253),
.A2(n_254),
.B1(n_256),
.B2(n_257),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_257),
.C(n_259),
.Y(n_283)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_260),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_264),
.B(n_265),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_283),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_276),
.B2(n_277),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_267),
.B(n_277),
.C(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_269),
.B(n_273),
.C(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_271),
.A2(n_273),
.B1(n_274),
.B2(n_275),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_271),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g273 ( 
.A(n_274),
.Y(n_273)
);

CKINVDCx14_ASAP7_75t_R g276 ( 
.A(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_279),
.B1(n_281),
.B2(n_282),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_278),
.A2(n_279),
.B1(n_300),
.B2(n_302),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_278),
.A2(n_296),
.B(n_300),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_279),
.B(n_281),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_281),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_286),
.B(n_287),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_289),
.B1(n_303),
.B2(n_304),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_290),
.B(n_295),
.C(n_304),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_292),
.B(n_294),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_291),
.B(n_292),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_293),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_308),
.C(n_317),
.Y(n_307)
);

FAx1_ASAP7_75t_SL g327 ( 
.A(n_294),
.B(n_308),
.CI(n_317),
.CON(n_327),
.SN(n_327)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_297),
.B1(n_298),
.B2(n_299),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_300),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_303),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_318),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_307),
.B(n_318),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_309),
.A2(n_310),
.B1(n_320),
.B2(n_323),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_310),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_310),
.B(n_313),
.C(n_315),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_310),
.B(n_323),
.C(n_324),
.Y(n_331)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_324),
.Y(n_318)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_320),
.Y(n_323)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_326),
.B(n_327),
.Y(n_328)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_327),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_331),
.B(n_332),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

CKINVDCx14_ASAP7_75t_R g335 ( 
.A(n_333),
.Y(n_335)
);


endmodule