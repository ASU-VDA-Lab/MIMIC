module fake_jpeg_29212_n_125 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_125);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_125;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_5),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_34),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_14),
.Y(n_49)
);

BUFx16f_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g51 ( 
.A(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_16),
.B(n_3),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_23),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_20),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_54),
.B(n_45),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_57),
.B1(n_59),
.B2(n_53),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_49),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_56),
.B(n_42),
.Y(n_64)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_48),
.A2(n_21),
.B1(n_39),
.B2(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_4),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_43),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_45),
.B1(n_50),
.B2(n_43),
.Y(n_70)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_61),
.Y(n_68)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_64),
.B(n_26),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_54),
.B(n_47),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_69),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_53),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_70),
.A2(n_72),
.B1(n_9),
.B2(n_10),
.Y(n_83)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_71),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_62),
.A2(n_50),
.B(n_51),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_7),
.B(n_8),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_74),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_6),
.Y(n_77)
);

A2O1A1Ixp33_ASAP7_75t_L g76 ( 
.A1(n_75),
.A2(n_50),
.B(n_52),
.C(n_8),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_76),
.B(n_77),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_46),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_78),
.B(n_85),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g100 ( 
.A1(n_80),
.A2(n_82),
.B(n_28),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_9),
.B(n_10),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_84),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_72),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_11),
.Y(n_85)
);

BUFx12f_ASAP7_75t_SL g87 ( 
.A(n_63),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_40),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_17),
.C(n_18),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_89),
.B(n_31),
.C(n_33),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_19),
.B1(n_22),
.B2(n_25),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_66),
.B1(n_29),
.B2(n_30),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_91),
.B(n_27),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_93),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_71),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_79),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_66),
.Y(n_97)
);

NAND3xp33_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_100),
.C(n_105),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_86),
.B1(n_102),
.B2(n_101),
.Y(n_115)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_87),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_99),
.A2(n_104),
.B(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_35),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_36),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_76),
.C(n_89),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_102),
.B1(n_94),
.B2(n_103),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_109),
.A2(n_115),
.B1(n_99),
.B2(n_104),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_112),
.B(n_114),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_106),
.C(n_100),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_116),
.B(n_118),
.C(n_112),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_117),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_116),
.C(n_119),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_121),
.B(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_123),
.A2(n_108),
.B(n_113),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_124),
.B(n_108),
.Y(n_125)
);


endmodule