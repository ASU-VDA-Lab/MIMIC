module fake_jpeg_27897_n_145 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_145);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_145;

wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_103;
wire n_50;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx10_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_21),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_22),
.B(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_11),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_29),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_2),
.B(n_8),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_8),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_46),
.A2(n_48),
.B1(n_43),
.B2(n_59),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_63),
.A2(n_42),
.B1(n_60),
.B2(n_58),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_0),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_64),
.B(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_55),
.B(n_0),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_56),
.Y(n_67)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_67),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_67),
.B(n_51),
.Y(n_72)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_72),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_76),
.A2(n_83),
.B1(n_1),
.B2(n_2),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_61),
.Y(n_77)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_77),
.Y(n_96)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_78),
.B(n_81),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_52),
.B1(n_49),
.B2(n_53),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_80),
.A2(n_45),
.B1(n_58),
.B2(n_4),
.Y(n_92)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_82),
.Y(n_99)
);

HAxp5_ASAP7_75t_SL g83 ( 
.A(n_62),
.B(n_45),
.CON(n_83),
.SN(n_83)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_60),
.C(n_42),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_84),
.B(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_57),
.C(n_50),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_89),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_80),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_97),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_92),
.A2(n_93),
.B1(n_94),
.B2(n_98),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g94 ( 
.A1(n_74),
.A2(n_26),
.B1(n_41),
.B2(n_40),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_69),
.A2(n_81),
.B1(n_83),
.B2(n_28),
.Y(n_98)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_69),
.Y(n_100)
);

INVx13_ASAP7_75t_L g102 ( 
.A(n_100),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_96),
.B(n_23),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_103),
.B(n_105),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_24),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_92),
.A2(n_20),
.B1(n_39),
.B2(n_38),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_108),
.A2(n_91),
.B1(n_87),
.B2(n_99),
.Y(n_115)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_106),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_114),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_103),
.B(n_107),
.Y(n_112)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_93),
.B1(n_98),
.B2(n_100),
.Y(n_113)
);

OA22x2_ASAP7_75t_L g128 ( 
.A1(n_113),
.A2(n_115),
.B1(n_5),
.B2(n_6),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_101),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_85),
.Y(n_116)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_95),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_1),
.B(n_4),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_110),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g129 ( 
.A(n_118),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_114),
.A2(n_105),
.B(n_104),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_120),
.B(n_122),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_117),
.A2(n_108),
.B(n_102),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_116),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_124),
.B(n_127),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_125),
.A2(n_128),
.B1(n_119),
.B2(n_121),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_116),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_102),
.Y(n_127)
);

INVxp33_ASAP7_75t_SL g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_130),
.Y(n_135)
);

AOI221xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_132),
.B1(n_128),
.B2(n_127),
.C(n_123),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_133),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_134),
.C(n_135),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_129),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_139),
.B(n_130),
.C(n_32),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_30),
.C(n_36),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_18),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_13),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_143),
.A2(n_33),
.B(n_35),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_144),
.B(n_12),
.Y(n_145)
);


endmodule