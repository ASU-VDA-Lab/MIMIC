module real_jpeg_1193_n_15 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_15);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_104;
wire n_153;
wire n_161;
wire n_64;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_173;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_164;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_175;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_30;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_167;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g51 ( 
.A(n_0),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_1),
.A2(n_50),
.B1(n_52),
.B2(n_58),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_1),
.Y(n_58)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_3),
.A2(n_25),
.B1(n_26),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_3),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_3),
.A2(n_30),
.B1(n_32),
.B2(n_67),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_3),
.A2(n_50),
.B1(n_52),
.B2(n_67),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_4),
.B(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_4),
.B(n_24),
.C(n_26),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_4),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_4),
.B(n_23),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_4),
.B(n_52),
.C(n_62),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_4),
.A2(n_25),
.B1(n_26),
.B2(n_90),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_4),
.B(n_56),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_70),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_4),
.A2(n_30),
.B1(n_32),
.B2(n_90),
.Y(n_165)
);

OAI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_5),
.A2(n_30),
.B1(n_32),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_5),
.A2(n_25),
.B1(n_26),
.B2(n_36),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_5),
.A2(n_36),
.B1(n_50),
.B2(n_52),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_5),
.A2(n_36),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_50),
.B1(n_52),
.B2(n_114),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_8),
.Y(n_114)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_11),
.A2(n_25),
.B1(n_26),
.B2(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_30),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_13),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_33),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_33),
.B1(n_50),
.B2(n_52),
.Y(n_150)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_117),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_116),
.Y(n_16)
);

INVxp67_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_19),
.B(n_80),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_59),
.C(n_72),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_20),
.B(n_173),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_39),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_21),
.B(n_40),
.C(n_48),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_29),
.B(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_22),
.A2(n_29),
.B1(n_97),
.B2(n_98),
.Y(n_96)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_23),
.B(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_23),
.B(n_35),
.Y(n_166)
);

AO22x2_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_23)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g38 ( 
.A1(n_24),
.A2(n_28),
.B1(n_30),
.B2(n_32),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_26),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_26),
.B(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_30),
.A2(n_32),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AOI32xp33_ASAP7_75t_L g107 ( 
.A1(n_30),
.A2(n_44),
.A3(n_87),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_32),
.B(n_75),
.Y(n_74)
);

NAND2xp33_ASAP7_75t_SL g109 ( 
.A(n_32),
.B(n_45),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_47),
.B2(n_48),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_85),
.Y(n_84)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_43),
.B(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_44),
.A2(n_45),
.B1(n_86),
.B2(n_87),
.Y(n_94)
);

INVx6_ASAP7_75t_SL g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_54),
.B1(n_55),
.B2(n_57),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_55),
.B(n_77),
.Y(n_76)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_50),
.A2(n_52),
.B1(n_62),
.B2(n_63),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_52),
.B(n_145),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_54),
.A2(n_55),
.B1(n_57),
.B2(n_112),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_54),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_54),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_54),
.A2(n_55),
.B1(n_123),
.B2(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_79),
.Y(n_125)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_78),
.B(n_150),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_59),
.B(n_72),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_60),
.A2(n_65),
.B(n_68),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_71),
.Y(n_102)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_60),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.Y(n_60)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_64),
.A2(n_100),
.B(n_102),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_64),
.A2(n_102),
.B(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_64),
.A2(n_66),
.B1(n_131),
.B2(n_139),
.Y(n_167)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_69),
.A2(n_139),
.B(n_140),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_71),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_76),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_73),
.A2(n_74),
.B1(n_76),
.B2(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_76),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_104),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_95),
.B2(n_103),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_90),
.B(n_91),
.C(n_92),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_90),
.Y(n_91)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI21xp5_ASAP7_75t_L g146 ( 
.A1(n_90),
.A2(n_125),
.B(n_147),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_91),
.Y(n_108)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_95),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_97),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_111),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_118),
.A2(n_171),
.B(n_175),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_160),
.B(n_170),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_120),
.A2(n_141),
.B(n_159),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_121),
.B(n_134),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_121),
.B(n_134),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_126),
.B1(n_132),
.B2(n_133),
.Y(n_121)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_129),
.C(n_132),
.Y(n_161)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_138),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_153),
.B(n_158),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_148),
.B(n_152),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_151),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_151),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_150),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_156),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_162),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_168),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_167),
.C(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_174),
.Y(n_175)
);


endmodule