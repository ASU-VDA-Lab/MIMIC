module fake_jpeg_24708_n_284 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_21;
wire n_57;
wire n_187;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx3_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx8_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx6f_ASAP7_75t_SL g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g30 ( 
.A(n_24),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_30),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_17),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_32),
.B(n_34),
.Y(n_51)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g56 ( 
.A(n_36),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_40),
.B(n_42),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_33),
.A2(n_15),
.B1(n_14),
.B2(n_27),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_43),
.A2(n_35),
.B1(n_18),
.B2(n_21),
.Y(n_72)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_44),
.Y(n_66)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_45),
.B(n_49),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_55),
.Y(n_60)
);

NAND2x1_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_24),
.Y(n_48)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_50),
.B(n_28),
.C(n_22),
.Y(n_73)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_37),
.A2(n_14),
.B1(n_15),
.B2(n_22),
.Y(n_50)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_34),
.B(n_18),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_37),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_57),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_33),
.A2(n_15),
.B1(n_14),
.B2(n_24),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_35),
.B1(n_38),
.B2(n_24),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_33),
.B1(n_35),
.B2(n_49),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_61),
.A2(n_65),
.B1(n_73),
.B2(n_44),
.Y(n_100)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_56),
.Y(n_64)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_68),
.B(n_69),
.Y(n_103)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_70),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_76),
.Y(n_94)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_72),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_58),
.B(n_29),
.Y(n_84)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_56),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_39),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_77),
.B(n_17),
.Y(n_93)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_59),
.Y(n_79)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_84),
.A2(n_21),
.B(n_74),
.Y(n_108)
);

OAI32xp33_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_51),
.A3(n_50),
.B1(n_43),
.B2(n_32),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_85),
.B(n_92),
.Y(n_111)
);

AO22x2_ASAP7_75t_L g86 ( 
.A1(n_82),
.A2(n_47),
.B1(n_52),
.B2(n_29),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_86),
.A2(n_98),
.B1(n_100),
.B2(n_72),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_60),
.B(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_93),
.B(n_17),
.Y(n_121)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_95),
.B(n_96),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_52),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_52),
.Y(n_97)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_79),
.A2(n_47),
.B1(n_21),
.B2(n_39),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_76),
.B(n_47),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_30),
.Y(n_102)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_SL g105 ( 
.A(n_67),
.B(n_23),
.C(n_16),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_77),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_86),
.B1(n_98),
.B2(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_107),
.B(n_113),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_108),
.A2(n_110),
.B(n_128),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_78),
.B(n_67),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_112),
.B(n_115),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_75),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_83),
.A2(n_40),
.B1(n_54),
.B2(n_53),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_116),
.A2(n_119),
.B1(n_89),
.B2(n_86),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_87),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_120),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_83),
.A2(n_64),
.B1(n_80),
.B2(n_66),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_121),
.B(n_125),
.Y(n_147)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_104),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_122),
.Y(n_130)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_99),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_127),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_101),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_91),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_126),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_94),
.B(n_23),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_63),
.B(n_66),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_101),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_125),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_131),
.B(n_152),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_88),
.B1(n_90),
.B2(n_86),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_132),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_100),
.B1(n_89),
.B2(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_123),
.B1(n_86),
.B2(n_109),
.Y(n_135)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_119),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_141),
.B(n_145),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_109),
.A2(n_86),
.B1(n_85),
.B2(n_98),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_144),
.B1(n_146),
.B2(n_148),
.Y(n_167)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_143),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_120),
.A2(n_98),
.B1(n_94),
.B2(n_103),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_98),
.B1(n_102),
.B2(n_103),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_92),
.B1(n_91),
.B2(n_95),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_118),
.A2(n_104),
.B1(n_80),
.B2(n_62),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_149),
.A2(n_153),
.B1(n_132),
.B2(n_134),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_111),
.B(n_70),
.C(n_25),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_150),
.B(n_126),
.C(n_26),
.Y(n_170)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_108),
.A2(n_70),
.B1(n_19),
.B2(n_28),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_143),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_154),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_140),
.A2(n_110),
.B(n_111),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_174),
.B(n_165),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_156),
.B(n_164),
.Y(n_182)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_151),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_158),
.B(n_160),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_138),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_159),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_149),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_139),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_142),
.A2(n_128),
.B1(n_129),
.B2(n_117),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_136),
.B1(n_137),
.B2(n_147),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g164 ( 
.A(n_147),
.B(n_121),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_165),
.B(n_172),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_122),
.Y(n_166)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_166),
.Y(n_185)
);

NAND3xp33_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_127),
.C(n_112),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_168),
.B(n_176),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_170),
.B(n_175),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g171 ( 
.A(n_130),
.Y(n_171)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_171),
.Y(n_187)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

BUFx5_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

AND2x4_ASAP7_75t_L g174 ( 
.A(n_140),
.B(n_26),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_25),
.Y(n_175)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_26),
.CI(n_25),
.CON(n_176),
.SN(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_145),
.B(n_25),
.C(n_26),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_175),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_172),
.A2(n_141),
.B1(n_152),
.B2(n_146),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_179),
.A2(n_176),
.B1(n_178),
.B2(n_19),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g180 ( 
.A(n_173),
.Y(n_180)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_180),
.Y(n_205)
);

OAI21xp33_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_133),
.B(n_153),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_183),
.A2(n_192),
.B(n_20),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_174),
.B(n_163),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_169),
.B(n_144),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_190),
.B(n_198),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_174),
.B(n_156),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_195),
.A2(n_190),
.B1(n_188),
.B2(n_184),
.Y(n_216)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_196),
.B(n_197),
.Y(n_211)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_199),
.B(n_200),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_155),
.B(n_22),
.Y(n_200)
);

NOR3xp33_ASAP7_75t_SL g201 ( 
.A(n_186),
.B(n_176),
.C(n_167),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_215),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g202 ( 
.A(n_191),
.Y(n_202)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_202),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_161),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_217),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_191),
.A2(n_160),
.B1(n_158),
.B2(n_170),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_185),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_189),
.B(n_199),
.C(n_181),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_209),
.B(n_182),
.C(n_188),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_181),
.A2(n_19),
.B1(n_1),
.B2(n_2),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_193),
.Y(n_212)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_212),
.Y(n_234)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_20),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_213),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_20),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_189),
.B(n_20),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_223),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_222),
.B(n_229),
.C(n_232),
.Y(n_243)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_209),
.B(n_183),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_225),
.B(n_208),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_211),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_227),
.B(n_233),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_204),
.Y(n_228)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_228),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_214),
.B(n_187),
.C(n_192),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_218),
.A2(n_192),
.B1(n_8),
.B2(n_9),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_230),
.A2(n_6),
.B1(n_13),
.B2(n_12),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_202),
.B(n_20),
.C(n_1),
.Y(n_232)
);

INVx13_ASAP7_75t_L g233 ( 
.A(n_205),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_236),
.B(n_220),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_235),
.A2(n_201),
.B1(n_203),
.B2(n_208),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_238),
.A2(n_245),
.B1(n_243),
.B2(n_237),
.Y(n_255)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_240),
.B(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_228),
.A2(n_217),
.B1(n_7),
.B2(n_10),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_11),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_222),
.B(n_6),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_226),
.Y(n_250)
);

AO22x2_ASAP7_75t_L g245 ( 
.A1(n_229),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_245),
.A2(n_246),
.B(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

NOR2xp67_ASAP7_75t_SL g249 ( 
.A(n_245),
.B(n_224),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_250),
.B(n_251),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_248),
.B(n_223),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_247),
.B(n_234),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_252),
.B(n_254),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_255),
.C(n_245),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_243),
.B(n_233),
.Y(n_256)
);

OR2x2_ASAP7_75t_L g263 ( 
.A(n_256),
.B(n_259),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_239),
.A2(n_11),
.B(n_4),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_258),
.A2(n_4),
.B(n_5),
.Y(n_268)
);

INVxp33_ASAP7_75t_L g260 ( 
.A(n_257),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_268),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_241),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_264),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_236),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_267),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_269),
.B(n_272),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_4),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_273),
.B(n_10),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_261),
.C(n_263),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.C(n_277),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_271),
.B(n_263),
.Y(n_276)
);

AOI311xp33_ASAP7_75t_L g280 ( 
.A1(n_276),
.A2(n_270),
.A3(n_12),
.B(n_13),
.C(n_3),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_281),
.B(n_279),
.C(n_278),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_3),
.C(n_20),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_3),
.Y(n_284)
);


endmodule