module fake_aes_1052_n_889 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_99, n_93, n_51, n_96, n_39, n_889);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_99;
input n_93;
input n_51;
input n_96;
input n_39;
output n_889;
wire n_117;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_125;
wire n_431;
wire n_484;
wire n_862;
wire n_852;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_152;
wire n_113;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_157;
wire n_765;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_789;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_860;
wire n_401;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_830;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_780;
wire n_726;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_171;
wire n_567;
wire n_809;
wire n_888;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_490;
wire n_247;
wire n_393;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_107;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_622;
wire n_549;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_799;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_716;
wire n_653;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_754;
wire n_775;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_870;
wire n_148;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_168;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_782;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_763;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_837;
wire n_128;
wire n_129;
wire n_410;
wire n_774;
wire n_867;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_785;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_781;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g106 ( .A(n_105), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_75), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_22), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_83), .Y(n_109) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_25), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_7), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_77), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_43), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_45), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_36), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_60), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_59), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_74), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_19), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_81), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_24), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_51), .Y(n_123) );
INVxp67_ASAP7_75t_L g124 ( .A(n_96), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_54), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_12), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_6), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_47), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_66), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_20), .Y(n_131) );
BUFx6f_ASAP7_75t_L g132 ( .A(n_40), .Y(n_132) );
INVx1_ASAP7_75t_SL g133 ( .A(n_78), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_57), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_62), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_11), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_52), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_95), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_28), .Y(n_139) );
INVxp67_ASAP7_75t_SL g140 ( .A(n_0), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_69), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_20), .Y(n_142) );
INVx1_ASAP7_75t_SL g143 ( .A(n_85), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_61), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_137), .Y(n_145) );
INVx6_ASAP7_75t_L g146 ( .A(n_132), .Y(n_146) );
INVx3_ASAP7_75t_L g147 ( .A(n_122), .Y(n_147) );
BUFx12f_ASAP7_75t_L g148 ( .A(n_107), .Y(n_148) );
NOR2xp33_ASAP7_75t_L g149 ( .A(n_123), .B(n_0), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_122), .B(n_1), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_106), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_108), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_137), .B(n_1), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_108), .Y(n_155) );
AND2x4_ASAP7_75t_L g156 ( .A(n_136), .B(n_2), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_141), .Y(n_157) );
INVx5_ASAP7_75t_L g158 ( .A(n_132), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_126), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_115), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_115), .Y(n_161) );
INVx3_ASAP7_75t_L g162 ( .A(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_141), .B(n_3), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_117), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_118), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_118), .Y(n_167) );
INVx6_ASAP7_75t_L g168 ( .A(n_132), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_132), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_120), .Y(n_170) );
AOI22xp33_ASAP7_75t_L g171 ( .A1(n_156), .A2(n_131), .B1(n_119), .B2(n_142), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_150), .B(n_110), .Y(n_172) );
NAND2xp33_ASAP7_75t_SL g173 ( .A(n_156), .B(n_112), .Y(n_173) );
NAND2xp33_ASAP7_75t_L g174 ( .A(n_150), .B(n_132), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_156), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_152), .B(n_124), .Y(n_176) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_156), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_152), .B(n_113), .Y(n_179) );
INVx2_ASAP7_75t_SL g180 ( .A(n_147), .Y(n_180) );
CKINVDCx6p67_ASAP7_75t_R g181 ( .A(n_148), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
BUFx10_ASAP7_75t_L g183 ( .A(n_153), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_147), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_153), .Y(n_185) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_155), .B(n_109), .Y(n_186) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_155), .B(n_114), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_160), .B(n_116), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_158), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_165), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_165), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_166), .Y(n_192) );
INVx2_ASAP7_75t_L g193 ( .A(n_158), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_148), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_160), .B(n_161), .Y(n_195) );
AND3x2_ASAP7_75t_L g196 ( .A(n_149), .B(n_140), .C(n_111), .Y(n_196) );
INVxp33_ASAP7_75t_SL g197 ( .A(n_159), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_161), .B(n_135), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_164), .B(n_113), .Y(n_199) );
AND2x2_ASAP7_75t_L g200 ( .A(n_164), .B(n_111), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_166), .Y(n_201) );
CKINVDCx5p33_ASAP7_75t_R g202 ( .A(n_159), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_167), .B(n_144), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_158), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_167), .B(n_147), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_147), .Y(n_206) );
OR2x6_ASAP7_75t_L g207 ( .A(n_154), .B(n_119), .Y(n_207) );
INVx1_ASAP7_75t_SL g208 ( .A(n_170), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_170), .B(n_162), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g210 ( .A(n_163), .Y(n_210) );
AND2x4_ASAP7_75t_L g211 ( .A(n_162), .B(n_131), .Y(n_211) );
XOR2xp5_ASAP7_75t_L g212 ( .A(n_145), .B(n_127), .Y(n_212) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_157), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_157), .Y(n_216) );
OR2x2_ASAP7_75t_L g217 ( .A(n_162), .B(n_142), .Y(n_217) );
INVx1_ASAP7_75t_SL g218 ( .A(n_162), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_158), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_158), .Y(n_220) );
AOI22xp5_ASAP7_75t_L g221 ( .A1(n_173), .A2(n_120), .B1(n_121), .B2(n_125), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_184), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_185), .B(n_208), .Y(n_223) );
INVx1_ASAP7_75t_L g224 ( .A(n_218), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_182), .B(n_133), .Y(n_226) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_183), .B(n_121), .Y(n_227) );
O2A1O1Ixp5_ASAP7_75t_L g228 ( .A1(n_195), .A2(n_138), .B(n_128), .C(n_129), .Y(n_228) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_172), .B(n_143), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_183), .B(n_125), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_210), .B(n_128), .Y(n_231) );
BUFx3_ASAP7_75t_L g232 ( .A(n_184), .Y(n_232) );
NOR2xp67_ASAP7_75t_L g233 ( .A(n_217), .B(n_4), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_209), .Y(n_234) );
INVx3_ASAP7_75t_L g235 ( .A(n_184), .Y(n_235) );
AND2x4_ASAP7_75t_SL g236 ( .A(n_181), .B(n_129), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_210), .B(n_130), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_175), .A2(n_139), .B1(n_138), .B2(n_130), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g239 ( .A(n_217), .B(n_5), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_211), .Y(n_240) );
NAND2x1p5_ASAP7_75t_L g241 ( .A(n_211), .B(n_139), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_188), .B(n_134), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_198), .B(n_134), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_203), .B(n_146), .Y(n_244) );
INVx2_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
BUFx4f_ASAP7_75t_L g246 ( .A(n_181), .Y(n_246) );
AND2x4_ASAP7_75t_SL g247 ( .A(n_194), .B(n_169), .Y(n_247) );
NAND2xp5_ASAP7_75t_SL g248 ( .A(n_178), .B(n_169), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_206), .Y(n_249) );
NOR3xp33_ASAP7_75t_L g250 ( .A(n_173), .B(n_6), .C(n_7), .Y(n_250) );
OR2x2_ASAP7_75t_L g251 ( .A(n_212), .B(n_8), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_211), .Y(n_252) );
NAND2xp33_ASAP7_75t_L g253 ( .A(n_171), .B(n_169), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_207), .B(n_146), .Y(n_254) );
AND2x2_ASAP7_75t_L g255 ( .A(n_207), .B(n_8), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_205), .Y(n_256) );
OAI22xp5_ASAP7_75t_L g257 ( .A1(n_207), .A2(n_168), .B1(n_146), .B2(n_169), .Y(n_257) );
AOI221x1_ASAP7_75t_L g258 ( .A1(n_206), .A2(n_168), .B1(n_146), .B2(n_56), .C(n_58), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_213), .A2(n_168), .B1(n_10), .B2(n_11), .Y(n_259) );
AND2x6_ASAP7_75t_SL g260 ( .A(n_194), .B(n_9), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_215), .Y(n_261) );
INVx2_ASAP7_75t_SL g262 ( .A(n_207), .Y(n_262) );
BUFx3_ASAP7_75t_L g263 ( .A(n_180), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_180), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g265 ( .A1(n_179), .A2(n_168), .B(n_55), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_200), .B(n_9), .Y(n_266) );
NAND3xp33_ASAP7_75t_L g267 ( .A(n_196), .B(n_10), .C(n_12), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_213), .A2(n_13), .B1(n_14), .B2(n_15), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_186), .B(n_63), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_216), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_200), .B(n_13), .Y(n_271) );
NOR2xp33_ASAP7_75t_R g272 ( .A(n_202), .B(n_14), .Y(n_272) );
O2A1O1Ixp33_ASAP7_75t_L g273 ( .A1(n_190), .A2(n_15), .B(n_16), .C(n_17), .Y(n_273) );
BUFx6f_ASAP7_75t_L g274 ( .A(n_232), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_271), .A2(n_197), .B1(n_202), .B2(n_192), .Y(n_275) );
OAI22x1_ASAP7_75t_L g276 ( .A1(n_268), .A2(n_197), .B1(n_176), .B2(n_187), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_232), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_227), .A2(n_174), .B(n_199), .Y(n_278) );
OAI21xp5_ASAP7_75t_L g279 ( .A1(n_256), .A2(n_191), .B(n_201), .Y(n_279) );
AOI33xp33_ASAP7_75t_L g280 ( .A1(n_238), .A2(n_220), .A3(n_214), .B1(n_204), .B2(n_193), .B3(n_189), .Y(n_280) );
NAND2xp5_ASAP7_75t_SL g281 ( .A(n_262), .B(n_220), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_234), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_273), .A2(n_174), .B(n_214), .C(n_204), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_223), .B(n_219), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_240), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_231), .B(n_219), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_236), .B(n_16), .Y(n_287) );
AOI21xp33_ASAP7_75t_L g288 ( .A1(n_262), .A2(n_193), .B(n_189), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_236), .B(n_17), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_252), .Y(n_290) );
OR2x2_ASAP7_75t_L g291 ( .A(n_251), .B(n_18), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_271), .Y(n_292) );
AOI21xp5_ASAP7_75t_L g293 ( .A1(n_227), .A2(n_177), .B(n_68), .Y(n_293) );
AO21x1_ASAP7_75t_L g294 ( .A1(n_265), .A2(n_18), .B(n_19), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_233), .A2(n_177), .B(n_23), .C(n_26), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_230), .A2(n_177), .B(n_27), .Y(n_296) );
OR2x4_ASAP7_75t_L g297 ( .A(n_246), .B(n_177), .Y(n_297) );
AOI21x1_ASAP7_75t_L g298 ( .A1(n_248), .A2(n_177), .B(n_29), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_271), .B(n_21), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_248), .A2(n_30), .B(n_31), .Y(n_300) );
NAND2x1p5_ASAP7_75t_L g301 ( .A(n_246), .B(n_32), .Y(n_301) );
INVx5_ASAP7_75t_L g302 ( .A(n_235), .Y(n_302) );
OAI22xp5_ASAP7_75t_L g303 ( .A1(n_241), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_303) );
O2A1O1Ixp5_ASAP7_75t_L g304 ( .A1(n_242), .A2(n_103), .B(n_38), .C(n_39), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_237), .B(n_37), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_235), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_241), .A2(n_41), .B1(n_42), .B2(n_44), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_235), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_225), .A2(n_46), .B(n_48), .Y(n_309) );
INVx5_ASAP7_75t_L g310 ( .A(n_255), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_239), .Y(n_311) );
INVx6_ASAP7_75t_L g312 ( .A(n_263), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_226), .B(n_49), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g314 ( .A1(n_275), .A2(n_224), .B1(n_238), .B2(n_266), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_282), .Y(n_315) );
OAI21xp5_ASAP7_75t_L g316 ( .A1(n_278), .A2(n_253), .B(n_228), .Y(n_316) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_287), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_285), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_290), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_275), .B(n_221), .Y(n_320) );
AOI21xp5_ASAP7_75t_L g321 ( .A1(n_305), .A2(n_243), .B(n_253), .Y(n_321) );
AOI21xp5_ASAP7_75t_L g322 ( .A1(n_286), .A2(n_264), .B(n_222), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_291), .B(n_229), .Y(n_323) );
NOR2xp33_ASAP7_75t_R g324 ( .A(n_289), .B(n_260), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_279), .Y(n_325) );
OAI21xp5_ASAP7_75t_SL g326 ( .A1(n_301), .A2(n_247), .B(n_259), .Y(n_326) );
OAI21x1_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_304), .B(n_296), .Y(n_327) );
AOI21xp5_ASAP7_75t_L g328 ( .A1(n_284), .A2(n_264), .B(n_245), .Y(n_328) );
INVx4_ASAP7_75t_L g329 ( .A(n_312), .Y(n_329) );
O2A1O1Ixp5_ASAP7_75t_SL g330 ( .A1(n_311), .A2(n_257), .B(n_270), .C(n_261), .Y(n_330) );
OA21x2_ASAP7_75t_L g331 ( .A1(n_304), .A2(n_258), .B(n_244), .Y(n_331) );
OAI21x1_ASAP7_75t_L g332 ( .A1(n_309), .A2(n_254), .B(n_245), .Y(n_332) );
AOI221x1_ASAP7_75t_L g333 ( .A1(n_295), .A2(n_250), .B1(n_269), .B2(n_267), .C(n_222), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_293), .A2(n_249), .B(n_269), .Y(n_334) );
INVx3_ASAP7_75t_L g335 ( .A(n_274), .Y(n_335) );
BUFx2_ASAP7_75t_L g336 ( .A(n_312), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_306), .Y(n_337) );
BUFx12f_ASAP7_75t_L g338 ( .A(n_301), .Y(n_338) );
OAI21x1_ASAP7_75t_L g339 ( .A1(n_294), .A2(n_249), .B(n_263), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_281), .A2(n_247), .B(n_53), .Y(n_340) );
INVx3_ASAP7_75t_L g341 ( .A(n_335), .Y(n_341) );
INVx4_ASAP7_75t_L g342 ( .A(n_338), .Y(n_342) );
CKINVDCx6p67_ASAP7_75t_R g343 ( .A(n_338), .Y(n_343) );
OAI21x1_ASAP7_75t_L g344 ( .A1(n_327), .A2(n_300), .B(n_307), .Y(n_344) );
INVx1_ASAP7_75t_L g345 ( .A(n_318), .Y(n_345) );
AO21x2_ASAP7_75t_L g346 ( .A1(n_339), .A2(n_295), .B(n_283), .Y(n_346) );
OAI21x1_ASAP7_75t_L g347 ( .A1(n_327), .A2(n_303), .B(n_299), .Y(n_347) );
AOI21xp5_ASAP7_75t_L g348 ( .A1(n_321), .A2(n_292), .B(n_311), .Y(n_348) );
OAI21x1_ASAP7_75t_L g349 ( .A1(n_339), .A2(n_313), .B(n_281), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_315), .B(n_310), .Y(n_350) );
AO21x2_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_283), .B(n_288), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_318), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_325), .A2(n_308), .B(n_280), .Y(n_353) );
OAI21xp5_ASAP7_75t_L g354 ( .A1(n_330), .A2(n_280), .B(n_302), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_325), .B(n_276), .Y(n_355) );
OR2x2_ASAP7_75t_L g356 ( .A(n_320), .B(n_310), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_319), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_315), .Y(n_358) );
OAI21x1_ASAP7_75t_L g359 ( .A1(n_330), .A2(n_297), .B(n_302), .Y(n_359) );
OAI21x1_ASAP7_75t_L g360 ( .A1(n_334), .A2(n_297), .B(n_302), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_323), .B(n_310), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_319), .B(n_310), .Y(n_362) );
OA21x2_ASAP7_75t_L g363 ( .A1(n_334), .A2(n_302), .B(n_277), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_332), .A2(n_312), .B(n_277), .Y(n_364) );
A2O1A1Ixp33_ASAP7_75t_L g365 ( .A1(n_326), .A2(n_277), .B(n_274), .C(n_272), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_335), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_337), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_317), .B(n_277), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_314), .B(n_274), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_337), .B(n_274), .Y(n_370) );
AOI21x1_ASAP7_75t_L g371 ( .A1(n_364), .A2(n_331), .B(n_333), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_345), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_363), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_363), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_345), .Y(n_375) );
AND2x2_ASAP7_75t_L g376 ( .A(n_352), .B(n_335), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_352), .Y(n_377) );
BUFx4f_ASAP7_75t_SL g378 ( .A(n_343), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_363), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_357), .Y(n_380) );
INVxp67_ASAP7_75t_SL g381 ( .A(n_369), .Y(n_381) );
OA21x2_ASAP7_75t_L g382 ( .A1(n_364), .A2(n_333), .B(n_332), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_363), .Y(n_383) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_358), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_357), .B(n_331), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_363), .Y(n_386) );
OR2x2_ASAP7_75t_L g387 ( .A(n_355), .B(n_336), .Y(n_387) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_367), .B(n_331), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_367), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_364), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_370), .B(n_331), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_353), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_355), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_353), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_353), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_353), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_346), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_360), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_346), .Y(n_401) );
OAI21x1_ASAP7_75t_L g402 ( .A1(n_344), .A2(n_340), .B(n_322), .Y(n_402) );
BUFx2_ASAP7_75t_L g403 ( .A(n_369), .Y(n_403) );
AOI21x1_ASAP7_75t_L g404 ( .A1(n_344), .A2(n_328), .B(n_336), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_346), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_369), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_370), .B(n_329), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_360), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_370), .B(n_329), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_356), .B(n_329), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_362), .B(n_272), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_354), .A2(n_50), .B(n_64), .Y(n_414) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_361), .B(n_324), .Y(n_415) );
BUFx3_ASAP7_75t_L g416 ( .A(n_350), .Y(n_416) );
OAI21x1_ASAP7_75t_L g417 ( .A1(n_344), .A2(n_65), .B(n_67), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_341), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_341), .Y(n_419) );
OA21x2_ASAP7_75t_L g420 ( .A1(n_354), .A2(n_70), .B(n_71), .Y(n_420) );
OR2x6_ASAP7_75t_L g421 ( .A(n_365), .B(n_72), .Y(n_421) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_356), .Y(n_422) );
OR2x2_ASAP7_75t_L g423 ( .A(n_422), .B(n_356), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_408), .B(n_351), .Y(n_424) );
BUFx8_ASAP7_75t_L g425 ( .A(n_388), .Y(n_425) );
OA21x2_ASAP7_75t_L g426 ( .A1(n_402), .A2(n_347), .B(n_349), .Y(n_426) );
AOI22xp33_ASAP7_75t_SL g427 ( .A1(n_378), .A2(n_342), .B1(n_350), .B2(n_361), .Y(n_427) );
HB1xp67_ASAP7_75t_L g428 ( .A(n_384), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_416), .B(n_343), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_390), .B(n_362), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_390), .B(n_362), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_413), .A2(n_350), .B1(n_368), .B2(n_342), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_413), .B(n_342), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_379), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_372), .B(n_368), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_372), .Y(n_436) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_384), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_422), .B(n_351), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_375), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_375), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_377), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_379), .Y(n_442) );
AOI22xp5_ASAP7_75t_L g443 ( .A1(n_413), .A2(n_343), .B1(n_342), .B2(n_341), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_379), .Y(n_445) );
OR2x2_ASAP7_75t_L g446 ( .A(n_416), .B(n_366), .Y(n_446) );
AO31x2_ASAP7_75t_L g447 ( .A1(n_399), .A2(n_348), .A3(n_351), .B(n_347), .Y(n_447) );
INVx3_ASAP7_75t_SL g448 ( .A(n_378), .Y(n_448) );
INVx3_ASAP7_75t_L g449 ( .A(n_373), .Y(n_449) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_402), .A2(n_347), .B(n_349), .Y(n_450) );
AND2x6_ASAP7_75t_L g451 ( .A(n_373), .B(n_366), .Y(n_451) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_409), .B(n_411), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_373), .Y(n_453) );
OR2x2_ASAP7_75t_L g454 ( .A(n_394), .B(n_351), .Y(n_454) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_394), .Y(n_455) );
AOI22xp5_ASAP7_75t_L g456 ( .A1(n_415), .A2(n_366), .B1(n_341), .B2(n_348), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_408), .B(n_341), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_377), .B(n_366), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_374), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_408), .B(n_366), .Y(n_460) );
INVx2_ASAP7_75t_SL g461 ( .A(n_388), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_374), .Y(n_462) );
INVx2_ASAP7_75t_SL g463 ( .A(n_388), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_416), .B(n_359), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_403), .B(n_359), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_380), .B(n_359), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_374), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_383), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_383), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_403), .B(n_349), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_383), .Y(n_471) );
HB1xp67_ASAP7_75t_L g472 ( .A(n_394), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_386), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_403), .B(n_73), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g475 ( .A1(n_416), .A2(n_76), .B1(n_79), .B2(n_80), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_386), .Y(n_476) );
INVx2_ASAP7_75t_L g477 ( .A(n_386), .Y(n_477) );
A2O1A1Ixp33_ASAP7_75t_L g478 ( .A1(n_412), .A2(n_82), .B(n_84), .C(n_86), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_380), .B(n_87), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_392), .B(n_88), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_392), .Y(n_481) );
INVxp67_ASAP7_75t_L g482 ( .A(n_415), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_395), .B(n_89), .Y(n_483) );
INVx3_ASAP7_75t_L g484 ( .A(n_421), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_392), .B(n_90), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_389), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_381), .B(n_91), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_376), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_376), .Y(n_489) );
BUFx2_ASAP7_75t_L g490 ( .A(n_409), .Y(n_490) );
AND2x4_ASAP7_75t_L g491 ( .A(n_419), .B(n_92), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_381), .B(n_93), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_385), .B(n_94), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_385), .B(n_97), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_395), .B(n_102), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_376), .Y(n_496) );
AND2x4_ASAP7_75t_L g497 ( .A(n_419), .B(n_98), .Y(n_497) );
OA21x2_ASAP7_75t_L g498 ( .A1(n_402), .A2(n_391), .B(n_398), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_387), .B(n_101), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_387), .B(n_99), .Y(n_500) );
INVx3_ASAP7_75t_L g501 ( .A(n_421), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_385), .B(n_100), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_387), .Y(n_503) );
BUFx2_ASAP7_75t_L g504 ( .A(n_409), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_411), .B(n_389), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_389), .B(n_411), .Y(n_506) );
OR2x2_ASAP7_75t_L g507 ( .A(n_412), .B(n_399), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_412), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_399), .B(n_406), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_399), .B(n_418), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_418), .Y(n_511) );
AOI221xp5_ASAP7_75t_L g512 ( .A1(n_401), .A2(n_405), .B1(n_406), .B2(n_407), .C(n_410), .Y(n_512) );
HB1xp67_ASAP7_75t_L g513 ( .A(n_418), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_418), .B(n_410), .Y(n_514) );
AND2x2_ASAP7_75t_L g515 ( .A(n_506), .B(n_406), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_434), .Y(n_516) );
OR2x2_ASAP7_75t_L g517 ( .A(n_505), .B(n_418), .Y(n_517) );
INVx4_ASAP7_75t_L g518 ( .A(n_448), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_436), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_439), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_434), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_490), .B(n_407), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g523 ( .A(n_503), .B(n_405), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_442), .Y(n_524) );
AND2x4_ASAP7_75t_L g525 ( .A(n_484), .B(n_400), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_504), .B(n_400), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_440), .Y(n_527) );
NOR2xp67_ASAP7_75t_L g528 ( .A(n_461), .B(n_401), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_506), .B(n_401), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_441), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_428), .Y(n_531) );
NOR2xp33_ASAP7_75t_L g532 ( .A(n_482), .B(n_421), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_508), .B(n_405), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_442), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_488), .B(n_398), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_452), .B(n_421), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_452), .B(n_421), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_444), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_423), .B(n_391), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_433), .B(n_421), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_437), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_489), .B(n_496), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_435), .Y(n_543) );
HB1xp67_ASAP7_75t_L g544 ( .A(n_449), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_481), .B(n_382), .Y(n_545) );
AND2x4_ASAP7_75t_SL g546 ( .A(n_461), .B(n_421), .Y(n_546) );
INVx3_ASAP7_75t_L g547 ( .A(n_451), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_423), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_444), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_481), .B(n_382), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_486), .B(n_382), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_486), .B(n_470), .Y(n_552) );
INVx1_ASAP7_75t_SL g553 ( .A(n_448), .Y(n_553) );
OR2x2_ASAP7_75t_L g554 ( .A(n_507), .B(n_391), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_507), .B(n_398), .Y(n_555) );
INVx2_ASAP7_75t_L g556 ( .A(n_445), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_430), .B(n_398), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_470), .B(n_382), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_431), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_455), .B(n_397), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_458), .Y(n_561) );
AND2x4_ASAP7_75t_L g562 ( .A(n_484), .B(n_404), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_433), .B(n_397), .Y(n_563) );
INVx3_ASAP7_75t_L g564 ( .A(n_451), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_472), .Y(n_565) );
NOR2xp67_ASAP7_75t_L g566 ( .A(n_463), .B(n_397), .Y(n_566) );
HB1xp67_ASAP7_75t_L g567 ( .A(n_449), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_463), .B(n_397), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_453), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_453), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_425), .Y(n_571) );
HB1xp67_ASAP7_75t_L g572 ( .A(n_449), .Y(n_572) );
BUFx2_ASAP7_75t_L g573 ( .A(n_425), .Y(n_573) );
NAND4xp25_ASAP7_75t_L g574 ( .A(n_432), .B(n_396), .C(n_393), .D(n_414), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_480), .B(n_420), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_493), .B(n_396), .Y(n_576) );
BUFx2_ASAP7_75t_L g577 ( .A(n_425), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_445), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_446), .B(n_396), .Y(n_579) );
INVx2_ASAP7_75t_L g580 ( .A(n_459), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_493), .B(n_396), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_459), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_462), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_424), .B(n_382), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_424), .B(n_382), .Y(n_585) );
INVx2_ASAP7_75t_L g586 ( .A(n_462), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_467), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_467), .B(n_393), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_494), .B(n_393), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_468), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_480), .B(n_414), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_494), .B(n_414), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_429), .B(n_414), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_468), .Y(n_594) );
BUFx3_ASAP7_75t_L g595 ( .A(n_451), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_484), .B(n_404), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_469), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_485), .B(n_414), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g599 ( .A(n_443), .B(n_414), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_485), .B(n_420), .Y(n_600) );
NAND2xp5_ASAP7_75t_SL g601 ( .A(n_501), .B(n_417), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_469), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_474), .B(n_420), .Y(n_603) );
HB1xp67_ASAP7_75t_L g604 ( .A(n_471), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_471), .B(n_420), .Y(n_605) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_473), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_473), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_476), .Y(n_608) );
INVxp67_ASAP7_75t_R g609 ( .A(n_474), .Y(n_609) );
INVx1_ASAP7_75t_SL g610 ( .A(n_502), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_457), .B(n_371), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_476), .B(n_420), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_427), .B(n_420), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_477), .B(n_417), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_457), .B(n_371), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_477), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_460), .B(n_371), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_509), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_451), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_460), .B(n_404), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_502), .B(n_417), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_509), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_513), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_502), .B(n_487), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_511), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_510), .Y(n_626) );
CKINVDCx16_ASAP7_75t_R g627 ( .A(n_487), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_466), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_465), .B(n_514), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_438), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_438), .Y(n_631) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_492), .B(n_497), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_465), .B(n_492), .Y(n_633) );
O2A1O1Ixp5_ASAP7_75t_SL g634 ( .A1(n_531), .A2(n_501), .B(n_495), .C(n_483), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_548), .B(n_454), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_630), .B(n_454), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_629), .B(n_514), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_541), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_519), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_520), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_618), .B(n_464), .Y(n_641) );
NOR2x1_ASAP7_75t_L g642 ( .A(n_518), .B(n_501), .Y(n_642) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_532), .A2(n_478), .B(n_500), .C(n_499), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_527), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_629), .B(n_514), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_631), .B(n_512), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_626), .B(n_447), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_628), .B(n_447), .Y(n_648) );
INVx2_ASAP7_75t_L g649 ( .A(n_604), .Y(n_649) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_604), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_553), .B(n_456), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_618), .B(n_447), .Y(n_652) );
AND2x4_ASAP7_75t_L g653 ( .A(n_595), .B(n_451), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_530), .Y(n_654) );
NOR2xp33_ASAP7_75t_L g655 ( .A(n_573), .B(n_479), .Y(n_655) );
INVx1_ASAP7_75t_L g656 ( .A(n_543), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g657 ( .A1(n_577), .A2(n_478), .B(n_475), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_532), .A2(n_451), .B1(n_491), .B2(n_497), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_552), .B(n_491), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_552), .B(n_491), .Y(n_660) );
AOI221xp5_ASAP7_75t_L g661 ( .A1(n_559), .A2(n_497), .B1(n_447), .B2(n_498), .C(n_426), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_561), .B(n_498), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_565), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_625), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_622), .B(n_563), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_516), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_542), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_595), .B(n_498), .Y(n_668) );
OR2x2_ASAP7_75t_L g669 ( .A(n_622), .B(n_426), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_516), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_623), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_584), .B(n_426), .Y(n_672) );
INVx2_ASAP7_75t_L g673 ( .A(n_521), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_609), .B(n_450), .Y(n_674) );
AND2x2_ASAP7_75t_L g675 ( .A(n_515), .B(n_450), .Y(n_675) );
INVx1_ASAP7_75t_SL g676 ( .A(n_544), .Y(n_676) );
AND2x2_ASAP7_75t_L g677 ( .A(n_515), .B(n_450), .Y(n_677) );
NAND2x1p5_ASAP7_75t_L g678 ( .A(n_518), .B(n_571), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_533), .Y(n_679) );
INVx2_ASAP7_75t_L g680 ( .A(n_521), .Y(n_680) );
AND2x2_ASAP7_75t_L g681 ( .A(n_529), .B(n_627), .Y(n_681) );
NOR2x1_ASAP7_75t_L g682 ( .A(n_518), .B(n_528), .Y(n_682) );
OR2x2_ASAP7_75t_L g683 ( .A(n_529), .B(n_517), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_522), .B(n_526), .Y(n_684) );
AND2x4_ASAP7_75t_L g685 ( .A(n_547), .B(n_564), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_523), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_584), .B(n_585), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_624), .B(n_540), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_568), .Y(n_689) );
INVx1_ASAP7_75t_SL g690 ( .A(n_544), .Y(n_690) );
AND2x2_ASAP7_75t_L g691 ( .A(n_558), .B(n_610), .Y(n_691) );
INVx2_ASAP7_75t_L g692 ( .A(n_524), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_585), .B(n_557), .Y(n_693) );
OR2x2_ASAP7_75t_L g694 ( .A(n_539), .B(n_606), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_606), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g696 ( .A(n_558), .B(n_535), .Y(n_696) );
INVx3_ASAP7_75t_L g697 ( .A(n_547), .Y(n_697) );
AND2x2_ASAP7_75t_L g698 ( .A(n_633), .B(n_536), .Y(n_698) );
INVx4_ASAP7_75t_L g699 ( .A(n_571), .Y(n_699) );
AND2x2_ASAP7_75t_L g700 ( .A(n_537), .B(n_611), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_611), .B(n_615), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_524), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_569), .Y(n_703) );
AND2x2_ASAP7_75t_L g704 ( .A(n_615), .B(n_617), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_570), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_551), .B(n_550), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_617), .B(n_550), .Y(n_707) );
INVx1_ASAP7_75t_SL g708 ( .A(n_567), .Y(n_708) );
OR2x6_ASAP7_75t_L g709 ( .A(n_632), .B(n_619), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_582), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_545), .B(n_551), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_534), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_579), .B(n_554), .Y(n_713) );
INVx1_ASAP7_75t_SL g714 ( .A(n_567), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_545), .B(n_590), .Y(n_715) );
OR2x2_ASAP7_75t_L g716 ( .A(n_555), .B(n_560), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_583), .B(n_597), .Y(n_717) );
OR2x2_ASAP7_75t_L g718 ( .A(n_594), .B(n_616), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g719 ( .A(n_608), .B(n_620), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_534), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_538), .Y(n_721) );
AND2x2_ASAP7_75t_L g722 ( .A(n_632), .B(n_525), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_538), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_549), .Y(n_724) );
NAND2x1p5_ASAP7_75t_L g725 ( .A(n_566), .B(n_564), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_549), .Y(n_726) );
OR2x2_ASAP7_75t_L g727 ( .A(n_556), .B(n_578), .Y(n_727) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_546), .B(n_564), .Y(n_728) );
HB1xp67_ASAP7_75t_L g729 ( .A(n_572), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_556), .B(n_578), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_580), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_525), .B(n_621), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_525), .B(n_572), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_580), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_586), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_593), .B(n_602), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_546), .A2(n_613), .B1(n_599), .B2(n_593), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_586), .B(n_607), .Y(n_738) );
INVxp67_ASAP7_75t_L g739 ( .A(n_650), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_639), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_699), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_640), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_679), .B(n_587), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_681), .B(n_547), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_644), .Y(n_745) );
NAND2x1_ASAP7_75t_L g746 ( .A(n_699), .B(n_562), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_654), .Y(n_747) );
OR2x2_ASAP7_75t_L g748 ( .A(n_687), .B(n_581), .Y(n_748) );
INVx1_ASAP7_75t_L g749 ( .A(n_656), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_664), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_671), .Y(n_751) );
OR2x6_ASAP7_75t_L g752 ( .A(n_709), .B(n_562), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_732), .B(n_599), .Y(n_753) );
INVx1_ASAP7_75t_L g754 ( .A(n_665), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_689), .Y(n_755) );
INVx1_ASAP7_75t_L g756 ( .A(n_638), .Y(n_756) );
NOR3xp33_ASAP7_75t_L g757 ( .A(n_657), .B(n_574), .C(n_613), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_684), .B(n_562), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_719), .Y(n_759) );
INVx2_ASAP7_75t_SL g760 ( .A(n_678), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_719), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_686), .B(n_607), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_687), .B(n_576), .Y(n_763) );
INVx2_ASAP7_75t_L g764 ( .A(n_650), .Y(n_764) );
AND2x2_ASAP7_75t_L g765 ( .A(n_700), .B(n_596), .Y(n_765) );
NOR2xp33_ASAP7_75t_L g766 ( .A(n_667), .B(n_589), .Y(n_766) );
AND2x2_ASAP7_75t_L g767 ( .A(n_637), .B(n_596), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g768 ( .A(n_646), .B(n_587), .Y(n_768) );
INVx1_ASAP7_75t_SL g769 ( .A(n_676), .Y(n_769) );
AOI32xp33_ASAP7_75t_L g770 ( .A1(n_682), .A2(n_603), .A3(n_600), .B1(n_591), .B2(n_598), .Y(n_770) );
INVx1_ASAP7_75t_L g771 ( .A(n_663), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_717), .Y(n_772) );
AND2x2_ASAP7_75t_L g773 ( .A(n_645), .B(n_596), .Y(n_773) );
INVxp67_ASAP7_75t_L g774 ( .A(n_651), .Y(n_774) );
INVx1_ASAP7_75t_L g775 ( .A(n_717), .Y(n_775) );
INVx1_ASAP7_75t_L g776 ( .A(n_683), .Y(n_776) );
INVx1_ASAP7_75t_L g777 ( .A(n_718), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_701), .B(n_575), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_703), .Y(n_779) );
NAND2xp33_ASAP7_75t_L g780 ( .A(n_678), .B(n_642), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_704), .B(n_602), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_655), .B(n_588), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_705), .Y(n_783) );
OR2x2_ASAP7_75t_L g784 ( .A(n_693), .B(n_696), .Y(n_784) );
INVx2_ASAP7_75t_L g785 ( .A(n_694), .Y(n_785) );
NAND2xp5_ASAP7_75t_SL g786 ( .A(n_668), .B(n_592), .Y(n_786) );
HB1xp67_ASAP7_75t_L g787 ( .A(n_729), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_646), .B(n_605), .Y(n_788) );
INVx2_ASAP7_75t_L g789 ( .A(n_735), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_647), .B(n_612), .Y(n_790) );
NOR5xp2_ASAP7_75t_L g791 ( .A(n_657), .B(n_601), .C(n_614), .D(n_729), .E(n_735), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_710), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_715), .Y(n_793) );
O2A1O1Ixp33_ASAP7_75t_L g794 ( .A1(n_643), .A2(n_601), .B(n_647), .C(n_648), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_715), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_716), .Y(n_796) );
AND2x2_ASAP7_75t_L g797 ( .A(n_707), .B(n_691), .Y(n_797) );
INVx2_ASAP7_75t_L g798 ( .A(n_649), .Y(n_798) );
AND2x4_ASAP7_75t_L g799 ( .A(n_685), .B(n_697), .Y(n_799) );
INVx2_ASAP7_75t_SL g800 ( .A(n_713), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_693), .B(n_672), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_672), .B(n_648), .Y(n_802) );
OR2x2_ASAP7_75t_L g803 ( .A(n_696), .B(n_706), .Y(n_803) );
AOI222xp33_ASAP7_75t_L g804 ( .A1(n_774), .A2(n_737), .B1(n_736), .B2(n_677), .C1(n_675), .C2(n_636), .Y(n_804) );
NOR2xp67_ASAP7_75t_L g805 ( .A(n_760), .B(n_697), .Y(n_805) );
AOI21xp33_ASAP7_75t_L g806 ( .A1(n_794), .A2(n_737), .B(n_662), .Y(n_806) );
XNOR2xp5_ASAP7_75t_L g807 ( .A(n_741), .B(n_698), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_772), .Y(n_808) );
NOR2xp33_ASAP7_75t_L g809 ( .A(n_800), .B(n_688), .Y(n_809) );
OAI31xp33_ASAP7_75t_L g810 ( .A1(n_757), .A2(n_674), .A3(n_725), .B(n_668), .Y(n_810) );
OAI21xp33_ASAP7_75t_SL g811 ( .A1(n_752), .A2(n_709), .B(n_728), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_752), .A2(n_658), .B1(n_709), .B2(n_725), .Y(n_812) );
NOR2xp67_ASAP7_75t_SL g813 ( .A(n_780), .B(n_722), .Y(n_813) );
INVx1_ASAP7_75t_SL g814 ( .A(n_797), .Y(n_814) );
INVxp67_ASAP7_75t_L g815 ( .A(n_787), .Y(n_815) );
HB1xp67_ASAP7_75t_L g816 ( .A(n_739), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g817 ( .A(n_788), .B(n_711), .Y(n_817) );
NAND2xp5_ASAP7_75t_L g818 ( .A(n_802), .B(n_662), .Y(n_818) );
HB1xp67_ASAP7_75t_L g819 ( .A(n_739), .Y(n_819) );
INVx2_ASAP7_75t_L g820 ( .A(n_789), .Y(n_820) );
AO22x1_ASAP7_75t_L g821 ( .A1(n_799), .A2(n_653), .B1(n_685), .B2(n_660), .Y(n_821) );
NAND2xp5_ASAP7_75t_SL g822 ( .A(n_794), .B(n_653), .Y(n_822) );
OAI33xp33_ASAP7_75t_L g823 ( .A1(n_802), .A2(n_636), .A3(n_635), .B1(n_706), .B2(n_652), .B3(n_669), .Y(n_823) );
INVx1_ASAP7_75t_L g824 ( .A(n_775), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g825 ( .A(n_788), .B(n_733), .Y(n_825) );
OR2x2_ASAP7_75t_L g826 ( .A(n_801), .B(n_641), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g827 ( .A1(n_752), .A2(n_659), .B1(n_708), .B2(n_714), .Y(n_827) );
INVx2_ASAP7_75t_L g828 ( .A(n_764), .Y(n_828) );
NAND3xp33_ASAP7_75t_L g829 ( .A(n_791), .B(n_634), .C(n_661), .Y(n_829) );
INVx1_ASAP7_75t_L g830 ( .A(n_759), .Y(n_830) );
AOI32xp33_ASAP7_75t_L g831 ( .A1(n_758), .A2(n_714), .A3(n_708), .B1(n_676), .B2(n_690), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_761), .Y(n_832) );
NOR4xp25_ASAP7_75t_L g833 ( .A(n_769), .B(n_661), .C(n_690), .D(n_695), .Y(n_833) );
NAND3xp33_ASAP7_75t_L g834 ( .A(n_791), .B(n_726), .C(n_723), .Y(n_834) );
OR2x2_ASAP7_75t_L g835 ( .A(n_801), .B(n_730), .Y(n_835) );
O2A1O1Ixp33_ASAP7_75t_SL g836 ( .A1(n_746), .A2(n_727), .B(n_720), .C(n_724), .Y(n_836) );
OA21x2_ASAP7_75t_L g837 ( .A1(n_768), .A2(n_731), .B(n_670), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_768), .Y(n_838) );
OAI22xp33_ASAP7_75t_L g839 ( .A1(n_784), .A2(n_666), .B1(n_673), .B2(n_680), .Y(n_839) );
AOI221xp5_ASAP7_75t_L g840 ( .A1(n_823), .A2(n_766), .B1(n_782), .B2(n_796), .C(n_755), .Y(n_840) );
OAI21x1_ASAP7_75t_L g841 ( .A1(n_822), .A2(n_786), .B(n_756), .Y(n_841) );
AOI21xp33_ASAP7_75t_SL g842 ( .A1(n_811), .A2(n_770), .B(n_799), .Y(n_842) );
AOI22xp5_ASAP7_75t_L g843 ( .A1(n_804), .A2(n_753), .B1(n_754), .B2(n_793), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g844 ( .A(n_838), .B(n_795), .Y(n_844) );
AOI21xp5_ASAP7_75t_L g845 ( .A1(n_836), .A2(n_762), .B(n_743), .Y(n_845) );
AOI22xp5_ASAP7_75t_L g846 ( .A1(n_812), .A2(n_777), .B1(n_776), .B2(n_744), .Y(n_846) );
AOI21xp5_ASAP7_75t_SL g847 ( .A1(n_812), .A2(n_749), .B(n_792), .Y(n_847) );
AOI221xp5_ASAP7_75t_L g848 ( .A1(n_806), .A2(n_751), .B1(n_771), .B2(n_750), .C(n_742), .Y(n_848) );
AND2x2_ASAP7_75t_L g849 ( .A(n_821), .B(n_765), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_806), .B(n_803), .Y(n_850) );
INVxp67_ASAP7_75t_L g851 ( .A(n_816), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_819), .B(n_790), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_835), .Y(n_853) );
INVx2_ASAP7_75t_L g854 ( .A(n_837), .Y(n_854) );
INVx1_ASAP7_75t_L g855 ( .A(n_808), .Y(n_855) );
NAND2xp5_ASAP7_75t_SL g856 ( .A(n_833), .B(n_769), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g857 ( .A1(n_810), .A2(n_740), .B1(n_747), .B2(n_745), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_824), .Y(n_858) );
AOI322xp5_ASAP7_75t_L g859 ( .A1(n_850), .A2(n_814), .A3(n_809), .B1(n_817), .B2(n_825), .C1(n_839), .C2(n_815), .Y(n_859) );
NAND2xp5_ASAP7_75t_L g860 ( .A(n_848), .B(n_832), .Y(n_860) );
AOI211xp5_ASAP7_75t_L g861 ( .A1(n_847), .A2(n_813), .B(n_829), .C(n_827), .Y(n_861) );
AOI321xp33_ASAP7_75t_L g862 ( .A1(n_856), .A2(n_827), .A3(n_818), .B1(n_830), .B2(n_785), .C(n_790), .Y(n_862) );
OAI21xp33_ASAP7_75t_L g863 ( .A1(n_846), .A2(n_831), .B(n_818), .Y(n_863) );
AOI211x1_ASAP7_75t_L g864 ( .A1(n_856), .A2(n_834), .B(n_767), .C(n_773), .Y(n_864) );
OAI21xp33_ASAP7_75t_L g865 ( .A1(n_857), .A2(n_807), .B(n_826), .Y(n_865) );
NAND2xp5_ASAP7_75t_L g866 ( .A(n_840), .B(n_837), .Y(n_866) );
OAI211xp5_ASAP7_75t_L g867 ( .A1(n_842), .A2(n_805), .B(n_762), .C(n_743), .Y(n_867) );
NAND4xp75_ASAP7_75t_L g868 ( .A(n_843), .B(n_779), .C(n_783), .D(n_778), .Y(n_868) );
INVx1_ASAP7_75t_SL g869 ( .A(n_866), .Y(n_869) );
NOR2xp33_ASAP7_75t_SL g870 ( .A(n_865), .B(n_849), .Y(n_870) );
NAND2xp5_ASAP7_75t_SL g871 ( .A(n_861), .B(n_857), .Y(n_871) );
NOR2xp33_ASAP7_75t_L g872 ( .A(n_867), .B(n_851), .Y(n_872) );
NOR2x1_ASAP7_75t_L g873 ( .A(n_868), .B(n_854), .Y(n_873) );
OAI221xp5_ASAP7_75t_L g874 ( .A1(n_870), .A2(n_862), .B1(n_859), .B2(n_863), .C(n_860), .Y(n_874) );
NAND4xp75_ASAP7_75t_L g875 ( .A(n_871), .B(n_864), .C(n_845), .D(n_854), .Y(n_875) );
NOR3xp33_ASAP7_75t_L g876 ( .A(n_869), .B(n_841), .C(n_852), .Y(n_876) );
NAND2x1p5_ASAP7_75t_L g877 ( .A(n_875), .B(n_873), .Y(n_877) );
OAI31xp33_ASAP7_75t_L g878 ( .A1(n_874), .A2(n_872), .A3(n_853), .B(n_855), .Y(n_878) );
AOI21xp5_ASAP7_75t_L g879 ( .A1(n_876), .A2(n_844), .B(n_858), .Y(n_879) );
XOR2xp5_ASAP7_75t_L g880 ( .A(n_877), .B(n_748), .Y(n_880) );
XNOR2x1_ASAP7_75t_L g881 ( .A(n_878), .B(n_828), .Y(n_881) );
AND2x2_ASAP7_75t_L g882 ( .A(n_881), .B(n_879), .Y(n_882) );
NAND2xp5_ASAP7_75t_L g883 ( .A(n_880), .B(n_820), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_882), .B(n_798), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_884), .A2(n_883), .B(n_763), .Y(n_885) );
OAI21xp5_ASAP7_75t_L g886 ( .A1(n_885), .A2(n_781), .B(n_738), .Y(n_886) );
OR2x6_ASAP7_75t_L g887 ( .A(n_886), .B(n_734), .Y(n_887) );
OR2x6_ASAP7_75t_L g888 ( .A(n_887), .B(n_692), .Y(n_888) );
AOI22xp33_ASAP7_75t_L g889 ( .A1(n_888), .A2(n_702), .B1(n_712), .B2(n_721), .Y(n_889) );
endmodule