module fake_ariane_1014_n_1041 (n_83, n_8, n_56, n_60, n_170, n_190, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_195, n_38, n_213, n_47, n_110, n_153, n_18, n_197, n_221, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_203, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_205, n_71, n_24, n_7, n_109, n_208, n_96, n_156, n_209, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_210, n_147, n_204, n_200, n_51, n_166, n_76, n_218, n_103, n_79, n_26, n_3, n_46, n_220, n_0, n_84, n_36, n_199, n_91, n_159, n_107, n_189, n_72, n_105, n_128, n_217, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_201, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_214, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_212, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_198, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_196, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_206, n_13, n_27, n_207, n_29, n_41, n_219, n_140, n_55, n_191, n_151, n_136, n_192, n_28, n_80, n_146, n_211, n_194, n_97, n_154, n_215, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_202, n_145, n_78, n_193, n_39, n_59, n_63, n_99, n_216, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1041);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_190;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_195;
input n_38;
input n_213;
input n_47;
input n_110;
input n_153;
input n_18;
input n_197;
input n_221;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_203;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_205;
input n_71;
input n_24;
input n_7;
input n_109;
input n_208;
input n_96;
input n_156;
input n_209;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_210;
input n_147;
input n_204;
input n_200;
input n_51;
input n_166;
input n_76;
input n_218;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_220;
input n_0;
input n_84;
input n_36;
input n_199;
input n_91;
input n_159;
input n_107;
input n_189;
input n_72;
input n_105;
input n_128;
input n_217;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_201;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_214;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_198;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_196;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_206;
input n_13;
input n_27;
input n_207;
input n_29;
input n_41;
input n_219;
input n_140;
input n_55;
input n_191;
input n_151;
input n_136;
input n_192;
input n_28;
input n_80;
input n_146;
input n_211;
input n_194;
input n_97;
input n_154;
input n_215;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_202;
input n_145;
input n_78;
input n_193;
input n_39;
input n_59;
input n_63;
input n_99;
input n_216;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1041;

wire n_295;
wire n_356;
wire n_556;
wire n_698;
wire n_695;
wire n_913;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_1008;
wire n_581;
wire n_294;
wire n_1020;
wire n_646;
wire n_640;
wire n_463;
wire n_1024;
wire n_830;
wire n_691;
wire n_404;
wire n_943;
wire n_678;
wire n_651;
wire n_987;
wire n_936;
wire n_347;
wire n_423;
wire n_961;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_1036;
wire n_564;
wire n_610;
wire n_752;
wire n_341;
wire n_1029;
wire n_985;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_969;
wire n_283;
wire n_919;
wire n_525;
wire n_806;
wire n_367;
wire n_970;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_952;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_940;
wire n_346;
wire n_1016;
wire n_764;
wire n_979;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_949;
wire n_956;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_232;
wire n_441;
wire n_568;
wire n_1032;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_960;
wire n_520;
wire n_980;
wire n_870;
wire n_714;
wire n_279;
wire n_958;
wire n_702;
wire n_905;
wire n_945;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_968;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_1009;
wire n_230;
wire n_270;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_995;
wire n_285;
wire n_473;
wire n_801;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_1018;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_953;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_1003;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_989;
wire n_331;
wire n_320;
wire n_309;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_1035;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_840;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_795;
wire n_398;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_507;
wire n_486;
wire n_465;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_971;
wire n_369;
wire n_240;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_323;
wire n_550;
wire n_1023;
wire n_988;
wire n_635;
wire n_707;
wire n_997;
wire n_330;
wire n_914;
wire n_400;
wire n_694;
wire n_689;
wire n_884;
wire n_983;
wire n_282;
wire n_328;
wire n_368;
wire n_1034;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_301;
wire n_248;
wire n_467;
wire n_432;
wire n_545;
wire n_1015;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_352;
wire n_538;
wire n_920;
wire n_899;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_1013;
wire n_986;
wire n_638;
wire n_334;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_1039;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_612;
wire n_449;
wire n_413;
wire n_392;
wire n_376;
wire n_957;
wire n_977;
wire n_512;
wire n_715;
wire n_889;
wire n_935;
wire n_579;
wire n_844;
wire n_1012;
wire n_459;
wire n_685;
wire n_321;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_950;
wire n_1017;
wire n_711;
wire n_877;
wire n_1021;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_617;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_942;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_490;
wire n_262;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_1006;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_1019;
wire n_297;
wire n_962;
wire n_662;
wire n_641;
wire n_1005;
wire n_503;
wire n_941;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_772;
wire n_747;
wire n_741;
wire n_847;
wire n_939;
wire n_371;
wire n_845;
wire n_888;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_676;
wire n_708;
wire n_551;
wire n_308;
wire n_417;
wire n_1038;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_993;
wire n_380;
wire n_948;
wire n_582;
wire n_284;
wire n_922;
wire n_1004;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_1022;
wire n_1033;
wire n_896;
wire n_409;
wire n_947;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_1031;
wire n_468;
wire n_853;
wire n_526;
wire n_742;
wire n_716;
wire n_696;
wire n_1040;
wire n_674;
wire n_482;
wire n_316;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_954;
wire n_912;
wire n_476;
wire n_460;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_762;
wire n_744;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_982;
wire n_915;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_966;
wire n_992;
wire n_298;
wire n_955;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_984;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_991;
wire n_389;
wire n_1007;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_606;
wire n_951;
wire n_1026;
wire n_938;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_509;
wire n_583;
wire n_1014;
wire n_724;
wire n_306;
wire n_666;
wire n_1000;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_378;
wire n_436;
wire n_946;
wire n_757;
wire n_375;
wire n_324;
wire n_1030;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_967;
wire n_998;
wire n_999;
wire n_472;
wire n_937;
wire n_296;
wire n_265;
wire n_746;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_751;
wire n_615;
wire n_1027;
wire n_996;
wire n_521;
wire n_963;
wire n_873;
wire n_496;
wire n_739;
wire n_1028;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_1001;
wire n_824;
wire n_428;
wire n_1002;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_959;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_975;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_1037;
wire n_981;
wire n_1010;
wire n_882;
wire n_990;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_944;
wire n_749;
wire n_994;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_973;
wire n_523;
wire n_268;
wire n_972;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_876;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_976;
wire n_353;
wire n_767;
wire n_736;
wire n_1025;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_964;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_978;
wire n_642;
wire n_1011;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_974;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_965;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_934;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g222 ( 
.A(n_7),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g223 ( 
.A(n_87),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_203),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_215),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_113),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_56),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_193),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_79),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_43),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_186),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_33),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_96),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_14),
.Y(n_235)
);

INVxp67_ASAP7_75t_SL g236 ( 
.A(n_154),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_64),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_46),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_149),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_135),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_107),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_108),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_125),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_72),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_75),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_38),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_208),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_77),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_67),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_73),
.Y(n_253)
);

BUFx5_ASAP7_75t_L g254 ( 
.A(n_98),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_51),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_30),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_153),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_70),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_83),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_148),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_204),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_117),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_205),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_30),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_189),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_27),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_168),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_90),
.Y(n_272)
);

BUFx10_ASAP7_75t_L g273 ( 
.A(n_185),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_88),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_167),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_176),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_170),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_3),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_171),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_210),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_211),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_158),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_196),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_38),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_44),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_60),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_220),
.Y(n_287)
);

INVx2_ASAP7_75t_SL g288 ( 
.A(n_18),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_213),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g290 ( 
.A(n_40),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_146),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_78),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_155),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_28),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_99),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_198),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_104),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_18),
.Y(n_298)
);

BUFx8_ASAP7_75t_SL g299 ( 
.A(n_54),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_80),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_2),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_207),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_136),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_201),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_0),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_97),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_82),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_53),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_48),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_95),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_165),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_36),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_214),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_23),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g315 ( 
.A(n_124),
.Y(n_315)
);

BUFx10_ASAP7_75t_L g316 ( 
.A(n_157),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_6),
.Y(n_317)
);

BUFx3_ASAP7_75t_L g318 ( 
.A(n_20),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_132),
.Y(n_319)
);

NAND2xp33_ASAP7_75t_R g320 ( 
.A(n_228),
.B(n_45),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_223),
.B(n_0),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_284),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_266),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_266),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_269),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_318),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_269),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_283),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_318),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_222),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_247),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_227),
.Y(n_333)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_312),
.Y(n_334)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_224),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_315),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_258),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_277),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_278),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_299),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_299),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_241),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_235),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_241),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_294),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_277),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_301),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_224),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g350 ( 
.A(n_249),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_229),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_224),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_225),
.B(n_231),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_238),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_233),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_232),
.B(n_1),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_226),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g359 ( 
.A(n_300),
.B(n_1),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_226),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_226),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_273),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_273),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_273),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_316),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_316),
.Y(n_366)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_267),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_316),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_270),
.Y(n_369)
);

XNOR2x1_ASAP7_75t_L g370 ( 
.A(n_290),
.B(n_298),
.Y(n_370)
);

NOR2xp67_ASAP7_75t_L g371 ( 
.A(n_305),
.B(n_2),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_243),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_317),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_250),
.Y(n_374)
);

INVxp33_ASAP7_75t_L g375 ( 
.A(n_227),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_256),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_324),
.B(n_3),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_342),
.B(n_260),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_333),
.Y(n_381)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_372),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_325),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_374),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_376),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_326),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_335),
.B(n_375),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_359),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_357),
.Y(n_389)
);

HB1xp67_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_340),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_331),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_332),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_359),
.B(n_260),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_353),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_340),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_335),
.B(n_263),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_341),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_345),
.Y(n_401)
);

BUFx8_ASAP7_75t_L g402 ( 
.A(n_358),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_341),
.Y(n_403)
);

XNOR2x2_ASAP7_75t_L g404 ( 
.A(n_370),
.B(n_293),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_328),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_351),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_354),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_349),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_321),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_323),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_338),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_327),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_330),
.Y(n_415)
);

INVxp33_ASAP7_75t_L g416 ( 
.A(n_343),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_377),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_369),
.Y(n_418)
);

BUFx3_ASAP7_75t_L g419 ( 
.A(n_360),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_R g420 ( 
.A(n_342),
.B(n_319),
.Y(n_420)
);

NOR2xp67_ASAP7_75t_L g421 ( 
.A(n_362),
.B(n_234),
.Y(n_421)
);

AND2x4_ASAP7_75t_L g422 ( 
.A(n_363),
.B(n_264),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_355),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_322),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_364),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_365),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_346),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_366),
.B(n_271),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_346),
.Y(n_429)
);

AND2x2_ASAP7_75t_L g430 ( 
.A(n_368),
.B(n_276),
.Y(n_430)
);

HB1xp67_ASAP7_75t_L g431 ( 
.A(n_369),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_356),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_329),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_371),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_344),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_423),
.Y(n_437)
);

INVx1_ASAP7_75t_SL g438 ( 
.A(n_383),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_414),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_387),
.B(n_344),
.Y(n_440)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_425),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_410),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_414),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_412),
.Y(n_444)
);

NAND2x1p5_ASAP7_75t_L g445 ( 
.A(n_436),
.B(n_292),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_386),
.Y(n_446)
);

NOR2x1p5_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_329),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_348),
.Y(n_448)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_425),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_411),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_389),
.B(n_336),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_395),
.B(n_348),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_411),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_410),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_395),
.B(n_352),
.Y(n_455)
);

INVx4_ASAP7_75t_SL g456 ( 
.A(n_394),
.Y(n_456)
);

INVx4_ASAP7_75t_L g457 ( 
.A(n_425),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_425),
.B(n_336),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_381),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_381),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_415),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_415),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g463 ( 
.A(n_425),
.B(n_350),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_392),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_412),
.Y(n_465)
);

AO21x2_ASAP7_75t_L g466 ( 
.A1(n_380),
.A2(n_308),
.B(n_303),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_388),
.B(n_352),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_392),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_419),
.B(n_361),
.Y(n_471)
);

INVx6_ASAP7_75t_L g472 ( 
.A(n_412),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_436),
.B(n_350),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_412),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_381),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_393),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_381),
.Y(n_477)
);

BUFx8_ASAP7_75t_SL g478 ( 
.A(n_405),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_378),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_384),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_436),
.B(n_361),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_413),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_378),
.Y(n_483)
);

AND2x4_ASAP7_75t_L g484 ( 
.A(n_419),
.B(n_334),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_406),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_426),
.B(n_373),
.Y(n_486)
);

OR2x2_ASAP7_75t_L g487 ( 
.A(n_417),
.B(n_373),
.Y(n_487)
);

INVx3_ASAP7_75t_L g488 ( 
.A(n_382),
.Y(n_488)
);

INVx4_ASAP7_75t_SL g489 ( 
.A(n_394),
.Y(n_489)
);

AND2x6_ASAP7_75t_L g490 ( 
.A(n_394),
.B(n_320),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_408),
.Y(n_491)
);

INVx4_ASAP7_75t_L g492 ( 
.A(n_388),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_382),
.Y(n_494)
);

AOI22xp33_ASAP7_75t_L g495 ( 
.A1(n_394),
.A2(n_236),
.B1(n_254),
.B2(n_310),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_385),
.Y(n_496)
);

NAND2x1p5_ASAP7_75t_L g497 ( 
.A(n_388),
.B(n_230),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

AND2x6_ASAP7_75t_L g499 ( 
.A(n_388),
.B(n_254),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_426),
.B(n_424),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_424),
.B(n_237),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_396),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_385),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_400),
.Y(n_504)
);

INVx4_ASAP7_75t_L g505 ( 
.A(n_422),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_398),
.B(n_239),
.Y(n_506)
);

INVx2_ASAP7_75t_SL g507 ( 
.A(n_417),
.Y(n_507)
);

BUFx3_ASAP7_75t_L g508 ( 
.A(n_400),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_422),
.B(n_240),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_422),
.B(n_4),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_434),
.B(n_313),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_401),
.Y(n_512)
);

INVx4_ASAP7_75t_L g513 ( 
.A(n_422),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_471),
.B(n_418),
.Y(n_514)
);

INVx2_ASAP7_75t_SL g515 ( 
.A(n_471),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_505),
.B(n_431),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_500),
.B(n_428),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g518 ( 
.A(n_478),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_500),
.B(n_428),
.Y(n_519)
);

INVxp67_ASAP7_75t_L g520 ( 
.A(n_478),
.Y(n_520)
);

INVx2_ASAP7_75t_L g521 ( 
.A(n_496),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_492),
.B(n_430),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_452),
.B(n_416),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_496),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_484),
.B(n_435),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_492),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_456),
.B(n_430),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_463),
.B(n_435),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_491),
.B(n_391),
.Y(n_529)
);

AND2x4_ASAP7_75t_L g530 ( 
.A(n_456),
.B(n_401),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_463),
.B(n_421),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_455),
.B(n_421),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_459),
.B(n_407),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_482),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_480),
.B(n_420),
.Y(n_535)
);

INVx8_ASAP7_75t_L g536 ( 
.A(n_490),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_459),
.B(n_407),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_496),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_484),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g540 ( 
.A(n_448),
.B(n_427),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_473),
.B(n_429),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_482),
.Y(n_542)
);

OAI22xp5_ASAP7_75t_L g543 ( 
.A1(n_510),
.A2(n_409),
.B1(n_434),
.B2(n_390),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_473),
.B(n_481),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_481),
.B(n_397),
.Y(n_545)
);

AOI21xp5_ASAP7_75t_L g546 ( 
.A1(n_468),
.A2(n_409),
.B(n_244),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_460),
.B(n_402),
.Y(n_547)
);

AOI22xp33_ASAP7_75t_L g548 ( 
.A1(n_490),
.A2(n_495),
.B1(n_404),
.B2(n_493),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_485),
.Y(n_549)
);

NOR2xp33_ASAP7_75t_L g550 ( 
.A(n_451),
.B(n_399),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_456),
.B(n_403),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_483),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g553 ( 
.A1(n_490),
.A2(n_404),
.B1(n_402),
.B2(n_379),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_480),
.B(n_402),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_496),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_505),
.B(n_432),
.Y(n_556)
);

OR2x2_ASAP7_75t_L g557 ( 
.A(n_438),
.B(n_432),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_513),
.B(n_402),
.Y(n_559)
);

AOI22xp5_ASAP7_75t_L g560 ( 
.A1(n_490),
.A2(n_279),
.B1(n_311),
.B2(n_309),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_460),
.B(n_254),
.Y(n_561)
);

AND2x6_ASAP7_75t_L g562 ( 
.A(n_510),
.B(n_254),
.Y(n_562)
);

A2O1A1Ixp33_ASAP7_75t_SL g563 ( 
.A1(n_486),
.A2(n_242),
.B(n_245),
.C(n_246),
.Y(n_563)
);

O2A1O1Ixp33_ASAP7_75t_L g564 ( 
.A1(n_504),
.A2(n_4),
.B(n_5),
.C(n_7),
.Y(n_564)
);

AOI22xp5_ASAP7_75t_L g565 ( 
.A1(n_490),
.A2(n_280),
.B1(n_307),
.B2(n_306),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_451),
.B(n_379),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_488),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_513),
.B(n_248),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_475),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_L g570 ( 
.A(n_440),
.B(n_251),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_493),
.B(n_252),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_508),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_487),
.B(n_5),
.Y(n_573)
);

A2O1A1Ixp33_ASAP7_75t_L g574 ( 
.A1(n_486),
.A2(n_304),
.B(n_302),
.C(n_297),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_446),
.Y(n_575)
);

INVx2_ASAP7_75t_SL g576 ( 
.A(n_437),
.Y(n_576)
);

AND2x4_ASAP7_75t_L g577 ( 
.A(n_489),
.B(n_8),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_508),
.B(n_253),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_501),
.B(n_255),
.Y(n_579)
);

HB1xp67_ASAP7_75t_SL g580 ( 
.A(n_507),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_450),
.Y(n_581)
);

OR2x6_ASAP7_75t_L g582 ( 
.A(n_447),
.B(n_445),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_495),
.A2(n_296),
.B1(n_295),
.B2(n_291),
.Y(n_584)
);

NOR2x2_ASAP7_75t_L g585 ( 
.A(n_479),
.B(n_8),
.Y(n_585)
);

AOI21xp5_ASAP7_75t_L g586 ( 
.A1(n_477),
.A2(n_259),
.B(n_257),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g587 ( 
.A(n_489),
.B(n_9),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_445),
.B(n_261),
.Y(n_588)
);

AOI22xp5_ASAP7_75t_L g589 ( 
.A1(n_458),
.A2(n_289),
.B1(n_287),
.B2(n_286),
.Y(n_589)
);

O2A1O1Ixp5_ASAP7_75t_L g590 ( 
.A1(n_441),
.A2(n_285),
.B(n_282),
.C(n_281),
.Y(n_590)
);

AOI22xp33_ASAP7_75t_L g591 ( 
.A1(n_494),
.A2(n_254),
.B1(n_274),
.B2(n_272),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_494),
.A2(n_254),
.B1(n_268),
.B2(n_265),
.Y(n_592)
);

OAI22xp5_ASAP7_75t_L g593 ( 
.A1(n_497),
.A2(n_275),
.B1(n_262),
.B2(n_11),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_475),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_458),
.A2(n_254),
.B1(n_10),
.B2(n_11),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_503),
.A2(n_9),
.B1(n_10),
.B2(n_12),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_512),
.B(n_12),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_489),
.B(n_13),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_453),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_L g600 ( 
.A(n_540),
.B(n_550),
.C(n_541),
.Y(n_600)
);

CKINVDCx8_ASAP7_75t_R g601 ( 
.A(n_534),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_533),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_R g603 ( 
.A(n_549),
.B(n_442),
.Y(n_603)
);

BUFx6f_ASAP7_75t_L g604 ( 
.A(n_569),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_R g605 ( 
.A(n_542),
.B(n_580),
.Y(n_605)
);

OR2x6_ASAP7_75t_L g606 ( 
.A(n_539),
.B(n_497),
.Y(n_606)
);

OR2x6_ASAP7_75t_L g607 ( 
.A(n_576),
.B(n_442),
.Y(n_607)
);

INVx5_ASAP7_75t_L g608 ( 
.A(n_551),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_517),
.B(n_511),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_552),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_551),
.B(n_527),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_523),
.A2(n_511),
.B1(n_499),
.B2(n_509),
.Y(n_612)
);

AND2x4_ASAP7_75t_L g613 ( 
.A(n_527),
.B(n_454),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_517),
.B(n_499),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_525),
.B(n_461),
.Y(n_615)
);

INVx1_ASAP7_75t_SL g616 ( 
.A(n_575),
.Y(n_616)
);

BUFx4f_ASAP7_75t_L g617 ( 
.A(n_582),
.Y(n_617)
);

NOR2x1_ASAP7_75t_L g618 ( 
.A(n_529),
.B(n_454),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_530),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_533),
.Y(n_620)
);

NOR2xp67_ASAP7_75t_L g621 ( 
.A(n_520),
.B(n_462),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_537),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_557),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_537),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_581),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_519),
.B(n_499),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_519),
.B(n_528),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_582),
.B(n_464),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_544),
.B(n_499),
.Y(n_629)
);

A2O1A1Ixp33_ASAP7_75t_L g630 ( 
.A1(n_545),
.A2(n_469),
.B(n_470),
.C(n_502),
.Y(n_630)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_577),
.Y(n_631)
);

AND3x1_ASAP7_75t_SL g632 ( 
.A(n_585),
.B(n_13),
.C(n_14),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_577),
.B(n_475),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_566),
.B(n_506),
.Y(n_635)
);

INVx3_ASAP7_75t_L g636 ( 
.A(n_530),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_518),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_522),
.B(n_499),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_548),
.B(n_503),
.Y(n_639)
);

AO22x1_ASAP7_75t_L g640 ( 
.A1(n_593),
.A2(n_498),
.B1(n_476),
.B2(n_439),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_582),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_587),
.B(n_475),
.Y(n_642)
);

INVxp67_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_599),
.Y(n_644)
);

BUFx6f_ASAP7_75t_L g645 ( 
.A(n_569),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_558),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_572),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_583),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_536),
.Y(n_650)
);

BUFx2_ASAP7_75t_SL g651 ( 
.A(n_562),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_R g652 ( 
.A(n_556),
.B(n_443),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_570),
.B(n_466),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_593),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_569),
.Y(n_655)
);

BUFx8_ASAP7_75t_L g656 ( 
.A(n_573),
.Y(n_656)
);

BUFx2_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_543),
.Y(n_658)
);

HB1xp67_ASAP7_75t_L g659 ( 
.A(n_543),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_535),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_521),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_561),
.Y(n_663)
);

NOR2x2_ASAP7_75t_L g664 ( 
.A(n_553),
.B(n_467),
.Y(n_664)
);

HB1xp67_ASAP7_75t_L g665 ( 
.A(n_562),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_635),
.B(n_532),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_627),
.B(n_531),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_L g668 ( 
.A1(n_627),
.A2(n_526),
.B1(n_579),
.B2(n_571),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_625),
.Y(n_669)
);

BUFx2_ASAP7_75t_L g670 ( 
.A(n_603),
.Y(n_670)
);

BUFx2_ASAP7_75t_L g671 ( 
.A(n_605),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_653),
.A2(n_561),
.B(n_546),
.Y(n_672)
);

AND2x2_ASAP7_75t_L g673 ( 
.A(n_658),
.B(n_516),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_608),
.Y(n_674)
);

AOI21x1_ASAP7_75t_L g675 ( 
.A1(n_629),
.A2(n_547),
.B(n_474),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_SL g676 ( 
.A(n_629),
.B(n_600),
.Y(n_676)
);

OAI21xp5_ASAP7_75t_L g677 ( 
.A1(n_614),
.A2(n_590),
.B(n_574),
.Y(n_677)
);

NAND3xp33_ASAP7_75t_L g678 ( 
.A(n_654),
.B(n_595),
.C(n_596),
.Y(n_678)
);

AND2x4_ASAP7_75t_L g679 ( 
.A(n_611),
.B(n_608),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_659),
.A2(n_554),
.B1(n_562),
.B2(n_559),
.Y(n_680)
);

CKINVDCx8_ASAP7_75t_R g681 ( 
.A(n_637),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_615),
.B(n_588),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g683 ( 
.A1(n_609),
.A2(n_526),
.B(n_536),
.Y(n_683)
);

INVx2_ASAP7_75t_SL g684 ( 
.A(n_617),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_638),
.A2(n_538),
.B(n_524),
.Y(n_685)
);

OAI21x1_ASAP7_75t_L g686 ( 
.A1(n_638),
.A2(n_555),
.B(n_547),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_608),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_610),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_650),
.Y(n_689)
);

AOI21xp5_ASAP7_75t_L g690 ( 
.A1(n_614),
.A2(n_626),
.B(n_620),
.Y(n_690)
);

AOI21xp5_ASAP7_75t_L g691 ( 
.A1(n_626),
.A2(n_536),
.B(n_568),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_612),
.A2(n_565),
.B(n_560),
.Y(n_692)
);

OAI22xp5_ASAP7_75t_L g693 ( 
.A1(n_602),
.A2(n_578),
.B1(n_594),
.B2(n_584),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_L g694 ( 
.A1(n_622),
.A2(n_562),
.B(n_586),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_611),
.B(n_594),
.Y(n_695)
);

AO21x2_ASAP7_75t_L g696 ( 
.A1(n_639),
.A2(n_563),
.B(n_466),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_663),
.A2(n_564),
.B(n_591),
.Y(n_697)
);

BUFx3_ASAP7_75t_L g698 ( 
.A(n_613),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_SL g699 ( 
.A(n_601),
.B(n_441),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_623),
.B(n_589),
.Y(n_700)
);

AOI21x1_ASAP7_75t_L g701 ( 
.A1(n_640),
.A2(n_465),
.B(n_444),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_639),
.A2(n_592),
.B(n_457),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_623),
.B(n_594),
.Y(n_703)
);

AO31x2_ASAP7_75t_L g704 ( 
.A1(n_630),
.A2(n_457),
.A3(n_449),
.B(n_465),
.Y(n_704)
);

AOI21xp5_ASAP7_75t_L g705 ( 
.A1(n_624),
.A2(n_449),
.B(n_444),
.Y(n_705)
);

OAI21x1_ASAP7_75t_L g706 ( 
.A1(n_662),
.A2(n_465),
.B(n_444),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_660),
.B(n_444),
.Y(n_707)
);

NOR2xp67_ASAP7_75t_SL g708 ( 
.A(n_651),
.B(n_465),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_644),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_646),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_648),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_634),
.A2(n_472),
.B(n_49),
.Y(n_712)
);

OAI21x1_ASAP7_75t_L g713 ( 
.A1(n_661),
.A2(n_618),
.B(n_647),
.Y(n_713)
);

OAI22x1_ASAP7_75t_L g714 ( 
.A1(n_631),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_714)
);

AO21x2_ASAP7_75t_L g715 ( 
.A1(n_652),
.A2(n_472),
.B(n_50),
.Y(n_715)
);

OAI21x1_ASAP7_75t_L g716 ( 
.A1(n_649),
.A2(n_665),
.B(n_636),
.Y(n_716)
);

BUFx6f_ASAP7_75t_L g717 ( 
.A(n_604),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_619),
.Y(n_718)
);

AOI21xp5_ASAP7_75t_L g719 ( 
.A1(n_642),
.A2(n_472),
.B(n_55),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_616),
.B(n_15),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_613),
.Y(n_721)
);

A2O1A1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_642),
.A2(n_16),
.B(n_17),
.C(n_19),
.Y(n_722)
);

INVx3_ASAP7_75t_L g723 ( 
.A(n_717),
.Y(n_723)
);

A2O1A1Ixp33_ASAP7_75t_L g724 ( 
.A1(n_666),
.A2(n_636),
.B(n_619),
.C(n_621),
.Y(n_724)
);

OAI21x1_ASAP7_75t_L g725 ( 
.A1(n_685),
.A2(n_645),
.B(n_604),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_688),
.Y(n_726)
);

OAI21x1_ASAP7_75t_L g727 ( 
.A1(n_685),
.A2(n_645),
.B(n_604),
.Y(n_727)
);

AOI21x1_ASAP7_75t_L g728 ( 
.A1(n_701),
.A2(n_606),
.B(n_657),
.Y(n_728)
);

INVx5_ASAP7_75t_L g729 ( 
.A(n_674),
.Y(n_729)
);

A2O1A1Ixp33_ASAP7_75t_L g730 ( 
.A1(n_666),
.A2(n_617),
.B(n_628),
.C(n_643),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_669),
.Y(n_731)
);

OAI21xp5_ASAP7_75t_L g732 ( 
.A1(n_678),
.A2(n_606),
.B(n_633),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_667),
.A2(n_656),
.B1(n_606),
.B2(n_664),
.Y(n_733)
);

OAI21x1_ASAP7_75t_L g734 ( 
.A1(n_686),
.A2(n_655),
.B(n_645),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_681),
.Y(n_735)
);

INVx5_ASAP7_75t_L g736 ( 
.A(n_674),
.Y(n_736)
);

AO21x1_ASAP7_75t_L g737 ( 
.A1(n_692),
.A2(n_628),
.B(n_650),
.Y(n_737)
);

NOR2xp33_ASAP7_75t_L g738 ( 
.A(n_700),
.B(n_616),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_709),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_681),
.Y(n_740)
);

OAI21x1_ASAP7_75t_L g741 ( 
.A1(n_686),
.A2(n_655),
.B(n_607),
.Y(n_741)
);

INVx3_ASAP7_75t_L g742 ( 
.A(n_717),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_688),
.Y(n_743)
);

OAI21x1_ASAP7_75t_L g744 ( 
.A1(n_672),
.A2(n_655),
.B(n_607),
.Y(n_744)
);

A2O1A1Ixp33_ASAP7_75t_L g745 ( 
.A1(n_722),
.A2(n_641),
.B(n_632),
.C(n_656),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_711),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_703),
.B(n_607),
.Y(n_747)
);

AOI221x1_ASAP7_75t_L g748 ( 
.A1(n_722),
.A2(n_19),
.B1(n_20),
.B2(n_21),
.C(n_22),
.Y(n_748)
);

OAI21x1_ASAP7_75t_SL g749 ( 
.A1(n_690),
.A2(n_694),
.B(n_677),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_SL g750 ( 
.A(n_699),
.B(n_21),
.C(n_22),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_670),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_682),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_752)
);

BUFx2_ASAP7_75t_L g753 ( 
.A(n_698),
.Y(n_753)
);

INVx4_ASAP7_75t_SL g754 ( 
.A(n_679),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_680),
.B(n_24),
.Y(n_755)
);

INVx2_ASAP7_75t_L g756 ( 
.A(n_710),
.Y(n_756)
);

NAND2x1p5_ASAP7_75t_L g757 ( 
.A(n_687),
.B(n_47),
.Y(n_757)
);

AO31x2_ASAP7_75t_L g758 ( 
.A1(n_668),
.A2(n_693),
.A3(n_683),
.B(n_691),
.Y(n_758)
);

INVx1_ASAP7_75t_SL g759 ( 
.A(n_671),
.Y(n_759)
);

OAI21x1_ASAP7_75t_L g760 ( 
.A1(n_672),
.A2(n_131),
.B(n_219),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_710),
.Y(n_761)
);

OAI21xp5_ASAP7_75t_L g762 ( 
.A1(n_676),
.A2(n_25),
.B(n_26),
.Y(n_762)
);

OAI21x1_ASAP7_75t_L g763 ( 
.A1(n_675),
.A2(n_130),
.B(n_218),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_720),
.B(n_26),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_698),
.B(n_27),
.Y(n_765)
);

BUFx12f_ASAP7_75t_L g766 ( 
.A(n_687),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_707),
.Y(n_767)
);

OAI22xp5_ASAP7_75t_L g768 ( 
.A1(n_676),
.A2(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_768)
);

INVx3_ASAP7_75t_SL g769 ( 
.A(n_721),
.Y(n_769)
);

BUFx2_ASAP7_75t_L g770 ( 
.A(n_721),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_673),
.A2(n_29),
.B1(n_31),
.B2(n_32),
.Y(n_771)
);

AO21x1_ASAP7_75t_L g772 ( 
.A1(n_719),
.A2(n_32),
.B(n_33),
.Y(n_772)
);

OAI21x1_ASAP7_75t_L g773 ( 
.A1(n_702),
.A2(n_138),
.B(n_217),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_735),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_756),
.B(n_718),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_764),
.B(n_714),
.Y(n_776)
);

OR2x6_ASAP7_75t_L g777 ( 
.A(n_730),
.B(n_716),
.Y(n_777)
);

AOI22xp33_ASAP7_75t_L g778 ( 
.A1(n_733),
.A2(n_684),
.B1(n_696),
.B2(n_679),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_SL g779 ( 
.A1(n_762),
.A2(n_715),
.B1(n_697),
.B2(n_679),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_731),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_739),
.Y(n_781)
);

OAI22xp5_ASAP7_75t_L g782 ( 
.A1(n_745),
.A2(n_718),
.B1(n_695),
.B2(n_689),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_730),
.B(n_717),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_746),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_756),
.Y(n_785)
);

NAND3xp33_ASAP7_75t_SL g786 ( 
.A(n_745),
.B(n_712),
.C(n_705),
.Y(n_786)
);

OA21x2_ASAP7_75t_L g787 ( 
.A1(n_725),
.A2(n_702),
.B(n_706),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_752),
.A2(n_695),
.B1(n_689),
.B2(n_717),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_761),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_755),
.A2(n_695),
.B1(n_697),
.B2(n_715),
.Y(n_790)
);

BUFx6f_ASAP7_75t_L g791 ( 
.A(n_769),
.Y(n_791)
);

NAND3xp33_ASAP7_75t_SL g792 ( 
.A(n_733),
.B(n_724),
.C(n_771),
.Y(n_792)
);

INVxp33_ASAP7_75t_L g793 ( 
.A(n_738),
.Y(n_793)
);

NAND2xp33_ASAP7_75t_R g794 ( 
.A(n_735),
.B(n_713),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_754),
.B(n_713),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_761),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_726),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_726),
.Y(n_798)
);

AOI222xp33_ASAP7_75t_L g799 ( 
.A1(n_755),
.A2(n_708),
.B1(n_35),
.B2(n_36),
.C1(n_37),
.C2(n_34),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_751),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_743),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_740),
.Y(n_802)
);

INVx5_ASAP7_75t_L g803 ( 
.A(n_766),
.Y(n_803)
);

INVx2_ASAP7_75t_SL g804 ( 
.A(n_751),
.Y(n_804)
);

INVx2_ASAP7_75t_SL g805 ( 
.A(n_740),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_754),
.B(n_716),
.Y(n_806)
);

BUFx2_ASAP7_75t_L g807 ( 
.A(n_753),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_743),
.Y(n_808)
);

AND2x4_ASAP7_75t_L g809 ( 
.A(n_754),
.B(n_706),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_729),
.B(n_704),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_738),
.A2(n_696),
.B1(n_704),
.B2(n_37),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_732),
.A2(n_750),
.B1(n_772),
.B2(n_767),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_747),
.B(n_704),
.Y(n_813)
);

CKINVDCx20_ASAP7_75t_R g814 ( 
.A(n_759),
.Y(n_814)
);

INVx3_ASAP7_75t_L g815 ( 
.A(n_766),
.Y(n_815)
);

AOI21xp5_ASAP7_75t_L g816 ( 
.A1(n_749),
.A2(n_704),
.B(n_35),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_728),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_723),
.Y(n_818)
);

OR2x2_ASAP7_75t_L g819 ( 
.A(n_765),
.B(n_34),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_742),
.Y(n_820)
);

NAND3xp33_ASAP7_75t_SL g821 ( 
.A(n_724),
.B(n_39),
.C(n_40),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_768),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_R g823 ( 
.A(n_769),
.B(n_57),
.Y(n_823)
);

OAI21x1_ASAP7_75t_L g824 ( 
.A1(n_773),
.A2(n_141),
.B(n_216),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_742),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_729),
.B(n_41),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_742),
.Y(n_827)
);

AND2x4_ASAP7_75t_L g828 ( 
.A(n_729),
.B(n_42),
.Y(n_828)
);

OAI22xp5_ASAP7_75t_L g829 ( 
.A1(n_770),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_822),
.A2(n_748),
.B1(n_757),
.B2(n_723),
.Y(n_830)
);

OAI211xp5_ASAP7_75t_L g831 ( 
.A1(n_799),
.A2(n_760),
.B(n_744),
.C(n_736),
.Y(n_831)
);

OAI222xp33_ASAP7_75t_L g832 ( 
.A1(n_788),
.A2(n_757),
.B1(n_736),
.B2(n_729),
.C1(n_737),
.C2(n_758),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_780),
.Y(n_833)
);

AOI22xp33_ASAP7_75t_L g834 ( 
.A1(n_792),
.A2(n_741),
.B1(n_744),
.B2(n_736),
.Y(n_834)
);

CKINVDCx11_ASAP7_75t_R g835 ( 
.A(n_814),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_781),
.Y(n_836)
);

AO21x2_ASAP7_75t_L g837 ( 
.A1(n_816),
.A2(n_773),
.B(n_763),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_800),
.B(n_741),
.Y(n_838)
);

AOI22xp33_ASAP7_75t_SL g839 ( 
.A1(n_788),
.A2(n_763),
.B1(n_760),
.B2(n_736),
.Y(n_839)
);

OAI211xp5_ASAP7_75t_L g840 ( 
.A1(n_799),
.A2(n_734),
.B(n_727),
.C(n_725),
.Y(n_840)
);

INVx3_ASAP7_75t_L g841 ( 
.A(n_810),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_786),
.A2(n_734),
.B(n_727),
.Y(n_842)
);

OR2x6_ASAP7_75t_L g843 ( 
.A(n_777),
.B(n_758),
.Y(n_843)
);

AOI22xp33_ASAP7_75t_L g844 ( 
.A1(n_776),
.A2(n_758),
.B1(n_63),
.B2(n_65),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_784),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_822),
.A2(n_758),
.B1(n_66),
.B2(n_68),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_SL g847 ( 
.A1(n_782),
.A2(n_62),
.B1(n_69),
.B2(n_71),
.Y(n_847)
);

AOI221xp5_ASAP7_75t_L g848 ( 
.A1(n_821),
.A2(n_74),
.B1(n_76),
.B2(n_81),
.C(n_84),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_789),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_785),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_807),
.B(n_793),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_804),
.B(n_85),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_824),
.A2(n_86),
.B(n_89),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_778),
.A2(n_91),
.B1(n_93),
.B2(n_94),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_774),
.Y(n_855)
);

A2O1A1Ixp33_ASAP7_75t_L g856 ( 
.A1(n_790),
.A2(n_100),
.B(n_101),
.C(n_102),
.Y(n_856)
);

AOI21xp33_ASAP7_75t_SL g857 ( 
.A1(n_802),
.A2(n_103),
.B(n_105),
.Y(n_857)
);

AOI221xp5_ASAP7_75t_L g858 ( 
.A1(n_812),
.A2(n_106),
.B1(n_109),
.B2(n_110),
.C(n_111),
.Y(n_858)
);

OAI22xp5_ASAP7_75t_L g859 ( 
.A1(n_779),
.A2(n_112),
.B1(n_114),
.B2(n_115),
.Y(n_859)
);

AOI221x1_ASAP7_75t_SL g860 ( 
.A1(n_829),
.A2(n_828),
.B1(n_826),
.B2(n_782),
.C(n_825),
.Y(n_860)
);

OAI22xp33_ASAP7_75t_L g861 ( 
.A1(n_819),
.A2(n_116),
.B1(n_118),
.B2(n_119),
.Y(n_861)
);

AO31x2_ASAP7_75t_L g862 ( 
.A1(n_817),
.A2(n_120),
.A3(n_121),
.B(n_122),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_818),
.B(n_123),
.Y(n_863)
);

OAI22xp33_ASAP7_75t_L g864 ( 
.A1(n_790),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_813),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_796),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_775),
.B(n_797),
.Y(n_867)
);

OAI33xp33_ASAP7_75t_L g868 ( 
.A1(n_829),
.A2(n_129),
.A3(n_133),
.B1(n_134),
.B2(n_137),
.B3(n_139),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_808),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_775),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_798),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_805),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_801),
.Y(n_873)
);

AOI22xp33_ASAP7_75t_L g874 ( 
.A1(n_811),
.A2(n_140),
.B1(n_142),
.B2(n_143),
.Y(n_874)
);

OAI221xp5_ASAP7_75t_L g875 ( 
.A1(n_783),
.A2(n_144),
.B1(n_145),
.B2(n_147),
.C(n_150),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_803),
.B(n_151),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_849),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_841),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_870),
.B(n_810),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_833),
.B(n_777),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_866),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_835),
.B(n_815),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_838),
.B(n_843),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_836),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_869),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_851),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_845),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_843),
.B(n_787),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_865),
.Y(n_889)
);

AND2x2_ASAP7_75t_L g890 ( 
.A(n_843),
.B(n_787),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_867),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_841),
.B(n_827),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_867),
.Y(n_893)
);

AND2x2_ASAP7_75t_L g894 ( 
.A(n_840),
.B(n_820),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_871),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_850),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_837),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_842),
.B(n_777),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_873),
.Y(n_899)
);

AND2x2_ASAP7_75t_L g900 ( 
.A(n_839),
.B(n_809),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_834),
.B(n_809),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_846),
.B(n_844),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_837),
.Y(n_903)
);

INVx2_ASAP7_75t_L g904 ( 
.A(n_862),
.Y(n_904)
);

OR2x2_ASAP7_75t_L g905 ( 
.A(n_831),
.B(n_815),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_862),
.Y(n_906)
);

AND2x2_ASAP7_75t_L g907 ( 
.A(n_830),
.B(n_826),
.Y(n_907)
);

INVxp67_ASAP7_75t_L g908 ( 
.A(n_830),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_860),
.B(n_828),
.Y(n_909)
);

INVx2_ASAP7_75t_SL g910 ( 
.A(n_876),
.Y(n_910)
);

OAI221xp5_ASAP7_75t_L g911 ( 
.A1(n_908),
.A2(n_859),
.B1(n_858),
.B2(n_856),
.C(n_848),
.Y(n_911)
);

HB1xp67_ASAP7_75t_L g912 ( 
.A(n_889),
.Y(n_912)
);

OR2x2_ASAP7_75t_L g913 ( 
.A(n_889),
.B(n_859),
.Y(n_913)
);

BUFx2_ASAP7_75t_L g914 ( 
.A(n_878),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_884),
.Y(n_915)
);

NAND3xp33_ASAP7_75t_L g916 ( 
.A(n_908),
.B(n_858),
.C(n_848),
.Y(n_916)
);

OAI33xp33_ASAP7_75t_L g917 ( 
.A1(n_893),
.A2(n_861),
.A3(n_864),
.B1(n_794),
.B2(n_868),
.B3(n_832),
.Y(n_917)
);

AO21x2_ASAP7_75t_L g918 ( 
.A1(n_906),
.A2(n_853),
.B(n_875),
.Y(n_918)
);

AOI221xp5_ASAP7_75t_L g919 ( 
.A1(n_894),
.A2(n_875),
.B1(n_857),
.B2(n_874),
.C(n_852),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_882),
.B(n_872),
.Y(n_920)
);

OR2x2_ASAP7_75t_L g921 ( 
.A(n_886),
.B(n_852),
.Y(n_921)
);

BUFx2_ASAP7_75t_L g922 ( 
.A(n_878),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_884),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_909),
.A2(n_847),
.B1(n_854),
.B2(n_791),
.Y(n_924)
);

AOI22xp33_ASAP7_75t_SL g925 ( 
.A1(n_902),
.A2(n_823),
.B1(n_876),
.B2(n_806),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_SL g926 ( 
.A1(n_902),
.A2(n_806),
.B1(n_795),
.B2(n_863),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_891),
.Y(n_927)
);

HB1xp67_ASAP7_75t_L g928 ( 
.A(n_891),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_887),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_886),
.B(n_791),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_930),
.B(n_898),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_930),
.B(n_898),
.Y(n_932)
);

OR2x2_ASAP7_75t_L g933 ( 
.A(n_928),
.B(n_893),
.Y(n_933)
);

NAND2x1_ASAP7_75t_L g934 ( 
.A(n_914),
.B(n_888),
.Y(n_934)
);

AND2x2_ASAP7_75t_L g935 ( 
.A(n_914),
.B(n_922),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_922),
.B(n_888),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_929),
.Y(n_937)
);

AND2x4_ASAP7_75t_L g938 ( 
.A(n_927),
.B(n_888),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_915),
.Y(n_939)
);

AOI221xp5_ASAP7_75t_L g940 ( 
.A1(n_917),
.A2(n_894),
.B1(n_909),
.B2(n_887),
.C(n_903),
.Y(n_940)
);

INVx2_ASAP7_75t_SL g941 ( 
.A(n_912),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_923),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_913),
.B(n_890),
.Y(n_943)
);

AND3x2_ASAP7_75t_L g944 ( 
.A(n_920),
.B(n_907),
.C(n_900),
.Y(n_944)
);

INVx2_ASAP7_75t_SL g945 ( 
.A(n_921),
.Y(n_945)
);

NAND4xp25_ASAP7_75t_L g946 ( 
.A(n_940),
.B(n_916),
.C(n_913),
.D(n_911),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_937),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_937),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_943),
.B(n_907),
.Y(n_949)
);

AOI22xp5_ASAP7_75t_L g950 ( 
.A1(n_944),
.A2(n_919),
.B1(n_924),
.B2(n_925),
.Y(n_950)
);

INVx3_ASAP7_75t_L g951 ( 
.A(n_934),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_941),
.B(n_877),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_933),
.Y(n_953)
);

OR2x2_ASAP7_75t_L g954 ( 
.A(n_953),
.B(n_933),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_947),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_951),
.B(n_949),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_951),
.B(n_943),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_952),
.Y(n_958)
);

INVx3_ASAP7_75t_SL g959 ( 
.A(n_948),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_950),
.Y(n_960)
);

OR2x2_ASAP7_75t_L g961 ( 
.A(n_946),
.B(n_941),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_950),
.B(n_936),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_958),
.B(n_939),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_961),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_954),
.Y(n_965)
);

OAI21xp5_ASAP7_75t_L g966 ( 
.A1(n_962),
.A2(n_905),
.B(n_934),
.Y(n_966)
);

A2O1A1Ixp33_ASAP7_75t_L g967 ( 
.A1(n_960),
.A2(n_905),
.B(n_956),
.C(n_955),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_965),
.B(n_959),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_967),
.A2(n_960),
.B(n_956),
.Y(n_969)
);

AOI221xp5_ASAP7_75t_L g970 ( 
.A1(n_964),
.A2(n_959),
.B1(n_955),
.B2(n_903),
.C(n_897),
.Y(n_970)
);

INVx2_ASAP7_75t_L g971 ( 
.A(n_963),
.Y(n_971)
);

OR2x2_ASAP7_75t_L g972 ( 
.A(n_966),
.B(n_956),
.Y(n_972)
);

OR2x2_ASAP7_75t_L g973 ( 
.A(n_968),
.B(n_957),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_971),
.B(n_939),
.Y(n_974)
);

CKINVDCx20_ASAP7_75t_L g975 ( 
.A(n_969),
.Y(n_975)
);

OAI32xp33_ASAP7_75t_L g976 ( 
.A1(n_972),
.A2(n_939),
.A3(n_936),
.B1(n_921),
.B2(n_935),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_970),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_977),
.B(n_910),
.C(n_897),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_973),
.B(n_855),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_974),
.Y(n_980)
);

NOR3xp33_ASAP7_75t_L g981 ( 
.A(n_975),
.B(n_910),
.C(n_897),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_976),
.B(n_939),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_977),
.B(n_942),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_SL g984 ( 
.A(n_973),
.B(n_935),
.Y(n_984)
);

NOR4xp25_ASAP7_75t_L g985 ( 
.A(n_977),
.B(n_942),
.C(n_945),
.D(n_931),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_980),
.Y(n_986)
);

OAI21xp33_ASAP7_75t_L g987 ( 
.A1(n_985),
.A2(n_938),
.B(n_945),
.Y(n_987)
);

AOI221xp5_ASAP7_75t_L g988 ( 
.A1(n_983),
.A2(n_981),
.B1(n_978),
.B2(n_982),
.C(n_984),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_979),
.A2(n_918),
.B1(n_910),
.B2(n_938),
.Y(n_989)
);

NAND4xp25_ASAP7_75t_L g990 ( 
.A(n_979),
.B(n_938),
.C(n_926),
.D(n_931),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_985),
.B(n_938),
.Y(n_991)
);

AOI22xp5_ASAP7_75t_L g992 ( 
.A1(n_981),
.A2(n_918),
.B1(n_903),
.B2(n_932),
.Y(n_992)
);

AOI211xp5_ASAP7_75t_L g993 ( 
.A1(n_985),
.A2(n_791),
.B(n_903),
.C(n_932),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_986),
.B(n_877),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_991),
.Y(n_995)
);

NOR2x1_ASAP7_75t_L g996 ( 
.A(n_990),
.B(n_803),
.Y(n_996)
);

AOI21xp33_ASAP7_75t_SL g997 ( 
.A1(n_987),
.A2(n_803),
.B(n_918),
.Y(n_997)
);

OAI211xp5_ASAP7_75t_L g998 ( 
.A1(n_988),
.A2(n_903),
.B(n_890),
.C(n_900),
.Y(n_998)
);

AOI221xp5_ASAP7_75t_L g999 ( 
.A1(n_993),
.A2(n_903),
.B1(n_906),
.B2(n_904),
.C(n_890),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_989),
.B(n_881),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_992),
.B(n_903),
.Y(n_1001)
);

AOI22xp5_ASAP7_75t_L g1002 ( 
.A1(n_988),
.A2(n_900),
.B1(n_881),
.B2(n_880),
.Y(n_1002)
);

OAI211xp5_ASAP7_75t_SL g1003 ( 
.A1(n_995),
.A2(n_880),
.B(n_879),
.C(n_904),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_994),
.Y(n_1004)
);

AND2x2_ASAP7_75t_L g1005 ( 
.A(n_996),
.B(n_892),
.Y(n_1005)
);

AND2x2_ASAP7_75t_L g1006 ( 
.A(n_997),
.B(n_892),
.Y(n_1006)
);

AOI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_998),
.A2(n_904),
.B1(n_901),
.B2(n_883),
.Y(n_1007)
);

OR2x2_ASAP7_75t_L g1008 ( 
.A(n_1000),
.B(n_885),
.Y(n_1008)
);

OR2x2_ASAP7_75t_L g1009 ( 
.A(n_1002),
.B(n_1001),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_999),
.B(n_885),
.Y(n_1010)
);

OAI22xp5_ASAP7_75t_SL g1011 ( 
.A1(n_995),
.A2(n_878),
.B1(n_879),
.B2(n_885),
.Y(n_1011)
);

OAI22xp33_ASAP7_75t_SL g1012 ( 
.A1(n_1009),
.A2(n_895),
.B1(n_896),
.B2(n_899),
.Y(n_1012)
);

NOR3xp33_ASAP7_75t_L g1013 ( 
.A(n_1004),
.B(n_901),
.C(n_883),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_1005),
.B(n_895),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_1008),
.B(n_895),
.C(n_896),
.Y(n_1015)
);

OAI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_1006),
.A2(n_795),
.B(n_899),
.Y(n_1016)
);

AOI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_1011),
.A2(n_899),
.B1(n_862),
.B2(n_159),
.Y(n_1017)
);

AOI22xp5_ASAP7_75t_L g1018 ( 
.A1(n_1010),
.A2(n_152),
.B1(n_156),
.B2(n_160),
.Y(n_1018)
);

NOR2xp33_ASAP7_75t_L g1019 ( 
.A(n_1003),
.B(n_161),
.Y(n_1019)
);

NAND4xp25_ASAP7_75t_L g1020 ( 
.A(n_1018),
.B(n_1007),
.C(n_163),
.D(n_164),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_1013),
.B(n_162),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_1014),
.B(n_166),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_1017),
.A2(n_1019),
.B1(n_1016),
.B2(n_1015),
.Y(n_1023)
);

AND2x4_ASAP7_75t_L g1024 ( 
.A(n_1012),
.B(n_169),
.Y(n_1024)
);

INVx1_ASAP7_75t_SL g1025 ( 
.A(n_1018),
.Y(n_1025)
);

AOI211xp5_ASAP7_75t_L g1026 ( 
.A1(n_1025),
.A2(n_172),
.B(n_174),
.C(n_175),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_1022),
.B(n_221),
.Y(n_1027)
);

BUFx2_ASAP7_75t_L g1028 ( 
.A(n_1024),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_1021),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_1028),
.B(n_1029),
.Y(n_1030)
);

NAND3xp33_ASAP7_75t_SL g1031 ( 
.A(n_1026),
.B(n_1023),
.C(n_1020),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_1030),
.Y(n_1032)
);

HB1xp67_ASAP7_75t_L g1033 ( 
.A(n_1031),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_L g1034 ( 
.A1(n_1032),
.A2(n_1027),
.B1(n_178),
.B2(n_179),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_1033),
.A2(n_177),
.B(n_180),
.Y(n_1035)
);

AOI22xp33_ASAP7_75t_L g1036 ( 
.A1(n_1035),
.A2(n_181),
.B1(n_182),
.B2(n_183),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_1034),
.Y(n_1037)
);

XOR2xp5_ASAP7_75t_L g1038 ( 
.A(n_1037),
.B(n_184),
.Y(n_1038)
);

OAI221xp5_ASAP7_75t_R g1039 ( 
.A1(n_1036),
.A2(n_188),
.B1(n_190),
.B2(n_192),
.C(n_194),
.Y(n_1039)
);

OAI221xp5_ASAP7_75t_R g1040 ( 
.A1(n_1038),
.A2(n_195),
.B1(n_197),
.B2(n_199),
.C(n_200),
.Y(n_1040)
);

AOI211xp5_ASAP7_75t_L g1041 ( 
.A1(n_1040),
.A2(n_1039),
.B(n_202),
.C(n_206),
.Y(n_1041)
);


endmodule