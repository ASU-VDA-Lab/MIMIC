module fake_netlist_6_4088_n_1271 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_235, n_256, n_18, n_21, n_193, n_147, n_269, n_258, n_154, n_191, n_88, n_3, n_209, n_98, n_260, n_265, n_113, n_39, n_63, n_223, n_270, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_226, n_228, n_252, n_266, n_166, n_28, n_184, n_212, n_268, n_271, n_50, n_158, n_49, n_7, n_210, n_216, n_83, n_206, n_217, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_215, n_178, n_247, n_225, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_227, n_132, n_188, n_102, n_186, n_204, n_245, n_0, n_87, n_195, n_261, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_213, n_164, n_257, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_254, n_142, n_20, n_143, n_207, n_2, n_242, n_180, n_19, n_47, n_62, n_29, n_155, n_219, n_75, n_109, n_150, n_233, n_263, n_122, n_264, n_45, n_255, n_205, n_34, n_140, n_218, n_70, n_120, n_234, n_251, n_214, n_274, n_37, n_15, n_67, n_33, n_82, n_27, n_236, n_246, n_38, n_110, n_151, n_61, n_112, n_172, n_237, n_81, n_59, n_244, n_181, n_76, n_36, n_182, n_26, n_124, n_238, n_239, n_55, n_126, n_202, n_94, n_97, n_108, n_267, n_58, n_116, n_211, n_64, n_220, n_117, n_118, n_175, n_224, n_48, n_231, n_65, n_230, n_25, n_40, n_93, n_80, n_141, n_240, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_259, n_177, n_176, n_273, n_114, n_86, n_198, n_104, n_222, n_95, n_179, n_243, n_9, n_248, n_107, n_10, n_71, n_74, n_229, n_253, n_6, n_190, n_14, n_123, n_262, n_136, n_72, n_187, n_89, n_249, n_173, n_201, n_250, n_103, n_111, n_60, n_159, n_272, n_157, n_162, n_170, n_185, n_35, n_183, n_232, n_115, n_12, n_69, n_128, n_241, n_30, n_79, n_275, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_221, n_1271);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_235;
input n_256;
input n_18;
input n_21;
input n_193;
input n_147;
input n_269;
input n_258;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_260;
input n_265;
input n_113;
input n_39;
input n_63;
input n_223;
input n_270;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_226;
input n_228;
input n_252;
input n_266;
input n_166;
input n_28;
input n_184;
input n_212;
input n_268;
input n_271;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_216;
input n_83;
input n_206;
input n_217;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_215;
input n_178;
input n_247;
input n_225;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_227;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_245;
input n_0;
input n_87;
input n_195;
input n_261;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_213;
input n_164;
input n_257;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_254;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_242;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_219;
input n_75;
input n_109;
input n_150;
input n_233;
input n_263;
input n_122;
input n_264;
input n_45;
input n_255;
input n_205;
input n_34;
input n_140;
input n_218;
input n_70;
input n_120;
input n_234;
input n_251;
input n_214;
input n_274;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_236;
input n_246;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_237;
input n_81;
input n_59;
input n_244;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_238;
input n_239;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_267;
input n_58;
input n_116;
input n_211;
input n_64;
input n_220;
input n_117;
input n_118;
input n_175;
input n_224;
input n_48;
input n_231;
input n_65;
input n_230;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_240;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_259;
input n_177;
input n_176;
input n_273;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_95;
input n_179;
input n_243;
input n_9;
input n_248;
input n_107;
input n_10;
input n_71;
input n_74;
input n_229;
input n_253;
input n_6;
input n_190;
input n_14;
input n_123;
input n_262;
input n_136;
input n_72;
input n_187;
input n_89;
input n_249;
input n_173;
input n_201;
input n_250;
input n_103;
input n_111;
input n_60;
input n_159;
input n_272;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_232;
input n_115;
input n_12;
input n_69;
input n_128;
input n_241;
input n_30;
input n_79;
input n_275;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;
input n_221;

output n_1271;

wire n_992;
wire n_801;
wire n_1234;
wire n_1199;
wire n_741;
wire n_1027;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_700;
wire n_1038;
wire n_578;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_783;
wire n_798;
wire n_509;
wire n_1209;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_442;
wire n_480;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_461;
wire n_873;
wire n_383;
wire n_447;
wire n_1172;
wire n_852;
wire n_1078;
wire n_544;
wire n_1140;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1143;
wire n_1232;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_641;
wire n_822;
wire n_693;
wire n_1056;
wire n_758;
wire n_516;
wire n_1163;
wire n_1180;
wire n_943;
wire n_491;
wire n_772;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_538;
wire n_1106;
wire n_886;
wire n_343;
wire n_953;
wire n_1094;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_638;
wire n_1211;
wire n_381;
wire n_887;
wire n_713;
wire n_976;
wire n_734;
wire n_1088;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_659;
wire n_407;
wire n_913;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_577;
wire n_619;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_323;
wire n_606;
wire n_818;
wire n_1123;
wire n_513;
wire n_645;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1162;
wire n_860;
wire n_788;
wire n_939;
wire n_821;
wire n_938;
wire n_1068;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_979;
wire n_905;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_547;
wire n_558;
wire n_1064;
wire n_634;
wire n_966;
wire n_764;
wire n_692;
wire n_733;
wire n_1233;
wire n_487;
wire n_1107;
wire n_1014;
wire n_882;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_277;
wire n_618;
wire n_1167;
wire n_674;
wire n_871;
wire n_922;
wire n_1069;
wire n_612;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_429;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_286;
wire n_928;
wire n_1214;
wire n_835;
wire n_690;
wire n_850;
wire n_816;
wire n_1157;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1124;
wire n_515;
wire n_598;
wire n_696;
wire n_961;
wire n_437;
wire n_1082;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_484;
wire n_891;
wire n_949;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_881;
wire n_1008;
wire n_760;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_304;
wire n_694;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_1044;
wire n_449;
wire n_1208;
wire n_1164;
wire n_1072;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_898;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_615;
wire n_1249;
wire n_1127;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_826;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_631;
wire n_720;
wire n_842;
wire n_843;
wire n_656;
wire n_989;
wire n_797;
wire n_1246;
wire n_899;
wire n_738;
wire n_1035;
wire n_294;
wire n_499;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_648;
wire n_657;
wire n_1049;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_777;
wire n_526;
wire n_1183;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1178;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_552;
wire n_912;
wire n_745;
wire n_1142;
wire n_716;
wire n_623;
wire n_1048;
wire n_1201;
wire n_884;
wire n_731;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_527;
wire n_312;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_589;
wire n_819;
wire n_767;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_399;
wire n_505;
wire n_319;
wire n_537;
wire n_311;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_1053;
wire n_416;
wire n_520;
wire n_418;
wire n_1093;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_518;
wire n_1185;
wire n_453;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1224;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_335;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_1096;
wire n_1091;
wire n_1267;
wire n_983;
wire n_427;
wire n_496;
wire n_906;
wire n_688;
wire n_1077;
wire n_351;
wire n_385;
wire n_858;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_664;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_485;
wire n_443;
wire n_892;
wire n_768;
wire n_421;
wire n_1095;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1024;
wire n_517;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1115;
wire n_750;
wire n_901;
wire n_468;
wire n_923;
wire n_504;
wire n_1015;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_785;
wire n_746;
wire n_609;
wire n_1168;
wire n_1216;
wire n_302;
wire n_380;
wire n_1190;
wire n_397;
wire n_1262;
wire n_1213;
wire n_782;
wire n_490;
wire n_809;
wire n_1043;
wire n_986;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_921;
wire n_711;
wire n_579;
wire n_937;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_456;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_936;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_482;
wire n_934;
wire n_420;
wire n_394;
wire n_942;
wire n_543;
wire n_1225;
wire n_325;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_548;
wire n_282;
wire n_833;
wire n_523;
wire n_707;
wire n_345;
wire n_799;
wire n_1155;
wire n_787;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_550;
wire n_652;
wire n_560;
wire n_1241;
wire n_569;
wire n_737;
wire n_1235;
wire n_1229;
wire n_306;
wire n_346;
wire n_1029;
wire n_790;
wire n_1210;
wire n_299;
wire n_1248;
wire n_902;
wire n_333;
wire n_1047;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_655;
wire n_706;
wire n_1045;
wire n_786;
wire n_1236;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1002;
wire n_545;
wire n_489;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_660;
wire n_438;
wire n_1200;
wire n_479;
wire n_869;
wire n_1154;
wire n_1113;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_817;
wire n_897;
wire n_846;
wire n_841;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1177;
wire n_332;
wire n_1150;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_1007;
wire n_855;
wire n_591;
wire n_853;
wire n_440;
wire n_695;
wire n_875;
wire n_367;
wire n_680;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_969;
wire n_988;
wire n_1065;
wire n_1255;
wire n_568;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_698;
wire n_1074;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1130;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_555;
wire n_389;
wire n_814;
wire n_669;
wire n_300;
wire n_747;
wire n_1105;
wire n_721;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_378;
wire n_1196;
wire n_377;
wire n_863;
wire n_601;
wire n_338;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1205;
wire n_1258;
wire n_1173;
wire n_525;
wire n_1116;
wire n_611;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_795;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_930;
wire n_888;
wire n_1112;
wire n_910;
wire n_911;
wire n_653;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_414;
wire n_563;
wire n_1011;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_779;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1109;
wire n_712;
wire n_348;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_1239;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_1149;
wire n_1184;
wire n_719;
wire n_455;
wire n_363;
wire n_1090;
wire n_592;
wire n_829;
wire n_1156;
wire n_393;
wire n_984;
wire n_503;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_981;
wire n_714;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_802;
wire n_561;
wire n_980;
wire n_1198;
wire n_436;
wire n_409;
wire n_1244;
wire n_756;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_583;
wire n_1039;
wire n_1034;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_359;
wire n_973;
wire n_1055;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_588;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1006;
wire n_373;
wire n_730;
wire n_670;
wire n_1089;
wire n_1242;
wire n_681;
wire n_1226;
wire n_412;
wire n_640;
wire n_965;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_457;
wire n_364;
wire n_629;
wire n_900;
wire n_827;
wire n_531;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_649;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_216),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_177),
.Y(n_277)
);

BUFx2_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_6),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_238),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_57),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_53),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_97),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_48),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_150),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_204),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_211),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_102),
.Y(n_288)
);

BUFx5_ASAP7_75t_L g289 ( 
.A(n_241),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_263),
.Y(n_291)
);

BUFx10_ASAP7_75t_L g292 ( 
.A(n_178),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_92),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g294 ( 
.A(n_228),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_234),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_268),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_30),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_219),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_98),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_53),
.Y(n_300)
);

CKINVDCx16_ASAP7_75t_R g301 ( 
.A(n_139),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_256),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g303 ( 
.A(n_265),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_84),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_227),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_17),
.Y(n_307)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_249),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_169),
.Y(n_309)
);

HB1xp67_ASAP7_75t_SL g310 ( 
.A(n_262),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_20),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_100),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_140),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_16),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_28),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_62),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_80),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g318 ( 
.A(n_225),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_213),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_64),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_240),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_275),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_215),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_13),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_131),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_25),
.Y(n_326)
);

INVx1_ASAP7_75t_SL g327 ( 
.A(n_171),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_235),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_185),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_172),
.Y(n_330)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_144),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_195),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_230),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_82),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_106),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_148),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_68),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_18),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_59),
.Y(n_339)
);

BUFx10_ASAP7_75t_L g340 ( 
.A(n_246),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_266),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_5),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_72),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_32),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_267),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_1),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_42),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_125),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_61),
.Y(n_349)
);

BUFx8_ASAP7_75t_SL g350 ( 
.A(n_118),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_52),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_87),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_104),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_174),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_126),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_37),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_168),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_224),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_114),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_271),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_161),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_41),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_207),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_146),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_56),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_2),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_189),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_194),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_180),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_105),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_72),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_274),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_221),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_202),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_160),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_75),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_138),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_242),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_115),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_4),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_101),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_162),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_20),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_21),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_264),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_203),
.Y(n_386)
);

BUFx10_ASAP7_75t_L g387 ( 
.A(n_127),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_152),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_47),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_210),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_233),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_151),
.Y(n_392)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_226),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_6),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_40),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_111),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_269),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_143),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_87),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_90),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_154),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_43),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_261),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_193),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_77),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_149),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_67),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_129),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_245),
.Y(n_410)
);

INVxp33_ASAP7_75t_SL g411 ( 
.A(n_229),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_85),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_29),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_1),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_92),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_22),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_76),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_198),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_0),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_173),
.Y(n_420)
);

INVx1_ASAP7_75t_SL g421 ( 
.A(n_103),
.Y(n_421)
);

BUFx3_ASAP7_75t_L g422 ( 
.A(n_14),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_170),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_273),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_116),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_236),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_10),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_255),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_179),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_110),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_252),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_159),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_41),
.Y(n_433)
);

BUFx3_ASAP7_75t_L g434 ( 
.A(n_119),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g435 ( 
.A(n_214),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_137),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_208),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_220),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_157),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_62),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_247),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_113),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_212),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_65),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_65),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_94),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_45),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g448 ( 
.A(n_250),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_89),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_132),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_258),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_190),
.Y(n_452)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_84),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_68),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_222),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_109),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_248),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_71),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_278),
.B(n_0),
.Y(n_459)
);

BUFx8_ASAP7_75t_SL g460 ( 
.A(n_366),
.Y(n_460)
);

BUFx2_ASAP7_75t_L g461 ( 
.A(n_412),
.Y(n_461)
);

BUFx8_ASAP7_75t_L g462 ( 
.A(n_288),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_297),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_294),
.Y(n_464)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_294),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_309),
.B(n_2),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_309),
.B(n_3),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_297),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_319),
.B(n_3),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_297),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_297),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_319),
.B(n_4),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_330),
.B(n_5),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_294),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_7),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_348),
.B(n_8),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_348),
.B(n_8),
.Y(n_477)
);

AND2x4_ASAP7_75t_L g478 ( 
.A(n_434),
.B(n_9),
.Y(n_478)
);

BUFx3_ASAP7_75t_L g479 ( 
.A(n_286),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_363),
.B(n_9),
.Y(n_480)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_394),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_412),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_422),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_276),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_301),
.B(n_11),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_277),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

BUFx12f_ASAP7_75t_L g489 ( 
.A(n_286),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_363),
.B(n_12),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_379),
.B(n_12),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_294),
.Y(n_492)
);

BUFx6f_ASAP7_75t_L g493 ( 
.A(n_318),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_318),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_379),
.B(n_14),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_318),
.Y(n_496)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_303),
.B(n_15),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g498 ( 
.A(n_316),
.Y(n_498)
);

BUFx12f_ASAP7_75t_L g499 ( 
.A(n_286),
.Y(n_499)
);

INVx5_ASAP7_75t_L g500 ( 
.A(n_318),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_427),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_279),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g503 ( 
.A(n_316),
.Y(n_503)
);

HB1xp67_ASAP7_75t_L g504 ( 
.A(n_352),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_427),
.Y(n_505)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_427),
.B(n_16),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_453),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_359),
.Y(n_508)
);

INVx5_ASAP7_75t_L g509 ( 
.A(n_359),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_453),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_281),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_359),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_423),
.B(n_17),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_453),
.Y(n_514)
);

BUFx2_ASAP7_75t_L g515 ( 
.A(n_284),
.Y(n_515)
);

BUFx12f_ASAP7_75t_L g516 ( 
.A(n_292),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g517 ( 
.A(n_359),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_423),
.B(n_19),
.Y(n_518)
);

BUFx6f_ASAP7_75t_L g519 ( 
.A(n_457),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_428),
.B(n_19),
.Y(n_520)
);

BUFx2_ASAP7_75t_L g521 ( 
.A(n_293),
.Y(n_521)
);

AND2x4_ASAP7_75t_L g522 ( 
.A(n_428),
.B(n_23),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g523 ( 
.A(n_292),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_457),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_457),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_308),
.B(n_24),
.Y(n_526)
);

INVx5_ASAP7_75t_L g527 ( 
.A(n_457),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_340),
.Y(n_528)
);

AND2x6_ASAP7_75t_L g529 ( 
.A(n_280),
.B(n_95),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_340),
.B(n_24),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_282),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_289),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_289),
.Y(n_533)
);

AND2x4_ASAP7_75t_L g534 ( 
.A(n_331),
.B(n_290),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_352),
.B(n_383),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_291),
.B(n_26),
.Y(n_536)
);

INVx5_ASAP7_75t_L g537 ( 
.A(n_340),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_298),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_327),
.B(n_27),
.Y(n_539)
);

INVxp67_ASAP7_75t_L g540 ( 
.A(n_305),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_383),
.B(n_27),
.Y(n_541)
);

BUFx2_ASAP7_75t_L g542 ( 
.A(n_324),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_307),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_302),
.Y(n_544)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_387),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_387),
.B(n_28),
.Y(n_546)
);

AND2x6_ASAP7_75t_L g547 ( 
.A(n_306),
.B(n_96),
.Y(n_547)
);

BUFx8_ASAP7_75t_SL g548 ( 
.A(n_300),
.Y(n_548)
);

BUFx12f_ASAP7_75t_L g549 ( 
.A(n_326),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_311),
.B(n_29),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_314),
.B(n_30),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_313),
.B(n_31),
.Y(n_552)
);

HB1xp67_ASAP7_75t_L g553 ( 
.A(n_315),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g554 ( 
.A(n_317),
.B(n_32),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_320),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_289),
.Y(n_556)
);

BUFx3_ASAP7_75t_L g557 ( 
.A(n_350),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_334),
.B(n_33),
.Y(n_558)
);

AND2x4_ASAP7_75t_L g559 ( 
.A(n_322),
.B(n_33),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g560 ( 
.A(n_339),
.Y(n_560)
);

INVx5_ASAP7_75t_L g561 ( 
.A(n_289),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_325),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_289),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_356),
.B(n_34),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_344),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_346),
.B(n_349),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_421),
.B(n_435),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_336),
.B(n_34),
.Y(n_568)
);

INVx5_ASAP7_75t_L g569 ( 
.A(n_289),
.Y(n_569)
);

INVx3_ASAP7_75t_L g570 ( 
.A(n_365),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_448),
.B(n_35),
.Y(n_571)
);

AND2x4_ASAP7_75t_L g572 ( 
.A(n_357),
.B(n_35),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_393),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_361),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_395),
.B(n_36),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_411),
.B(n_36),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_393),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_364),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_369),
.B(n_374),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_399),
.B(n_402),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_283),
.Y(n_581)
);

BUFx8_ASAP7_75t_L g582 ( 
.A(n_406),
.Y(n_582)
);

HB1xp67_ASAP7_75t_L g583 ( 
.A(n_408),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_393),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g585 ( 
.A(n_433),
.B(n_37),
.Y(n_585)
);

BUFx3_ASAP7_75t_L g586 ( 
.A(n_285),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_414),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_393),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_419),
.B(n_38),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_446),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_454),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_375),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_377),
.B(n_39),
.Y(n_593)
);

AND2x6_ASAP7_75t_L g594 ( 
.A(n_382),
.B(n_99),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_386),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_337),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_445),
.B(n_40),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_287),
.Y(n_598)
);

OAI22xp33_ASAP7_75t_L g599 ( 
.A1(n_575),
.A2(n_342),
.B1(n_343),
.B2(n_338),
.Y(n_599)
);

AO22x2_ASAP7_75t_L g600 ( 
.A1(n_530),
.A2(n_392),
.B1(n_398),
.B2(n_397),
.Y(n_600)
);

AOI22x1_ASAP7_75t_L g601 ( 
.A1(n_513),
.A2(n_351),
.B1(n_362),
.B2(n_347),
.Y(n_601)
);

AO22x2_ASAP7_75t_L g602 ( 
.A1(n_530),
.A2(n_401),
.B1(n_418),
.B2(n_404),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_507),
.Y(n_603)
);

OAI22xp33_ASAP7_75t_L g604 ( 
.A1(n_575),
.A2(n_376),
.B1(n_380),
.B2(n_371),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_463),
.Y(n_605)
);

BUFx10_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_468),
.Y(n_607)
);

OR2x6_ASAP7_75t_L g608 ( 
.A(n_557),
.B(n_420),
.Y(n_608)
);

OAI22xp33_ASAP7_75t_L g609 ( 
.A1(n_585),
.A2(n_389),
.B1(n_400),
.B2(n_384),
.Y(n_609)
);

OR2x2_ASAP7_75t_L g610 ( 
.A(n_461),
.B(n_413),
.Y(n_610)
);

AND2x4_ASAP7_75t_L g611 ( 
.A(n_473),
.B(n_424),
.Y(n_611)
);

OAI22xp33_ASAP7_75t_SL g612 ( 
.A1(n_486),
.A2(n_310),
.B1(n_416),
.B2(n_415),
.Y(n_612)
);

AO22x2_ASAP7_75t_L g613 ( 
.A1(n_486),
.A2(n_431),
.B1(n_437),
.B2(n_430),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_528),
.B(n_409),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_481),
.A2(n_440),
.B1(n_444),
.B2(n_417),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_567),
.B(n_441),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_470),
.Y(n_617)
);

OAI22xp33_ASAP7_75t_L g618 ( 
.A1(n_585),
.A2(n_449),
.B1(n_458),
.B2(n_447),
.Y(n_618)
);

OAI22xp33_ASAP7_75t_SL g619 ( 
.A1(n_545),
.A2(n_456),
.B1(n_295),
.B2(n_296),
.Y(n_619)
);

INVx1_ASAP7_75t_SL g620 ( 
.A(n_548),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_502),
.B(n_299),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_511),
.B(n_304),
.Y(n_622)
);

AOI22xp5_ASAP7_75t_L g623 ( 
.A1(n_576),
.A2(n_321),
.B1(n_333),
.B2(n_312),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_576),
.A2(n_353),
.B1(n_373),
.B2(n_341),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_471),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_485),
.Y(n_626)
);

AO22x2_ASAP7_75t_L g627 ( 
.A1(n_546),
.A2(n_44),
.B1(n_42),
.B2(n_43),
.Y(n_627)
);

AO22x2_ASAP7_75t_L g628 ( 
.A1(n_475),
.A2(n_46),
.B1(n_44),
.B2(n_45),
.Y(n_628)
);

INVx2_ASAP7_75t_SL g629 ( 
.A(n_479),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_505),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_497),
.A2(n_328),
.B1(n_329),
.B2(n_323),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_510),
.Y(n_633)
);

OAI22xp33_ASAP7_75t_R g634 ( 
.A1(n_526),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_515),
.B(n_332),
.Y(n_635)
);

OAI22xp33_ASAP7_75t_R g636 ( 
.A1(n_526),
.A2(n_51),
.B1(n_49),
.B2(n_50),
.Y(n_636)
);

AND2x2_ASAP7_75t_L g637 ( 
.A(n_521),
.B(n_335),
.Y(n_637)
);

AO22x2_ASAP7_75t_L g638 ( 
.A1(n_475),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_638)
);

INVx3_ASAP7_75t_L g639 ( 
.A(n_464),
.Y(n_639)
);

INVx1_ASAP7_75t_SL g640 ( 
.A(n_548),
.Y(n_640)
);

AND2x4_ASAP7_75t_L g641 ( 
.A(n_586),
.B(n_345),
.Y(n_641)
);

AO22x2_ASAP7_75t_L g642 ( 
.A1(n_478),
.A2(n_56),
.B1(n_54),
.B2(n_55),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_514),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_464),
.Y(n_644)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_542),
.B(n_354),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_539),
.A2(n_358),
.B1(n_360),
.B2(n_355),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_592),
.Y(n_647)
);

AO22x2_ASAP7_75t_L g648 ( 
.A1(n_478),
.A2(n_57),
.B1(n_54),
.B2(n_55),
.Y(n_648)
);

AO22x2_ASAP7_75t_L g649 ( 
.A1(n_459),
.A2(n_60),
.B1(n_58),
.B2(n_59),
.Y(n_649)
);

INVx4_ASAP7_75t_L g650 ( 
.A(n_484),
.Y(n_650)
);

OAI22xp33_ASAP7_75t_L g651 ( 
.A1(n_593),
.A2(n_467),
.B1(n_469),
.B2(n_466),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_596),
.B(n_367),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_523),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_595),
.Y(n_654)
);

OAI22xp5_ASAP7_75t_SL g655 ( 
.A1(n_539),
.A2(n_455),
.B1(n_452),
.B2(n_451),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_SL g656 ( 
.A1(n_528),
.A2(n_450),
.B1(n_443),
.B2(n_442),
.Y(n_656)
);

OAI22xp5_ASAP7_75t_L g657 ( 
.A1(n_571),
.A2(n_439),
.B1(n_438),
.B2(n_436),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_528),
.B(n_368),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_SL g659 ( 
.A1(n_537),
.A2(n_432),
.B1(n_429),
.B2(n_426),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_498),
.Y(n_660)
);

AOI22xp5_ASAP7_75t_L g661 ( 
.A1(n_571),
.A2(n_549),
.B1(n_564),
.B2(n_554),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_465),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_474),
.Y(n_663)
);

INVx1_ASAP7_75t_SL g664 ( 
.A(n_537),
.Y(n_664)
);

OAI22xp33_ASAP7_75t_SL g665 ( 
.A1(n_537),
.A2(n_467),
.B1(n_469),
.B2(n_466),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_482),
.B(n_370),
.Y(n_666)
);

BUFx10_ASAP7_75t_L g667 ( 
.A(n_487),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_474),
.Y(n_668)
);

INVx3_ASAP7_75t_L g669 ( 
.A(n_474),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_492),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_492),
.Y(n_671)
);

AOI22xp5_ASAP7_75t_L g672 ( 
.A1(n_597),
.A2(n_372),
.B1(n_410),
.B2(n_407),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_498),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_593),
.A2(n_425),
.B1(n_405),
.B2(n_403),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_493),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_493),
.Y(n_676)
);

OAI22xp5_ASAP7_75t_SL g677 ( 
.A1(n_550),
.A2(n_396),
.B1(n_391),
.B2(n_390),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_489),
.A2(n_388),
.B1(n_385),
.B2(n_381),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_L g679 ( 
.A1(n_472),
.A2(n_378),
.B1(n_60),
.B2(n_61),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_493),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_494),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_647),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_654),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_616),
.B(n_598),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_617),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_644),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_662),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_625),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_676),
.Y(n_689)
);

INVxp67_ASAP7_75t_L g690 ( 
.A(n_610),
.Y(n_690)
);

AND2x4_ASAP7_75t_SL g691 ( 
.A(n_667),
.B(n_536),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_626),
.Y(n_692)
);

AND2x2_ASAP7_75t_L g693 ( 
.A(n_606),
.B(n_581),
.Y(n_693)
);

AND2x4_ASAP7_75t_SL g694 ( 
.A(n_667),
.B(n_536),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_633),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_605),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_639),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_639),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_605),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_669),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_664),
.B(n_534),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_666),
.B(n_534),
.Y(n_702)
);

AND2x2_ASAP7_75t_L g703 ( 
.A(n_629),
.B(n_483),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_663),
.Y(n_704)
);

XNOR2x2_ASAP7_75t_L g705 ( 
.A(n_649),
.B(n_627),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_668),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_651),
.B(n_579),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_660),
.B(n_488),
.Y(n_708)
);

XOR2xp5_ASAP7_75t_L g709 ( 
.A(n_623),
.B(n_553),
.Y(n_709)
);

INVx4_ASAP7_75t_L g710 ( 
.A(n_662),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_653),
.B(n_503),
.Y(n_711)
);

NOR2xp33_ASAP7_75t_L g712 ( 
.A(n_665),
.B(n_579),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_673),
.Y(n_713)
);

NAND2x1p5_ASAP7_75t_L g714 ( 
.A(n_650),
.B(n_552),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_599),
.B(n_499),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_671),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_604),
.B(n_609),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_675),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_680),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_641),
.B(n_552),
.Y(n_720)
);

AND2x4_ASAP7_75t_L g721 ( 
.A(n_641),
.B(n_559),
.Y(n_721)
);

BUFx6f_ASAP7_75t_L g722 ( 
.A(n_662),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_681),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_670),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_670),
.Y(n_725)
);

NAND2x1p5_ASAP7_75t_L g726 ( 
.A(n_650),
.B(n_559),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_603),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_630),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_603),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_607),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_631),
.Y(n_731)
);

AND2x2_ASAP7_75t_L g732 ( 
.A(n_621),
.B(n_503),
.Y(n_732)
);

XOR2xp5_ASAP7_75t_L g733 ( 
.A(n_624),
.B(n_560),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_643),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_618),
.B(n_516),
.Y(n_735)
);

BUFx2_ASAP7_75t_L g736 ( 
.A(n_622),
.Y(n_736)
);

OAI21xp5_ASAP7_75t_L g737 ( 
.A1(n_611),
.A2(n_547),
.B(n_529),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_R g738 ( 
.A(n_635),
.B(n_568),
.Y(n_738)
);

INVxp33_ASAP7_75t_SL g739 ( 
.A(n_655),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_600),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_637),
.B(n_504),
.Y(n_741)
);

AOI21xp5_ASAP7_75t_L g742 ( 
.A1(n_613),
.A2(n_477),
.B(n_476),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_602),
.Y(n_743)
);

INVx4_ASAP7_75t_L g744 ( 
.A(n_608),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_658),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_602),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_645),
.B(n_652),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_613),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_657),
.B(n_538),
.Y(n_749)
);

AND2x6_ASAP7_75t_L g750 ( 
.A(n_658),
.B(n_513),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_601),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_628),
.Y(n_752)
);

OR2x6_ASAP7_75t_L g753 ( 
.A(n_649),
.B(n_550),
.Y(n_753)
);

INVxp67_ASAP7_75t_SL g754 ( 
.A(n_679),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_638),
.Y(n_755)
);

NAND2x1p5_ASAP7_75t_L g756 ( 
.A(n_614),
.B(n_568),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_SL g757 ( 
.A(n_612),
.B(n_460),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_745),
.B(n_608),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_745),
.B(n_572),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_708),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_684),
.B(n_632),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_747),
.B(n_674),
.Y(n_762)
);

AND2x2_ASAP7_75t_SL g763 ( 
.A(n_717),
.B(n_522),
.Y(n_763)
);

AND2x2_ASAP7_75t_SL g764 ( 
.A(n_717),
.B(n_522),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_684),
.B(n_646),
.Y(n_765)
);

AND2x2_ASAP7_75t_L g766 ( 
.A(n_732),
.B(n_642),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_696),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_682),
.Y(n_768)
);

HB1xp67_ASAP7_75t_L g769 ( 
.A(n_711),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_696),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_741),
.B(n_642),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_751),
.B(n_672),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_683),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_699),
.Y(n_774)
);

INVxp67_ASAP7_75t_SL g775 ( 
.A(n_722),
.Y(n_775)
);

INVx3_ASAP7_75t_L g776 ( 
.A(n_699),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_750),
.B(n_707),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_702),
.B(n_648),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_707),
.A2(n_661),
.B(n_547),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_701),
.B(n_648),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_720),
.B(n_721),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_720),
.B(n_627),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_721),
.B(n_712),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_737),
.A2(n_547),
.B(n_529),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_712),
.B(n_504),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_750),
.B(n_742),
.Y(n_786)
);

INVxp67_ASAP7_75t_SL g787 ( 
.A(n_722),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_728),
.Y(n_788)
);

INVx4_ASAP7_75t_L g789 ( 
.A(n_750),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_728),
.Y(n_790)
);

AND2x2_ASAP7_75t_SL g791 ( 
.A(n_748),
.B(n_572),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_748),
.B(n_583),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_740),
.B(n_583),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_727),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_685),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_743),
.B(n_540),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_729),
.Y(n_797)
);

BUFx3_ASAP7_75t_L g798 ( 
.A(n_708),
.Y(n_798)
);

AND2x2_ASAP7_75t_L g799 ( 
.A(n_746),
.B(n_591),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_685),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_688),
.Y(n_801)
);

INVx3_ASAP7_75t_L g802 ( 
.A(n_688),
.Y(n_802)
);

INVx2_ASAP7_75t_SL g803 ( 
.A(n_703),
.Y(n_803)
);

BUFx6f_ASAP7_75t_L g804 ( 
.A(n_722),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_692),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_736),
.Y(n_806)
);

BUFx6f_ASAP7_75t_L g807 ( 
.A(n_722),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_749),
.B(n_547),
.Y(n_808)
);

CKINVDCx12_ASAP7_75t_R g809 ( 
.A(n_753),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_692),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_695),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_695),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_704),
.Y(n_813)
);

BUFx5_ASAP7_75t_L g814 ( 
.A(n_686),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_713),
.B(n_594),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_SL g816 ( 
.A(n_693),
.B(n_619),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_713),
.B(n_591),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_689),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_730),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_714),
.B(n_726),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_754),
.B(n_714),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_731),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_756),
.Y(n_823)
);

INVx2_ASAP7_75t_L g824 ( 
.A(n_734),
.Y(n_824)
);

INVx4_ASAP7_75t_L g825 ( 
.A(n_687),
.Y(n_825)
);

INVx1_ASAP7_75t_SL g826 ( 
.A(n_691),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_754),
.B(n_615),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_726),
.B(n_570),
.Y(n_828)
);

HB1xp67_ASAP7_75t_L g829 ( 
.A(n_738),
.Y(n_829)
);

AND2x2_ASAP7_75t_L g830 ( 
.A(n_756),
.B(n_570),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_691),
.B(n_694),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_706),
.B(n_594),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_687),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_694),
.B(n_590),
.Y(n_834)
);

BUFx6f_ASAP7_75t_L g835 ( 
.A(n_710),
.Y(n_835)
);

AND2x2_ASAP7_75t_SL g836 ( 
.A(n_715),
.B(n_476),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_690),
.B(n_753),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_715),
.B(n_656),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_716),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_753),
.B(n_590),
.Y(n_840)
);

INVxp67_ASAP7_75t_SL g841 ( 
.A(n_724),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_718),
.A2(n_509),
.B(n_500),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_817),
.B(n_735),
.Y(n_843)
);

BUFx2_ASAP7_75t_L g844 ( 
.A(n_806),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_804),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_770),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_774),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_781),
.B(n_744),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_821),
.Y(n_849)
);

OR2x6_ASAP7_75t_L g850 ( 
.A(n_831),
.B(n_744),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_765),
.B(n_735),
.Y(n_851)
);

BUFx2_ASAP7_75t_L g852 ( 
.A(n_783),
.Y(n_852)
);

BUFx6f_ASAP7_75t_L g853 ( 
.A(n_804),
.Y(n_853)
);

OR2x6_ASAP7_75t_L g854 ( 
.A(n_831),
.B(n_752),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_770),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_761),
.B(n_739),
.Y(n_857)
);

INVx4_ASAP7_75t_L g858 ( 
.A(n_804),
.Y(n_858)
);

INVx6_ASAP7_75t_L g859 ( 
.A(n_758),
.Y(n_859)
);

INVx2_ASAP7_75t_SL g860 ( 
.A(n_834),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_767),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_770),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_817),
.B(n_755),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_777),
.B(n_719),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_785),
.B(n_723),
.Y(n_865)
);

BUFx12f_ASAP7_75t_L g866 ( 
.A(n_758),
.Y(n_866)
);

INVxp67_ASAP7_75t_L g867 ( 
.A(n_769),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_785),
.B(n_709),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_776),
.Y(n_869)
);

BUFx2_ASAP7_75t_L g870 ( 
.A(n_783),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_763),
.B(n_733),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_SL g872 ( 
.A(n_764),
.B(n_757),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_764),
.B(n_827),
.Y(n_873)
);

AND2x2_ASAP7_75t_L g874 ( 
.A(n_803),
.B(n_829),
.Y(n_874)
);

BUFx2_ASAP7_75t_L g875 ( 
.A(n_837),
.Y(n_875)
);

AND2x4_ASAP7_75t_L g876 ( 
.A(n_781),
.B(n_697),
.Y(n_876)
);

INVx4_ASAP7_75t_L g877 ( 
.A(n_804),
.Y(n_877)
);

OR2x6_ASAP7_75t_L g878 ( 
.A(n_782),
.B(n_677),
.Y(n_878)
);

BUFx2_ASAP7_75t_L g879 ( 
.A(n_821),
.Y(n_879)
);

INVx3_ASAP7_75t_L g880 ( 
.A(n_776),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_776),
.Y(n_881)
);

NAND2x1_ASAP7_75t_SL g882 ( 
.A(n_766),
.B(n_678),
.Y(n_882)
);

NOR2xp67_ASAP7_75t_L g883 ( 
.A(n_772),
.B(n_698),
.Y(n_883)
);

INVx3_ASAP7_75t_L g884 ( 
.A(n_804),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_807),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_SL g886 ( 
.A(n_836),
.B(n_620),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_788),
.Y(n_887)
);

BUFx3_ASAP7_75t_L g888 ( 
.A(n_798),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_790),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_836),
.B(n_762),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_827),
.B(n_791),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_823),
.B(n_551),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_807),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_791),
.B(n_700),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_797),
.B(n_779),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_800),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_797),
.B(n_725),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_840),
.Y(n_898)
);

NOR2xp33_ASAP7_75t_SL g899 ( 
.A(n_789),
.B(n_640),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_814),
.B(n_532),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_814),
.B(n_533),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_807),
.Y(n_902)
);

NOR2xp33_ASAP7_75t_SL g903 ( 
.A(n_789),
.B(n_705),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_800),
.Y(n_904)
);

AND2x4_ASAP7_75t_L g905 ( 
.A(n_759),
.B(n_531),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_807),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_801),
.Y(n_907)
);

NAND2xp33_ASAP7_75t_L g908 ( 
.A(n_823),
.B(n_393),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_805),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_814),
.B(n_556),
.Y(n_910)
);

AND2x4_ASAP7_75t_L g911 ( 
.A(n_898),
.B(n_759),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_866),
.Y(n_912)
);

BUFx2_ASAP7_75t_L g913 ( 
.A(n_844),
.Y(n_913)
);

INVx5_ASAP7_75t_L g914 ( 
.A(n_845),
.Y(n_914)
);

INVx4_ASAP7_75t_L g915 ( 
.A(n_845),
.Y(n_915)
);

BUFx12f_ASAP7_75t_L g916 ( 
.A(n_850),
.Y(n_916)
);

BUFx6f_ASAP7_75t_L g917 ( 
.A(n_845),
.Y(n_917)
);

AND2x4_ASAP7_75t_L g918 ( 
.A(n_848),
.B(n_822),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_L g919 ( 
.A(n_851),
.B(n_838),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_853),
.Y(n_920)
);

NAND2x1p5_ASAP7_75t_L g921 ( 
.A(n_858),
.B(n_825),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_859),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_847),
.Y(n_923)
);

AND2x2_ASAP7_75t_L g924 ( 
.A(n_843),
.B(n_766),
.Y(n_924)
);

INVx1_ASAP7_75t_SL g925 ( 
.A(n_849),
.Y(n_925)
);

INVx6_ASAP7_75t_L g926 ( 
.A(n_859),
.Y(n_926)
);

BUFx2_ASAP7_75t_R g927 ( 
.A(n_868),
.Y(n_927)
);

INVx1_ASAP7_75t_SL g928 ( 
.A(n_849),
.Y(n_928)
);

NOR2xp33_ASAP7_75t_L g929 ( 
.A(n_857),
.B(n_780),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_896),
.Y(n_930)
);

BUFx12f_ASAP7_75t_L g931 ( 
.A(n_850),
.Y(n_931)
);

BUFx3_ASAP7_75t_L g932 ( 
.A(n_855),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_891),
.B(n_771),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_888),
.Y(n_934)
);

INVx1_ASAP7_75t_SL g935 ( 
.A(n_874),
.Y(n_935)
);

HB1xp67_ASAP7_75t_L g936 ( 
.A(n_879),
.Y(n_936)
);

BUFx2_ASAP7_75t_R g937 ( 
.A(n_868),
.Y(n_937)
);

BUFx2_ASAP7_75t_SL g938 ( 
.A(n_848),
.Y(n_938)
);

BUFx6f_ASAP7_75t_SL g939 ( 
.A(n_878),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_873),
.B(n_771),
.Y(n_940)
);

INVx1_ASAP7_75t_SL g941 ( 
.A(n_852),
.Y(n_941)
);

BUFx4f_ASAP7_75t_SL g942 ( 
.A(n_875),
.Y(n_942)
);

INVx5_ASAP7_75t_L g943 ( 
.A(n_853),
.Y(n_943)
);

INVx1_ASAP7_75t_SL g944 ( 
.A(n_870),
.Y(n_944)
);

BUFx2_ASAP7_75t_SL g945 ( 
.A(n_860),
.Y(n_945)
);

BUFx4_ASAP7_75t_SL g946 ( 
.A(n_878),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_904),
.Y(n_947)
);

INVx6_ASAP7_75t_L g948 ( 
.A(n_854),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_907),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_909),
.Y(n_950)
);

CKINVDCx11_ASAP7_75t_R g951 ( 
.A(n_878),
.Y(n_951)
);

INVx5_ASAP7_75t_L g952 ( 
.A(n_853),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_861),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_905),
.Y(n_954)
);

BUFx6f_ASAP7_75t_L g955 ( 
.A(n_906),
.Y(n_955)
);

INVx1_ASAP7_75t_SL g956 ( 
.A(n_863),
.Y(n_956)
);

BUFx6f_ASAP7_75t_L g957 ( 
.A(n_906),
.Y(n_957)
);

BUFx6f_ASAP7_75t_L g958 ( 
.A(n_906),
.Y(n_958)
);

BUFx6f_ASAP7_75t_L g959 ( 
.A(n_858),
.Y(n_959)
);

NAND2x1p5_ASAP7_75t_L g960 ( 
.A(n_877),
.B(n_825),
.Y(n_960)
);

CKINVDCx6p67_ASAP7_75t_R g961 ( 
.A(n_892),
.Y(n_961)
);

BUFx3_ASAP7_75t_L g962 ( 
.A(n_876),
.Y(n_962)
);

CKINVDCx20_ASAP7_75t_R g963 ( 
.A(n_871),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_887),
.Y(n_964)
);

INVxp67_ASAP7_75t_SL g965 ( 
.A(n_884),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_889),
.Y(n_966)
);

INVxp67_ASAP7_75t_L g967 ( 
.A(n_936),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_953),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_923),
.Y(n_969)
);

AOI22xp33_ASAP7_75t_L g970 ( 
.A1(n_919),
.A2(n_872),
.B1(n_890),
.B2(n_873),
.Y(n_970)
);

BUFx2_ASAP7_75t_L g971 ( 
.A(n_913),
.Y(n_971)
);

BUFx8_ASAP7_75t_SL g972 ( 
.A(n_963),
.Y(n_972)
);

INVx6_ASAP7_75t_L g973 ( 
.A(n_926),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_925),
.Y(n_974)
);

AND2x2_ASAP7_75t_L g975 ( 
.A(n_924),
.B(n_778),
.Y(n_975)
);

INVx4_ASAP7_75t_L g976 ( 
.A(n_914),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_932),
.Y(n_977)
);

AOI22xp33_ASAP7_75t_L g978 ( 
.A1(n_929),
.A2(n_903),
.B1(n_778),
.B2(n_816),
.Y(n_978)
);

INVx6_ASAP7_75t_L g979 ( 
.A(n_926),
.Y(n_979)
);

AOI22xp33_ASAP7_75t_SL g980 ( 
.A1(n_939),
.A2(n_886),
.B1(n_899),
.B2(n_634),
.Y(n_980)
);

INVx2_ASAP7_75t_L g981 ( 
.A(n_930),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_947),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_939),
.A2(n_886),
.B1(n_899),
.B2(n_636),
.Y(n_983)
);

AOI22xp33_ASAP7_75t_SL g984 ( 
.A1(n_940),
.A2(n_462),
.B1(n_786),
.B2(n_895),
.Y(n_984)
);

BUFx6f_ASAP7_75t_L g985 ( 
.A(n_914),
.Y(n_985)
);

BUFx10_ASAP7_75t_L g986 ( 
.A(n_912),
.Y(n_986)
);

INVxp67_ASAP7_75t_SL g987 ( 
.A(n_965),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_933),
.A2(n_956),
.B1(n_865),
.B2(n_506),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_SL g989 ( 
.A1(n_956),
.A2(n_462),
.B1(n_865),
.B2(n_823),
.Y(n_989)
);

INVx2_ASAP7_75t_L g990 ( 
.A(n_949),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_950),
.Y(n_991)
);

OAI22xp33_ASAP7_75t_L g992 ( 
.A1(n_935),
.A2(n_738),
.B1(n_897),
.B2(n_823),
.Y(n_992)
);

BUFx12f_ASAP7_75t_L g993 ( 
.A(n_951),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_964),
.Y(n_994)
);

AOI22xp33_ASAP7_75t_L g995 ( 
.A1(n_918),
.A2(n_954),
.B1(n_911),
.B2(n_948),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_928),
.B(n_792),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_966),
.A2(n_506),
.B1(n_558),
.B2(n_551),
.Y(n_997)
);

NAND2x1p5_ASAP7_75t_L g998 ( 
.A(n_914),
.B(n_877),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_L g999 ( 
.A1(n_961),
.A2(n_589),
.B1(n_558),
.B2(n_480),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_918),
.A2(n_589),
.B1(n_480),
.B2(n_490),
.Y(n_1000)
);

AOI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_911),
.A2(n_809),
.B1(n_867),
.B2(n_826),
.Y(n_1001)
);

CKINVDCx11_ASAP7_75t_R g1002 ( 
.A(n_916),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_SL g1003 ( 
.A1(n_946),
.A2(n_773),
.B1(n_768),
.B2(n_819),
.Y(n_1003)
);

OAI22xp33_ASAP7_75t_L g1004 ( 
.A1(n_941),
.A2(n_897),
.B1(n_894),
.B2(n_892),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_SL g1005 ( 
.A(n_934),
.Y(n_1005)
);

INVx6_ASAP7_75t_L g1006 ( 
.A(n_926),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_942),
.Y(n_1007)
);

BUFx10_ASAP7_75t_L g1008 ( 
.A(n_948),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_941),
.Y(n_1009)
);

BUFx8_ASAP7_75t_L g1010 ( 
.A(n_931),
.Y(n_1010)
);

INVx6_ASAP7_75t_L g1011 ( 
.A(n_914),
.Y(n_1011)
);

INVx2_ASAP7_75t_L g1012 ( 
.A(n_959),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_959),
.Y(n_1013)
);

OAI22xp5_ASAP7_75t_L g1014 ( 
.A1(n_938),
.A2(n_808),
.B1(n_883),
.B2(n_820),
.Y(n_1014)
);

CKINVDCx6p67_ASAP7_75t_R g1015 ( 
.A(n_922),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_946),
.Y(n_1016)
);

NAND3xp33_ASAP7_75t_L g1017 ( 
.A(n_984),
.B(n_582),
.C(n_830),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_972),
.Y(n_1018)
);

AOI22xp33_ASAP7_75t_L g1019 ( 
.A1(n_980),
.A2(n_828),
.B1(n_822),
.B2(n_824),
.Y(n_1019)
);

HB1xp67_ASAP7_75t_L g1020 ( 
.A(n_974),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_980),
.A2(n_828),
.B1(n_824),
.B2(n_944),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_983),
.A2(n_944),
.B1(n_819),
.B2(n_794),
.Y(n_1022)
);

BUFx8_ASAP7_75t_SL g1023 ( 
.A(n_993),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_981),
.Y(n_1024)
);

INVx2_ASAP7_75t_L g1025 ( 
.A(n_990),
.Y(n_1025)
);

AOI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_970),
.A2(n_818),
.B1(n_962),
.B2(n_659),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_999),
.A2(n_839),
.B1(n_908),
.B2(n_864),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_969),
.Y(n_1028)
);

CKINVDCx20_ASAP7_75t_R g1029 ( 
.A(n_1002),
.Y(n_1029)
);

NOR2xp33_ASAP7_75t_L g1030 ( 
.A(n_1009),
.B(n_927),
.Y(n_1030)
);

BUFx6f_ASAP7_75t_L g1031 ( 
.A(n_985),
.Y(n_1031)
);

INVx2_ASAP7_75t_SL g1032 ( 
.A(n_1011),
.Y(n_1032)
);

AOI22xp5_ASAP7_75t_L g1033 ( 
.A1(n_989),
.A2(n_945),
.B1(n_796),
.B2(n_799),
.Y(n_1033)
);

OAI22xp33_ASAP7_75t_L g1034 ( 
.A1(n_1001),
.A2(n_815),
.B1(n_784),
.B2(n_927),
.Y(n_1034)
);

HB1xp67_ASAP7_75t_L g1035 ( 
.A(n_974),
.Y(n_1035)
);

BUFx4f_ASAP7_75t_SL g1036 ( 
.A(n_1015),
.Y(n_1036)
);

INVx1_ASAP7_75t_SL g1037 ( 
.A(n_971),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_1016),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_988),
.B(n_975),
.Y(n_1039)
);

OR2x2_ASAP7_75t_L g1040 ( 
.A(n_996),
.B(n_793),
.Y(n_1040)
);

HB1xp67_ASAP7_75t_L g1041 ( 
.A(n_967),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_982),
.Y(n_1042)
);

OAI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_978),
.A2(n_937),
.B1(n_960),
.B2(n_921),
.Y(n_1043)
);

AOI22xp33_ASAP7_75t_SL g1044 ( 
.A1(n_1010),
.A2(n_541),
.B1(n_491),
.B2(n_495),
.Y(n_1044)
);

AOI22xp33_ASAP7_75t_L g1045 ( 
.A1(n_1000),
.A2(n_810),
.B1(n_812),
.B2(n_811),
.Y(n_1045)
);

BUFx12f_ASAP7_75t_L g1046 ( 
.A(n_986),
.Y(n_1046)
);

AOI222xp33_ASAP7_75t_L g1047 ( 
.A1(n_1003),
.A2(n_580),
.B1(n_566),
.B2(n_520),
.C1(n_518),
.C2(n_535),
.Y(n_1047)
);

AOI22xp33_ASAP7_75t_SL g1048 ( 
.A1(n_1010),
.A2(n_520),
.B1(n_882),
.B2(n_943),
.Y(n_1048)
);

CKINVDCx6p67_ASAP7_75t_R g1049 ( 
.A(n_1005),
.Y(n_1049)
);

AOI222xp33_ASAP7_75t_L g1050 ( 
.A1(n_997),
.A2(n_580),
.B1(n_566),
.B2(n_535),
.C1(n_543),
.C2(n_587),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_1000),
.A2(n_812),
.B1(n_813),
.B2(n_841),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_991),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_994),
.Y(n_1053)
);

AOI22xp33_ASAP7_75t_L g1054 ( 
.A1(n_1004),
.A2(n_813),
.B1(n_795),
.B2(n_802),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_968),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_L g1056 ( 
.A1(n_1004),
.A2(n_813),
.B1(n_795),
.B2(n_802),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_SL g1057 ( 
.A1(n_1005),
.A2(n_952),
.B1(n_943),
.B2(n_959),
.Y(n_1057)
);

OAI22xp33_ASAP7_75t_L g1058 ( 
.A1(n_1007),
.A2(n_952),
.B1(n_943),
.B2(n_880),
.Y(n_1058)
);

HB1xp67_ASAP7_75t_L g1059 ( 
.A(n_977),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_986),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_985),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_1053),
.Y(n_1062)
);

AOI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1017),
.A2(n_992),
.B1(n_995),
.B2(n_1014),
.Y(n_1063)
);

AOI22xp33_ASAP7_75t_L g1064 ( 
.A1(n_1044),
.A2(n_565),
.B1(n_555),
.B2(n_813),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_1022),
.A2(n_987),
.B1(n_1011),
.B2(n_973),
.Y(n_1065)
);

AOI22xp33_ASAP7_75t_L g1066 ( 
.A1(n_1047),
.A2(n_813),
.B1(n_1013),
.B2(n_1012),
.Y(n_1066)
);

AND2x2_ASAP7_75t_L g1067 ( 
.A(n_1039),
.B(n_1008),
.Y(n_1067)
);

AND2x2_ASAP7_75t_L g1068 ( 
.A(n_1053),
.B(n_846),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1021),
.A2(n_1006),
.B1(n_973),
.B2(n_979),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_1034),
.A2(n_856),
.B1(n_869),
.B2(n_862),
.Y(n_1070)
);

OAI222xp33_ASAP7_75t_L g1071 ( 
.A1(n_1033),
.A2(n_976),
.B1(n_998),
.B2(n_915),
.C1(n_880),
.C2(n_881),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1048),
.A2(n_814),
.B1(n_881),
.B2(n_832),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_SL g1073 ( 
.A1(n_1043),
.A2(n_985),
.B1(n_976),
.B2(n_998),
.Y(n_1073)
);

OAI222xp33_ASAP7_75t_L g1074 ( 
.A1(n_1019),
.A2(n_915),
.B1(n_910),
.B2(n_901),
.C1(n_900),
.C2(n_563),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_1020),
.B(n_917),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1028),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1024),
.Y(n_1077)
);

OAI222xp33_ASAP7_75t_L g1078 ( 
.A1(n_1026),
.A2(n_910),
.B1(n_584),
.B2(n_588),
.C1(n_577),
.C2(n_573),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_1035),
.B(n_958),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1030),
.A2(n_814),
.B1(n_574),
.B2(n_544),
.Y(n_1080)
);

HB1xp67_ASAP7_75t_L g1081 ( 
.A(n_1041),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_1024),
.B(n_958),
.Y(n_1082)
);

AND2x2_ASAP7_75t_L g1083 ( 
.A(n_1025),
.B(n_920),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_1050),
.A2(n_814),
.B1(n_832),
.B2(n_578),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_1037),
.A2(n_1027),
.B1(n_1046),
.B2(n_1040),
.Y(n_1085)
);

OAI22xp5_ASAP7_75t_L g1086 ( 
.A1(n_1060),
.A2(n_957),
.B1(n_955),
.B2(n_885),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1025),
.B(n_562),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_SL g1088 ( 
.A1(n_1060),
.A2(n_58),
.B1(n_63),
.B2(n_66),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_1055),
.B(n_63),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_1059),
.A2(n_885),
.B1(n_893),
.B2(n_902),
.Y(n_1090)
);

AOI22xp5_ASAP7_75t_L g1091 ( 
.A1(n_1049),
.A2(n_787),
.B1(n_775),
.B2(n_825),
.Y(n_1091)
);

OAI22xp5_ASAP7_75t_L g1092 ( 
.A1(n_1057),
.A2(n_835),
.B1(n_833),
.B2(n_512),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_1042),
.B(n_67),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_1052),
.A2(n_835),
.B1(n_833),
.B2(n_561),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1054),
.B(n_494),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1061),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_1045),
.A2(n_561),
.B1(n_569),
.B2(n_519),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_1032),
.A2(n_561),
.B1(n_569),
.B2(n_519),
.Y(n_1098)
);

NAND3xp33_ASAP7_75t_L g1099 ( 
.A(n_1056),
.B(n_1051),
.C(n_1018),
.Y(n_1099)
);

OAI222xp33_ASAP7_75t_L g1100 ( 
.A1(n_1018),
.A2(n_69),
.B1(n_70),
.B2(n_71),
.C1(n_73),
.C2(n_74),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_L g1101 ( 
.A1(n_1029),
.A2(n_1058),
.B1(n_1023),
.B2(n_1061),
.Y(n_1101)
);

OAI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1061),
.A2(n_842),
.B1(n_525),
.B2(n_524),
.C(n_519),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_L g1103 ( 
.A1(n_1023),
.A2(n_508),
.B1(n_524),
.B2(n_517),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_1081),
.B(n_1031),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_1076),
.Y(n_1105)
);

NAND3xp33_ASAP7_75t_L g1106 ( 
.A(n_1064),
.B(n_1031),
.C(n_1038),
.Y(n_1106)
);

NOR3xp33_ASAP7_75t_L g1107 ( 
.A(n_1100),
.B(n_1036),
.C(n_69),
.Y(n_1107)
);

NAND3xp33_ASAP7_75t_L g1108 ( 
.A(n_1063),
.B(n_1031),
.C(n_496),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1066),
.A2(n_524),
.B1(n_508),
.B2(n_494),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_1076),
.B(n_77),
.Y(n_1110)
);

NOR2xp33_ASAP7_75t_L g1111 ( 
.A(n_1067),
.B(n_78),
.Y(n_1111)
);

AOI221xp5_ASAP7_75t_L g1112 ( 
.A1(n_1088),
.A2(n_508),
.B1(n_79),
.B2(n_80),
.C(n_81),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1067),
.B(n_78),
.Y(n_1113)
);

NAND3xp33_ASAP7_75t_L g1114 ( 
.A(n_1085),
.B(n_527),
.C(n_509),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_SL g1115 ( 
.A1(n_1073),
.A2(n_82),
.B(n_83),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_1062),
.B(n_83),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1077),
.B(n_85),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1077),
.B(n_86),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1093),
.B(n_86),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_1096),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_1080),
.B(n_527),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1093),
.B(n_88),
.Y(n_1122)
);

OAI21xp5_ASAP7_75t_SL g1123 ( 
.A1(n_1099),
.A2(n_88),
.B(n_89),
.Y(n_1123)
);

AND2x2_ASAP7_75t_L g1124 ( 
.A(n_1096),
.B(n_90),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_1083),
.B(n_91),
.Y(n_1125)
);

OR2x2_ASAP7_75t_L g1126 ( 
.A(n_1075),
.B(n_91),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_1068),
.B(n_93),
.Y(n_1127)
);

OAI21xp5_ASAP7_75t_SL g1128 ( 
.A1(n_1101),
.A2(n_107),
.B(n_108),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_1068),
.B(n_1079),
.Y(n_1129)
);

NAND2xp5_ASAP7_75t_L g1130 ( 
.A(n_1083),
.B(n_112),
.Y(n_1130)
);

AND2x2_ASAP7_75t_L g1131 ( 
.A(n_1089),
.B(n_117),
.Y(n_1131)
);

AOI22xp33_ASAP7_75t_L g1132 ( 
.A1(n_1084),
.A2(n_120),
.B1(n_121),
.B2(n_122),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1082),
.B(n_123),
.Y(n_1133)
);

AND2x2_ASAP7_75t_L g1134 ( 
.A(n_1069),
.B(n_124),
.Y(n_1134)
);

OAI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_1103),
.A2(n_128),
.B(n_130),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_1065),
.B(n_133),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_L g1137 ( 
.A(n_1087),
.B(n_134),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1071),
.B(n_135),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1072),
.B(n_136),
.Y(n_1139)
);

OAI21xp5_ASAP7_75t_SL g1140 ( 
.A1(n_1078),
.A2(n_141),
.B(n_142),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1074),
.A2(n_145),
.B(n_147),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_1105),
.Y(n_1142)
);

INVx2_ASAP7_75t_SL g1143 ( 
.A(n_1104),
.Y(n_1143)
);

OR2x2_ASAP7_75t_L g1144 ( 
.A(n_1129),
.B(n_1095),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_1113),
.B(n_1086),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_1120),
.B(n_1110),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1110),
.B(n_1091),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1125),
.B(n_1091),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_1111),
.B(n_1070),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1125),
.B(n_1095),
.Y(n_1150)
);

AND2x2_ASAP7_75t_L g1151 ( 
.A(n_1124),
.B(n_1094),
.Y(n_1151)
);

NAND3xp33_ASAP7_75t_L g1152 ( 
.A(n_1112),
.B(n_1107),
.C(n_1123),
.Y(n_1152)
);

OR2x2_ASAP7_75t_L g1153 ( 
.A(n_1126),
.B(n_1090),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1128),
.A2(n_1092),
.B1(n_1102),
.B2(n_1097),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1124),
.Y(n_1155)
);

AO21x2_ASAP7_75t_L g1156 ( 
.A1(n_1121),
.A2(n_1098),
.B(n_155),
.Y(n_1156)
);

NOR3xp33_ASAP7_75t_L g1157 ( 
.A(n_1115),
.B(n_153),
.C(n_156),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1127),
.B(n_158),
.Y(n_1158)
);

AO21x2_ASAP7_75t_L g1159 ( 
.A1(n_1121),
.A2(n_163),
.B(n_164),
.Y(n_1159)
);

NAND4xp75_ASAP7_75t_L g1160 ( 
.A(n_1138),
.B(n_165),
.C(n_166),
.D(n_167),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1116),
.Y(n_1161)
);

NOR3xp33_ASAP7_75t_SL g1162 ( 
.A(n_1114),
.B(n_175),
.C(n_176),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_1117),
.Y(n_1163)
);

INVx2_ASAP7_75t_L g1164 ( 
.A(n_1118),
.Y(n_1164)
);

BUFx2_ASAP7_75t_SL g1165 ( 
.A(n_1161),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1142),
.Y(n_1166)
);

NAND4xp75_ASAP7_75t_L g1167 ( 
.A(n_1162),
.B(n_1141),
.C(n_1134),
.D(n_1136),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_1142),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1155),
.Y(n_1169)
);

AND2x2_ASAP7_75t_L g1170 ( 
.A(n_1143),
.B(n_1119),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1161),
.B(n_1164),
.Y(n_1171)
);

INVx2_ASAP7_75t_SL g1172 ( 
.A(n_1143),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1164),
.B(n_1122),
.Y(n_1173)
);

INVx3_ASAP7_75t_L g1174 ( 
.A(n_1155),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1146),
.Y(n_1175)
);

XNOR2x1_ASAP7_75t_L g1176 ( 
.A(n_1152),
.B(n_1106),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1146),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1163),
.Y(n_1178)
);

INVx3_ASAP7_75t_L g1179 ( 
.A(n_1150),
.Y(n_1179)
);

AND2x2_ASAP7_75t_L g1180 ( 
.A(n_1147),
.B(n_1148),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1144),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_1144),
.Y(n_1182)
);

INVx3_ASAP7_75t_L g1183 ( 
.A(n_1150),
.Y(n_1183)
);

AND2x2_ASAP7_75t_L g1184 ( 
.A(n_1147),
.B(n_1131),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1148),
.B(n_1108),
.Y(n_1185)
);

OR2x2_ASAP7_75t_L g1186 ( 
.A(n_1153),
.B(n_1130),
.Y(n_1186)
);

NOR2xp67_ASAP7_75t_L g1187 ( 
.A(n_1178),
.B(n_1145),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1166),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1166),
.Y(n_1189)
);

INVx1_ASAP7_75t_SL g1190 ( 
.A(n_1165),
.Y(n_1190)
);

XNOR2x1_ASAP7_75t_L g1191 ( 
.A(n_1176),
.B(n_1149),
.Y(n_1191)
);

NOR2xp33_ASAP7_75t_L g1192 ( 
.A(n_1176),
.B(n_1158),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1168),
.Y(n_1193)
);

INVx1_ASAP7_75t_SL g1194 ( 
.A(n_1165),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1178),
.Y(n_1195)
);

INVx1_ASAP7_75t_SL g1196 ( 
.A(n_1172),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_1172),
.Y(n_1197)
);

XOR2x2_ASAP7_75t_L g1198 ( 
.A(n_1184),
.B(n_1157),
.Y(n_1198)
);

OA22x2_ASAP7_75t_L g1199 ( 
.A1(n_1173),
.A2(n_1135),
.B1(n_1140),
.B2(n_1154),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1169),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1188),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1189),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1193),
.Y(n_1203)
);

OA22x2_ASAP7_75t_L g1204 ( 
.A1(n_1190),
.A2(n_1170),
.B1(n_1183),
.B2(n_1179),
.Y(n_1204)
);

INVxp67_ASAP7_75t_L g1205 ( 
.A(n_1191),
.Y(n_1205)
);

XOR2x2_ASAP7_75t_L g1206 ( 
.A(n_1198),
.B(n_1167),
.Y(n_1206)
);

OAI22x1_ASAP7_75t_L g1207 ( 
.A1(n_1192),
.A2(n_1183),
.B1(n_1179),
.B2(n_1170),
.Y(n_1207)
);

OA22x2_ASAP7_75t_L g1208 ( 
.A1(n_1194),
.A2(n_1183),
.B1(n_1182),
.B2(n_1181),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1195),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1187),
.Y(n_1210)
);

BUFx3_ASAP7_75t_L g1211 ( 
.A(n_1196),
.Y(n_1211)
);

OA22x2_ASAP7_75t_L g1212 ( 
.A1(n_1197),
.A2(n_1182),
.B1(n_1181),
.B2(n_1185),
.Y(n_1212)
);

BUFx2_ASAP7_75t_SL g1213 ( 
.A(n_1199),
.Y(n_1213)
);

INVx2_ASAP7_75t_L g1214 ( 
.A(n_1211),
.Y(n_1214)
);

NOR2x1_ASAP7_75t_SL g1215 ( 
.A(n_1211),
.B(n_1180),
.Y(n_1215)
);

OAI322xp33_ASAP7_75t_L g1216 ( 
.A1(n_1205),
.A2(n_1199),
.A3(n_1186),
.B1(n_1171),
.B2(n_1200),
.C1(n_1153),
.C2(n_1177),
.Y(n_1216)
);

AOI22x1_ASAP7_75t_L g1217 ( 
.A1(n_1213),
.A2(n_1186),
.B1(n_1151),
.B2(n_1180),
.Y(n_1217)
);

INVx2_ASAP7_75t_L g1218 ( 
.A(n_1208),
.Y(n_1218)
);

INVxp67_ASAP7_75t_SL g1219 ( 
.A(n_1210),
.Y(n_1219)
);

INVx2_ASAP7_75t_L g1220 ( 
.A(n_1208),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1201),
.Y(n_1221)
);

OA22x2_ASAP7_75t_L g1222 ( 
.A1(n_1218),
.A2(n_1210),
.B1(n_1207),
.B2(n_1206),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1219),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1219),
.Y(n_1224)
);

OA22x2_ASAP7_75t_L g1225 ( 
.A1(n_1220),
.A2(n_1202),
.B1(n_1203),
.B2(n_1209),
.Y(n_1225)
);

AOI22xp5_ASAP7_75t_L g1226 ( 
.A1(n_1214),
.A2(n_1212),
.B1(n_1204),
.B2(n_1167),
.Y(n_1226)
);

AOI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1222),
.A2(n_1220),
.B1(n_1221),
.B2(n_1160),
.Y(n_1227)
);

HB1xp67_ASAP7_75t_L g1228 ( 
.A(n_1223),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1224),
.Y(n_1229)
);

HB1xp67_ASAP7_75t_L g1230 ( 
.A(n_1225),
.Y(n_1230)
);

OAI22xp5_ASAP7_75t_L g1231 ( 
.A1(n_1226),
.A2(n_1217),
.B1(n_1216),
.B2(n_1215),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1230),
.B(n_1174),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1228),
.Y(n_1233)
);

NOR4xp25_ASAP7_75t_L g1234 ( 
.A(n_1229),
.B(n_1132),
.C(n_1133),
.D(n_1139),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1227),
.Y(n_1235)
);

AO22x2_ASAP7_75t_L g1236 ( 
.A1(n_1231),
.A2(n_1169),
.B1(n_1175),
.B2(n_1109),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1233),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_SL g1238 ( 
.A(n_1234),
.B(n_1151),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1232),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1235),
.B(n_1159),
.Y(n_1240)
);

AOI22xp5_ASAP7_75t_L g1241 ( 
.A1(n_1236),
.A2(n_1159),
.B1(n_1156),
.B2(n_1137),
.Y(n_1241)
);

HB1xp67_ASAP7_75t_L g1242 ( 
.A(n_1239),
.Y(n_1242)
);

OAI22x1_ASAP7_75t_L g1243 ( 
.A1(n_1238),
.A2(n_1236),
.B1(n_1159),
.B2(n_1156),
.Y(n_1243)
);

OR3x2_ASAP7_75t_L g1244 ( 
.A(n_1240),
.B(n_1156),
.C(n_182),
.Y(n_1244)
);

NOR3xp33_ASAP7_75t_L g1245 ( 
.A(n_1241),
.B(n_181),
.C(n_183),
.Y(n_1245)
);

INVx2_ASAP7_75t_L g1246 ( 
.A(n_1237),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1246),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1244),
.Y(n_1248)
);

INVxp67_ASAP7_75t_SL g1249 ( 
.A(n_1243),
.Y(n_1249)
);

AOI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1245),
.A2(n_184),
.B1(n_186),
.B2(n_187),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1242),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1242),
.Y(n_1252)
);

AO22x2_ASAP7_75t_L g1253 ( 
.A1(n_1249),
.A2(n_188),
.B1(n_191),
.B2(n_192),
.Y(n_1253)
);

OAI22x1_ASAP7_75t_L g1254 ( 
.A1(n_1251),
.A2(n_196),
.B1(n_197),
.B2(n_199),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1252),
.Y(n_1255)
);

OAI22xp5_ASAP7_75t_L g1256 ( 
.A1(n_1248),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1247),
.Y(n_1257)
);

INVx1_ASAP7_75t_L g1258 ( 
.A(n_1255),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1257),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1253),
.Y(n_1260)
);

AO22x2_ASAP7_75t_L g1261 ( 
.A1(n_1260),
.A2(n_1256),
.B1(n_1254),
.B2(n_1250),
.Y(n_1261)
);

OAI22xp5_ASAP7_75t_L g1262 ( 
.A1(n_1258),
.A2(n_217),
.B1(n_218),
.B2(n_223),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1261),
.Y(n_1263)
);

HB1xp67_ASAP7_75t_L g1264 ( 
.A(n_1262),
.Y(n_1264)
);

AOI22xp5_ASAP7_75t_SL g1265 ( 
.A1(n_1263),
.A2(n_1259),
.B1(n_231),
.B2(n_232),
.Y(n_1265)
);

OAI22xp33_ASAP7_75t_L g1266 ( 
.A1(n_1264),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_1266)
);

AOI22xp5_ASAP7_75t_L g1267 ( 
.A1(n_1263),
.A2(n_251),
.B1(n_253),
.B2(n_254),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1265),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1267),
.Y(n_1269)
);

AOI221xp5_ASAP7_75t_L g1270 ( 
.A1(n_1268),
.A2(n_1266),
.B1(n_257),
.B2(n_259),
.C(n_260),
.Y(n_1270)
);

AOI211xp5_ASAP7_75t_L g1271 ( 
.A1(n_1270),
.A2(n_1269),
.B(n_270),
.C(n_272),
.Y(n_1271)
);


endmodule