module fake_jpeg_3278_n_177 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_177);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_177;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx5_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_12),
.B(n_14),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_9),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_16),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_38),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_30),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_29),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_31),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_13),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_44),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_67),
.Y(n_72)
);

INVx11_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

BUFx2_ASAP7_75t_SL g78 ( 
.A(n_65),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_51),
.B(n_42),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_66),
.B(n_68),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_48),
.B(n_0),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_60),
.Y(n_69)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_60),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_70),
.Y(n_73)
);

CKINVDCx12_ASAP7_75t_R g71 ( 
.A(n_65),
.Y(n_71)
);

BUFx2_ASAP7_75t_SL g93 ( 
.A(n_71),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_69),
.Y(n_75)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_75),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_67),
.A2(n_49),
.B1(n_46),
.B2(n_58),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_80),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_50),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_49),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_83),
.B(n_84),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_64),
.B1(n_70),
.B2(n_69),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_85),
.A2(n_88),
.B1(n_91),
.B2(n_62),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_73),
.Y(n_86)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_86),
.B(n_98),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_87),
.B(n_94),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_55),
.B1(n_59),
.B2(n_45),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_89),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_77),
.A2(n_50),
.B1(n_57),
.B2(n_62),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_68),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_L g95 ( 
.A1(n_74),
.A2(n_52),
.B(n_54),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_56),
.B(n_61),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_77),
.B(n_46),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_79),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_86),
.B(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_112),
.Y(n_122)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_95),
.B(n_57),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_103),
.B(n_104),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_2),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_96),
.B1(n_86),
.B2(n_98),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_40),
.B1(n_39),
.B2(n_37),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_97),
.Y(n_109)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_109),
.Y(n_123)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_111),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_91),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_96),
.A2(n_52),
.B(n_54),
.C(n_53),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_97),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_118),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_92),
.A2(n_58),
.B(n_47),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_78),
.B(n_65),
.C(n_41),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_135)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_90),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_90),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_120),
.B(n_134),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_101),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_126),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_125),
.B(n_131),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_101),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_133),
.B1(n_136),
.B2(n_132),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_130),
.A2(n_4),
.B1(n_7),
.B2(n_8),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_35),
.C(n_33),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_136),
.C(n_137),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_106),
.B(n_3),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_135),
.A2(n_117),
.B1(n_109),
.B2(n_118),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_32),
.C(n_28),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_107),
.B(n_27),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_113),
.B(n_26),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_138),
.B(n_7),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_139),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_140),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_108),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_141),
.B(n_145),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_122),
.A2(n_116),
.B1(n_5),
.B2(n_6),
.Y(n_143)
);

AND2x2_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_129),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_146),
.B(n_149),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_150),
.B(n_151),
.C(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_123),
.Y(n_151)
);

AOI321xp33_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_153),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C(n_13),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_127),
.B(n_9),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_156),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_159),
.B(n_143),
.Y(n_165)
);

AOI221xp5_ASAP7_75t_L g161 ( 
.A1(n_141),
.A2(n_124),
.B1(n_135),
.B2(n_15),
.C(n_16),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_161),
.A2(n_149),
.B(n_139),
.Y(n_164)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_163),
.B(n_164),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_165),
.A2(n_144),
.B1(n_155),
.B2(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_168),
.B(n_140),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_154),
.B1(n_166),
.B2(n_163),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_170),
.A2(n_171),
.B1(n_168),
.B2(n_167),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_170),
.C(n_161),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_173),
.A2(n_147),
.B1(n_135),
.B2(n_23),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g175 ( 
.A1(n_174),
.A2(n_21),
.A3(n_25),
.B1(n_24),
.B2(n_20),
.C1(n_10),
.C2(n_17),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_175),
.A2(n_142),
.B1(n_14),
.B2(n_17),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_176),
.B(n_142),
.Y(n_177)
);


endmodule