module real_aes_6877_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_281;
wire n_496;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g112 ( .A(n_0), .Y(n_112) );
A2O1A1Ixp33_ASAP7_75t_L g459 ( .A1(n_1), .A2(n_137), .B(n_140), .C(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g144 ( .A(n_2), .Y(n_144) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_3), .A2(n_160), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_4), .B(n_172), .Y(n_485) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_5), .A2(n_15), .B1(n_695), .B2(n_696), .Y(n_694) );
CKINVDCx20_ASAP7_75t_R g696 ( .A(n_5), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g176 ( .A1(n_6), .A2(n_160), .B(n_177), .Y(n_176) );
AND2x6_ASAP7_75t_L g137 ( .A(n_7), .B(n_138), .Y(n_137) );
AOI21xp5_ASAP7_75t_L g246 ( .A1(n_8), .A2(n_247), .B(n_248), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_9), .B(n_43), .Y(n_113) );
INVx1_ASAP7_75t_L g452 ( .A(n_10), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g463 ( .A(n_11), .B(n_148), .Y(n_463) );
INVx1_ASAP7_75t_L g182 ( .A(n_12), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_13), .B(n_239), .Y(n_238) );
INVx1_ASAP7_75t_L g129 ( .A(n_14), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g695 ( .A(n_15), .Y(n_695) );
INVx1_ASAP7_75t_L g253 ( .A(n_16), .Y(n_253) );
A2O1A1Ixp33_ASAP7_75t_L g470 ( .A1(n_17), .A2(n_146), .B(n_254), .C(n_471), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_18), .B(n_172), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_19), .B(n_165), .Y(n_227) );
AOI222xp33_ASAP7_75t_L g115 ( .A1(n_20), .A2(n_116), .B1(n_694), .B2(n_697), .C1(n_700), .C2(n_705), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_21), .B(n_160), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_22), .B(n_522), .Y(n_521) );
A2O1A1Ixp33_ASAP7_75t_L g442 ( .A1(n_23), .A2(n_150), .B(n_239), .C(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_24), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g492 ( .A(n_25), .B(n_148), .Y(n_492) );
A2O1A1Ixp33_ASAP7_75t_L g250 ( .A1(n_26), .A2(n_251), .B(n_252), .C(n_254), .Y(n_250) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_27), .B(n_148), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g488 ( .A(n_28), .Y(n_488) );
INVx1_ASAP7_75t_L g501 ( .A(n_29), .Y(n_501) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_30), .Y(n_136) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_31), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_32), .B(n_148), .Y(n_147) );
INVx1_ASAP7_75t_L g519 ( .A(n_33), .Y(n_519) );
INVx1_ASAP7_75t_L g197 ( .A(n_34), .Y(n_197) );
INVx2_ASAP7_75t_L g135 ( .A(n_35), .Y(n_135) );
CKINVDCx20_ASAP7_75t_R g465 ( .A(n_36), .Y(n_465) );
A2O1A1Ixp33_ASAP7_75t_L g482 ( .A1(n_37), .A2(n_168), .B(n_239), .C(n_483), .Y(n_482) );
INVxp67_ASAP7_75t_L g520 ( .A(n_38), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_39), .A2(n_137), .B(n_140), .C(n_212), .Y(n_211) );
CKINVDCx14_ASAP7_75t_R g481 ( .A(n_40), .Y(n_481) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_41), .A2(n_140), .B(n_500), .C(n_505), .Y(n_499) );
OAI22xp5_ASAP7_75t_SL g713 ( .A1(n_42), .A2(n_89), .B1(n_714), .B2(n_715), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_42), .Y(n_715) );
INVx1_ASAP7_75t_L g195 ( .A(n_44), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g450 ( .A1(n_45), .A2(n_180), .B(n_216), .C(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_46), .B(n_148), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_47), .B(n_108), .Y(n_720) );
CKINVDCx20_ASAP7_75t_R g507 ( .A(n_48), .Y(n_507) );
CKINVDCx20_ASAP7_75t_R g516 ( .A(n_49), .Y(n_516) );
INVx1_ASAP7_75t_L g441 ( .A(n_50), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g198 ( .A(n_51), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_52), .B(n_160), .Y(n_241) );
AOI22xp5_ASAP7_75t_L g192 ( .A1(n_53), .A2(n_140), .B1(n_150), .B2(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g220 ( .A(n_54), .Y(n_220) );
CKINVDCx16_ASAP7_75t_R g131 ( .A(n_55), .Y(n_131) );
A2O1A1Ixp33_ASAP7_75t_L g179 ( .A1(n_56), .A2(n_168), .B(n_180), .C(n_181), .Y(n_179) );
CKINVDCx14_ASAP7_75t_R g449 ( .A(n_57), .Y(n_449) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_58), .Y(n_230) );
INVx1_ASAP7_75t_L g178 ( .A(n_59), .Y(n_178) );
INVx1_ASAP7_75t_L g138 ( .A(n_60), .Y(n_138) );
INVx1_ASAP7_75t_L g128 ( .A(n_61), .Y(n_128) );
INVx1_ASAP7_75t_SL g484 ( .A(n_62), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_63), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_64), .B(n_172), .Y(n_445) );
INVx1_ASAP7_75t_L g491 ( .A(n_65), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_SL g164 ( .A1(n_66), .A2(n_165), .B(n_166), .C(n_168), .Y(n_164) );
INVxp67_ASAP7_75t_L g167 ( .A(n_67), .Y(n_167) );
INVx1_ASAP7_75t_L g105 ( .A(n_68), .Y(n_105) );
AOI21xp5_ASAP7_75t_L g447 ( .A1(n_69), .A2(n_160), .B(n_448), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_70), .Y(n_495) );
CKINVDCx20_ASAP7_75t_R g200 ( .A(n_71), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_72), .A2(n_160), .B(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g223 ( .A(n_73), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_74), .A2(n_247), .B(n_515), .Y(n_514) );
INVx1_ASAP7_75t_L g469 ( .A(n_75), .Y(n_469) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_76), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g224 ( .A1(n_77), .A2(n_137), .B(n_140), .C(n_225), .Y(n_224) );
AOI21xp5_ASAP7_75t_L g439 ( .A1(n_78), .A2(n_160), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g472 ( .A(n_79), .Y(n_472) );
NAND2xp5_ASAP7_75t_SL g213 ( .A(n_80), .B(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g126 ( .A(n_81), .Y(n_126) );
INVx1_ASAP7_75t_L g461 ( .A(n_82), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_83), .B(n_165), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g139 ( .A1(n_84), .A2(n_137), .B(n_140), .C(n_143), .Y(n_139) );
OR2x2_ASAP7_75t_L g109 ( .A(n_85), .B(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g430 ( .A(n_85), .Y(n_430) );
OR2x2_ASAP7_75t_L g693 ( .A(n_85), .B(n_111), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_L g489 ( .A1(n_86), .A2(n_140), .B(n_490), .C(n_493), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_87), .B(n_155), .Y(n_183) );
CKINVDCx20_ASAP7_75t_R g153 ( .A(n_88), .Y(n_153) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_89), .A2(n_101), .B1(n_114), .B2(n_706), .C1(n_711), .C2(n_721), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g714 ( .A(n_89), .Y(n_714) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_90), .A2(n_137), .B(n_140), .C(n_236), .Y(n_235) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_91), .Y(n_243) );
INVx1_ASAP7_75t_L g163 ( .A(n_92), .Y(n_163) );
CKINVDCx16_ASAP7_75t_R g249 ( .A(n_93), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g237 ( .A(n_94), .B(n_145), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_95), .B(n_158), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_96), .B(n_158), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_97), .B(n_105), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g159 ( .A1(n_98), .A2(n_160), .B(n_161), .Y(n_159) );
INVx2_ASAP7_75t_L g444 ( .A(n_99), .Y(n_444) );
INVx1_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
NAND2xp33_ASAP7_75t_L g102 ( .A(n_103), .B(n_107), .Y(n_102) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_104), .B(n_106), .Y(n_103) );
INVx1_ASAP7_75t_SL g710 ( .A(n_104), .Y(n_710) );
INVx1_ASAP7_75t_L g709 ( .A(n_106), .Y(n_709) );
OA21x2_ASAP7_75t_L g722 ( .A1(n_106), .A2(n_710), .B(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g719 ( .A(n_109), .Y(n_719) );
BUFx2_ASAP7_75t_L g723 ( .A(n_109), .Y(n_723) );
NOR2x2_ASAP7_75t_L g699 ( .A(n_110), .B(n_430), .Y(n_699) );
INVx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g429 ( .A(n_111), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
OAI22xp5_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_429), .B1(n_431), .B2(n_693), .Y(n_116) );
INVx1_ASAP7_75t_L g701 ( .A(n_117), .Y(n_701) );
NAND2x1_ASAP7_75t_L g117 ( .A(n_118), .B(n_345), .Y(n_117) );
NOR5xp2_ASAP7_75t_L g118 ( .A(n_119), .B(n_268), .C(n_300), .D(n_315), .E(n_332), .Y(n_118) );
A2O1A1Ixp33_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_184), .B(n_205), .C(n_256), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_156), .Y(n_120) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_121), .B(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_121), .B(n_320), .Y(n_383) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_122), .B(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_122), .B(n_202), .Y(n_269) );
AND2x2_ASAP7_75t_L g310 ( .A(n_122), .B(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_122), .B(n_279), .Y(n_314) );
OR2x2_ASAP7_75t_L g351 ( .A(n_122), .B(n_190), .Y(n_351) );
INVx3_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x2_ASAP7_75t_L g189 ( .A(n_123), .B(n_190), .Y(n_189) );
INVx3_ASAP7_75t_L g259 ( .A(n_123), .Y(n_259) );
OR2x2_ASAP7_75t_L g422 ( .A(n_123), .B(n_262), .Y(n_422) );
AO21x2_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_130), .B(n_152), .Y(n_123) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_124), .A2(n_191), .B(n_199), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_124), .B(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g218 ( .A(n_124), .Y(n_218) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_125), .Y(n_158) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_127), .Y(n_125) );
AND2x2_ASAP7_75t_SL g155 ( .A(n_126), .B(n_127), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
OAI21xp5_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_132), .B(n_139), .Y(n_130) );
OAI22xp33_ASAP7_75t_L g191 ( .A1(n_132), .A2(n_170), .B1(n_192), .B2(n_198), .Y(n_191) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_132), .A2(n_223), .B(n_224), .Y(n_222) );
OAI21xp5_ASAP7_75t_L g457 ( .A1(n_132), .A2(n_458), .B(n_459), .Y(n_457) );
OAI21xp5_ASAP7_75t_L g487 ( .A1(n_132), .A2(n_488), .B(n_489), .Y(n_487) );
O2A1O1Ixp33_ASAP7_75t_L g497 ( .A1(n_132), .A2(n_155), .B(n_498), .C(n_499), .Y(n_497) );
NAND2x1p5_ASAP7_75t_L g132 ( .A(n_133), .B(n_137), .Y(n_132) );
AND2x4_ASAP7_75t_L g160 ( .A(n_133), .B(n_137), .Y(n_160) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx1_ASAP7_75t_L g504 ( .A(n_134), .Y(n_504) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g141 ( .A(n_135), .Y(n_141) );
INVx1_ASAP7_75t_L g151 ( .A(n_135), .Y(n_151) );
INVx1_ASAP7_75t_L g142 ( .A(n_136), .Y(n_142) );
INVx3_ASAP7_75t_L g146 ( .A(n_136), .Y(n_146) );
BUFx6f_ASAP7_75t_L g148 ( .A(n_136), .Y(n_148) );
INVx1_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_136), .Y(n_194) );
INVx4_ASAP7_75t_SL g170 ( .A(n_137), .Y(n_170) );
BUFx3_ASAP7_75t_L g505 ( .A(n_137), .Y(n_505) );
INVx5_ASAP7_75t_L g162 ( .A(n_140), .Y(n_162) );
AND2x6_ASAP7_75t_L g140 ( .A(n_141), .B(n_142), .Y(n_140) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
BUFx3_ASAP7_75t_L g217 ( .A(n_141), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g143 ( .A1(n_144), .A2(n_145), .B(n_147), .C(n_149), .Y(n_143) );
O2A1O1Ixp33_ASAP7_75t_L g500 ( .A1(n_145), .A2(n_501), .B(n_502), .C(n_503), .Y(n_500) );
OAI22xp33_ASAP7_75t_L g518 ( .A1(n_145), .A2(n_251), .B1(n_519), .B2(n_520), .Y(n_518) );
INVx5_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_146), .B(n_167), .Y(n_166) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_146), .B(n_182), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_146), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g180 ( .A(n_148), .Y(n_180) );
INVx4_ASAP7_75t_L g239 ( .A(n_148), .Y(n_239) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_154), .B(n_230), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g242 ( .A(n_154), .B(n_243), .Y(n_242) );
AO21x2_ASAP7_75t_L g456 ( .A1(n_154), .A2(n_457), .B(n_464), .Y(n_456) );
INVx1_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g233 ( .A(n_155), .Y(n_233) );
OA21x2_ASAP7_75t_L g245 ( .A1(n_155), .A2(n_246), .B(n_255), .Y(n_245) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_155), .A2(n_447), .B(n_453), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_156), .A2(n_325), .B1(n_326), .B2(n_329), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_156), .B(n_259), .Y(n_408) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_174), .Y(n_156) );
AND2x2_ASAP7_75t_L g204 ( .A(n_157), .B(n_190), .Y(n_204) );
AND2x2_ASAP7_75t_L g261 ( .A(n_157), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g266 ( .A(n_157), .Y(n_266) );
INVx3_ASAP7_75t_L g279 ( .A(n_157), .Y(n_279) );
OR2x2_ASAP7_75t_L g299 ( .A(n_157), .B(n_262), .Y(n_299) );
AND2x2_ASAP7_75t_L g318 ( .A(n_157), .B(n_175), .Y(n_318) );
BUFx2_ASAP7_75t_L g350 ( .A(n_157), .Y(n_350) );
OA21x2_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_171), .Y(n_157) );
INVx4_ASAP7_75t_L g173 ( .A(n_158), .Y(n_173) );
HB1xp67_ASAP7_75t_L g438 ( .A(n_158), .Y(n_438) );
BUFx2_ASAP7_75t_L g247 ( .A(n_160), .Y(n_247) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_163), .B(n_164), .C(n_170), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g177 ( .A1(n_162), .A2(n_170), .B(n_178), .C(n_179), .Y(n_177) );
O2A1O1Ixp33_ASAP7_75t_L g248 ( .A1(n_162), .A2(n_170), .B(n_249), .C(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g440 ( .A1(n_162), .A2(n_170), .B(n_441), .C(n_442), .Y(n_440) );
O2A1O1Ixp33_ASAP7_75t_SL g448 ( .A1(n_162), .A2(n_170), .B(n_449), .C(n_450), .Y(n_448) );
O2A1O1Ixp33_ASAP7_75t_SL g468 ( .A1(n_162), .A2(n_170), .B(n_469), .C(n_470), .Y(n_468) );
O2A1O1Ixp33_ASAP7_75t_L g480 ( .A1(n_162), .A2(n_170), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_SL g515 ( .A1(n_162), .A2(n_170), .B(n_516), .C(n_517), .Y(n_515) );
INVx3_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
HB1xp67_ASAP7_75t_L g240 ( .A(n_169), .Y(n_240) );
INVx1_ASAP7_75t_L g493 ( .A(n_170), .Y(n_493) );
OA21x2_ASAP7_75t_L g175 ( .A1(n_172), .A2(n_176), .B(n_183), .Y(n_175) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_SL g219 ( .A(n_173), .B(n_220), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g464 ( .A(n_173), .B(n_465), .Y(n_464) );
AO21x2_ASAP7_75t_L g486 ( .A1(n_173), .A2(n_487), .B(n_494), .Y(n_486) );
NOR2xp33_ASAP7_75t_L g506 ( .A(n_173), .B(n_507), .Y(n_506) );
AND2x4_ASAP7_75t_L g265 ( .A(n_174), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_SL g174 ( .A(n_175), .Y(n_174) );
BUFx2_ASAP7_75t_L g188 ( .A(n_175), .Y(n_188) );
INVx2_ASAP7_75t_L g203 ( .A(n_175), .Y(n_203) );
OR2x2_ASAP7_75t_L g281 ( .A(n_175), .B(n_262), .Y(n_281) );
AND2x2_ASAP7_75t_L g311 ( .A(n_175), .B(n_190), .Y(n_311) );
AND2x2_ASAP7_75t_L g328 ( .A(n_175), .B(n_259), .Y(n_328) );
AND2x2_ASAP7_75t_L g368 ( .A(n_175), .B(n_279), .Y(n_368) );
AND2x2_ASAP7_75t_SL g404 ( .A(n_175), .B(n_204), .Y(n_404) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp33_ASAP7_75t_SL g185 ( .A(n_186), .B(n_201), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_187), .B(n_189), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_187), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_SL g187 ( .A(n_188), .Y(n_187) );
OAI21xp33_ASAP7_75t_L g342 ( .A1(n_188), .A2(n_204), .B(n_343), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g398 ( .A(n_188), .B(n_190), .Y(n_398) );
AND2x2_ASAP7_75t_L g334 ( .A(n_189), .B(n_335), .Y(n_334) );
INVx3_ASAP7_75t_L g262 ( .A(n_190), .Y(n_262) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_190), .Y(n_360) );
OAI22xp5_ASAP7_75t_SL g193 ( .A1(n_194), .A2(n_195), .B1(n_196), .B2(n_197), .Y(n_193) );
INVx2_ASAP7_75t_L g196 ( .A(n_194), .Y(n_196) );
INVx4_ASAP7_75t_L g251 ( .A(n_194), .Y(n_251) );
INVx2_ASAP7_75t_L g462 ( .A(n_196), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_201), .B(n_259), .Y(n_427) );
INVx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
AOI22xp33_ASAP7_75t_L g369 ( .A1(n_202), .A2(n_370), .B1(n_371), .B2(n_376), .Y(n_369) );
AND2x2_ASAP7_75t_L g202 ( .A(n_203), .B(n_204), .Y(n_202) );
AND2x2_ASAP7_75t_L g260 ( .A(n_203), .B(n_261), .Y(n_260) );
OR2x2_ASAP7_75t_L g298 ( .A(n_203), .B(n_299), .Y(n_298) );
INVx1_ASAP7_75t_SL g335 ( .A(n_203), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_204), .B(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g389 ( .A(n_204), .Y(n_389) );
CKINVDCx16_ASAP7_75t_R g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_231), .Y(n_206) );
INVx4_ASAP7_75t_L g275 ( .A(n_207), .Y(n_275) );
AND2x2_ASAP7_75t_L g353 ( .A(n_207), .B(n_320), .Y(n_353) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_221), .Y(n_207) );
INVx3_ASAP7_75t_L g272 ( .A(n_208), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_287), .Y(n_286) );
INVx1_ASAP7_75t_L g290 ( .A(n_208), .Y(n_290) );
INVx2_ASAP7_75t_L g304 ( .A(n_208), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_208), .B(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g361 ( .A(n_208), .B(n_356), .Y(n_361) );
AND2x2_ASAP7_75t_L g426 ( .A(n_208), .B(n_396), .Y(n_426) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_219), .Y(n_208) );
AOI21xp5_ASAP7_75t_SL g209 ( .A1(n_210), .A2(n_211), .B(n_218), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_214), .B(n_215), .Y(n_212) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_215), .A2(n_226), .B(n_227), .Y(n_225) );
O2A1O1Ixp5_ASAP7_75t_L g460 ( .A1(n_215), .A2(n_461), .B(n_462), .C(n_463), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_215), .A2(n_462), .B(n_491), .C(n_492), .Y(n_490) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g254 ( .A(n_217), .Y(n_254) );
INVx1_ASAP7_75t_L g228 ( .A(n_218), .Y(n_228) );
AND2x2_ASAP7_75t_L g267 ( .A(n_221), .B(n_245), .Y(n_267) );
INVx2_ASAP7_75t_L g287 ( .A(n_221), .Y(n_287) );
AO21x2_ASAP7_75t_L g221 ( .A1(n_222), .A2(n_228), .B(n_229), .Y(n_221) );
INVx1_ASAP7_75t_L g513 ( .A(n_228), .Y(n_513) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_228), .A2(n_529), .B(n_530), .Y(n_528) );
INVx1_ASAP7_75t_L g292 ( .A(n_231), .Y(n_292) );
AND2x2_ASAP7_75t_L g338 ( .A(n_231), .B(n_286), .Y(n_338) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_244), .Y(n_231) );
INVx2_ASAP7_75t_L g277 ( .A(n_232), .Y(n_277) );
INVx1_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
AND2x2_ASAP7_75t_L g303 ( .A(n_232), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_232), .B(n_287), .Y(n_341) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_234), .B(n_242), .Y(n_232) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_233), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_L g522 ( .A(n_233), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_241), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_237), .A2(n_238), .B(n_240), .Y(n_236) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_239), .B(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g320 ( .A(n_244), .B(n_277), .Y(n_320) );
INVx1_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g273 ( .A(n_245), .Y(n_273) );
AND2x2_ASAP7_75t_L g356 ( .A(n_245), .B(n_287), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_251), .B(n_253), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_251), .B(n_444), .Y(n_443) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_251), .B(n_472), .Y(n_471) );
OAI21xp5_ASAP7_75t_SL g256 ( .A1(n_257), .A2(n_263), .B(n_267), .Y(n_256) );
INVx1_ASAP7_75t_SL g301 ( .A(n_257), .Y(n_301) );
AND2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_260), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_258), .B(n_265), .Y(n_358) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g307 ( .A(n_259), .B(n_262), .Y(n_307) );
AND2x2_ASAP7_75t_L g336 ( .A(n_259), .B(n_280), .Y(n_336) );
OR2x2_ASAP7_75t_L g339 ( .A(n_259), .B(n_299), .Y(n_339) );
AOI222xp33_ASAP7_75t_L g403 ( .A1(n_260), .A2(n_352), .B1(n_404), .B2(n_405), .C1(n_407), .C2(n_409), .Y(n_403) );
BUFx2_ASAP7_75t_L g317 ( .A(n_262), .Y(n_317) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g306 ( .A(n_265), .B(n_307), .Y(n_306) );
INVx3_ASAP7_75t_SL g323 ( .A(n_265), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_265), .B(n_317), .Y(n_377) );
AND2x2_ASAP7_75t_L g312 ( .A(n_267), .B(n_272), .Y(n_312) );
INVx1_ASAP7_75t_L g331 ( .A(n_267), .Y(n_331) );
OAI221xp5_ASAP7_75t_SL g268 ( .A1(n_269), .A2(n_270), .B1(n_274), .B2(n_278), .C(n_282), .Y(n_268) );
OR2x2_ASAP7_75t_L g340 ( .A(n_270), .B(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
AND2x2_ASAP7_75t_L g325 ( .A(n_272), .B(n_295), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_272), .B(n_285), .Y(n_365) );
AND2x2_ASAP7_75t_L g370 ( .A(n_272), .B(n_320), .Y(n_370) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_272), .Y(n_380) );
NAND2x1_ASAP7_75t_SL g391 ( .A(n_272), .B(n_392), .Y(n_391) );
OR2x2_ASAP7_75t_L g276 ( .A(n_273), .B(n_277), .Y(n_276) );
INVx2_ASAP7_75t_L g296 ( .A(n_273), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_273), .B(n_291), .Y(n_322) );
INVx1_ASAP7_75t_L g388 ( .A(n_273), .Y(n_388) );
INVx1_ASAP7_75t_L g363 ( .A(n_274), .Y(n_363) );
OR2x2_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx1_ASAP7_75t_L g375 ( .A(n_275), .Y(n_375) );
NOR2xp67_ASAP7_75t_L g387 ( .A(n_275), .B(n_388), .Y(n_387) );
INVx2_ASAP7_75t_L g392 ( .A(n_276), .Y(n_392) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_276), .B(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g295 ( .A(n_277), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_277), .B(n_287), .Y(n_308) );
INVx1_ASAP7_75t_L g374 ( .A(n_277), .Y(n_374) );
INVx1_ASAP7_75t_L g395 ( .A(n_278), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_283), .A2(n_288), .B(n_297), .Y(n_282) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
AND2x2_ASAP7_75t_L g428 ( .A(n_284), .B(n_361), .Y(n_428) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g396 ( .A(n_285), .B(n_356), .Y(n_396) );
AOI32xp33_ASAP7_75t_L g309 ( .A1(n_286), .A2(n_292), .A3(n_310), .B1(n_312), .B2(n_313), .Y(n_309) );
AOI322xp5_ASAP7_75t_L g411 ( .A1(n_286), .A2(n_318), .A3(n_401), .B1(n_412), .B2(n_413), .C1(n_414), .C2(n_416), .Y(n_411) );
INVx2_ASAP7_75t_L g291 ( .A(n_287), .Y(n_291) );
INVx1_ASAP7_75t_L g401 ( .A(n_287), .Y(n_401) );
OAI22xp5_ASAP7_75t_L g288 ( .A1(n_289), .A2(n_292), .B1(n_293), .B2(n_294), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_289), .B(n_295), .Y(n_344) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_291), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_290), .B(n_356), .Y(n_406) );
INVx1_ASAP7_75t_L g293 ( .A(n_291), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g410 ( .A(n_291), .B(n_320), .Y(n_410) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_SL g297 ( .A(n_298), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g393 ( .A(n_299), .B(n_394), .Y(n_393) );
OAI221xp5_ASAP7_75t_SL g300 ( .A1(n_301), .A2(n_302), .B1(n_305), .B2(n_308), .C(n_309), .Y(n_300) );
OR2x2_ASAP7_75t_L g321 ( .A(n_302), .B(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g330 ( .A(n_302), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g355 ( .A(n_303), .B(n_356), .Y(n_355) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
AND2x2_ASAP7_75t_L g359 ( .A(n_313), .B(n_360), .Y(n_359) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI221xp5_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_319), .B1(n_321), .B2(n_323), .C(n_324), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_317), .A2(n_348), .B1(n_352), .B2(n_353), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_318), .B(n_419), .Y(n_418) );
INVx1_ASAP7_75t_L g423 ( .A(n_318), .Y(n_423) );
INVx1_ASAP7_75t_L g417 ( .A(n_320), .Y(n_417) );
INVx1_ASAP7_75t_SL g352 ( .A(n_321), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_323), .B(n_351), .Y(n_413) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_328), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_SL g394 ( .A(n_328), .Y(n_394) );
INVx1_ASAP7_75t_SL g329 ( .A(n_330), .Y(n_329) );
OAI221xp5_ASAP7_75t_SL g332 ( .A1(n_333), .A2(n_337), .B1(n_339), .B2(n_340), .C(n_342), .Y(n_332) );
NOR2xp33_ASAP7_75t_SL g333 ( .A(n_334), .B(n_336), .Y(n_333) );
AOI22xp5_ASAP7_75t_L g397 ( .A1(n_334), .A2(n_352), .B1(n_398), .B2(n_399), .Y(n_397) );
CKINVDCx14_ASAP7_75t_R g337 ( .A(n_338), .Y(n_337) );
OAI21xp33_ASAP7_75t_L g416 ( .A1(n_339), .A2(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
NOR3xp33_ASAP7_75t_SL g345 ( .A(n_346), .B(n_378), .C(n_402), .Y(n_345) );
NAND4xp25_ASAP7_75t_L g346 ( .A(n_347), .B(n_354), .C(n_362), .D(n_369), .Y(n_346) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
OR2x2_ASAP7_75t_L g349 ( .A(n_350), .B(n_351), .Y(n_349) );
INVx1_ASAP7_75t_L g425 ( .A(n_350), .Y(n_425) );
INVx3_ASAP7_75t_SL g419 ( .A(n_351), .Y(n_419) );
OR2x2_ASAP7_75t_L g424 ( .A(n_351), .B(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_357), .B1(n_359), .B2(n_361), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_356), .B(n_374), .Y(n_415) );
INVxp67_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
OAI21xp5_ASAP7_75t_SL g362 ( .A1(n_363), .A2(n_364), .B(n_366), .Y(n_362) );
INVxp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVxp67_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_379), .A2(n_381), .B(n_384), .C(n_397), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g412 ( .A(n_383), .Y(n_412) );
AOI222xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_389), .B1(n_390), .B2(n_393), .C1(n_395), .C2(n_396), .Y(n_384) );
INVxp67_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NAND4xp25_ASAP7_75t_SL g421 ( .A(n_394), .B(n_422), .C(n_423), .D(n_424), .Y(n_421) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NAND3xp33_ASAP7_75t_SL g402 ( .A(n_403), .B(n_411), .C(n_420), .Y(n_402) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_426), .B1(n_427), .B2(n_428), .Y(n_420) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_429), .A2(n_701), .B1(n_702), .B2(n_704), .Y(n_700) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_431), .A2(n_704), .B1(n_713), .B2(n_716), .Y(n_712) );
INVx1_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx2_ASAP7_75t_L g704 ( .A(n_432), .Y(n_704) );
AND2x2_ASAP7_75t_L g432 ( .A(n_433), .B(n_619), .Y(n_432) );
NOR4xp25_ASAP7_75t_L g433 ( .A(n_434), .B(n_561), .C(n_591), .D(n_601), .Y(n_433) );
OAI211xp5_ASAP7_75t_L g434 ( .A1(n_435), .A2(n_474), .B(n_524), .C(n_551), .Y(n_434) );
OAI222xp33_ASAP7_75t_L g646 ( .A1(n_435), .A2(n_566), .B1(n_647), .B2(n_648), .C1(n_649), .C2(n_650), .Y(n_646) );
OR2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_454), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g572 ( .A1(n_436), .A2(n_559), .A3(n_560), .B1(n_573), .B2(n_578), .B3(n_580), .Y(n_572) );
OAI211xp5_ASAP7_75t_SL g629 ( .A1(n_436), .A2(n_630), .B(n_632), .C(n_634), .Y(n_629) );
OR2x2_ASAP7_75t_L g645 ( .A(n_436), .B(n_631), .Y(n_645) );
INVx1_ASAP7_75t_L g678 ( .A(n_436), .Y(n_678) );
OR2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_446), .Y(n_436) );
INVx2_ASAP7_75t_L g555 ( .A(n_437), .Y(n_555) );
AND2x2_ASAP7_75t_L g571 ( .A(n_437), .B(n_466), .Y(n_571) );
HB1xp67_ASAP7_75t_L g606 ( .A(n_437), .Y(n_606) );
AND2x2_ASAP7_75t_L g635 ( .A(n_437), .B(n_446), .Y(n_635) );
OA21x2_ASAP7_75t_L g437 ( .A1(n_438), .A2(n_439), .B(n_445), .Y(n_437) );
OA21x2_ASAP7_75t_L g466 ( .A1(n_438), .A2(n_467), .B(n_473), .Y(n_466) );
OA21x2_ASAP7_75t_L g478 ( .A1(n_438), .A2(n_479), .B(n_485), .Y(n_478) );
INVx2_ASAP7_75t_L g535 ( .A(n_446), .Y(n_535) );
BUFx3_ASAP7_75t_L g543 ( .A(n_446), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_446), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g554 ( .A(n_446), .B(n_555), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g583 ( .A(n_446), .B(n_455), .Y(n_583) );
AND2x2_ASAP7_75t_L g652 ( .A(n_446), .B(n_586), .Y(n_652) );
INVx2_ASAP7_75t_SL g546 ( .A(n_454), .Y(n_546) );
OR2x2_ASAP7_75t_L g454 ( .A(n_455), .B(n_466), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_455), .B(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g588 ( .A(n_455), .Y(n_588) );
AND2x2_ASAP7_75t_L g599 ( .A(n_455), .B(n_555), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_455), .B(n_584), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_455), .B(n_586), .Y(n_631) );
AND2x2_ASAP7_75t_L g690 ( .A(n_455), .B(n_635), .Y(n_690) );
INVx4_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g560 ( .A(n_456), .B(n_466), .Y(n_560) );
AND2x2_ASAP7_75t_L g570 ( .A(n_456), .B(n_571), .Y(n_570) );
BUFx3_ASAP7_75t_L g592 ( .A(n_456), .Y(n_592) );
AND3x2_ASAP7_75t_L g651 ( .A(n_456), .B(n_652), .C(n_653), .Y(n_651) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_466), .Y(n_542) );
INVx1_ASAP7_75t_SL g586 ( .A(n_466), .Y(n_586) );
NAND3xp33_ASAP7_75t_L g598 ( .A(n_466), .B(n_535), .C(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_508), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g621 ( .A1(n_475), .A2(n_570), .B(n_622), .C(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_477), .B(n_496), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_477), .B(n_628), .Y(n_627) );
INVx2_ASAP7_75t_SL g638 ( .A(n_477), .Y(n_638) );
AND2x2_ASAP7_75t_L g659 ( .A(n_477), .B(n_510), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g687 ( .A(n_477), .B(n_568), .Y(n_687) );
AND2x2_ASAP7_75t_L g477 ( .A(n_478), .B(n_486), .Y(n_477) );
AND2x2_ASAP7_75t_L g532 ( .A(n_478), .B(n_523), .Y(n_532) );
INVx2_ASAP7_75t_L g539 ( .A(n_478), .Y(n_539) );
AND2x2_ASAP7_75t_L g559 ( .A(n_478), .B(n_510), .Y(n_559) );
AND2x2_ASAP7_75t_L g609 ( .A(n_478), .B(n_496), .Y(n_609) );
INVx1_ASAP7_75t_L g613 ( .A(n_478), .Y(n_613) );
INVx2_ASAP7_75t_SL g523 ( .A(n_486), .Y(n_523) );
BUFx2_ASAP7_75t_L g549 ( .A(n_486), .Y(n_549) );
AND2x2_ASAP7_75t_L g676 ( .A(n_486), .B(n_496), .Y(n_676) );
INVx3_ASAP7_75t_SL g510 ( .A(n_496), .Y(n_510) );
AND2x2_ASAP7_75t_L g531 ( .A(n_496), .B(n_532), .Y(n_531) );
AND2x4_ASAP7_75t_L g538 ( .A(n_496), .B(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g568 ( .A(n_496), .B(n_528), .Y(n_568) );
OR2x2_ASAP7_75t_L g577 ( .A(n_496), .B(n_523), .Y(n_577) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_496), .Y(n_595) );
AND2x2_ASAP7_75t_L g600 ( .A(n_496), .B(n_553), .Y(n_600) );
AND2x2_ASAP7_75t_L g628 ( .A(n_496), .B(n_512), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_496), .B(n_664), .Y(n_663) );
OR2x2_ASAP7_75t_L g666 ( .A(n_496), .B(n_511), .Y(n_666) );
OR2x6_ASAP7_75t_L g496 ( .A(n_497), .B(n_506), .Y(n_496) );
INVx2_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g517 ( .A(n_504), .B(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x2_ASAP7_75t_L g509 ( .A(n_510), .B(n_511), .Y(n_509) );
AND2x2_ASAP7_75t_L g590 ( .A(n_510), .B(n_539), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_510), .B(n_532), .Y(n_618) );
AND2x2_ASAP7_75t_L g636 ( .A(n_510), .B(n_553), .Y(n_636) );
OR2x2_ASAP7_75t_L g511 ( .A(n_512), .B(n_523), .Y(n_511) );
AND2x2_ASAP7_75t_L g537 ( .A(n_512), .B(n_523), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_512), .B(n_566), .Y(n_565) );
BUFx3_ASAP7_75t_L g575 ( .A(n_512), .Y(n_575) );
OR2x2_ASAP7_75t_L g623 ( .A(n_512), .B(n_543), .Y(n_623) );
OA21x2_ASAP7_75t_L g512 ( .A1(n_513), .A2(n_514), .B(n_521), .Y(n_512) );
INVx1_ASAP7_75t_L g529 ( .A(n_514), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_521), .Y(n_530) );
AND2x2_ASAP7_75t_L g558 ( .A(n_523), .B(n_528), .Y(n_558) );
INVx1_ASAP7_75t_L g566 ( .A(n_523), .Y(n_566) );
AND2x2_ASAP7_75t_L g661 ( .A(n_523), .B(n_539), .Y(n_661) );
AOI222xp33_ASAP7_75t_L g524 ( .A1(n_525), .A2(n_533), .B1(n_536), .B2(n_540), .C1(n_544), .C2(n_547), .Y(n_524) );
INVx1_ASAP7_75t_L g656 ( .A(n_525), .Y(n_656) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_531), .Y(n_525) );
AND2x2_ASAP7_75t_L g552 ( .A(n_526), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_L g563 ( .A(n_526), .B(n_532), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_526), .B(n_554), .Y(n_579) );
OAI222xp33_ASAP7_75t_L g601 ( .A1(n_526), .A2(n_602), .B1(n_607), .B2(n_608), .C1(n_616), .C2(n_618), .Y(n_601) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx1_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g589 ( .A(n_528), .B(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_528), .B(n_609), .Y(n_649) );
AND2x2_ASAP7_75t_L g660 ( .A(n_528), .B(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g668 ( .A(n_531), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g647 ( .A(n_533), .B(n_584), .Y(n_647) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_535), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g605 ( .A(n_535), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_538), .Y(n_536) );
INVx3_ASAP7_75t_L g550 ( .A(n_538), .Y(n_550) );
O2A1O1Ixp33_ASAP7_75t_L g640 ( .A1(n_538), .A2(n_641), .B(n_644), .C(n_646), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_538), .B(n_575), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_538), .B(n_558), .Y(n_680) );
AND2x2_ASAP7_75t_L g553 ( .A(n_539), .B(n_549), .Y(n_553) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .Y(n_541) );
INVx1_ASAP7_75t_L g580 ( .A(n_542), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_543), .B(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g632 ( .A(n_543), .B(n_633), .Y(n_632) );
AND2x2_ASAP7_75t_L g671 ( .A(n_543), .B(n_571), .Y(n_671) );
INVx1_ASAP7_75t_L g683 ( .A(n_543), .Y(n_683) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_546), .B(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g547 ( .A(n_548), .Y(n_547) );
OR2x2_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .Y(n_548) );
INVx1_ASAP7_75t_L g664 ( .A(n_549), .Y(n_664) );
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_552), .A2(n_554), .B(n_556), .C(n_560), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g596 ( .A1(n_552), .A2(n_582), .B1(n_597), .B2(n_600), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_553), .B(n_567), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_553), .B(n_575), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_554), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_SL g617 ( .A(n_554), .Y(n_617) );
AND2x2_ASAP7_75t_L g624 ( .A(n_554), .B(n_604), .Y(n_624) );
INVx2_ASAP7_75t_L g585 ( .A(n_555), .Y(n_585) );
INVxp67_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NOR4xp25_ASAP7_75t_L g562 ( .A(n_559), .B(n_563), .C(n_564), .D(n_567), .Y(n_562) );
INVx1_ASAP7_75t_SL g633 ( .A(n_560), .Y(n_633) );
AND2x2_ASAP7_75t_L g677 ( .A(n_560), .B(n_678), .Y(n_677) );
OAI211xp5_ASAP7_75t_SL g561 ( .A1(n_562), .A2(n_569), .B(n_572), .C(n_581), .Y(n_561) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_SL g567 ( .A(n_568), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_568), .B(n_638), .Y(n_689) );
AOI22xp5_ASAP7_75t_L g688 ( .A1(n_570), .A2(n_689), .B1(n_690), .B2(n_691), .Y(n_688) );
INVx1_ASAP7_75t_SL g643 ( .A(n_571), .Y(n_643) );
AND2x2_ASAP7_75t_L g682 ( .A(n_571), .B(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_576), .Y(n_574) );
NAND2xp5_ASAP7_75t_SL g675 ( .A(n_575), .B(n_676), .Y(n_675) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g594 ( .A(n_579), .B(n_595), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_580), .B(n_605), .Y(n_665) );
OAI21xp5_ASAP7_75t_SL g581 ( .A1(n_582), .A2(n_587), .B(n_589), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_583), .B(n_584), .Y(n_582) );
INVx1_ASAP7_75t_L g657 ( .A(n_584), .Y(n_657) );
AND2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g685 ( .A(n_585), .Y(n_685) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_586), .Y(n_612) );
OAI21xp33_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_593), .B(n_596), .Y(n_591) );
CKINVDCx16_ASAP7_75t_R g604 ( .A(n_592), .Y(n_604) );
OR2x2_ASAP7_75t_L g642 ( .A(n_592), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
AOI21xp33_ASAP7_75t_SL g637 ( .A1(n_595), .A2(n_638), .B(n_639), .Y(n_637) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_599), .A2(n_626), .B1(n_629), .B2(n_636), .C(n_637), .Y(n_625) );
INVx1_ASAP7_75t_SL g669 ( .A(n_600), .Y(n_669) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .Y(n_603) );
OR2x2_ASAP7_75t_L g616 ( .A(n_604), .B(n_617), .Y(n_616) );
INVxp67_ASAP7_75t_L g653 ( .A(n_606), .Y(n_653) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_613), .B2(n_614), .Y(n_608) );
INVx1_ASAP7_75t_L g648 ( .A(n_609), .Y(n_648) );
INVxp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_612), .B(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
NOR4xp25_ASAP7_75t_L g619 ( .A(n_620), .B(n_654), .C(n_667), .D(n_679), .Y(n_619) );
NAND3xp33_ASAP7_75t_SL g620 ( .A(n_621), .B(n_625), .C(n_640), .Y(n_620) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_623), .B(n_642), .Y(n_641) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_630), .B(n_635), .Y(n_639) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
OAI221xp5_ASAP7_75t_SL g667 ( .A1(n_642), .A2(n_668), .B1(n_669), .B2(n_670), .C(n_672), .Y(n_667) );
O2A1O1Ixp33_ASAP7_75t_L g658 ( .A1(n_644), .A2(n_659), .B(n_660), .C(n_662), .Y(n_658) );
INVx2_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_645), .A2(n_663), .B1(n_665), .B2(n_666), .Y(n_662) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_656), .B(n_657), .C(n_658), .Y(n_654) );
INVx1_ASAP7_75t_L g673 ( .A(n_666), .Y(n_673) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
OAI21xp5_ASAP7_75t_SL g672 ( .A1(n_673), .A2(n_674), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI221xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_681), .B1(n_684), .B2(n_686), .C(n_688), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVxp67_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g703 ( .A(n_693), .Y(n_703) );
INVx1_ASAP7_75t_L g705 ( .A(n_694), .Y(n_705) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx3_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g702 ( .A(n_703), .Y(n_702) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_708), .B(n_710), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
OAI21xp5_ASAP7_75t_SL g711 ( .A1(n_712), .A2(n_717), .B(n_720), .Y(n_711) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_713), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_SL g718 ( .A(n_719), .Y(n_718) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_722), .Y(n_721) );
endmodule