module fake_jpeg_31326_n_323 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_323);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_323;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_12),
.B(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_15),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_10),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_3),
.B(n_12),
.Y(n_40)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_48),
.Y(n_107)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_50),
.B(n_55),
.Y(n_118)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

INVx3_ASAP7_75t_SL g115 ( 
.A(n_52),
.Y(n_115)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_53),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_19),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_56),
.B(n_69),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

INVx6_ASAP7_75t_L g109 ( 
.A(n_57),
.Y(n_109)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_61),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_36),
.Y(n_63)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_63),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_23),
.B(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_64),
.B(n_67),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx6_ASAP7_75t_L g134 ( 
.A(n_65),
.Y(n_134)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_34),
.B(n_10),
.Y(n_67)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_68),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_26),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx13_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_28),
.B(n_11),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_71),
.B(n_73),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_26),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_72),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_36),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_31),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_75),
.Y(n_132)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_17),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_19),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_76),
.B(n_78),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_77),
.B(n_80),
.Y(n_130)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx11_ASAP7_75t_SL g79 ( 
.A(n_31),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_79),
.Y(n_108)
);

NAND2x1_ASAP7_75t_SL g80 ( 
.A(n_31),
.B(n_0),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_99)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_82),
.B(n_85),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_18),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_46),
.Y(n_84)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_37),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_93),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_30),
.B(n_11),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_92),
.Y(n_127)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_25),
.Y(n_89)
);

AOI21xp33_ASAP7_75t_L g126 ( 
.A1(n_89),
.A2(n_16),
.B(n_2),
.Y(n_126)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_33),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_22),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_25),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_35),
.B(n_12),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_94),
.B(n_95),
.Y(n_128)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_33),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_96),
.A2(n_42),
.B1(n_2),
.B2(n_1),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_24),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_94),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_47),
.B1(n_43),
.B2(n_29),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_98),
.A2(n_103),
.B1(n_104),
.B2(n_113),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_57),
.A2(n_47),
.B1(n_43),
.B2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_49),
.A2(n_24),
.B1(n_33),
.B2(n_42),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_77),
.A2(n_33),
.B1(n_42),
.B2(n_6),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_114),
.A2(n_116),
.B1(n_117),
.B2(n_119),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_54),
.A2(n_42),
.B1(n_13),
.B2(n_6),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_84),
.A2(n_6),
.B1(n_9),
.B2(n_14),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_81),
.A2(n_14),
.B1(n_16),
.B2(n_1),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_90),
.B1(n_70),
.B2(n_72),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_122),
.A2(n_124),
.B1(n_138),
.B2(n_140),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_79),
.A2(n_14),
.B1(n_16),
.B2(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_131),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_80),
.A2(n_62),
.B1(n_65),
.B2(n_67),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_71),
.A2(n_88),
.B1(n_64),
.B2(n_74),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_89),
.A2(n_44),
.B1(n_25),
.B2(n_45),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_146),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_49),
.A2(n_44),
.B1(n_25),
.B2(n_45),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_49),
.A2(n_44),
.B1(n_25),
.B2(n_45),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_49),
.A2(n_44),
.B1(n_25),
.B2(n_45),
.Y(n_146)
);

INVx5_ASAP7_75t_L g148 ( 
.A(n_142),
.Y(n_148)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_148),
.Y(n_191)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_121),
.Y(n_149)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_149),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_127),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_150),
.B(n_152),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_133),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_154),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_133),
.B(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_155),
.B(n_156),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_128),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_128),
.B(n_136),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_158),
.B(n_159),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_118),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_139),
.B(n_125),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_162),
.B(n_169),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_163),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_115),
.A2(n_107),
.B1(n_101),
.B2(n_100),
.Y(n_164)
);

INVx13_ASAP7_75t_L g183 ( 
.A(n_164),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_112),
.Y(n_165)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_165),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_129),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_166),
.B(n_167),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_123),
.Y(n_167)
);

INVx13_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_130),
.B(n_123),
.Y(n_169)
);

CKINVDCx12_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_174),
.Y(n_182)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_109),
.Y(n_171)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_171),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_137),
.B(n_103),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_172),
.B(n_120),
.C(n_106),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_132),
.B(n_115),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_173),
.B(n_176),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx14_ASAP7_75t_R g175 ( 
.A(n_135),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_177),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_115),
.B(n_108),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g178 ( 
.A(n_126),
.B(n_101),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_178),
.B(n_111),
.Y(n_201)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_179),
.B(n_180),
.Y(n_189)
);

INVx13_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_169),
.A2(n_102),
.B(n_99),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_186),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_178),
.A2(n_113),
.B(n_104),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_152),
.B(n_156),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_196),
.B(n_200),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_155),
.B(n_108),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_207),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_157),
.A2(n_105),
.B1(n_112),
.B2(n_134),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_161),
.B1(n_160),
.B2(n_147),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_162),
.B(n_110),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_173),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_167),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_207),
.A2(n_157),
.B1(n_166),
.B2(n_172),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_208),
.A2(n_203),
.B1(n_206),
.B2(n_205),
.Y(n_230)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_194),
.Y(n_209)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_209),
.Y(n_229)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g242 ( 
.A(n_211),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_150),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_212),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_195),
.Y(n_213)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_213),
.Y(n_235)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_195),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_215),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_184),
.B(n_158),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_220),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_184),
.B(n_197),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_188),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_181),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_198),
.B(n_151),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_222),
.B(n_223),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_181),
.B(n_159),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_224),
.A2(n_183),
.B1(n_188),
.B2(n_189),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_151),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_225),
.B(n_227),
.Y(n_239)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_199),
.Y(n_227)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_200),
.B(n_196),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g236 ( 
.A(n_228),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_231),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_208),
.A2(n_190),
.B1(n_205),
.B2(n_186),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_237),
.A2(n_238),
.B1(n_246),
.B2(n_215),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_226),
.A2(n_186),
.B1(n_201),
.B2(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_219),
.B(n_192),
.C(n_204),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_244),
.C(n_225),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_192),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_221),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_199),
.C(n_153),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_209),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_238),
.A2(n_216),
.B(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_247),
.B(n_249),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_228),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_251),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_252),
.B(n_257),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_236),
.A2(n_216),
.B(n_218),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_253),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_233),
.B(n_223),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_255),
.A2(n_256),
.B1(n_261),
.B2(n_257),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_233),
.B(n_239),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_239),
.B(n_210),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_212),
.C(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_259),
.C(n_244),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_222),
.C(n_217),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_260),
.A2(n_213),
.B1(n_214),
.B2(n_242),
.Y(n_275)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_235),
.Y(n_261)
);

AO21x2_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_183),
.B(n_224),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_262),
.A2(n_234),
.B1(n_237),
.B2(n_189),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_263),
.B(n_266),
.C(n_269),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_264),
.B(n_262),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_254),
.A2(n_262),
.B1(n_253),
.B2(n_250),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_265),
.B(n_271),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_241),
.C(n_232),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_258),
.B(n_232),
.C(n_230),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_259),
.B(n_210),
.C(n_227),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_270),
.B(n_182),
.C(n_248),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_275),
.A2(n_262),
.B1(n_229),
.B2(n_211),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_254),
.A2(n_242),
.B1(n_229),
.B2(n_187),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_276),
.B(n_187),
.Y(n_287)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_274),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_277),
.B(n_282),
.Y(n_296)
);

OAI322xp33_ASAP7_75t_L g278 ( 
.A1(n_272),
.A2(n_255),
.A3(n_247),
.B1(n_260),
.B2(n_262),
.C1(n_251),
.C2(n_261),
.Y(n_278)
);

BUFx24_ASAP7_75t_SL g289 ( 
.A(n_278),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_281),
.B(n_283),
.C(n_288),
.Y(n_294)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_274),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_248),
.C(n_262),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_284),
.A2(n_286),
.B1(n_276),
.B2(n_268),
.Y(n_293)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_272),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_285),
.B(n_287),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_182),
.C(n_202),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_273),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_279),
.C(n_288),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_265),
.B(n_264),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_292),
.B(n_295),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_297),
.B1(n_194),
.B2(n_191),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_269),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_267),
.B1(n_275),
.B2(n_270),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_289),
.A2(n_284),
.B1(n_281),
.B2(n_266),
.Y(n_300)
);

OR2x2_ASAP7_75t_L g307 ( 
.A(n_300),
.B(n_290),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_295),
.B(n_202),
.C(n_193),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_296),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_303),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_294),
.B(n_185),
.C(n_177),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_304),
.B(n_294),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_299),
.B(n_291),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g311 ( 
.A1(n_305),
.A2(n_298),
.B(n_163),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_307),
.Y(n_313)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_308),
.B(n_191),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_309),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_313),
.A3(n_148),
.B1(n_180),
.B2(n_170),
.C1(n_168),
.C2(n_171),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_314),
.B1(n_179),
.B2(n_154),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_305),
.A2(n_187),
.B1(n_154),
.B2(n_171),
.Y(n_314)
);

AOI21xp33_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_310),
.B(n_306),
.Y(n_316)
);

AOI21x1_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_317),
.B(n_180),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g320 ( 
.A(n_318),
.B(n_179),
.CI(n_193),
.CON(n_320),
.SN(n_320)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_319),
.Y(n_321)
);

NOR3xp33_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_320),
.C(n_174),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_322),
.B(n_148),
.Y(n_323)
);


endmodule