module real_jpeg_33980_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_578;
wire n_328;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_546;
wire n_285;
wire n_172;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx2_ASAP7_75t_L g112 ( 
.A(n_0),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_0),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g258 ( 
.A(n_0),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_0),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g412 ( 
.A(n_0),
.Y(n_412)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_1),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_41),
.Y(n_40)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_2),
.B(n_55),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g94 ( 
.A(n_2),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_2),
.B(n_208),
.Y(n_207)
);

NAND2x1_ASAP7_75t_L g255 ( 
.A(n_2),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_2),
.B(n_346),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_2),
.B(n_510),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_3),
.B(n_35),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_3),
.B(n_89),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_3),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g173 ( 
.A(n_3),
.B(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_3),
.B(n_236),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_3),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

AND2x2_ASAP7_75t_L g458 ( 
.A(n_3),
.B(n_459),
.Y(n_458)
);

AND2x4_ASAP7_75t_SL g166 ( 
.A(n_4),
.B(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_4),
.B(n_178),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_4),
.B(n_170),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g314 ( 
.A(n_4),
.B(n_315),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g341 ( 
.A(n_4),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_4),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_4),
.B(n_236),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_4),
.B(n_453),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_5),
.B(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_5),
.B(n_263),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_5),
.B(n_289),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_5),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_5),
.B(n_402),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_5),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_5),
.B(n_426),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_6),
.B(n_77),
.Y(n_76)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_6),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_6),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_6),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_6),
.B(n_63),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_7),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g157 ( 
.A(n_7),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_7),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_8),
.Y(n_44)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_8),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_9),
.Y(n_82)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_9),
.Y(n_151)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_9),
.Y(n_324)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_9),
.Y(n_347)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_10),
.Y(n_274)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_10),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_11),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_11),
.B(n_89),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_11),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_11),
.B(n_268),
.Y(n_267)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_11),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_11),
.B(n_236),
.Y(n_349)
);

AND2x4_ASAP7_75t_SL g463 ( 
.A(n_11),
.B(n_464),
.Y(n_463)
);

AND2x4_ASAP7_75t_SL g507 ( 
.A(n_11),
.B(n_508),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_12),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_12),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_12),
.B(n_245),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_12),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_12),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_12),
.B(n_232),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_12),
.B(n_474),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_13),
.A2(n_15),
.B1(n_21),
.B2(n_24),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_14),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_14),
.B(n_252),
.Y(n_251)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_14),
.B(n_101),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_14),
.B(n_297),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_14),
.B(n_366),
.Y(n_365)
);

AND2x2_ASAP7_75t_L g377 ( 
.A(n_14),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_14),
.B(n_411),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_14),
.B(n_245),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_16),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_16),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_16),
.Y(n_134)
);

NAND2x1_ASAP7_75t_L g169 ( 
.A(n_16),
.B(n_170),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_16),
.B(n_200),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_16),
.B(n_302),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_16),
.B(n_321),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_16),
.B(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_17),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_17),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g270 ( 
.A(n_17),
.Y(n_270)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_18),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_18),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_18),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_19),
.B(n_46),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_19),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_19),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_19),
.B(n_479),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

BUFx12f_ASAP7_75t_SL g22 ( 
.A(n_23),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_219),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_R g25 ( 
.A(n_26),
.B(n_217),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_183),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_27),
.B(n_183),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_120),
.C(n_138),
.Y(n_27)
);

HB1xp67_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_29),
.B(n_120),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_84),
.B1(n_85),
.B2(n_119),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_30),
.B(n_105),
.C(n_185),
.Y(n_184)
);

MAJx2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_50),
.C(n_67),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_50),
.C(n_67),
.Y(n_119)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

XNOR2xp5_ASAP7_75t_L g531 ( 
.A(n_32),
.B(n_51),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_34),
.B(n_124),
.C(n_125),
.Y(n_123)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_38),
.Y(n_137)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_38),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_45),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_40),
.Y(n_124)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_44),
.Y(n_317)
);

BUFx6f_ASAP7_75t_L g465 ( 
.A(n_44),
.Y(n_465)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_45),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_49),
.Y(n_299)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_61),
.B(n_66),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_56),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_56),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_53),
.A2(n_54),
.B1(n_62),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_58),
.Y(n_56)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_59),
.Y(n_286)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_59),
.Y(n_342)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_59),
.Y(n_399)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_60),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g175 ( 
.A(n_65),
.Y(n_175)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_67),
.Y(n_532)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_74),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_68),
.B(n_75),
.C(n_83),
.Y(n_122)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g70 ( 
.A(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_76),
.B1(n_79),
.B2(n_83),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_76),
.B1(n_128),
.B2(n_132),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_76),
.B(n_192),
.C(n_193),
.Y(n_191)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_79),
.B(n_107),
.C(n_110),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_79),
.A2(n_83),
.B1(n_110),
.B2(n_152),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_79),
.B(n_107),
.C(n_110),
.Y(n_182)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx6_ASAP7_75t_L g309 ( 
.A(n_82),
.Y(n_309)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_104),
.B2(n_105),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g185 ( 
.A(n_86),
.Y(n_185)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

XOR2x1_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_93),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_88),
.B(n_94),
.C(n_100),
.Y(n_205)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

XNOR2x1_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_100),
.Y(n_93)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_99),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_99),
.Y(n_290)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

MAJx2_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_113),
.C(n_117),
.Y(n_105)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_109),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_110),
.B(n_148),
.Y(n_495)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_111),
.Y(n_427)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_164),
.C(n_176),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_113),
.B(n_118),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_113),
.A2(n_176),
.B1(n_177),
.B2(n_546),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_113),
.Y(n_546)
);

INVx3_ASAP7_75t_SL g114 ( 
.A(n_115),
.Y(n_114)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_115),
.Y(n_453)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx8_ASAP7_75t_L g254 ( 
.A(n_116),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_126),
.Y(n_120)
);

XNOR2xp5_ASAP7_75t_L g121 ( 
.A(n_122),
.B(n_123),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_122),
.B(n_123),
.C(n_126),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_127),
.B(n_133),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_128),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_128),
.A2(n_132),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_133),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_138),
.B(n_577),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_161),
.C(n_179),
.Y(n_138)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_140),
.B(n_528),
.Y(n_527)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_146),
.C(n_158),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_142),
.B(n_554),
.Y(n_553)
);

XNOR2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_146),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.C(n_153),
.Y(n_146)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_150),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

OA22x2_ASAP7_75t_L g494 ( 
.A1(n_153),
.A2(n_495),
.B1(n_496),
.B2(n_497),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_153),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g541 ( 
.A(n_153),
.B(n_496),
.Y(n_541)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx4_ASAP7_75t_SL g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_157),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_158),
.B(n_553),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_160),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g528 ( 
.A1(n_162),
.A2(n_163),
.B1(n_180),
.B2(n_529),
.Y(n_528)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_169),
.C(n_172),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_165),
.B(n_169),
.C(n_172),
.Y(n_547)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_166),
.B(n_173),
.Y(n_491)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_169),
.B(n_491),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_169),
.B(n_491),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_171),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g172 ( 
.A(n_173),
.Y(n_172)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_180),
.Y(n_529)
);

XOR2x1_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_182),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

XNOR2x1_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_188),
.Y(n_186)
);

XNOR2x1_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_204),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_195),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

XOR2x2_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_203),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g474 ( 
.A(n_203),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.Y(n_206)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx8_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g508 ( 
.A(n_216),
.Y(n_508)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_578),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_570),
.Y(n_220)
);

OAI21x1_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_523),
.B(n_567),
.Y(n_221)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_439),
.B(n_521),
.Y(n_222)
);

OAI21x1_ASAP7_75t_SL g223 ( 
.A1(n_224),
.A2(n_353),
.B(n_437),
.Y(n_223)
);

NOR3xp33_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_332),
.C(n_335),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_226),
.B(n_333),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_277),
.Y(n_226)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_227),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_227),
.B(n_519),
.C(n_520),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_249),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_228),
.B(n_250),
.C(n_260),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_238),
.C(n_243),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_229),
.B(n_352),
.Y(n_351)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_234),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_230),
.A2(n_231),
.B1(n_234),
.B2(n_235),
.Y(n_339)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_237),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_238),
.A2(n_239),
.B1(n_243),
.B2(n_244),
.Y(n_352)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_260),
.Y(n_249)
);

OA21x2_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_255),
.B(n_259),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_251),
.B(n_255),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx8_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g481 ( 
.A1(n_259),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.Y(n_481)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_259),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_SL g499 ( 
.A(n_259),
.B(n_472),
.C(n_483),
.Y(n_499)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_266),
.Y(n_260)
);

HB1xp67_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_262),
.Y(n_446)
);

BUFx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_271),
.B1(n_275),
.B2(n_276),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_267),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_267),
.B(n_275),
.C(n_446),
.Y(n_445)
);

INVx3_ASAP7_75t_SL g268 ( 
.A(n_269),
.Y(n_268)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_269),
.Y(n_402)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g363 ( 
.A(n_270),
.Y(n_363)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_271),
.Y(n_275)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_274),
.Y(n_451)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_278),
.B(n_334),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_311),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g519 ( 
.A(n_279),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_287),
.C(n_300),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_280),
.B(n_337),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJx2_ASAP7_75t_L g329 ( 
.A(n_281),
.B(n_283),
.C(n_284),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_287),
.B(n_300),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_291),
.C(n_296),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_288),
.B(n_291),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_295),
.Y(n_374)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_296),
.Y(n_391)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

BUFx3_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_305),
.B1(n_306),
.B2(n_310),
.Y(n_300)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_301),
.Y(n_310)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_310),
.Y(n_328)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

HB1xp67_ASAP7_75t_L g520 ( 
.A(n_311),
.Y(n_520)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_312),
.B(n_327),
.Y(n_311)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_312),
.B(n_328),
.C(n_331),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_318),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_314),
.B(n_320),
.C(n_325),
.Y(n_482)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_325),
.B2(n_326),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_322),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_330),
.B2(n_331),
.Y(n_327)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_329),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_335),
.B(n_438),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_338),
.C(n_350),
.Y(n_335)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_336),
.B(n_435),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_338),
.B(n_351),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.C(n_343),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_339),
.B(n_340),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_343),
.B(n_383),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_348),
.Y(n_343)
);

AO22x1_ASAP7_75t_SL g380 ( 
.A1(n_344),
.A2(n_345),
.B1(n_348),
.B2(n_349),
.Y(n_380)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_354),
.A2(n_432),
.B(n_436),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_355),
.A2(n_393),
.B(n_431),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_381),
.Y(n_355)
);

OR2x2_ASAP7_75t_L g431 ( 
.A(n_356),
.B(n_381),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_375),
.C(n_380),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_357),
.A2(n_358),
.B1(n_404),
.B2(n_406),
.Y(n_403)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_SL g358 ( 
.A(n_359),
.B(n_364),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_359),
.B(n_387),
.C(n_388),
.Y(n_386)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_370),
.Y(n_364)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_365),
.Y(n_388)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

BUFx3_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g513 ( 
.A(n_369),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_375),
.A2(n_376),
.B1(n_380),
.B2(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_379),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_377),
.B(n_379),
.Y(n_396)
);

INVx1_ASAP7_75t_SL g405 ( 
.A(n_380),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_382),
.A2(n_384),
.B1(n_385),
.B2(n_392),
.Y(n_381)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_382),
.Y(n_392)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_SL g385 ( 
.A(n_386),
.B(n_389),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_386),
.B(n_389),
.C(n_392),
.Y(n_433)
);

XOR2x1_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_391),
.Y(n_389)
);

AOI21x1_ASAP7_75t_SL g393 ( 
.A1(n_394),
.A2(n_407),
.B(n_430),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_403),
.Y(n_394)
);

NOR2xp67_ASAP7_75t_SL g430 ( 
.A(n_395),
.B(n_403),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_396),
.B(n_397),
.C(n_400),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_396),
.B(n_415),
.Y(n_414)
);

AOI22xp33_ASAP7_75t_L g415 ( 
.A1(n_397),
.A2(n_398),
.B1(n_400),
.B2(n_401),
.Y(n_415)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_404),
.Y(n_406)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_408),
.A2(n_416),
.B(n_429),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_414),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g429 ( 
.A(n_409),
.B(n_414),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_410),
.B(n_413),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_413),
.Y(n_423)
);

BUFx4f_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g424 ( 
.A(n_413),
.B(n_425),
.Y(n_424)
);

AOI21xp5_ASAP7_75t_L g416 ( 
.A1(n_417),
.A2(n_424),
.B(n_428),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_423),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_423),
.Y(n_428)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

NAND2xp33_ASAP7_75t_SL g432 ( 
.A(n_433),
.B(n_434),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_434),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_440),
.A2(n_485),
.B(n_515),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_440),
.B(n_485),
.C(n_522),
.Y(n_521)
);

MAJx2_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_468),
.C(n_470),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_441),
.B(n_517),
.Y(n_516)
);

XOR2xp5_ASAP7_75t_SL g441 ( 
.A(n_442),
.B(n_443),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_442),
.B(n_444),
.C(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_444),
.B(n_456),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_445),
.B(n_447),
.Y(n_444)
);

A2O1A1Ixp33_ASAP7_75t_L g501 ( 
.A1(n_445),
.A2(n_452),
.B(n_455),
.C(n_502),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_448),
.A2(n_452),
.B1(n_454),
.B2(n_455),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g455 ( 
.A(n_448),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_448),
.B(n_454),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g449 ( 
.A(n_450),
.Y(n_449)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_452),
.Y(n_454)
);

HB1xp67_ASAP7_75t_L g487 ( 
.A(n_456),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_461),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_SL g540 ( 
.A(n_457),
.B(n_462),
.C(n_466),
.Y(n_540)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

MAJx2_ASAP7_75t_L g493 ( 
.A(n_458),
.B(n_463),
.C(n_467),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_460),
.Y(n_459)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_462),
.A2(n_463),
.B1(n_466),
.B2(n_467),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_463),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_466),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XOR2xp5_ASAP7_75t_L g517 ( 
.A(n_469),
.B(n_471),
.Y(n_517)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_472),
.B(n_481),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_473),
.B(n_475),
.Y(n_472)
);

MAJx2_ASAP7_75t_L g504 ( 
.A(n_473),
.B(n_477),
.C(n_480),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_478),
.B2(n_480),
.Y(n_475)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_476),
.Y(n_480)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_482),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_488),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g561 ( 
.A(n_486),
.B(n_562),
.C(n_563),
.Y(n_561)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_498),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_489),
.Y(n_563)
);

XNOR2x1_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_492),
.Y(n_489)
);

XNOR2x1_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_494),
.Y(n_492)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_493),
.Y(n_543)
);

AO22x1_ASAP7_75t_L g537 ( 
.A1(n_494),
.A2(n_538),
.B1(n_539),
.B2(n_543),
.Y(n_537)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_495),
.B(n_497),
.Y(n_542)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_498),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_R g555 ( 
.A(n_499),
.B(n_556),
.C(n_557),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g566 ( 
.A(n_499),
.B(n_556),
.C(n_557),
.Y(n_566)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_501),
.B(n_503),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g556 ( 
.A(n_501),
.Y(n_556)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_503),
.Y(n_557)
);

XNOR2x1_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_505),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_507),
.C(n_550),
.Y(n_549)
);

OAI22x1_ASAP7_75t_L g505 ( 
.A1(n_506),
.A2(n_507),
.B1(n_509),
.B2(n_514),
.Y(n_505)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_507),
.Y(n_506)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_509),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g550 ( 
.A(n_509),
.Y(n_550)
);

INVx3_ASAP7_75t_L g510 ( 
.A(n_511),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_512),
.Y(n_511)
);

INVx3_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_516),
.B(n_518),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_516),
.B(n_518),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_560),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_524),
.A2(n_568),
.B(n_569),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_525),
.B(n_551),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_525),
.B(n_551),
.Y(n_569)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_535),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_530),
.B1(n_533),
.B2(n_534),
.Y(n_526)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_527),
.Y(n_534)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_530),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_530),
.Y(n_575)
);

XOR2x1_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g573 ( 
.A(n_534),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_535),
.Y(n_574)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_544),
.C(n_548),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_537),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_537),
.B(n_559),
.Y(n_558)
);

NAND3xp33_ASAP7_75t_L g539 ( 
.A(n_540),
.B(n_541),
.C(n_542),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_544),
.B(n_549),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_545),
.B(n_547),
.Y(n_544)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_552),
.B(n_555),
.C(n_558),
.Y(n_551)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_566),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_565),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_561),
.B(n_564),
.Y(n_560)
);

NOR2xp67_ASAP7_75t_L g568 ( 
.A(n_561),
.B(n_564),
.Y(n_568)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_572),
.B(n_576),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_L g580 ( 
.A(n_572),
.B(n_576),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_573),
.B(n_574),
.C(n_575),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

HB1xp67_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);


endmodule