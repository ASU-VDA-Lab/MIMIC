module fake_netlist_6_4221_n_603 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_186, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_603);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_186;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_603;

wire n_591;
wire n_435;
wire n_326;
wire n_256;
wire n_440;
wire n_587;
wire n_507;
wire n_580;
wire n_209;
wire n_367;
wire n_465;
wire n_590;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_208;
wire n_462;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_578;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_524;
wire n_342;
wire n_358;
wire n_449;
wire n_188;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_396;
wire n_495;
wire n_350;
wire n_585;
wire n_568;
wire n_392;
wire n_442;
wire n_480;
wire n_382;
wire n_557;
wire n_349;
wire n_233;
wire n_255;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_471;
wire n_289;
wire n_421;
wire n_424;
wire n_238;
wire n_573;
wire n_202;
wire n_320;
wire n_327;
wire n_369;
wire n_597;
wire n_280;
wire n_287;
wire n_353;
wire n_555;
wire n_389;
wire n_415;
wire n_230;
wire n_461;
wire n_383;
wire n_200;
wire n_447;
wire n_198;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_229;
wire n_542;
wire n_305;
wire n_532;
wire n_535;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_510;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_506;
wire n_360;
wire n_235;
wire n_536;
wire n_191;
wire n_340;
wire n_387;
wire n_452;
wire n_344;
wire n_581;
wire n_428;
wire n_432;
wire n_516;
wire n_525;
wire n_491;
wire n_371;
wire n_567;
wire n_189;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_197;
wire n_343;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_529;
wire n_445;
wire n_425;
wire n_454;
wire n_218;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_490;
wire n_290;
wire n_220;
wire n_224;
wire n_196;
wire n_402;
wire n_352;
wire n_478;
wire n_574;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_374;
wire n_366;
wire n_407;
wire n_450;
wire n_272;
wire n_526;
wire n_348;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_330;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_279;
wire n_252;
wire n_228;
wire n_565;
wire n_594;
wire n_356;
wire n_577;
wire n_552;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_592;
wire n_323;
wire n_393;
wire n_411;
wire n_503;
wire n_599;
wire n_513;
wire n_321;
wire n_331;
wire n_227;
wire n_570;
wire n_406;
wire n_483;
wire n_204;
wire n_482;
wire n_474;
wire n_527;
wire n_261;
wire n_420;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_476;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_325;
wire n_329;
wire n_464;
wire n_600;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_211;
wire n_523;
wire n_322;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_505;
wire n_240;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_311;
wire n_403;
wire n_253;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_556;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_560;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_444;
wire n_586;
wire n_423;
wire n_318;
wire n_303;
wire n_511;
wire n_467;
wire n_306;
wire n_269;
wire n_193;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_571;
wire n_268;
wire n_404;
wire n_271;
wire n_439;
wire n_217;
wire n_210;
wire n_518;
wire n_299;
wire n_206;
wire n_453;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_355;
wire n_426;
wire n_317;
wire n_431;
wire n_347;
wire n_459;
wire n_502;
wire n_328;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_257;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_242;
wire n_401;
wire n_324;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_251;
wire n_301;
wire n_274;
wire n_412;
wire n_267;
wire n_438;
wire n_339;
wire n_434;
wire n_515;
wire n_315;
wire n_427;
wire n_288;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_528;
wire n_391;
wire n_457;
wire n_364;
wire n_385;
wire n_295;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_501;
wire n_531;
wire n_361;
wire n_508;
wire n_379;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_192;
wire n_283;

INVx1_ASAP7_75t_L g188 ( 
.A(n_61),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_75),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_175),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_110),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_16),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_19),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_74),
.Y(n_194)
);

INVxp33_ASAP7_75t_SL g195 ( 
.A(n_122),
.Y(n_195)
);

INVxp33_ASAP7_75t_SL g196 ( 
.A(n_51),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_62),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_35),
.Y(n_198)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_162),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_31),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_154),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_106),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_84),
.Y(n_206)
);

INVxp67_ASAP7_75t_SL g207 ( 
.A(n_6),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_47),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVxp67_ASAP7_75t_SL g210 ( 
.A(n_83),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_96),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVxp67_ASAP7_75t_SL g213 ( 
.A(n_142),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_45),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_120),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_136),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_173),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_53),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_39),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_99),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_2),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_4),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_20),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_95),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_5),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_128),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_50),
.Y(n_227)
);

INVxp67_ASAP7_75t_SL g228 ( 
.A(n_42),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_68),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_121),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_135),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_43),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_87),
.Y(n_233)
);

BUFx2_ASAP7_75t_L g234 ( 
.A(n_151),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_181),
.Y(n_235)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_176),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_105),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_161),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_138),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_149),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_126),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_91),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_11),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_146),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_112),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_134),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_93),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_155),
.Y(n_248)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_0),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_30),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_103),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_69),
.Y(n_252)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_41),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_37),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_71),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_143),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_166),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_64),
.Y(n_258)
);

INVxp33_ASAP7_75t_L g259 ( 
.A(n_168),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_46),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_81),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_59),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_169),
.Y(n_263)
);

INVxp33_ASAP7_75t_SL g264 ( 
.A(n_66),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_3),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVxp33_ASAP7_75t_SL g268 ( 
.A(n_171),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_10),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_7),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_147),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_60),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_89),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_101),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_72),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_140),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_18),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_15),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_24),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_92),
.Y(n_280)
);

INVxp67_ASAP7_75t_SL g281 ( 
.A(n_139),
.Y(n_281)
);

CKINVDCx16_ASAP7_75t_R g282 ( 
.A(n_133),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_117),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_9),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_148),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_27),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_80),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_184),
.Y(n_289)
);

INVxp33_ASAP7_75t_L g290 ( 
.A(n_153),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_40),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_109),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_98),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_108),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_21),
.Y(n_295)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_13),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g298 ( 
.A(n_94),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_182),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g300 ( 
.A(n_107),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_152),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_88),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_125),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_179),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_79),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_67),
.Y(n_306)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_34),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_85),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_44),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_160),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_49),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_73),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_174),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_32),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_119),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g316 ( 
.A(n_159),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_158),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_123),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_102),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_23),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_167),
.Y(n_321)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_100),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_145),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_65),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_90),
.Y(n_325)
);

INVxp33_ASAP7_75t_L g326 ( 
.A(n_36),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_127),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_111),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_97),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_14),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_22),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_25),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_70),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_185),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_124),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_55),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_266),
.Y(n_337)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_221),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_227),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_188),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_191),
.Y(n_341)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_249),
.B(n_0),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_189),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_227),
.Y(n_345)
);

BUFx10_ASAP7_75t_L g346 ( 
.A(n_298),
.Y(n_346)
);

BUFx3_ASAP7_75t_L g347 ( 
.A(n_248),
.Y(n_347)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_227),
.Y(n_349)
);

AO21x2_ASAP7_75t_L g350 ( 
.A1(n_190),
.A2(n_205),
.B(n_203),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_333),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_327),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_206),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_209),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_192),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_211),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_197),
.B(n_1),
.Y(n_357)
);

INVx2_ASAP7_75t_SL g358 ( 
.A(n_194),
.Y(n_358)
);

INVx3_ASAP7_75t_L g359 ( 
.A(n_215),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_216),
.Y(n_360)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_282),
.Y(n_361)
);

AND2x4_ASAP7_75t_L g362 ( 
.A(n_199),
.B(n_1),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_217),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_306),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_218),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_220),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g367 ( 
.A1(n_259),
.A2(n_2),
.B1(n_3),
.B2(n_12),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_290),
.B(n_17),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_222),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_223),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_232),
.Y(n_371)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_236),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_198),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_225),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_226),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_230),
.Y(n_376)
);

INVx8_ASAP7_75t_L g377 ( 
.A(n_201),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_231),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_316),
.A2(n_26),
.B1(n_28),
.B2(n_33),
.Y(n_379)
);

INVx2_ASAP7_75t_SL g380 ( 
.A(n_204),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_238),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_253),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_239),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_241),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_208),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_254),
.Y(n_386)
);

BUFx4f_ASAP7_75t_L g387 ( 
.A(n_255),
.Y(n_387)
);

NAND2xp33_ASAP7_75t_L g388 ( 
.A(n_326),
.B(n_38),
.Y(n_388)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_256),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_219),
.Y(n_390)
);

BUFx10_ASAP7_75t_L g391 ( 
.A(n_258),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_261),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_265),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_267),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_260),
.B(n_52),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_269),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_270),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_273),
.Y(n_398)
);

BUFx3_ASAP7_75t_L g399 ( 
.A(n_224),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_274),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_195),
.B(n_196),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_212),
.B(n_54),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_275),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g404 ( 
.A(n_264),
.B(n_56),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_268),
.B(n_57),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_276),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_338),
.Y(n_407)
);

NAND4xp25_ASAP7_75t_SL g408 ( 
.A(n_351),
.B(n_367),
.C(n_342),
.D(n_337),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g409 ( 
.A(n_339),
.Y(n_409)
);

INVxp67_ASAP7_75t_SL g410 ( 
.A(n_347),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_339),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g412 ( 
.A(n_358),
.B(n_296),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_341),
.B(n_329),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_385),
.B(n_277),
.Y(n_414)
);

NAND2x1p5_ASAP7_75t_L g415 ( 
.A(n_395),
.B(n_237),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_345),
.Y(n_416)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_348),
.A2(n_322),
.B1(n_335),
.B2(n_235),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_348),
.Y(n_418)
);

INVx2_ASAP7_75t_SL g419 ( 
.A(n_346),
.Y(n_419)
);

BUFx2_ASAP7_75t_L g420 ( 
.A(n_355),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_345),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_401),
.B(n_212),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_399),
.Y(n_423)
);

BUFx6f_ASAP7_75t_L g424 ( 
.A(n_371),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_353),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g426 ( 
.A(n_352),
.B(n_279),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_380),
.Y(n_427)
);

O2A1O1Ixp33_ASAP7_75t_L g428 ( 
.A1(n_357),
.A2(n_233),
.B(n_257),
.C(n_250),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_354),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_390),
.B(n_402),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_350),
.B(n_280),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_361),
.B(n_233),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_344),
.B(n_285),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_360),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_371),
.Y(n_435)
);

AND2x6_ASAP7_75t_SL g436 ( 
.A(n_368),
.B(n_286),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_349),
.B(n_287),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_372),
.B(n_289),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

NAND2xp33_ASAP7_75t_SL g440 ( 
.A(n_364),
.B(n_193),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_372),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g442 ( 
.A(n_366),
.B(n_369),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_382),
.B(n_293),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_374),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_382),
.B(n_297),
.Y(n_445)
);

AND2x4_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_307),
.Y(n_446)
);

OAI21xp5_ASAP7_75t_L g447 ( 
.A1(n_387),
.A2(n_404),
.B(n_405),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_375),
.Y(n_449)
);

INVx5_ASAP7_75t_L g450 ( 
.A(n_391),
.Y(n_450)
);

BUFx3_ASAP7_75t_L g451 ( 
.A(n_356),
.Y(n_451)
);

NAND2x1_ASAP7_75t_L g452 ( 
.A(n_379),
.B(n_302),
.Y(n_452)
);

BUFx3_ASAP7_75t_L g453 ( 
.A(n_365),
.Y(n_453)
);

INVx2_ASAP7_75t_SL g454 ( 
.A(n_377),
.Y(n_454)
);

AOI21xp5_ASAP7_75t_L g455 ( 
.A1(n_431),
.A2(n_388),
.B(n_394),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_441),
.B(n_392),
.Y(n_456)
);

INVx2_ASAP7_75t_SL g457 ( 
.A(n_407),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_430),
.B(n_422),
.Y(n_458)
);

O2A1O1Ixp5_ASAP7_75t_L g459 ( 
.A1(n_452),
.A2(n_447),
.B(n_414),
.C(n_413),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_427),
.B(n_415),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_435),
.Y(n_461)
);

AND2x2_ASAP7_75t_L g462 ( 
.A(n_448),
.B(n_398),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g463 ( 
.A1(n_433),
.A2(n_443),
.B(n_438),
.Y(n_463)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_408),
.A2(n_384),
.B(n_370),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_442),
.Y(n_465)
);

O2A1O1Ixp33_ASAP7_75t_SL g466 ( 
.A1(n_428),
.A2(n_311),
.B(n_304),
.C(n_308),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g467 ( 
.A1(n_445),
.A2(n_376),
.B(n_381),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_412),
.A2(n_262),
.B1(n_284),
.B2(n_278),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g469 ( 
.A1(n_437),
.A2(n_378),
.B(n_389),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_453),
.Y(n_471)
);

OAI21x1_ASAP7_75t_L g472 ( 
.A1(n_432),
.A2(n_403),
.B(n_400),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_410),
.B(n_377),
.Y(n_473)
);

AO31x2_ASAP7_75t_L g474 ( 
.A1(n_425),
.A2(n_403),
.A3(n_400),
.B(n_397),
.Y(n_474)
);

OAI21x1_ASAP7_75t_L g475 ( 
.A1(n_426),
.A2(n_340),
.B(n_343),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_423),
.Y(n_476)
);

OAI21x1_ASAP7_75t_L g477 ( 
.A1(n_429),
.A2(n_397),
.B(n_396),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_446),
.B(n_383),
.Y(n_478)
);

AO31x2_ASAP7_75t_L g479 ( 
.A1(n_434),
.A2(n_396),
.A3(n_340),
.B(n_343),
.Y(n_479)
);

OAI21x1_ASAP7_75t_L g480 ( 
.A1(n_439),
.A2(n_319),
.B(n_309),
.Y(n_480)
);

INVx4_ASAP7_75t_L g481 ( 
.A(n_420),
.Y(n_481)
);

OAI21x1_ASAP7_75t_L g482 ( 
.A1(n_444),
.A2(n_313),
.B(n_321),
.Y(n_482)
);

BUFx3_ASAP7_75t_L g483 ( 
.A(n_424),
.Y(n_483)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_449),
.A2(n_393),
.B(n_386),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g485 ( 
.A(n_436),
.B(n_362),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_424),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_418),
.B(n_362),
.Y(n_487)
);

NOR4xp25_ASAP7_75t_L g488 ( 
.A(n_411),
.B(n_336),
.C(n_330),
.D(n_328),
.Y(n_488)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_416),
.A2(n_334),
.B(n_210),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_458),
.B(n_454),
.Y(n_490)
);

AOI21x1_ASAP7_75t_SL g491 ( 
.A1(n_485),
.A2(n_281),
.B(n_228),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_487),
.B(n_462),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_463),
.B(n_207),
.Y(n_493)
);

AOI221x1_ASAP7_75t_SL g494 ( 
.A1(n_468),
.A2(n_310),
.B1(n_323),
.B2(n_417),
.C(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_456),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_457),
.B(n_450),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_483),
.Y(n_497)
);

A2O1A1Ixp33_ASAP7_75t_L g498 ( 
.A1(n_459),
.A2(n_464),
.B(n_460),
.C(n_455),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_476),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_465),
.Y(n_500)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_450),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_477),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g503 ( 
.A1(n_470),
.A2(n_214),
.B1(n_200),
.B2(n_324),
.Y(n_503)
);

AOI21x1_ASAP7_75t_SL g504 ( 
.A1(n_478),
.A2(n_213),
.B(n_300),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g505 ( 
.A(n_471),
.B(n_419),
.Y(n_505)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_473),
.A2(n_202),
.B1(n_229),
.B2(n_245),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_472),
.B(n_450),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_488),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_409),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_461),
.B(n_409),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g511 ( 
.A1(n_475),
.A2(n_240),
.B(n_332),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_474),
.B(n_421),
.Y(n_512)
);

AOI221x1_ASAP7_75t_SL g513 ( 
.A1(n_466),
.A2(n_294),
.B1(n_251),
.B2(n_263),
.C(n_318),
.Y(n_513)
);

O2A1O1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_292),
.B(n_301),
.C(n_305),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_474),
.Y(n_515)
);

OR2x2_ASAP7_75t_L g516 ( 
.A(n_474),
.B(n_421),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_467),
.Y(n_517)
);

OA21x2_ASAP7_75t_L g518 ( 
.A1(n_469),
.A2(n_331),
.B(n_325),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g519 ( 
.A(n_492),
.B(n_479),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_500),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_516),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_512),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g523 ( 
.A(n_506),
.B(n_479),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_510),
.Y(n_524)
);

AND2x2_ASAP7_75t_L g525 ( 
.A(n_495),
.B(n_479),
.Y(n_525)
);

AO21x2_ASAP7_75t_L g526 ( 
.A1(n_498),
.A2(n_511),
.B(n_515),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_497),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_497),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g529 ( 
.A(n_496),
.B(n_484),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_509),
.Y(n_530)
);

INVx3_ASAP7_75t_L g531 ( 
.A(n_502),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_493),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_497),
.Y(n_533)
);

HB1xp67_ASAP7_75t_L g534 ( 
.A(n_499),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g535 ( 
.A(n_490),
.B(n_291),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_505),
.Y(n_536)
);

AND2x2_ASAP7_75t_L g537 ( 
.A(n_501),
.B(n_517),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_482),
.Y(n_538)
);

OAI31xp33_ASAP7_75t_L g539 ( 
.A1(n_514),
.A2(n_288),
.A3(n_320),
.B(n_317),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_494),
.B(n_480),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_503),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_522),
.B(n_513),
.Y(n_543)
);

OAI21x1_ASAP7_75t_L g544 ( 
.A1(n_538),
.A2(n_504),
.B(n_491),
.Y(n_544)
);

AND2x2_ASAP7_75t_L g545 ( 
.A(n_520),
.B(n_508),
.Y(n_545)
);

NOR2x1p5_ASAP7_75t_L g546 ( 
.A(n_536),
.B(n_283),
.Y(n_546)
);

HB1xp67_ASAP7_75t_L g547 ( 
.A(n_530),
.Y(n_547)
);

INVx2_ASAP7_75t_SL g548 ( 
.A(n_527),
.Y(n_548)
);

BUFx2_ASAP7_75t_L g549 ( 
.A(n_528),
.Y(n_549)
);

NAND3xp33_ASAP7_75t_SL g550 ( 
.A(n_539),
.B(n_272),
.C(n_315),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_519),
.Y(n_551)
);

AO21x1_ASAP7_75t_L g552 ( 
.A1(n_540),
.A2(n_518),
.B(n_63),
.Y(n_552)
);

OA21x2_ASAP7_75t_L g553 ( 
.A1(n_538),
.A2(n_518),
.B(n_314),
.Y(n_553)
);

BUFx2_ASAP7_75t_L g554 ( 
.A(n_533),
.Y(n_554)
);

OAI21xp5_ASAP7_75t_L g555 ( 
.A1(n_532),
.A2(n_312),
.B(n_303),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_556),
.B(n_541),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_545),
.B(n_524),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_551),
.B(n_537),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_551),
.B(n_535),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_547),
.B(n_525),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_543),
.B(n_529),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_549),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_555),
.B(n_539),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_554),
.Y(n_566)
);

OAI211xp5_ASAP7_75t_L g567 ( 
.A1(n_550),
.A2(n_523),
.B(n_242),
.C(n_252),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_548),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_557),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_559),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_561),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g572 ( 
.A(n_563),
.B(n_562),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_558),
.B(n_556),
.Y(n_573)
);

AND2x2_ASAP7_75t_L g574 ( 
.A(n_560),
.B(n_566),
.Y(n_574)
);

NAND3xp33_ASAP7_75t_L g575 ( 
.A(n_565),
.B(n_540),
.C(n_244),
.Y(n_575)
);

NOR3xp33_ASAP7_75t_L g576 ( 
.A(n_575),
.B(n_567),
.C(n_564),
.Y(n_576)
);

OAI322xp33_ASAP7_75t_L g577 ( 
.A1(n_572),
.A2(n_568),
.A3(n_299),
.B1(n_295),
.B2(n_271),
.C1(n_246),
.C2(n_243),
.Y(n_577)
);

AOI221xp5_ASAP7_75t_L g578 ( 
.A1(n_570),
.A2(n_567),
.B1(n_552),
.B2(n_526),
.C(n_531),
.Y(n_578)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_571),
.B(n_58),
.Y(n_579)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_573),
.A2(n_544),
.B(n_553),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_574),
.B(n_546),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_580),
.Y(n_582)
);

AND2x2_ASAP7_75t_L g583 ( 
.A(n_581),
.B(n_569),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_579),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_576),
.B(n_546),
.Y(n_585)
);

INVxp33_ASAP7_75t_L g586 ( 
.A(n_578),
.Y(n_586)
);

NAND4xp75_ASAP7_75t_L g587 ( 
.A(n_585),
.B(n_577),
.C(n_78),
.D(n_82),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_R g588 ( 
.A(n_583),
.B(n_77),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_584),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_582),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_590),
.Y(n_591)
);

NOR3xp33_ASAP7_75t_L g592 ( 
.A(n_587),
.B(n_586),
.C(n_86),
.Y(n_592)
);

NOR3xp33_ASAP7_75t_L g593 ( 
.A(n_589),
.B(n_586),
.C(n_104),
.Y(n_593)
);

AOI221xp5_ASAP7_75t_L g594 ( 
.A1(n_588),
.A2(n_114),
.B1(n_115),
.B2(n_116),
.C(n_118),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_591),
.B(n_129),
.Y(n_595)
);

AOI32xp33_ASAP7_75t_L g596 ( 
.A1(n_592),
.A2(n_130),
.A3(n_131),
.B1(n_132),
.B2(n_137),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_594),
.A2(n_141),
.B1(n_144),
.B2(n_150),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g598 ( 
.A(n_593),
.B(n_186),
.Y(n_598)
);

AOI221x1_ASAP7_75t_L g599 ( 
.A1(n_595),
.A2(n_156),
.B1(n_163),
.B2(n_164),
.C(n_165),
.Y(n_599)
);

CKINVDCx20_ASAP7_75t_R g600 ( 
.A(n_598),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_L g601 ( 
.A1(n_596),
.A2(n_597),
.B1(n_177),
.B2(n_178),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_601),
.B(n_180),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g603 ( 
.A1(n_602),
.A2(n_600),
.B1(n_599),
.B2(n_183),
.Y(n_603)
);


endmodule