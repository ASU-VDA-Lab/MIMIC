module fake_aes_2109_n_701 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_701);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_701;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_649;
wire n_276;
wire n_526;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_22), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_77), .Y(n_80) );
INVxp67_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
NOR2xp33_ASAP7_75t_L g82 ( .A(n_27), .B(n_76), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_43), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_71), .Y(n_84) );
CKINVDCx20_ASAP7_75t_R g85 ( .A(n_26), .Y(n_85) );
INVxp67_ASAP7_75t_SL g86 ( .A(n_74), .Y(n_86) );
INVx2_ASAP7_75t_SL g87 ( .A(n_45), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_72), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_62), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_61), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_29), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_46), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_66), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_32), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_39), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_56), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_14), .Y(n_98) );
INVx4_ASAP7_75t_R g99 ( .A(n_58), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_78), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_69), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_2), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_53), .Y(n_103) );
INVx2_ASAP7_75t_L g104 ( .A(n_44), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_20), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_65), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g107 ( .A(n_25), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_35), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_18), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g110 ( .A(n_13), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_40), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_70), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_19), .Y(n_113) );
INVxp33_ASAP7_75t_SL g114 ( .A(n_2), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_59), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_4), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g117 ( .A(n_24), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_33), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_7), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_8), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_4), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_28), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_11), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_48), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g125 ( .A(n_36), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_30), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_121), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_121), .B(n_0), .Y(n_128) );
INVx3_ASAP7_75t_L g129 ( .A(n_120), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_79), .Y(n_130) );
INVx6_ASAP7_75t_L g131 ( .A(n_120), .Y(n_131) );
OA21x2_ASAP7_75t_L g132 ( .A1(n_104), .A2(n_34), .B(n_73), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_87), .B(n_0), .Y(n_133) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_104), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_97), .B(n_1), .Y(n_135) );
CKINVDCx16_ASAP7_75t_R g136 ( .A(n_85), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_123), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
BUFx6f_ASAP7_75t_L g139 ( .A(n_120), .Y(n_139) );
BUFx2_ASAP7_75t_L g140 ( .A(n_115), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_116), .Y(n_141) );
OAI22xp5_ASAP7_75t_SL g142 ( .A1(n_102), .A2(n_1), .B1(n_3), .B2(n_5), .Y(n_142) );
INVx3_ASAP7_75t_L g143 ( .A(n_120), .Y(n_143) );
BUFx8_ASAP7_75t_L g144 ( .A(n_80), .Y(n_144) );
AND2x2_ASAP7_75t_L g145 ( .A(n_119), .B(n_3), .Y(n_145) );
NAND2xp33_ASAP7_75t_L g146 ( .A(n_115), .B(n_38), .Y(n_146) );
CKINVDCx20_ASAP7_75t_R g147 ( .A(n_102), .Y(n_147) );
AND2x4_ASAP7_75t_L g148 ( .A(n_83), .B(n_5), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_84), .Y(n_149) );
OAI22xp5_ASAP7_75t_L g150 ( .A1(n_98), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_90), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_91), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_126), .B(n_6), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_92), .Y(n_155) );
OA21x2_ASAP7_75t_L g156 ( .A1(n_93), .A2(n_42), .B(n_68), .Y(n_156) );
INVx3_ASAP7_75t_L g157 ( .A(n_94), .Y(n_157) );
NAND2xp5_ASAP7_75t_SL g158 ( .A(n_96), .B(n_9), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_100), .Y(n_159) );
AO22x1_ASAP7_75t_L g160 ( .A1(n_98), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_160) );
BUFx3_ASAP7_75t_L g161 ( .A(n_103), .Y(n_161) );
INVx4_ASAP7_75t_L g162 ( .A(n_125), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_108), .Y(n_163) );
OAI22xp5_ASAP7_75t_L g164 ( .A1(n_114), .A2(n_10), .B1(n_12), .B2(n_14), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_112), .B(n_12), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_113), .Y(n_166) );
AND2x6_ASAP7_75t_L g167 ( .A(n_118), .B(n_50), .Y(n_167) );
OAI22xp5_ASAP7_75t_L g168 ( .A1(n_114), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_82), .Y(n_169) );
INVx4_ASAP7_75t_L g170 ( .A(n_88), .Y(n_170) );
INVx1_ASAP7_75t_L g171 ( .A(n_128), .Y(n_171) );
NAND2xp5_ASAP7_75t_SL g172 ( .A(n_140), .B(n_81), .Y(n_172) );
AND2x2_ASAP7_75t_L g173 ( .A(n_140), .B(n_110), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_162), .B(n_101), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_134), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_167), .Y(n_176) );
OR2x6_ASAP7_75t_L g177 ( .A(n_160), .B(n_110), .Y(n_177) );
INVx2_ASAP7_75t_L g178 ( .A(n_134), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_162), .B(n_101), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_162), .B(n_86), .Y(n_180) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_162), .B(n_124), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_170), .B(n_122), .Y(n_182) );
INVx6_ASAP7_75t_L g183 ( .A(n_170), .Y(n_183) );
AOI22xp33_ASAP7_75t_L g184 ( .A1(n_128), .A2(n_148), .B1(n_167), .B2(n_145), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_128), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_170), .B(n_117), .Y(n_186) );
NOR2xp33_ASAP7_75t_L g187 ( .A(n_170), .B(n_106), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_130), .B(n_105), .Y(n_188) );
NAND2xp33_ASAP7_75t_SL g189 ( .A(n_137), .B(n_111), .Y(n_189) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_136), .Y(n_190) );
BUFx8_ASAP7_75t_SL g191 ( .A(n_147), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_144), .B(n_95), .Y(n_192) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_130), .B(n_111), .Y(n_193) );
AOI22xp33_ASAP7_75t_L g194 ( .A1(n_128), .A2(n_109), .B1(n_107), .B2(n_85), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_149), .B(n_109), .Y(n_195) );
INVx4_ASAP7_75t_SL g196 ( .A(n_167), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_134), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_134), .Y(n_198) );
INVx1_ASAP7_75t_L g199 ( .A(n_138), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_167), .Y(n_200) );
AND2x2_ASAP7_75t_L g201 ( .A(n_137), .B(n_107), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
NOR3xp33_ASAP7_75t_L g203 ( .A(n_142), .B(n_99), .C(n_16), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_149), .B(n_15), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_138), .Y(n_205) );
BUFx4f_ASAP7_75t_L g206 ( .A(n_167), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_153), .B(n_17), .Y(n_207) );
INVx4_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_153), .B(n_21), .Y(n_209) );
NOR2xp33_ASAP7_75t_SL g210 ( .A(n_144), .B(n_23), .Y(n_210) );
OR2x6_ASAP7_75t_L g211 ( .A(n_160), .B(n_31), .Y(n_211) );
BUFx10_ASAP7_75t_L g212 ( .A(n_148), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_155), .B(n_37), .Y(n_213) );
BUFx10_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_134), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_144), .Y(n_216) );
AOI22xp33_ASAP7_75t_L g217 ( .A1(n_148), .A2(n_41), .B1(n_47), .B2(n_49), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_155), .B(n_51), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_167), .Y(n_219) );
NAND2xp33_ASAP7_75t_SL g220 ( .A(n_154), .B(n_54), .Y(n_220) );
NAND2xp33_ASAP7_75t_R g221 ( .A(n_156), .B(n_75), .Y(n_221) );
BUFx3_ASAP7_75t_L g222 ( .A(n_167), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_135), .A2(n_145), .B1(n_166), .B2(n_152), .Y(n_223) );
BUFx10_ASAP7_75t_L g224 ( .A(n_133), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_154), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_163), .B(n_55), .Y(n_226) );
INVx4_ASAP7_75t_SL g227 ( .A(n_169), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_134), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_139), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_163), .B(n_57), .Y(n_230) );
BUFx2_ASAP7_75t_L g231 ( .A(n_144), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_154), .Y(n_232) );
NAND3xp33_ASAP7_75t_L g233 ( .A(n_141), .B(n_60), .C(n_63), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_139), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_224), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_227), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_184), .A2(n_159), .B(n_157), .C(n_152), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_227), .Y(n_238) );
CKINVDCx5p33_ASAP7_75t_R g239 ( .A(n_191), .Y(n_239) );
AO22x1_ASAP7_75t_L g240 ( .A1(n_203), .A2(n_150), .B1(n_168), .B2(n_164), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_216), .B(n_141), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_231), .B(n_145), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_223), .B(n_165), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_173), .B(n_136), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_225), .A2(n_135), .B(n_165), .C(n_151), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_201), .B(n_135), .Y(n_246) );
AOI22xp33_ASAP7_75t_L g247 ( .A1(n_171), .A2(n_151), .B1(n_166), .B2(n_152), .Y(n_247) );
INVx6_ASAP7_75t_L g248 ( .A(n_212), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_212), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_199), .Y(n_250) );
INVx6_ASAP7_75t_L g251 ( .A(n_214), .Y(n_251) );
A2O1A1Ixp33_ASAP7_75t_L g252 ( .A1(n_184), .A2(n_157), .B(n_159), .C(n_151), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_223), .B(n_165), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_232), .A2(n_150), .B(n_168), .C(n_164), .Y(n_254) );
OAI22xp5_ASAP7_75t_SL g255 ( .A1(n_177), .A2(n_142), .B1(n_127), .B2(n_156), .Y(n_255) );
INVxp67_ASAP7_75t_L g256 ( .A(n_193), .Y(n_256) );
NAND2xp5_ASAP7_75t_SL g257 ( .A(n_200), .B(n_169), .Y(n_257) );
INVx1_ASAP7_75t_L g258 ( .A(n_202), .Y(n_258) );
AOI22xp5_ASAP7_75t_L g259 ( .A1(n_193), .A2(n_195), .B1(n_177), .B2(n_172), .Y(n_259) );
CKINVDCx11_ASAP7_75t_R g260 ( .A(n_177), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_205), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_174), .B(n_161), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_185), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_179), .B(n_161), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_188), .B(n_161), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_227), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_211), .Y(n_267) );
INVx3_ASAP7_75t_L g268 ( .A(n_214), .Y(n_268) );
INVx2_ASAP7_75t_SL g269 ( .A(n_224), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_180), .B(n_169), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_180), .B(n_159), .Y(n_271) );
BUFx3_ASAP7_75t_L g272 ( .A(n_211), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_181), .B(n_159), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_181), .B(n_157), .Y(n_274) );
INVxp33_ASAP7_75t_L g275 ( .A(n_195), .Y(n_275) );
NAND2x1p5_ASAP7_75t_L g276 ( .A(n_192), .B(n_158), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_211), .A2(n_166), .B1(n_157), .B2(n_169), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_182), .B(n_169), .Y(n_278) );
AOI22xp33_ASAP7_75t_L g279 ( .A1(n_220), .A2(n_169), .B1(n_127), .B2(n_146), .Y(n_279) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_182), .B(n_132), .Y(n_280) );
NOR2xp33_ASAP7_75t_L g281 ( .A(n_186), .B(n_156), .Y(n_281) );
INVx4_ASAP7_75t_L g282 ( .A(n_183), .Y(n_282) );
INVx2_ASAP7_75t_SL g283 ( .A(n_190), .Y(n_283) );
INVx2_ASAP7_75t_SL g284 ( .A(n_204), .Y(n_284) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_187), .B(n_156), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_187), .B(n_132), .Y(n_286) );
AND2x2_ASAP7_75t_L g287 ( .A(n_194), .B(n_156), .Y(n_287) );
NAND2x1_ASAP7_75t_L g288 ( .A(n_183), .B(n_217), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g289 ( .A1(n_189), .A2(n_132), .B1(n_129), .B2(n_143), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_183), .B(n_132), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_200), .B(n_132), .Y(n_291) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_208), .B(n_139), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_207), .Y(n_293) );
OR2x2_ASAP7_75t_L g294 ( .A(n_194), .B(n_129), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_210), .B(n_196), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_209), .B(n_129), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_206), .A2(n_129), .B(n_143), .Y(n_297) );
OAI22xp5_ASAP7_75t_SL g298 ( .A1(n_217), .A2(n_131), .B1(n_143), .B2(n_139), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_196), .B(n_143), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_209), .B(n_131), .Y(n_300) );
BUFx6f_ASAP7_75t_L g301 ( .A(n_176), .Y(n_301) );
AOI21xp5_ASAP7_75t_L g302 ( .A1(n_206), .A2(n_139), .B(n_131), .Y(n_302) );
OAI21xp5_ASAP7_75t_L g303 ( .A1(n_281), .A2(n_219), .B(n_208), .Y(n_303) );
AOI21xp5_ASAP7_75t_L g304 ( .A1(n_290), .A2(n_219), .B(n_222), .Y(n_304) );
OR2x6_ASAP7_75t_L g305 ( .A(n_241), .B(n_176), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_263), .Y(n_306) );
AOI21xp5_ASAP7_75t_L g307 ( .A1(n_280), .A2(n_222), .B(n_218), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_250), .Y(n_308) );
OR2x2_ASAP7_75t_L g309 ( .A(n_244), .B(n_226), .Y(n_309) );
BUFx4f_ASAP7_75t_L g310 ( .A(n_241), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g311 ( .A(n_275), .B(n_230), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_286), .A2(n_213), .B(n_198), .Y(n_312) );
NAND2xp5_ASAP7_75t_SL g313 ( .A(n_249), .B(n_196), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_293), .B(n_213), .Y(n_314) );
OAI22xp5_ASAP7_75t_SL g315 ( .A1(n_239), .A2(n_233), .B1(n_221), .B2(n_131), .Y(n_315) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_242), .B(n_131), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_245), .B(n_198), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_277), .A2(n_221), .B1(n_139), .B2(n_228), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_242), .B(n_197), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_258), .Y(n_320) );
OAI221xp5_ASAP7_75t_L g321 ( .A1(n_256), .A2(n_259), .B1(n_254), .B2(n_253), .C(n_243), .Y(n_321) );
NOR3xp33_ASAP7_75t_SL g322 ( .A(n_255), .B(n_64), .C(n_67), .Y(n_322) );
NAND2xp33_ASAP7_75t_R g323 ( .A(n_287), .B(n_175), .Y(n_323) );
NAND2xp5_ASAP7_75t_SL g324 ( .A(n_249), .B(n_175), .Y(n_324) );
INVx6_ASAP7_75t_L g325 ( .A(n_248), .Y(n_325) );
OAI22x1_ASAP7_75t_L g326 ( .A1(n_267), .A2(n_256), .B1(n_260), .B2(n_283), .Y(n_326) );
BUFx3_ASAP7_75t_L g327 ( .A(n_235), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_261), .Y(n_328) );
BUFx3_ASAP7_75t_L g329 ( .A(n_269), .Y(n_329) );
INVx3_ASAP7_75t_SL g330 ( .A(n_248), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_268), .B(n_178), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_237), .A2(n_178), .B(n_197), .C(n_215), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_245), .B(n_215), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_301), .Y(n_334) );
NOR2xp33_ASAP7_75t_SL g335 ( .A(n_272), .B(n_228), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_252), .B(n_229), .Y(n_336) );
BUFx3_ASAP7_75t_L g337 ( .A(n_246), .Y(n_337) );
AOI21xp5_ASAP7_75t_L g338 ( .A1(n_291), .A2(n_229), .B(n_234), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_SL g339 ( .A1(n_288), .A2(n_234), .B(n_257), .C(n_278), .Y(n_339) );
OAI22xp5_ASAP7_75t_L g340 ( .A1(n_277), .A2(n_247), .B1(n_267), .B2(n_279), .Y(n_340) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_270), .A2(n_264), .B(n_262), .Y(n_341) );
AND2x2_ASAP7_75t_L g342 ( .A(n_240), .B(n_284), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_268), .B(n_301), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_291), .A2(n_281), .B(n_285), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_247), .B(n_271), .Y(n_345) );
AOI21xp5_ASAP7_75t_L g346 ( .A1(n_285), .A2(n_257), .B(n_292), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_294), .Y(n_347) );
O2A1O1Ixp33_ASAP7_75t_L g348 ( .A1(n_270), .A2(n_265), .B(n_274), .C(n_273), .Y(n_348) );
NOR2xp33_ASAP7_75t_L g349 ( .A(n_248), .B(n_251), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_L g350 ( .A1(n_276), .A2(n_296), .B(n_279), .C(n_292), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_251), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_276), .B(n_289), .Y(n_352) );
O2A1O1Ixp5_ASAP7_75t_L g353 ( .A1(n_302), .A2(n_297), .B(n_282), .C(n_300), .Y(n_353) );
AOI21xp5_ASAP7_75t_L g354 ( .A1(n_236), .A2(n_238), .B(n_266), .Y(n_354) );
NOR3xp33_ASAP7_75t_SL g355 ( .A(n_298), .B(n_251), .C(n_295), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_342), .B(n_299), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_303), .A2(n_301), .B(n_282), .Y(n_357) );
OAI21xp5_ASAP7_75t_L g358 ( .A1(n_346), .A2(n_301), .B(n_348), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_334), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_306), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g361 ( .A1(n_310), .A2(n_337), .B1(n_347), .B2(n_321), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_309), .B(n_328), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g363 ( .A1(n_310), .A2(n_305), .B1(n_314), .B2(n_318), .Y(n_363) );
OAI21xp5_ASAP7_75t_L g364 ( .A1(n_344), .A2(n_312), .B(n_304), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g365 ( .A1(n_307), .A2(n_314), .B(n_339), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_308), .B(n_320), .Y(n_366) );
OAI221xp5_ASAP7_75t_L g367 ( .A1(n_311), .A2(n_352), .B1(n_327), .B2(n_329), .C(n_340), .Y(n_367) );
O2A1O1Ixp33_ASAP7_75t_SL g368 ( .A1(n_352), .A2(n_317), .B(n_333), .C(n_336), .Y(n_368) );
O2A1O1Ixp33_ASAP7_75t_L g369 ( .A1(n_340), .A2(n_316), .B(n_350), .C(n_319), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
OAI21x1_ASAP7_75t_L g371 ( .A1(n_338), .A2(n_336), .B(n_318), .Y(n_371) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_334), .Y(n_372) );
AO31x2_ASAP7_75t_L g373 ( .A1(n_317), .A2(n_354), .A3(n_344), .B(n_323), .Y(n_373) );
INVx2_ASAP7_75t_L g374 ( .A(n_353), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_305), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_345), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_335), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_324), .Y(n_378) );
AOI21xp5_ASAP7_75t_L g379 ( .A1(n_341), .A2(n_332), .B(n_331), .Y(n_379) );
OAI21x1_ASAP7_75t_L g380 ( .A1(n_343), .A2(n_313), .B(n_349), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_305), .B(n_330), .Y(n_381) );
NAND3xp33_ASAP7_75t_L g382 ( .A(n_322), .B(n_355), .C(n_351), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_326), .B(n_325), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_315), .Y(n_384) );
O2A1O1Ixp33_ASAP7_75t_SL g385 ( .A1(n_325), .A2(n_252), .B(n_237), .C(n_288), .Y(n_385) );
O2A1O1Ixp33_ASAP7_75t_SL g386 ( .A1(n_325), .A2(n_252), .B(n_237), .C(n_288), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_330), .Y(n_387) );
BUFx6f_ASAP7_75t_L g388 ( .A(n_334), .Y(n_388) );
INVx1_ASAP7_75t_SL g389 ( .A(n_387), .Y(n_389) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_363), .A2(n_367), .B1(n_376), .B2(n_362), .Y(n_390) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_365), .A2(n_368), .B(n_364), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_387), .Y(n_392) );
AOI21xp5_ASAP7_75t_L g393 ( .A1(n_364), .A2(n_374), .B(n_386), .Y(n_393) );
AOI21xp5_ASAP7_75t_L g394 ( .A1(n_374), .A2(n_385), .B(n_379), .Y(n_394) );
AOI21xp5_ASAP7_75t_L g395 ( .A1(n_358), .A2(n_369), .B(n_371), .Y(n_395) );
OAI211xp5_ASAP7_75t_SL g396 ( .A1(n_361), .A2(n_383), .B(n_384), .C(n_381), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_384), .A2(n_382), .B1(n_376), .B2(n_356), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_371), .A2(n_357), .B(n_380), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_360), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_360), .B(n_366), .Y(n_400) );
AO21x2_ASAP7_75t_L g401 ( .A1(n_382), .A2(n_380), .B(n_359), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_356), .B(n_373), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_356), .B(n_375), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_375), .A2(n_378), .B1(n_377), .B2(n_370), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_373), .B(n_375), .Y(n_405) );
AO21x2_ASAP7_75t_L g406 ( .A1(n_359), .A2(n_370), .B(n_378), .Y(n_406) );
AOI21xp5_ASAP7_75t_L g407 ( .A1(n_372), .A2(n_388), .B(n_375), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_372), .Y(n_408) );
NAND2x1_ASAP7_75t_L g409 ( .A(n_372), .B(n_388), .Y(n_409) );
INVx5_ASAP7_75t_L g410 ( .A(n_375), .Y(n_410) );
INVx3_ASAP7_75t_L g411 ( .A(n_372), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_372), .A2(n_363), .B1(n_367), .B2(n_347), .Y(n_412) );
AOI221xp5_ASAP7_75t_L g413 ( .A1(n_388), .A2(n_254), .B1(n_240), .B2(n_321), .C(n_203), .Y(n_413) );
HB1xp67_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_373), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_388), .A2(n_255), .B1(n_384), .B2(n_260), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g417 ( .A1(n_390), .A2(n_373), .B1(n_388), .B2(n_397), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_400), .B(n_399), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_399), .Y(n_419) );
INVx2_ASAP7_75t_SL g420 ( .A(n_410), .Y(n_420) );
AOI22xp33_ASAP7_75t_L g421 ( .A1(n_396), .A2(n_416), .B1(n_413), .B2(n_412), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g422 ( .A(n_389), .B(n_392), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_400), .B(n_403), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_413), .A2(n_390), .B1(n_412), .B2(n_402), .Y(n_424) );
BUFx3_ASAP7_75t_L g425 ( .A(n_410), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_415), .Y(n_426) );
AO21x2_ASAP7_75t_L g427 ( .A1(n_391), .A2(n_395), .B(n_394), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_411), .Y(n_428) );
OR2x6_ASAP7_75t_L g429 ( .A(n_402), .B(n_405), .Y(n_429) );
AOI21xp5_ASAP7_75t_SL g430 ( .A1(n_405), .A2(n_415), .B(n_414), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_403), .B(n_410), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_389), .B(n_410), .Y(n_433) );
OR2x2_ASAP7_75t_L g434 ( .A(n_401), .B(n_406), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_393), .B(n_410), .Y(n_435) );
AO21x2_ASAP7_75t_L g436 ( .A1(n_407), .A2(n_401), .B(n_408), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_408), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_406), .Y(n_438) );
BUFx3_ASAP7_75t_L g439 ( .A(n_410), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_401), .Y(n_440) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_408), .B(n_411), .Y(n_441) );
NOR2xp67_ASAP7_75t_SL g442 ( .A(n_411), .B(n_398), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AO21x2_ASAP7_75t_L g444 ( .A1(n_398), .A2(n_409), .B(n_411), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_398), .Y(n_445) );
OA21x2_ASAP7_75t_L g446 ( .A1(n_404), .A2(n_391), .B(n_395), .Y(n_446) );
AO21x1_ASAP7_75t_SL g447 ( .A1(n_409), .A2(n_402), .B(n_405), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_399), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_408), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_408), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_399), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_410), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_426), .Y(n_453) );
INVx4_ASAP7_75t_L g454 ( .A(n_425), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_429), .B(n_426), .Y(n_455) );
INVx2_ASAP7_75t_SL g456 ( .A(n_425), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AOI322xp5_ASAP7_75t_L g458 ( .A1(n_418), .A2(n_451), .A3(n_421), .B1(n_448), .B2(n_419), .C1(n_424), .C2(n_423), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_423), .B(n_429), .Y(n_459) );
AND2x2_ASAP7_75t_L g460 ( .A(n_429), .B(n_447), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_448), .B(n_418), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_432), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_429), .Y(n_463) );
BUFx3_ASAP7_75t_L g464 ( .A(n_425), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_429), .Y(n_465) );
NOR3xp33_ASAP7_75t_L g466 ( .A(n_422), .B(n_433), .C(n_452), .Y(n_466) );
OR2x2_ASAP7_75t_L g467 ( .A(n_429), .B(n_451), .Y(n_467) );
INVx2_ASAP7_75t_L g468 ( .A(n_443), .Y(n_468) );
BUFx2_ASAP7_75t_L g469 ( .A(n_444), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_447), .B(n_437), .Y(n_470) );
AND2x2_ASAP7_75t_L g471 ( .A(n_437), .B(n_450), .Y(n_471) );
INVx1_ASAP7_75t_SL g472 ( .A(n_439), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_432), .Y(n_473) );
AND2x2_ASAP7_75t_SL g474 ( .A(n_430), .B(n_435), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_445), .Y(n_475) );
AO21x2_ASAP7_75t_L g476 ( .A1(n_427), .A2(n_440), .B(n_445), .Y(n_476) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_437), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_444), .B(n_435), .Y(n_478) );
AND2x4_ASAP7_75t_L g479 ( .A(n_444), .B(n_450), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_438), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_449), .B(n_431), .Y(n_481) );
OR2x6_ASAP7_75t_L g482 ( .A(n_430), .B(n_417), .Y(n_482) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
BUFx3_ASAP7_75t_L g484 ( .A(n_439), .Y(n_484) );
INVxp67_ASAP7_75t_SL g485 ( .A(n_442), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_438), .B(n_440), .Y(n_486) );
INVxp67_ASAP7_75t_SL g487 ( .A(n_442), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_431), .B(n_441), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_420), .B(n_452), .Y(n_489) );
INVx2_ASAP7_75t_L g490 ( .A(n_436), .Y(n_490) );
BUFx6f_ASAP7_75t_L g491 ( .A(n_446), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_417), .B(n_441), .Y(n_492) );
CKINVDCx20_ASAP7_75t_R g493 ( .A(n_439), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_420), .B(n_452), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_420), .A2(n_428), .B1(n_446), .B2(n_427), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_428), .B(n_427), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_434), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_436), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_427), .B(n_446), .Y(n_499) );
INVxp67_ASAP7_75t_L g500 ( .A(n_494), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_459), .B(n_434), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_453), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_459), .B(n_436), .Y(n_504) );
HB1xp67_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
AND2x2_ASAP7_75t_L g506 ( .A(n_488), .B(n_436), .Y(n_506) );
OAI31xp33_ASAP7_75t_L g507 ( .A1(n_489), .A2(n_428), .A3(n_446), .B(n_472), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_462), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_460), .B(n_428), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_457), .Y(n_510) );
INVx2_ASAP7_75t_L g511 ( .A(n_468), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_488), .B(n_446), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_462), .Y(n_513) );
NAND2x1p5_ASAP7_75t_L g514 ( .A(n_454), .B(n_464), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_467), .B(n_497), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_466), .A2(n_455), .B1(n_463), .B2(n_465), .Y(n_516) );
INVx2_ASAP7_75t_L g517 ( .A(n_468), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_455), .B(n_481), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_455), .B(n_481), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_468), .Y(n_520) );
AND2x2_ASAP7_75t_L g521 ( .A(n_470), .B(n_460), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_470), .B(n_460), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_473), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
INVxp67_ASAP7_75t_SL g525 ( .A(n_477), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_480), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_461), .B(n_458), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_470), .B(n_467), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_461), .B(n_458), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_480), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_457), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_466), .B(n_497), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_496), .B(n_486), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_493), .B(n_454), .Y(n_534) );
HB1xp67_ASAP7_75t_L g535 ( .A(n_477), .Y(n_535) );
INVx1_ASAP7_75t_SL g536 ( .A(n_472), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_486), .B(n_471), .Y(n_537) );
NAND2x1_ASAP7_75t_L g538 ( .A(n_454), .B(n_482), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_463), .B(n_465), .Y(n_539) );
OR2x2_ASAP7_75t_L g540 ( .A(n_486), .B(n_475), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_471), .B(n_496), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_471), .B(n_456), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_475), .B(n_499), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_475), .B(n_492), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_499), .B(n_479), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_499), .B(n_479), .Y(n_546) );
NOR2x1_ASAP7_75t_SL g547 ( .A(n_454), .B(n_464), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_456), .B(n_464), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_476), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_456), .B(n_484), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_545), .B(n_479), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_545), .B(n_478), .Y(n_552) );
INVx2_ASAP7_75t_L g553 ( .A(n_511), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_511), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_546), .B(n_478), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_508), .Y(n_556) );
OR2x2_ASAP7_75t_L g557 ( .A(n_515), .B(n_544), .Y(n_557) );
INVxp67_ASAP7_75t_SL g558 ( .A(n_547), .Y(n_558) );
INVx1_ASAP7_75t_SL g559 ( .A(n_536), .Y(n_559) );
AND2x2_ASAP7_75t_L g560 ( .A(n_546), .B(n_478), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_541), .B(n_478), .Y(n_561) );
INVxp67_ASAP7_75t_L g562 ( .A(n_547), .Y(n_562) );
INVx2_ASAP7_75t_SL g563 ( .A(n_514), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_502), .Y(n_564) );
INVx1_ASAP7_75t_L g565 ( .A(n_502), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_508), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_527), .B(n_492), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_529), .B(n_532), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_541), .B(n_469), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_513), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_517), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_533), .B(n_469), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_503), .Y(n_573) );
INVx2_ASAP7_75t_SL g574 ( .A(n_514), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_503), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_513), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_520), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_537), .B(n_484), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_531), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_531), .Y(n_581) );
AND2x4_ASAP7_75t_L g582 ( .A(n_521), .B(n_482), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_510), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_533), .B(n_483), .Y(n_584) );
CKINVDCx16_ASAP7_75t_R g585 ( .A(n_534), .Y(n_585) );
OR2x2_ASAP7_75t_L g586 ( .A(n_515), .B(n_476), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g587 ( .A(n_537), .B(n_484), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_500), .B(n_476), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_533), .B(n_483), .Y(n_589) );
INVxp67_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_512), .A2(n_482), .B1(n_474), .B2(n_491), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_505), .B(n_543), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_544), .B(n_476), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_523), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_535), .Y(n_595) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_516), .A2(n_474), .B1(n_482), .B2(n_485), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_506), .B(n_482), .Y(n_597) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_525), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_523), .Y(n_599) );
INVx4_ASAP7_75t_L g600 ( .A(n_514), .Y(n_600) );
OR2x2_ASAP7_75t_L g601 ( .A(n_540), .B(n_490), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_540), .B(n_490), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_543), .B(n_490), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_557), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_557), .B(n_506), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_595), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_567), .B(n_512), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_561), .B(n_504), .Y(n_608) );
INVx2_ASAP7_75t_SL g609 ( .A(n_600), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_568), .B(n_501), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_556), .Y(n_611) );
NOR2xp67_ASAP7_75t_SL g612 ( .A(n_600), .B(n_550), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_569), .B(n_501), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_556), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
AOI21xp33_ASAP7_75t_L g616 ( .A1(n_588), .A2(n_549), .B(n_507), .Y(n_616) );
BUFx2_ASAP7_75t_L g617 ( .A(n_558), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_566), .Y(n_618) );
INVx1_ASAP7_75t_L g619 ( .A(n_566), .Y(n_619) );
AND2x2_ASAP7_75t_L g620 ( .A(n_561), .B(n_504), .Y(n_620) );
OAI22xp5_ASAP7_75t_L g621 ( .A1(n_562), .A2(n_538), .B1(n_522), .B2(n_521), .Y(n_621) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_600), .B(n_538), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_570), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_570), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_577), .Y(n_625) );
INVx1_ASAP7_75t_L g626 ( .A(n_577), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_569), .B(n_519), .Y(n_627) );
INVx2_ASAP7_75t_L g628 ( .A(n_553), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_554), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_598), .B(n_519), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_599), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_599), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_563), .A2(n_522), .B(n_509), .C(n_474), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_551), .B(n_528), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_583), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_590), .B(n_518), .Y(n_636) );
INVx2_ASAP7_75t_L g637 ( .A(n_554), .Y(n_637) );
INVxp67_ASAP7_75t_L g638 ( .A(n_559), .Y(n_638) );
NAND2xp5_ASAP7_75t_SL g639 ( .A(n_585), .B(n_509), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_592), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_605), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_617), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_605), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_617), .B(n_560), .Y(n_644) );
INVx1_ASAP7_75t_L g645 ( .A(n_635), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_606), .Y(n_646) );
AOI322xp5_ASAP7_75t_L g647 ( .A1(n_639), .A2(n_582), .A3(n_597), .B1(n_560), .B2(n_552), .C1(n_555), .C2(n_587), .Y(n_647) );
INVx2_ASAP7_75t_L g648 ( .A(n_615), .Y(n_648) );
NAND2xp5_ASAP7_75t_SL g649 ( .A(n_609), .B(n_563), .Y(n_649) );
AOI31xp33_ASAP7_75t_L g650 ( .A1(n_622), .A2(n_574), .A3(n_591), .B(n_596), .Y(n_650) );
INVxp67_ASAP7_75t_L g651 ( .A(n_638), .Y(n_651) );
AOI21xp33_ASAP7_75t_SL g652 ( .A1(n_622), .A2(n_574), .B(n_582), .Y(n_652) );
OAI21xp33_ASAP7_75t_SL g653 ( .A1(n_639), .A2(n_552), .B(n_555), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_604), .B(n_586), .Y(n_654) );
INVx1_ASAP7_75t_SL g655 ( .A(n_609), .Y(n_655) );
INVxp67_ASAP7_75t_L g656 ( .A(n_612), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_608), .B(n_551), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_615), .Y(n_658) );
AOI21xp33_ASAP7_75t_L g659 ( .A1(n_616), .A2(n_549), .B(n_593), .Y(n_659) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_633), .A2(n_593), .B1(n_586), .B2(n_579), .C(n_601), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_607), .B(n_584), .Y(n_661) );
OAI22xp5_ASAP7_75t_L g662 ( .A1(n_633), .A2(n_582), .B1(n_597), .B2(n_528), .Y(n_662) );
NOR3xp33_ASAP7_75t_L g663 ( .A(n_621), .B(n_573), .C(n_565), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_642), .A2(n_630), .B1(n_627), .B2(n_613), .Y(n_664) );
AOI211xp5_ASAP7_75t_L g665 ( .A1(n_653), .A2(n_612), .B(n_610), .C(n_640), .Y(n_665) );
OAI21xp5_ASAP7_75t_L g666 ( .A1(n_642), .A2(n_636), .B(n_634), .Y(n_666) );
AOI21xp5_ASAP7_75t_L g667 ( .A1(n_649), .A2(n_542), .B(n_603), .Y(n_667) );
A2O1A1Ixp33_ASAP7_75t_L g668 ( .A1(n_652), .A2(n_634), .B(n_608), .C(n_620), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g669 ( .A1(n_656), .A2(n_620), .B1(n_572), .B2(n_584), .Y(n_669) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_662), .A2(n_589), .B1(n_572), .B2(n_509), .Y(n_670) );
O2A1O1Ixp5_ASAP7_75t_L g671 ( .A1(n_649), .A2(n_625), .B(n_632), .C(n_631), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_641), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_651), .Y(n_673) );
AOI322xp5_ASAP7_75t_L g674 ( .A1(n_643), .A2(n_589), .A3(n_518), .B1(n_624), .B2(n_623), .C1(n_619), .C2(n_618), .Y(n_674) );
OAI221xp5_ASAP7_75t_L g675 ( .A1(n_650), .A2(n_626), .B1(n_614), .B2(n_611), .C(n_602), .Y(n_675) );
AOI22xp5_ASAP7_75t_L g676 ( .A1(n_663), .A2(n_482), .B1(n_594), .B2(n_581), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g677 ( .A1(n_644), .A2(n_575), .A3(n_564), .B1(n_580), .B2(n_637), .C1(n_628), .C2(n_629), .Y(n_677) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_665), .B(n_655), .Y(n_678) );
OAI211xp5_ASAP7_75t_L g679 ( .A1(n_675), .A2(n_647), .B(n_659), .C(n_660), .Y(n_679) );
NAND3xp33_ASAP7_75t_L g680 ( .A(n_673), .B(n_646), .C(n_645), .Y(n_680) );
A2O1A1Ixp33_ASAP7_75t_L g681 ( .A1(n_668), .A2(n_644), .B(n_657), .C(n_654), .Y(n_681) );
NOR3xp33_ASAP7_75t_SL g682 ( .A(n_669), .B(n_661), .C(n_658), .Y(n_682) );
A2O1A1Ixp33_ASAP7_75t_L g683 ( .A1(n_671), .A2(n_657), .B(n_648), .C(n_658), .Y(n_683) );
AOI221xp5_ASAP7_75t_L g684 ( .A1(n_664), .A2(n_648), .B1(n_637), .B2(n_628), .C(n_629), .Y(n_684) );
NAND2xp5_ASAP7_75t_SL g685 ( .A(n_677), .B(n_674), .Y(n_685) );
O2A1O1Ixp33_ASAP7_75t_L g686 ( .A1(n_685), .A2(n_666), .B(n_672), .C(n_670), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_684), .B(n_667), .Y(n_687) );
OAI211xp5_ASAP7_75t_SL g688 ( .A1(n_678), .A2(n_676), .B(n_495), .C(n_539), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_680), .Y(n_689) );
NAND3xp33_ASAP7_75t_L g690 ( .A(n_682), .B(n_524), .C(n_530), .Y(n_690) );
AOI211xp5_ASAP7_75t_L g691 ( .A1(n_686), .A2(n_679), .B(n_681), .C(n_683), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g692 ( .A(n_689), .B(n_485), .C(n_487), .Y(n_692) );
NOR3xp33_ASAP7_75t_L g693 ( .A(n_688), .B(n_487), .C(n_530), .Y(n_693) );
INVx4_ASAP7_75t_L g694 ( .A(n_691), .Y(n_694) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_692), .B(n_687), .Y(n_695) );
INVx2_ASAP7_75t_SL g696 ( .A(n_695), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_696), .A2(n_694), .B1(n_693), .B2(n_690), .Y(n_697) );
AOI222xp33_ASAP7_75t_SL g698 ( .A1(n_697), .A2(n_526), .B1(n_524), .B2(n_578), .C1(n_571), .C2(n_576), .Y(n_698) );
OR2x2_ASAP7_75t_L g699 ( .A(n_698), .B(n_602), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_699), .A2(n_526), .B(n_498), .Y(n_700) );
AOI21xp33_ASAP7_75t_L g701 ( .A1(n_700), .A2(n_601), .B(n_539), .Y(n_701) );
endmodule