module real_aes_17183_n_376 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_375, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_376);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_375;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_376;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_2003;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1994;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1959;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_1966;
wire n_1346;
wire n_552;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1583;
wire n_1250;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1632;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_1648;
wire n_724;
wire n_1914;
wire n_1945;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_877;
wire n_424;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1973;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_948;
wire n_399;
wire n_1499;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1946;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_1971;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_1404;
wire n_602;
wire n_402;
wire n_733;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_1569;
wire n_895;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1580;
wire n_1000;
wire n_1187;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1474;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1185;
wire n_661;
wire n_1102;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_1175;
wire n_778;
wire n_1170;
wire n_522;
wire n_1475;
wire n_1928;
wire n_977;
wire n_943;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1939;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1671;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1802;
wire n_1855;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_524;
wire n_1496;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_1143;
wire n_929;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1457;
wire n_1343;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1931;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_423;
wire n_1969;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1584;
wire n_1277;
wire n_1049;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1352;
wire n_729;
wire n_1323;
wire n_1280;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g627 ( .A(n_0), .Y(n_627) );
OAI211xp5_ASAP7_75t_L g1515 ( .A1(n_1), .A2(n_772), .B(n_1512), .C(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1528 ( .A(n_1), .Y(n_1528) );
INVx1_ASAP7_75t_L g1594 ( .A(n_2), .Y(n_1594) );
OAI211xp5_ASAP7_75t_L g1620 ( .A1(n_2), .A2(n_1621), .B(n_1622), .C(n_1626), .Y(n_1620) );
INVx1_ASAP7_75t_L g391 ( .A(n_3), .Y(n_391) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_3), .B(n_401), .Y(n_542) );
AND2x2_ASAP7_75t_L g626 ( .A(n_3), .B(n_278), .Y(n_626) );
AND2x2_ASAP7_75t_L g642 ( .A(n_3), .B(n_433), .Y(n_642) );
INVx1_ASAP7_75t_L g1045 ( .A(n_4), .Y(n_1045) );
INVx1_ASAP7_75t_L g1665 ( .A(n_5), .Y(n_1665) );
OAI22xp5_ASAP7_75t_L g628 ( .A1(n_6), .A2(n_287), .B1(n_629), .B2(n_635), .Y(n_628) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_6), .A2(n_640), .B(n_643), .C(n_650), .Y(n_639) );
INVx1_ASAP7_75t_L g1447 ( .A(n_7), .Y(n_1447) );
INVx1_ASAP7_75t_L g1099 ( .A(n_8), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g851 ( .A1(n_9), .A2(n_299), .B1(n_489), .B2(n_775), .Y(n_851) );
OAI22xp33_ASAP7_75t_L g858 ( .A1(n_9), .A2(n_299), .B1(n_859), .B2(n_860), .Y(n_858) );
AOI22xp5_ASAP7_75t_L g1689 ( .A1(n_10), .A2(n_78), .B1(n_1690), .B2(n_1692), .Y(n_1689) );
XOR2x2_ASAP7_75t_L g1896 ( .A(n_10), .B(n_1897), .Y(n_1896) );
AOI22xp33_ASAP7_75t_L g1953 ( .A1(n_10), .A2(n_1954), .B1(n_1957), .B2(n_1999), .Y(n_1953) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_11), .A2(n_83), .B1(n_519), .B2(n_520), .Y(n_524) );
AOI22xp33_ASAP7_75t_L g567 ( .A1(n_11), .A2(n_246), .B1(n_544), .B2(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g966 ( .A(n_12), .Y(n_966) );
OAI211xp5_ASAP7_75t_L g1663 ( .A1(n_13), .A2(n_828), .B(n_1507), .C(n_1664), .Y(n_1663) );
INVx1_ASAP7_75t_L g1672 ( .A(n_13), .Y(n_1672) );
AOI22xp33_ASAP7_75t_L g1445 ( .A1(n_14), .A2(n_89), .B1(n_467), .B2(n_598), .Y(n_1445) );
AOI221xp5_ASAP7_75t_L g1462 ( .A1(n_14), .A2(n_28), .B1(n_657), .B2(n_1463), .C(n_1465), .Y(n_1462) );
INVx1_ASAP7_75t_L g1964 ( .A(n_15), .Y(n_1964) );
OAI22xp5_ASAP7_75t_L g994 ( .A1(n_16), .A2(n_54), .B1(n_925), .B2(n_995), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_16), .A2(n_54), .B1(n_921), .B2(n_1005), .Y(n_1004) );
INVx1_ASAP7_75t_L g1535 ( .A(n_17), .Y(n_1535) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_18), .A2(n_319), .B1(n_519), .B2(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_18), .A2(n_369), .B1(n_657), .B2(n_658), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g1612 ( .A1(n_19), .A2(n_198), .B1(n_596), .B2(n_1613), .Y(n_1612) );
INVx1_ASAP7_75t_L g1623 ( .A(n_19), .Y(n_1623) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_20), .A2(n_32), .B1(n_532), .B2(n_1310), .Y(n_1339) );
INVx1_ASAP7_75t_L g1378 ( .A(n_20), .Y(n_1378) );
INVx1_ASAP7_75t_L g697 ( .A(n_21), .Y(n_697) );
INVx1_ASAP7_75t_L g1131 ( .A(n_22), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g1137 ( .A1(n_22), .A2(n_772), .B(n_1138), .C(n_1140), .Y(n_1137) );
INVx1_ASAP7_75t_L g798 ( .A(n_23), .Y(n_798) );
INVx1_ASAP7_75t_L g917 ( .A(n_24), .Y(n_917) );
OAI22xp33_ASAP7_75t_L g1181 ( .A1(n_25), .A2(n_179), .B1(n_762), .B2(n_763), .Y(n_1181) );
OAI22xp33_ASAP7_75t_L g1183 ( .A1(n_25), .A2(n_179), .B1(n_393), .B2(n_1077), .Y(n_1183) );
INVx1_ASAP7_75t_L g1102 ( .A(n_26), .Y(n_1102) );
CKINVDCx5p33_ASAP7_75t_R g1203 ( .A(n_27), .Y(n_1203) );
AOI22xp33_ASAP7_75t_SL g1454 ( .A1(n_28), .A2(n_263), .B1(n_517), .B2(n_532), .Y(n_1454) );
INVx2_ASAP7_75t_L g478 ( .A(n_29), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_30), .A2(n_374), .B1(n_681), .B2(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1579 ( .A(n_30), .Y(n_1579) );
OAI22xp33_ASAP7_75t_L g743 ( .A1(n_31), .A2(n_303), .B1(n_393), .B2(n_744), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g761 ( .A1(n_31), .A2(n_303), .B1(n_762), .B2(n_763), .Y(n_761) );
AOI221xp5_ASAP7_75t_L g1356 ( .A1(n_32), .A2(n_53), .B1(n_681), .B2(n_1357), .C(n_1359), .Y(n_1356) );
INVx1_ASAP7_75t_L g886 ( .A(n_33), .Y(n_886) );
INVx1_ASAP7_75t_L g1451 ( .A(n_34), .Y(n_1451) );
INVx1_ASAP7_75t_L g1974 ( .A(n_35), .Y(n_1974) );
OAI22xp5_ASAP7_75t_L g1065 ( .A1(n_36), .A2(n_308), .B1(n_930), .B2(n_1066), .Y(n_1065) );
OAI22xp5_ASAP7_75t_L g1078 ( .A1(n_36), .A2(n_345), .B1(n_1079), .B2(n_1081), .Y(n_1078) );
INVx1_ASAP7_75t_L g430 ( .A(n_37), .Y(n_430) );
AOI22xp5_ASAP7_75t_L g1714 ( .A1(n_38), .A2(n_247), .B1(n_1682), .B2(n_1687), .Y(n_1714) );
INVx1_ASAP7_75t_L g1110 ( .A(n_39), .Y(n_1110) );
OA222x2_ASAP7_75t_L g1248 ( .A1(n_40), .A2(n_95), .B1(n_271), .B2(n_1249), .C1(n_1251), .C2(n_1257), .Y(n_1248) );
INVx1_ASAP7_75t_L g1307 ( .A(n_40), .Y(n_1307) );
HB1xp67_ASAP7_75t_L g386 ( .A(n_41), .Y(n_386) );
AND2x2_ASAP7_75t_L g1683 ( .A(n_41), .B(n_384), .Y(n_1683) );
AOI22xp5_ASAP7_75t_L g1681 ( .A1(n_42), .A2(n_221), .B1(n_1682), .B2(n_1687), .Y(n_1681) );
AOI22xp33_ASAP7_75t_L g1402 ( .A1(n_43), .A2(n_353), .B1(n_418), .B2(n_569), .Y(n_1402) );
INVxp67_ASAP7_75t_SL g1419 ( .A(n_43), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1559 ( .A1(n_44), .A2(n_228), .B1(n_548), .B2(n_1560), .Y(n_1559) );
AOI22xp33_ASAP7_75t_L g1585 ( .A1(n_44), .A2(n_289), .B1(n_607), .B2(n_1586), .Y(n_1585) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_45), .A2(n_240), .B1(n_519), .B2(n_1308), .Y(n_1340) );
INVx1_ASAP7_75t_L g1361 ( .A(n_45), .Y(n_1361) );
AOI22xp5_ASAP7_75t_L g1698 ( .A1(n_46), .A2(n_296), .B1(n_1682), .B2(n_1687), .Y(n_1698) );
INVx1_ASAP7_75t_L g1541 ( .A(n_47), .Y(n_1541) );
INVx1_ASAP7_75t_L g967 ( .A(n_48), .Y(n_967) );
INVx1_ASAP7_75t_L g710 ( .A(n_49), .Y(n_710) );
OAI22xp5_ASAP7_75t_L g919 ( .A1(n_50), .A2(n_293), .B1(n_920), .B2(n_921), .Y(n_919) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_50), .A2(n_209), .B1(n_489), .B2(n_930), .Y(n_929) );
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_51), .Y(n_1207) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_52), .A2(n_208), .B1(n_842), .B2(n_844), .Y(n_841) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_52), .A2(n_208), .B1(n_393), .B2(n_744), .Y(n_861) );
AOI22xp33_ASAP7_75t_SL g1345 ( .A1(n_53), .A2(n_341), .B1(n_532), .B2(n_1346), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g1450 ( .A(n_55), .Y(n_1450) );
OAI22xp5_ASAP7_75t_L g1471 ( .A1(n_55), .A2(n_197), .B1(n_870), .B2(n_1472), .Y(n_1471) );
AOI22xp5_ASAP7_75t_L g1710 ( .A1(n_56), .A2(n_128), .B1(n_1682), .B2(n_1687), .Y(n_1710) );
AOI22xp33_ASAP7_75t_SL g933 ( .A1(n_57), .A2(n_136), .B1(n_934), .B2(n_935), .Y(n_933) );
AOI22xp33_ASAP7_75t_SL g954 ( .A1(n_57), .A2(n_277), .B1(n_948), .B2(n_955), .Y(n_954) );
INVx1_ASAP7_75t_L g1644 ( .A(n_58), .Y(n_1644) );
INVx1_ASAP7_75t_L g1970 ( .A(n_59), .Y(n_1970) );
INVx1_ASAP7_75t_L g1158 ( .A(n_60), .Y(n_1158) );
INVx1_ASAP7_75t_L g792 ( .A(n_61), .Y(n_792) );
OAI211xp5_ASAP7_75t_L g745 ( .A1(n_62), .A2(n_746), .B(n_748), .C(n_749), .Y(n_745) );
INVx1_ASAP7_75t_L g771 ( .A(n_62), .Y(n_771) );
CKINVDCx5p33_ASAP7_75t_R g1273 ( .A(n_63), .Y(n_1273) );
INVx1_ASAP7_75t_L g1458 ( .A(n_64), .Y(n_1458) );
INVx1_ASAP7_75t_L g1038 ( .A(n_65), .Y(n_1038) );
INVx1_ASAP7_75t_L g1606 ( .A(n_66), .Y(n_1606) );
AOI21xp33_ASAP7_75t_L g1627 ( .A1(n_66), .A2(n_678), .B(n_941), .Y(n_1627) );
AOI22xp5_ASAP7_75t_L g1708 ( .A1(n_67), .A2(n_202), .B1(n_1690), .B2(n_1709), .Y(n_1708) );
INVx1_ASAP7_75t_L g1178 ( .A(n_68), .Y(n_1178) );
AOI22xp33_ASAP7_75t_SL g1407 ( .A1(n_69), .A2(n_286), .B1(n_418), .B2(n_1408), .Y(n_1407) );
AOI22xp33_ASAP7_75t_L g1420 ( .A1(n_69), .A2(n_268), .B1(n_955), .B2(n_1299), .Y(n_1420) );
OAI22xp33_ASAP7_75t_L g1667 ( .A1(n_70), .A2(n_152), .B1(n_774), .B2(n_833), .Y(n_1667) );
OAI22xp5_ASAP7_75t_L g1673 ( .A1(n_70), .A2(n_152), .B1(n_755), .B2(n_860), .Y(n_1673) );
CKINVDCx5p33_ASAP7_75t_R g1449 ( .A(n_71), .Y(n_1449) );
INVx1_ASAP7_75t_L g1482 ( .A(n_72), .Y(n_1482) );
BUFx6f_ASAP7_75t_L g398 ( .A(n_73), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g1341 ( .A1(n_74), .A2(n_84), .B1(n_1342), .B2(n_1344), .Y(n_1341) );
INVx1_ASAP7_75t_L g1360 ( .A(n_74), .Y(n_1360) );
INVx1_ASAP7_75t_L g1152 ( .A(n_75), .Y(n_1152) );
OAI22xp33_ASAP7_75t_SL g1397 ( .A1(n_76), .A2(n_274), .B1(n_877), .B2(n_882), .Y(n_1397) );
INVx1_ASAP7_75t_L g1433 ( .A(n_76), .Y(n_1433) );
INVx1_ASAP7_75t_L g1602 ( .A(n_77), .Y(n_1602) );
OAI22xp5_ASAP7_75t_L g1617 ( .A1(n_77), .A2(n_334), .B1(n_1618), .B2(n_1619), .Y(n_1617) );
CKINVDCx5p33_ASAP7_75t_R g1332 ( .A(n_79), .Y(n_1332) );
INVx1_ASAP7_75t_L g701 ( .A(n_80), .Y(n_701) );
OAI22xp33_ASAP7_75t_L g1220 ( .A1(n_81), .A2(n_131), .B1(n_393), .B2(n_1077), .Y(n_1220) );
OAI22xp33_ASAP7_75t_L g1229 ( .A1(n_81), .A2(n_131), .B1(n_844), .B2(n_930), .Y(n_1229) );
AOI21xp33_ASAP7_75t_L g1569 ( .A1(n_82), .A2(n_552), .B(n_1401), .Y(n_1569) );
AOI22xp33_ASAP7_75t_L g1580 ( .A1(n_82), .A2(n_228), .B1(n_1310), .B2(n_1581), .Y(n_1580) );
AOI22xp33_ASAP7_75t_SL g550 ( .A1(n_83), .A2(n_113), .B1(n_551), .B2(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g1382 ( .A(n_84), .Y(n_1382) );
AOI22xp33_ASAP7_75t_L g1768 ( .A1(n_85), .A2(n_266), .B1(n_1690), .B2(n_1692), .Y(n_1768) );
INVx1_ASAP7_75t_L g1991 ( .A(n_86), .Y(n_1991) );
OAI211xp5_ASAP7_75t_L g1996 ( .A1(n_86), .A2(n_748), .B(n_1186), .C(n_1997), .Y(n_1996) );
INVx1_ASAP7_75t_L g821 ( .A(n_87), .Y(n_821) );
OAI211xp5_ASAP7_75t_L g827 ( .A1(n_87), .A2(n_765), .B(n_828), .C(n_829), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g581 ( .A1(n_88), .A2(n_330), .B1(n_582), .B2(n_589), .Y(n_581) );
INVx1_ASAP7_75t_L g644 ( .A(n_88), .Y(n_644) );
INVx1_ASAP7_75t_L g1481 ( .A(n_89), .Y(n_1481) );
INVx1_ASAP7_75t_L g1906 ( .A(n_90), .Y(n_1906) );
INVx1_ASAP7_75t_L g1041 ( .A(n_91), .Y(n_1041) );
INVx1_ASAP7_75t_L g789 ( .A(n_92), .Y(n_789) );
CKINVDCx5p33_ASAP7_75t_R g1552 ( .A(n_93), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g1930 ( .A1(n_94), .A2(n_276), .B1(n_926), .B2(n_1136), .Y(n_1930) );
OAI22xp5_ASAP7_75t_L g1941 ( .A1(n_94), .A2(n_276), .B1(n_1942), .B2(n_1943), .Y(n_1941) );
OAI221xp5_ASAP7_75t_L g1292 ( .A1(n_95), .A2(n_216), .B1(n_1293), .B2(n_1295), .C(n_1297), .Y(n_1292) );
OAI22xp5_ASAP7_75t_L g1369 ( .A1(n_96), .A2(n_325), .B1(n_425), .B2(n_870), .Y(n_1369) );
INVx1_ASAP7_75t_L g1384 ( .A(n_96), .Y(n_1384) );
INVx1_ASAP7_75t_L g1265 ( .A(n_97), .Y(n_1265) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_97), .A2(n_149), .B1(n_522), .B2(n_607), .Y(n_1324) );
INVx1_ASAP7_75t_L g888 ( .A(n_98), .Y(n_888) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_99), .A2(n_195), .B1(n_755), .B2(n_757), .Y(n_754) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_99), .A2(n_195), .B1(n_774), .B2(n_775), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1725 ( .A1(n_100), .A2(n_203), .B1(n_1682), .B2(n_1690), .Y(n_1725) );
INVx1_ASAP7_75t_L g429 ( .A(n_101), .Y(n_429) );
AOI22xp33_ASAP7_75t_SL g531 ( .A1(n_102), .A2(n_191), .B1(n_532), .B2(n_534), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_102), .A2(n_253), .B1(n_544), .B2(n_546), .Y(n_543) );
XOR2x2_ASAP7_75t_L g1017 ( .A(n_103), .B(n_1018), .Y(n_1017) );
AOI22xp33_ASAP7_75t_L g1724 ( .A1(n_103), .A2(n_324), .B1(n_1687), .B2(n_1692), .Y(n_1724) );
INVx1_ASAP7_75t_L g1968 ( .A(n_104), .Y(n_1968) );
XNOR2xp5_ASAP7_75t_L g778 ( .A(n_105), .B(n_779), .Y(n_778) );
AOI22xp5_ASAP7_75t_L g1700 ( .A1(n_105), .A2(n_175), .B1(n_1690), .B2(n_1701), .Y(n_1700) );
XNOR2xp5_ASAP7_75t_L g1639 ( .A(n_106), .B(n_1640), .Y(n_1639) );
CKINVDCx5p33_ASAP7_75t_R g1457 ( .A(n_107), .Y(n_1457) );
AOI22xp33_ASAP7_75t_SL g606 ( .A1(n_108), .A2(n_279), .B1(n_535), .B2(n_607), .Y(n_606) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_108), .A2(n_331), .B1(n_652), .B2(n_654), .C(n_655), .Y(n_651) );
AOI22xp33_ASAP7_75t_L g1453 ( .A1(n_109), .A2(n_346), .B1(n_520), .B2(n_1342), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1478 ( .A1(n_109), .A2(n_236), .B1(n_418), .B2(n_681), .C(n_1479), .Y(n_1478) );
INVx1_ASAP7_75t_L g1905 ( .A(n_110), .Y(n_1905) );
INVx1_ASAP7_75t_L g1648 ( .A(n_111), .Y(n_1648) );
INVx1_ASAP7_75t_L g1153 ( .A(n_112), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_113), .A2(n_246), .B1(n_519), .B2(n_520), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g1769 ( .A1(n_114), .A2(n_359), .B1(n_1682), .B2(n_1687), .Y(n_1769) );
OAI22xp33_ASAP7_75t_L g1514 ( .A1(n_115), .A2(n_171), .B1(n_501), .B2(n_844), .Y(n_1514) );
OAI22xp33_ASAP7_75t_L g1522 ( .A1(n_115), .A2(n_171), .B1(n_393), .B2(n_744), .Y(n_1522) );
INVx1_ASAP7_75t_L g1387 ( .A(n_116), .Y(n_1387) );
INVx1_ASAP7_75t_L g1917 ( .A(n_117), .Y(n_1917) );
INVx1_ASAP7_75t_L g751 ( .A(n_118), .Y(n_751) );
OAI22xp33_ASAP7_75t_L g1126 ( .A1(n_119), .A2(n_125), .B1(n_1007), .B2(n_1077), .Y(n_1126) );
OAI22xp33_ASAP7_75t_L g1134 ( .A1(n_119), .A2(n_125), .B1(n_826), .B2(n_842), .Y(n_1134) );
INVx1_ASAP7_75t_L g1495 ( .A(n_120), .Y(n_1495) );
INVx1_ASAP7_75t_L g1611 ( .A(n_121), .Y(n_1611) );
AOI22xp33_ASAP7_75t_L g1625 ( .A1(n_121), .A2(n_281), .B1(n_418), .B2(n_569), .Y(n_1625) );
CKINVDCx5p33_ASAP7_75t_R g1551 ( .A(n_122), .Y(n_1551) );
INVx1_ASAP7_75t_L g384 ( .A(n_123), .Y(n_384) );
INVx1_ASAP7_75t_L g1967 ( .A(n_124), .Y(n_1967) );
XOR2x2_ASAP7_75t_L g838 ( .A(n_126), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g1024 ( .A(n_127), .Y(n_1024) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_129), .A2(n_170), .B1(n_755), .B2(n_757), .Y(n_822) );
OAI22xp33_ASAP7_75t_L g832 ( .A1(n_129), .A2(n_170), .B1(n_774), .B2(n_833), .Y(n_832) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_130), .A2(n_163), .B1(n_968), .B2(n_1266), .Y(n_1396) );
NOR2xp33_ASAP7_75t_L g1437 ( .A(n_130), .B(n_1438), .Y(n_1437) );
CKINVDCx5p33_ASAP7_75t_R g1352 ( .A(n_132), .Y(n_1352) );
INVx1_ASAP7_75t_L g1503 ( .A(n_133), .Y(n_1503) );
INVx1_ASAP7_75t_L g704 ( .A(n_134), .Y(n_704) );
XOR2xp5_ASAP7_75t_L g1958 ( .A(n_135), .B(n_1959), .Y(n_1958) );
AOI22xp33_ASAP7_75t_L g944 ( .A1(n_136), .A2(n_258), .B1(n_534), .B2(n_945), .Y(n_944) );
AOI22xp33_ASAP7_75t_L g599 ( .A1(n_137), .A2(n_369), .B1(n_519), .B2(n_600), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_137), .A2(n_676), .B(n_678), .Y(n_675) );
OAI22xp5_ASAP7_75t_L g1132 ( .A1(n_138), .A2(n_311), .B1(n_755), .B2(n_913), .Y(n_1132) );
OAI22xp5_ASAP7_75t_L g1135 ( .A1(n_138), .A2(n_311), .B1(n_833), .B2(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g881 ( .A(n_139), .Y(n_881) );
INVx1_ASAP7_75t_L g1130 ( .A(n_140), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1072 ( .A1(n_141), .A2(n_345), .B1(n_1073), .B2(n_1074), .Y(n_1072) );
OAI22xp33_ASAP7_75t_L g1076 ( .A1(n_141), .A2(n_308), .B1(n_393), .B2(n_1077), .Y(n_1076) );
INVx1_ASAP7_75t_L g1092 ( .A(n_142), .Y(n_1092) );
AOI22xp33_ASAP7_75t_SL g1697 ( .A1(n_142), .A2(n_239), .B1(n_1690), .B2(n_1692), .Y(n_1697) );
AOI22xp33_ASAP7_75t_SL g1608 ( .A1(n_143), .A2(n_297), .B1(n_467), .B2(n_948), .Y(n_1608) );
AOI21xp33_ASAP7_75t_L g1624 ( .A1(n_143), .A2(n_676), .B(n_1401), .Y(n_1624) );
INVx1_ASAP7_75t_L g1155 ( .A(n_144), .Y(n_1155) );
INVx1_ASAP7_75t_L g422 ( .A(n_145), .Y(n_422) );
INVx1_ASAP7_75t_L g820 ( .A(n_146), .Y(n_820) );
INVx1_ASAP7_75t_L g1000 ( .A(n_147), .Y(n_1000) );
OAI211xp5_ASAP7_75t_L g1008 ( .A1(n_147), .A2(n_1009), .B(n_1010), .C(n_1012), .Y(n_1008) );
OAI211xp5_ASAP7_75t_L g1174 ( .A1(n_148), .A2(n_828), .B(n_1175), .C(n_1177), .Y(n_1174) );
INVx1_ASAP7_75t_L g1189 ( .A(n_148), .Y(n_1189) );
AOI22xp33_ASAP7_75t_L g1274 ( .A1(n_149), .A2(n_205), .B1(n_1255), .B2(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g784 ( .A(n_150), .Y(n_784) );
INVx1_ASAP7_75t_L g1166 ( .A(n_151), .Y(n_1166) );
OAI22xp5_ASAP7_75t_L g1280 ( .A1(n_153), .A2(n_216), .B1(n_633), .B2(n_1281), .Y(n_1280) );
INVx1_ASAP7_75t_L g1309 ( .A(n_153), .Y(n_1309) );
INVx1_ASAP7_75t_L g1497 ( .A(n_154), .Y(n_1497) );
INVx1_ASAP7_75t_L g1498 ( .A(n_155), .Y(n_1498) );
OAI211xp5_ASAP7_75t_L g1221 ( .A1(n_156), .A2(n_450), .B(n_1222), .C(n_1224), .Y(n_1221) );
INVx1_ASAP7_75t_L g1233 ( .A(n_156), .Y(n_1233) );
INVx1_ASAP7_75t_L g974 ( .A(n_157), .Y(n_974) );
INVx1_ASAP7_75t_L g613 ( .A(n_158), .Y(n_613) );
OAI221xp5_ASAP7_75t_L g660 ( .A1(n_158), .A2(n_218), .B1(n_661), .B2(n_665), .C(n_669), .Y(n_660) );
OAI221xp5_ASAP7_75t_L g1411 ( .A1(n_159), .A2(n_356), .B1(n_1215), .B2(n_1412), .C(n_1414), .Y(n_1411) );
INVx1_ASAP7_75t_L g1430 ( .A(n_159), .Y(n_1430) );
INVx1_ASAP7_75t_L g1399 ( .A(n_160), .Y(n_1399) );
AOI22xp33_ASAP7_75t_L g1425 ( .A1(n_160), .A2(n_286), .B1(n_535), .B2(n_1299), .Y(n_1425) );
INVx1_ASAP7_75t_L g1655 ( .A(n_161), .Y(n_1655) );
CKINVDCx5p33_ASAP7_75t_R g1404 ( .A(n_162), .Y(n_1404) );
INVx1_ASAP7_75t_L g1432 ( .A(n_163), .Y(n_1432) );
INVx1_ASAP7_75t_L g1651 ( .A(n_164), .Y(n_1651) );
INVx1_ASAP7_75t_L g850 ( .A(n_165), .Y(n_850) );
OAI211xp5_ASAP7_75t_L g853 ( .A1(n_165), .A2(n_854), .B(n_855), .C(n_856), .Y(n_853) );
INVx1_ASAP7_75t_L g916 ( .A(n_166), .Y(n_916) );
OAI211xp5_ASAP7_75t_L g927 ( .A1(n_166), .A2(n_718), .B(n_828), .C(n_928), .Y(n_927) );
OAI211xp5_ASAP7_75t_L g1068 ( .A1(n_167), .A2(n_718), .B(n_772), .C(n_1069), .Y(n_1068) );
INVx1_ASAP7_75t_L g1088 ( .A(n_167), .Y(n_1088) );
INVx1_ASAP7_75t_L g1106 ( .A(n_168), .Y(n_1106) );
OAI22xp33_ASAP7_75t_L g1992 ( .A1(n_169), .A2(n_284), .B1(n_826), .B2(n_930), .Y(n_1992) );
OAI22xp5_ASAP7_75t_L g1994 ( .A1(n_169), .A2(n_284), .B1(n_920), .B2(n_921), .Y(n_1994) );
OAI22xp33_ASAP7_75t_L g1935 ( .A1(n_172), .A2(n_187), .B1(n_1073), .B2(n_1936), .Y(n_1935) );
OAI22xp33_ASAP7_75t_L g1939 ( .A1(n_172), .A2(n_187), .B1(n_921), .B2(n_1940), .Y(n_1939) );
INVx1_ASAP7_75t_L g878 ( .A(n_173), .Y(n_878) );
INVx1_ASAP7_75t_L g1965 ( .A(n_174), .Y(n_1965) );
INVx1_ASAP7_75t_L g1971 ( .A(n_176), .Y(n_1971) );
INVx1_ASAP7_75t_L g1517 ( .A(n_177), .Y(n_1517) );
INVx1_ASAP7_75t_L g1162 ( .A(n_178), .Y(n_1162) );
INVx1_ASAP7_75t_L g1652 ( .A(n_180), .Y(n_1652) );
OAI22xp33_ASAP7_75t_L g1662 ( .A1(n_181), .A2(n_364), .B1(n_844), .B2(n_995), .Y(n_1662) );
OAI22xp33_ASAP7_75t_L g1669 ( .A1(n_181), .A2(n_364), .B1(n_393), .B2(n_1077), .Y(n_1669) );
INVx1_ASAP7_75t_L g1933 ( .A(n_182), .Y(n_1933) );
INVx1_ASAP7_75t_L g717 ( .A(n_183), .Y(n_717) );
OAI211xp5_ASAP7_75t_L g1127 ( .A1(n_184), .A2(n_1009), .B(n_1128), .C(n_1129), .Y(n_1127) );
INVx1_ASAP7_75t_L g1141 ( .A(n_184), .Y(n_1141) );
INVx1_ASAP7_75t_L g802 ( .A(n_185), .Y(n_802) );
OAI22xp33_ASAP7_75t_L g1986 ( .A1(n_186), .A2(n_214), .B1(n_774), .B2(n_1074), .Y(n_1986) );
OAI22xp33_ASAP7_75t_L g1995 ( .A1(n_186), .A2(n_214), .B1(n_1079), .B2(n_1081), .Y(n_1995) );
XNOR2xp5_ASAP7_75t_L g410 ( .A(n_188), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g1646 ( .A(n_189), .Y(n_1646) );
INVx1_ASAP7_75t_L g883 ( .A(n_190), .Y(n_883) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_191), .A2(n_329), .B1(n_551), .B2(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g1500 ( .A(n_192), .Y(n_1500) );
INVx1_ASAP7_75t_L g1911 ( .A(n_193), .Y(n_1911) );
AOI221xp5_ASAP7_75t_L g1555 ( .A1(n_194), .A2(n_362), .B1(n_1263), .B2(n_1556), .C(n_1558), .Y(n_1555) );
AOI22xp33_ASAP7_75t_L g1584 ( .A1(n_194), .A2(n_374), .B1(n_602), .B2(n_796), .Y(n_1584) );
XOR2x2_ASAP7_75t_L g961 ( .A(n_196), .B(n_962), .Y(n_961) );
INVxp67_ASAP7_75t_SL g1460 ( .A(n_197), .Y(n_1460) );
AOI22xp33_ASAP7_75t_L g1628 ( .A1(n_198), .A2(n_297), .B1(n_418), .B2(n_569), .Y(n_1628) );
CKINVDCx5p33_ASAP7_75t_R g1272 ( .A(n_199), .Y(n_1272) );
INVx1_ASAP7_75t_L g999 ( .A(n_200), .Y(n_999) );
INVx1_ASAP7_75t_L g978 ( .A(n_201), .Y(n_978) );
INVx1_ASAP7_75t_L g1390 ( .A(n_202), .Y(n_1390) );
INVx1_ASAP7_75t_L g437 ( .A(n_204), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_204), .A2(n_317), .B1(n_474), .B2(n_481), .Y(n_473) );
INVx1_ASAP7_75t_L g1320 ( .A(n_205), .Y(n_1320) );
XNOR2xp5_ASAP7_75t_L g687 ( .A(n_206), .B(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g801 ( .A(n_207), .Y(n_801) );
INVx1_ASAP7_75t_L g914 ( .A(n_209), .Y(n_914) );
OAI22xp33_ASAP7_75t_L g1180 ( .A1(n_210), .A2(n_365), .B1(n_1066), .B2(n_1074), .Y(n_1180) );
OAI22xp33_ASAP7_75t_L g1184 ( .A1(n_210), .A2(n_365), .B1(n_1079), .B2(n_1081), .Y(n_1184) );
INVx1_ASAP7_75t_L g871 ( .A(n_211), .Y(n_871) );
INVx1_ASAP7_75t_L g1098 ( .A(n_212), .Y(n_1098) );
AOI221x1_ASAP7_75t_SL g1259 ( .A1(n_213), .A2(n_285), .B1(n_1260), .B2(n_1262), .C(n_1264), .Y(n_1259) );
AOI21xp33_ASAP7_75t_L g1322 ( .A1(n_213), .A2(n_592), .B(n_1323), .Y(n_1322) );
INVx2_ASAP7_75t_L g1685 ( .A(n_215), .Y(n_1685) );
AND2x2_ASAP7_75t_L g1688 ( .A(n_215), .B(n_1686), .Y(n_1688) );
AND2x2_ASAP7_75t_L g1693 ( .A(n_215), .B(n_320), .Y(n_1693) );
OAI22xp33_ASAP7_75t_L g1001 ( .A1(n_217), .A2(n_283), .B1(n_489), .B2(n_926), .Y(n_1001) );
OAI22xp33_ASAP7_75t_L g1014 ( .A1(n_217), .A2(n_283), .B1(n_755), .B2(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g609 ( .A(n_218), .Y(n_609) );
INVx1_ASAP7_75t_L g918 ( .A(n_219), .Y(n_918) );
AOI22xp5_ASAP7_75t_L g1716 ( .A1(n_220), .A2(n_275), .B1(n_1687), .B2(n_1690), .Y(n_1716) );
INVx1_ASAP7_75t_L g849 ( .A(n_222), .Y(n_849) );
INVx1_ASAP7_75t_L g1070 ( .A(n_223), .Y(n_1070) );
OAI22xp5_ASAP7_75t_L g1532 ( .A1(n_224), .A2(n_1533), .B1(n_1587), .B2(n_1588), .Y(n_1532) );
INVxp67_ASAP7_75t_L g1588 ( .A(n_224), .Y(n_1588) );
CKINVDCx5p33_ASAP7_75t_R g1267 ( .A(n_225), .Y(n_1267) );
AOI22xp33_ASAP7_75t_L g1717 ( .A1(n_226), .A2(n_229), .B1(n_1682), .B2(n_1701), .Y(n_1717) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_227), .A2(n_361), .B1(n_544), .B2(n_560), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g950 ( .A1(n_227), .A2(n_235), .B1(n_951), .B2(n_953), .Y(n_950) );
INVx1_ASAP7_75t_L g1518 ( .A(n_230), .Y(n_1518) );
OAI211xp5_ASAP7_75t_L g1523 ( .A1(n_230), .A2(n_1010), .B(n_1524), .C(n_1525), .Y(n_1523) );
XOR2x2_ASAP7_75t_L g1190 ( .A(n_231), .B(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g695 ( .A(n_232), .Y(n_695) );
OAI211xp5_ASAP7_75t_L g1931 ( .A1(n_233), .A2(n_828), .B(n_1028), .C(n_1932), .Y(n_1931) );
INVx1_ASAP7_75t_L g1946 ( .A(n_233), .Y(n_1946) );
OAI221xp5_ASAP7_75t_SL g1547 ( .A1(n_234), .A2(n_312), .B1(n_1548), .B2(n_1549), .C(n_1550), .Y(n_1547) );
INVx1_ASAP7_75t_L g1565 ( .A(n_234), .Y(n_1565) );
AOI22xp33_ASAP7_75t_SL g942 ( .A1(n_235), .A2(n_358), .B1(n_544), .B2(n_568), .Y(n_942) );
AOI22xp33_ASAP7_75t_L g1444 ( .A1(n_236), .A2(n_332), .B1(n_1157), .B2(n_1344), .Y(n_1444) );
INVx1_ASAP7_75t_L g971 ( .A(n_237), .Y(n_971) );
INVx1_ASAP7_75t_L g1046 ( .A(n_238), .Y(n_1046) );
INVx1_ASAP7_75t_L g1380 ( .A(n_240), .Y(n_1380) );
INVx1_ASAP7_75t_L g972 ( .A(n_241), .Y(n_972) );
INVx2_ASAP7_75t_L g461 ( .A(n_242), .Y(n_461) );
INVx1_ASAP7_75t_L g530 ( .A(n_242), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_242), .B(n_478), .Y(n_588) );
AOI22xp5_ASAP7_75t_L g1702 ( .A1(n_243), .A2(n_368), .B1(n_1682), .B2(n_1687), .Y(n_1702) );
INVx1_ASAP7_75t_L g1649 ( .A(n_244), .Y(n_1649) );
INVx1_ASAP7_75t_L g1111 ( .A(n_245), .Y(n_1111) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_248), .A2(n_254), .B1(n_859), .B2(n_860), .Y(n_1227) );
OAI22xp33_ASAP7_75t_L g1234 ( .A1(n_248), .A2(n_254), .B1(n_775), .B2(n_1066), .Y(n_1234) );
CKINVDCx5p33_ASAP7_75t_R g1201 ( .A(n_249), .Y(n_1201) );
XNOR2xp5_ASAP7_75t_L g570 ( .A(n_250), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g1916 ( .A(n_251), .Y(n_1916) );
INVx1_ASAP7_75t_L g1103 ( .A(n_252), .Y(n_1103) );
AOI22xp33_ASAP7_75t_SL g512 ( .A1(n_253), .A2(n_329), .B1(n_513), .B2(n_517), .Y(n_512) );
OAI22xp33_ASAP7_75t_L g817 ( .A1(n_255), .A2(n_282), .B1(n_393), .B2(n_744), .Y(n_817) );
OAI22xp5_ASAP7_75t_L g825 ( .A1(n_255), .A2(n_282), .B1(n_762), .B2(n_826), .Y(n_825) );
BUFx3_ASAP7_75t_L g472 ( .A(n_256), .Y(n_472) );
INVx1_ASAP7_75t_L g1538 ( .A(n_257), .Y(n_1538) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_258), .A2(n_277), .B1(n_554), .B2(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g980 ( .A(n_259), .Y(n_980) );
INVx1_ASAP7_75t_L g1179 ( .A(n_260), .Y(n_1179) );
OAI211xp5_ASAP7_75t_L g1185 ( .A1(n_260), .A2(n_748), .B(n_1186), .C(n_1188), .Y(n_1185) );
INVx1_ASAP7_75t_L g708 ( .A(n_261), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g595 ( .A1(n_262), .A2(n_331), .B1(n_517), .B2(n_596), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_262), .A2(n_279), .B1(n_657), .B2(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g1480 ( .A(n_263), .Y(n_1480) );
INVx1_ASAP7_75t_L g753 ( .A(n_264), .Y(n_753) );
OAI211xp5_ASAP7_75t_SL g764 ( .A1(n_264), .A2(n_765), .B(n_767), .C(n_772), .Y(n_764) );
INVx1_ASAP7_75t_L g868 ( .A(n_265), .Y(n_868) );
CKINVDCx5p33_ASAP7_75t_R g1198 ( .A(n_267), .Y(n_1198) );
AOI21xp33_ASAP7_75t_L g1400 ( .A1(n_268), .A2(n_552), .B(n_1401), .Y(n_1400) );
INVx1_ASAP7_75t_L g1034 ( .A(n_269), .Y(n_1034) );
INVx1_ASAP7_75t_L g874 ( .A(n_270), .Y(n_874) );
INVx1_ASAP7_75t_L g1298 ( .A(n_271), .Y(n_1298) );
INVx1_ASAP7_75t_L g1598 ( .A(n_272), .Y(n_1598) );
INVx1_ASAP7_75t_L g1973 ( .A(n_273), .Y(n_1973) );
INVx1_ASAP7_75t_L g1436 ( .A(n_274), .Y(n_1436) );
BUFx3_ASAP7_75t_L g401 ( .A(n_278), .Y(n_401) );
INVx1_ASAP7_75t_L g433 ( .A(n_278), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g1519 ( .A1(n_280), .A2(n_328), .B1(n_489), .B2(n_833), .Y(n_1519) );
OAI22xp5_ASAP7_75t_L g1529 ( .A1(n_280), .A2(n_328), .B1(n_755), .B2(n_757), .Y(n_1529) );
INVx1_ASAP7_75t_L g1607 ( .A(n_281), .Y(n_1607) );
INVx1_ASAP7_75t_L g1319 ( .A(n_285), .Y(n_1319) );
INVx1_ASAP7_75t_L g1246 ( .A(n_288), .Y(n_1246) );
INVx1_ASAP7_75t_L g1568 ( .A(n_289), .Y(n_1568) );
INVx1_ASAP7_75t_L g1027 ( .A(n_290), .Y(n_1027) );
INVx1_ASAP7_75t_L g794 ( .A(n_291), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_292), .Y(n_1204) );
OAI22xp5_ASAP7_75t_L g924 ( .A1(n_293), .A2(n_375), .B1(n_925), .B2(n_926), .Y(n_924) );
INVx1_ASAP7_75t_L g1501 ( .A(n_294), .Y(n_1501) );
CKINVDCx5p33_ASAP7_75t_R g1354 ( .A(n_295), .Y(n_1354) );
INVx1_ASAP7_75t_L g471 ( .A(n_298), .Y(n_471) );
INVx1_ASAP7_75t_L g494 ( .A(n_298), .Y(n_494) );
INVx1_ASAP7_75t_L g1666 ( .A(n_300), .Y(n_1666) );
OAI211xp5_ASAP7_75t_L g1670 ( .A1(n_300), .A2(n_855), .B(n_1186), .C(n_1671), .Y(n_1670) );
OAI22xp5_ASAP7_75t_L g1589 ( .A1(n_301), .A2(n_1590), .B1(n_1591), .B2(n_1634), .Y(n_1589) );
INVxp67_ASAP7_75t_L g1634 ( .A(n_301), .Y(n_1634) );
INVx1_ASAP7_75t_L g1160 ( .A(n_302), .Y(n_1160) );
CKINVDCx5p33_ASAP7_75t_R g1225 ( .A(n_304), .Y(n_1225) );
INVxp67_ASAP7_75t_SL g1595 ( .A(n_305), .Y(n_1595) );
OAI221xp5_ASAP7_75t_L g1630 ( .A1(n_305), .A2(n_363), .B1(n_625), .B2(n_1631), .C(n_1632), .Y(n_1630) );
INVx1_ASAP7_75t_L g1030 ( .A(n_306), .Y(n_1030) );
OAI211xp5_ASAP7_75t_L g818 ( .A1(n_307), .A2(n_746), .B(n_748), .C(n_819), .Y(n_818) );
INVx1_ASAP7_75t_L g831 ( .A(n_307), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g1200 ( .A(n_309), .Y(n_1200) );
INVx1_ASAP7_75t_L g1504 ( .A(n_310), .Y(n_1504) );
INVx1_ASAP7_75t_L g1574 ( .A(n_312), .Y(n_1574) );
CKINVDCx5p33_ASAP7_75t_R g1599 ( .A(n_313), .Y(n_1599) );
INVx1_ASAP7_75t_L g1990 ( .A(n_314), .Y(n_1990) );
INVx1_ASAP7_75t_L g976 ( .A(n_315), .Y(n_976) );
AOI22xp5_ASAP7_75t_SL g1713 ( .A1(n_316), .A2(n_372), .B1(n_1690), .B2(n_1701), .Y(n_1713) );
INVx1_ASAP7_75t_L g441 ( .A(n_317), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g1348 ( .A(n_318), .Y(n_1348) );
INVxp67_ASAP7_75t_SL g670 ( .A(n_319), .Y(n_670) );
INVx1_ASAP7_75t_L g1686 ( .A(n_320), .Y(n_1686) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_320), .B(n_1685), .Y(n_1691) );
CKINVDCx5p33_ASAP7_75t_R g1206 ( .A(n_321), .Y(n_1206) );
OAI211xp5_ASAP7_75t_SL g1987 ( .A1(n_322), .A2(n_828), .B(n_1988), .C(n_1989), .Y(n_1987) );
INVx1_ASAP7_75t_L g1998 ( .A(n_322), .Y(n_1998) );
INVx1_ASAP7_75t_L g444 ( .A(n_323), .Y(n_444) );
INVx1_ASAP7_75t_L g1335 ( .A(n_325), .Y(n_1335) );
INVx1_ASAP7_75t_L g1934 ( .A(n_326), .Y(n_1934) );
OAI211xp5_ASAP7_75t_L g1944 ( .A1(n_326), .A2(n_450), .B(n_1215), .C(n_1945), .Y(n_1944) );
OAI211xp5_ASAP7_75t_L g997 ( .A1(n_327), .A2(n_772), .B(n_847), .C(n_998), .Y(n_997) );
INVx1_ASAP7_75t_L g1013 ( .A(n_327), .Y(n_1013) );
INVx1_ASAP7_75t_L g647 ( .A(n_330), .Y(n_647) );
INVx1_ASAP7_75t_L g1467 ( .A(n_332), .Y(n_1467) );
INVx1_ASAP7_75t_L g1901 ( .A(n_333), .Y(n_1901) );
INVx1_ASAP7_75t_L g1603 ( .A(n_334), .Y(n_1603) );
INVx1_ASAP7_75t_L g1410 ( .A(n_335), .Y(n_1410) );
INVx1_ASAP7_75t_L g785 ( .A(n_336), .Y(n_785) );
INVx1_ASAP7_75t_L g1654 ( .A(n_337), .Y(n_1654) );
INVx1_ASAP7_75t_L g1226 ( .A(n_338), .Y(n_1226) );
OAI211xp5_ASAP7_75t_L g1230 ( .A1(n_338), .A2(n_772), .B(n_1231), .C(n_1232), .Y(n_1230) );
CKINVDCx5p33_ASAP7_75t_R g1610 ( .A(n_339), .Y(n_1610) );
OAI22xp5_ASAP7_75t_L g906 ( .A1(n_340), .A2(n_907), .B1(n_956), .B2(n_957), .Y(n_906) );
INVxp67_ASAP7_75t_SL g957 ( .A(n_340), .Y(n_957) );
AOI211xp5_ASAP7_75t_SL g1376 ( .A1(n_341), .A2(n_438), .B(n_1377), .C(n_1379), .Y(n_1376) );
INVx1_ASAP7_75t_L g1108 ( .A(n_342), .Y(n_1108) );
AOI21xp5_ASAP7_75t_SL g1405 ( .A1(n_343), .A2(n_552), .B(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1418 ( .A(n_343), .Y(n_1418) );
INVx1_ASAP7_75t_L g720 ( .A(n_344), .Y(n_720) );
INVx1_ASAP7_75t_L g1466 ( .A(n_346), .Y(n_1466) );
XNOR2xp5_ASAP7_75t_L g1147 ( .A(n_347), .B(n_1148), .Y(n_1147) );
INVx1_ASAP7_75t_L g1164 ( .A(n_348), .Y(n_1164) );
INVx1_ASAP7_75t_L g1910 ( .A(n_349), .Y(n_1910) );
INVx1_ASAP7_75t_L g1492 ( .A(n_350), .Y(n_1492) );
INVx1_ASAP7_75t_L g1902 ( .A(n_351), .Y(n_1902) );
XOR2x2_ASAP7_75t_L g1487 ( .A(n_352), .B(n_1488), .Y(n_1487) );
INVxp67_ASAP7_75t_L g1424 ( .A(n_353), .Y(n_1424) );
OAI211xp5_ASAP7_75t_L g845 ( .A1(n_354), .A2(n_772), .B(n_846), .C(n_848), .Y(n_845) );
INVx1_ASAP7_75t_L g857 ( .A(n_354), .Y(n_857) );
CKINVDCx5p33_ASAP7_75t_R g1195 ( .A(n_355), .Y(n_1195) );
INVxp67_ASAP7_75t_SL g1435 ( .A(n_356), .Y(n_1435) );
BUFx6f_ASAP7_75t_L g397 ( .A(n_357), .Y(n_397) );
AOI22xp33_ASAP7_75t_SL g947 ( .A1(n_358), .A2(n_361), .B1(n_520), .B2(n_948), .Y(n_947) );
CKINVDCx5p33_ASAP7_75t_R g1285 ( .A(n_360), .Y(n_1285) );
INVx1_ASAP7_75t_L g1578 ( .A(n_362), .Y(n_1578) );
INVx1_ASAP7_75t_L g1597 ( .A(n_363), .Y(n_1597) );
INVx1_ASAP7_75t_L g415 ( .A(n_366), .Y(n_415) );
INVx1_ASAP7_75t_L g1071 ( .A(n_367), .Y(n_1071) );
OAI211xp5_ASAP7_75t_L g1084 ( .A1(n_367), .A2(n_746), .B(n_748), .C(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g457 ( .A(n_370), .Y(n_457) );
INVx2_ASAP7_75t_L g511 ( .A(n_370), .Y(n_511) );
INVx1_ASAP7_75t_L g529 ( .A(n_370), .Y(n_529) );
CKINVDCx5p33_ASAP7_75t_R g1288 ( .A(n_371), .Y(n_1288) );
CKINVDCx5p33_ASAP7_75t_R g1337 ( .A(n_373), .Y(n_1337) );
INVx1_ASAP7_75t_L g911 ( .A(n_375), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_402), .B(n_1674), .Y(n_376) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx4f_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_387), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g1952 ( .A(n_381), .B(n_390), .Y(n_1952) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_383), .B(n_385), .Y(n_382) );
NOR2xp33_ASAP7_75t_L g1956 ( .A(n_383), .B(n_386), .Y(n_1956) );
INVx1_ASAP7_75t_L g2001 ( .A(n_383), .Y(n_2001) );
HB1xp67_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g2003 ( .A(n_386), .B(n_2001), .Y(n_2003) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_389), .B(n_392), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AND2x4_ASAP7_75t_L g453 ( .A(n_390), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AND2x4_ASAP7_75t_L g564 ( .A(n_391), .B(n_401), .Y(n_564) );
AND2x4_ASAP7_75t_L g679 ( .A(n_391), .B(n_400), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_392), .A2(n_429), .B1(n_430), .B2(n_431), .Y(n_428) );
INVxp67_ASAP7_75t_SL g920 ( .A(n_392), .Y(n_920) );
INVx1_ASAP7_75t_L g1940 ( .A(n_392), .Y(n_1940) );
AND2x4_ASAP7_75t_SL g1951 ( .A(n_392), .B(n_1952), .Y(n_1951) );
INVx3_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g393 ( .A(n_394), .B(n_399), .Y(n_393) );
OR2x6_ASAP7_75t_L g756 ( .A(n_394), .B(n_432), .Y(n_756) );
BUFx4f_ASAP7_75t_L g885 ( .A(n_394), .Y(n_885) );
INVx1_ASAP7_75t_L g1062 ( .A(n_394), .Y(n_1062) );
INVxp67_ASAP7_75t_L g1494 ( .A(n_394), .Y(n_1494) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx4f_ASAP7_75t_L g726 ( .A(n_395), .Y(n_726) );
INVx3_ASAP7_75t_L g870 ( .A(n_395), .Y(n_870) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_397), .B(n_398), .Y(n_396) );
INVx2_ASAP7_75t_L g420 ( .A(n_397), .Y(n_420) );
INVx2_ASAP7_75t_L g427 ( .A(n_397), .Y(n_427) );
AND2x2_ASAP7_75t_L g434 ( .A(n_397), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_L g440 ( .A(n_397), .B(n_398), .Y(n_440) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
NAND2x1_ASAP7_75t_L g674 ( .A(n_397), .B(n_398), .Y(n_674) );
INVx1_ASAP7_75t_L g421 ( .A(n_398), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_398), .B(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g435 ( .A(n_398), .Y(n_435) );
BUFx2_ASAP7_75t_L g443 ( .A(n_398), .Y(n_443) );
AND2x2_ASAP7_75t_L g549 ( .A(n_398), .B(n_427), .Y(n_549) );
OR2x2_ASAP7_75t_L g734 ( .A(n_398), .B(n_420), .Y(n_734) );
OR2x6_ASAP7_75t_L g1007 ( .A(n_399), .B(n_870), .Y(n_1007) );
INVxp67_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g452 ( .A(n_400), .Y(n_452) );
INVx2_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
BUFx2_ASAP7_75t_L g417 ( .A(n_401), .Y(n_417) );
AND2x4_ASAP7_75t_L g447 ( .A(n_401), .B(n_448), .Y(n_447) );
XNOR2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_1237), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_1143), .B1(n_1144), .B2(n_1236), .Y(n_403) );
INVx1_ASAP7_75t_L g1236 ( .A(n_404), .Y(n_1236) );
AOI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_1090), .B2(n_1142), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
XNOR2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_836), .Y(n_406) );
AOI22xp33_ASAP7_75t_SL g407 ( .A1(n_408), .A2(n_409), .B1(n_686), .B2(n_835), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
XNOR2x1_ASAP7_75t_L g409 ( .A(n_410), .B(n_570), .Y(n_409) );
NAND3x1_ASAP7_75t_L g411 ( .A(n_412), .B(n_507), .C(n_536), .Y(n_411) );
AOI22xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_453), .B1(n_458), .B2(n_465), .Y(n_412) );
NAND4xp25_ASAP7_75t_L g413 ( .A(n_414), .B(n_428), .C(n_436), .D(n_450), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_415), .A2(n_416), .B1(n_422), .B2(n_423), .Y(n_414) );
AOI22xp33_ASAP7_75t_L g487 ( .A1(n_415), .A2(n_422), .B1(n_488), .B2(n_495), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g910 ( .A1(n_416), .A2(n_911), .B1(n_912), .B2(n_914), .Y(n_910) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
OR2x2_ASAP7_75t_L g424 ( .A(n_417), .B(n_425), .Y(n_424) );
AND2x4_ASAP7_75t_L g442 ( .A(n_417), .B(n_443), .Y(n_442) );
AND2x2_ASAP7_75t_L g750 ( .A(n_417), .B(n_443), .Y(n_750) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_418), .Y(n_657) );
INVx3_ASAP7_75t_L g1358 ( .A(n_418), .Y(n_1358) );
A2O1A1Ixp33_ASAP7_75t_L g1370 ( .A1(n_418), .A2(n_1337), .B(n_1371), .C(n_1375), .Y(n_1370) );
A2O1A1Ixp33_ASAP7_75t_L g1473 ( .A1(n_418), .A2(n_1451), .B(n_1474), .C(n_1477), .Y(n_1473) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
INVx3_ASAP7_75t_L g545 ( .A(n_419), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_419), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g646 ( .A(n_419), .B(n_642), .Y(n_646) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
HB1xp67_ASAP7_75t_L g1374 ( .A(n_420), .Y(n_1374) );
INVx2_ASAP7_75t_L g913 ( .A(n_423), .Y(n_913) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx2_ASAP7_75t_L g758 ( .A(n_424), .Y(n_758) );
BUFx2_ASAP7_75t_L g1083 ( .A(n_424), .Y(n_1083) );
INVx8_ASAP7_75t_L g729 ( .A(n_425), .Y(n_729) );
BUFx2_ASAP7_75t_L g1121 ( .A(n_425), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_429), .A2(n_430), .B1(n_500), .B2(n_502), .Y(n_499) );
INVx4_ASAP7_75t_L g744 ( .A(n_431), .Y(n_744) );
INVx3_ASAP7_75t_SL g921 ( .A(n_431), .Y(n_921) );
CKINVDCx16_ASAP7_75t_R g1077 ( .A(n_431), .Y(n_1077) );
AND2x4_ASAP7_75t_L g431 ( .A(n_432), .B(n_434), .Y(n_431) );
HB1xp67_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx6f_ASAP7_75t_L g553 ( .A(n_434), .Y(n_553) );
BUFx3_ASAP7_75t_L g653 ( .A(n_434), .Y(n_653) );
INVx2_ASAP7_75t_L g677 ( .A(n_434), .Y(n_677) );
AOI222xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_438), .B1(n_441), .B2(n_442), .C1(n_444), .C2(n_445), .Y(n_436) );
BUFx3_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x2_ASAP7_75t_L g451 ( .A(n_439), .B(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g654 ( .A(n_439), .Y(n_654) );
AND2x6_ASAP7_75t_L g659 ( .A(n_439), .B(n_626), .Y(n_659) );
AND2x4_ASAP7_75t_SL g664 ( .A(n_439), .B(n_642), .Y(n_664) );
BUFx6f_ASAP7_75t_L g1263 ( .A(n_439), .Y(n_1263) );
BUFx6f_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g558 ( .A(n_440), .Y(n_558) );
AOI22xp33_ASAP7_75t_L g819 ( .A1(n_442), .A2(n_447), .B1(n_820), .B2(n_821), .Y(n_819) );
AOI22xp33_ASAP7_75t_L g1012 ( .A1(n_442), .A2(n_447), .B1(n_999), .B2(n_1013), .Y(n_1012) );
BUFx3_ASAP7_75t_L g1086 ( .A(n_442), .Y(n_1086) );
INVx1_ASAP7_75t_L g667 ( .A(n_443), .Y(n_667) );
INVx1_ASAP7_75t_L g1283 ( .A(n_443), .Y(n_1283) );
AOI22xp33_ASAP7_75t_L g1372 ( .A1(n_443), .A2(n_1332), .B1(n_1352), .B2(n_1373), .Y(n_1372) );
BUFx2_ASAP7_75t_L g1476 ( .A(n_443), .Y(n_1476) );
AOI211xp5_ASAP7_75t_L g466 ( .A1(n_444), .A2(n_467), .B(n_473), .C(n_485), .Y(n_466) );
AOI222xp33_ASAP7_75t_L g915 ( .A1(n_445), .A2(n_654), .B1(n_750), .B2(n_916), .C1(n_917), .C2(n_918), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g1129 ( .A1(n_445), .A2(n_750), .B1(n_1130), .B2(n_1131), .Y(n_1129) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
INVx2_ASAP7_75t_L g752 ( .A(n_446), .Y(n_752) );
INVx2_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
BUFx3_ASAP7_75t_L g1087 ( .A(n_447), .Y(n_1087) );
INVx2_ASAP7_75t_L g1527 ( .A(n_447), .Y(n_1527) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_448), .B(n_626), .Y(n_634) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND3xp33_ASAP7_75t_L g909 ( .A(n_450), .B(n_910), .C(n_915), .Y(n_909) );
INVx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g748 ( .A(n_451), .Y(n_748) );
INVx1_ASAP7_75t_L g855 ( .A(n_451), .Y(n_855) );
AND2x2_ASAP7_75t_L g1011 ( .A(n_452), .B(n_562), .Y(n_1011) );
BUFx3_ASAP7_75t_L g759 ( .A(n_453), .Y(n_759) );
BUFx2_ASAP7_75t_SL g823 ( .A(n_453), .Y(n_823) );
BUFx2_ASAP7_75t_L g922 ( .A(n_453), .Y(n_922) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x2_ASAP7_75t_L g633 ( .A(n_455), .B(n_634), .Y(n_633) );
INVxp67_ASAP7_75t_L g637 ( .A(n_455), .Y(n_637) );
INVx1_ASAP7_75t_L g1287 ( .A(n_455), .Y(n_1287) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g464 ( .A(n_456), .Y(n_464) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OAI31xp33_ASAP7_75t_L g840 ( .A1(n_458), .A2(n_841), .A3(n_845), .B(n_851), .Y(n_840) );
OAI31xp33_ASAP7_75t_L g923 ( .A1(n_458), .A2(n_924), .A3(n_927), .B(n_929), .Y(n_923) );
OAI31xp33_ASAP7_75t_L g1173 ( .A1(n_458), .A2(n_1174), .A3(n_1180), .B(n_1181), .Y(n_1173) );
OAI31xp33_ASAP7_75t_L g1228 ( .A1(n_458), .A2(n_1229), .A3(n_1230), .B(n_1234), .Y(n_1228) );
AOI211xp5_ASAP7_75t_L g1591 ( .A1(n_458), .A2(n_1592), .B(n_1604), .C(n_1615), .Y(n_1591) );
AND2x4_ASAP7_75t_L g458 ( .A(n_459), .B(n_462), .Y(n_458) );
AND2x2_ASAP7_75t_SL g777 ( .A(n_459), .B(n_462), .Y(n_777) );
AND2x2_ASAP7_75t_L g1002 ( .A(n_459), .B(n_462), .Y(n_1002) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_459), .B(n_462), .Y(n_1439) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_459), .B(n_462), .Y(n_1520) );
INVx1_ASAP7_75t_SL g459 ( .A(n_460), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
AND3x4_ASAP7_75t_L g509 ( .A(n_461), .B(n_477), .C(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g580 ( .A(n_461), .Y(n_580) );
NAND2xp33_ASAP7_75t_SL g693 ( .A(n_461), .B(n_478), .Y(n_693) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
INVx1_ASAP7_75t_L g566 ( .A(n_464), .Y(n_566) );
OR2x2_ASAP7_75t_L g587 ( .A(n_464), .B(n_588), .Y(n_587) );
OR2x2_ASAP7_75t_L g692 ( .A(n_464), .B(n_693), .Y(n_692) );
AND2x2_ASAP7_75t_SL g1123 ( .A(n_464), .B(n_564), .Y(n_1123) );
NAND3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_487), .C(n_499), .Y(n_465) );
INVx1_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx2_ASAP7_75t_L g955 ( .A(n_468), .Y(n_955) );
INVx1_ASAP7_75t_L g1346 ( .A(n_468), .Y(n_1346) );
INVx2_ASAP7_75t_L g1586 ( .A(n_468), .Y(n_1586) );
INVx2_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
AND2x4_ASAP7_75t_L g485 ( .A(n_469), .B(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g517 ( .A(n_469), .Y(n_517) );
BUFx2_ASAP7_75t_L g535 ( .A(n_469), .Y(n_535) );
BUFx2_ASAP7_75t_L g576 ( .A(n_469), .Y(n_576) );
BUFx3_ASAP7_75t_L g1300 ( .A(n_469), .Y(n_1300) );
BUFx2_ASAP7_75t_L g1310 ( .A(n_469), .Y(n_1310) );
BUFx2_ASAP7_75t_L g1600 ( .A(n_469), .Y(n_1600) );
AND2x4_ASAP7_75t_L g469 ( .A(n_470), .B(n_472), .Y(n_469) );
INVx1_ASAP7_75t_L g523 ( .A(n_470), .Y(n_523) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g484 ( .A(n_471), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_471), .B(n_472), .Y(n_498) );
BUFx6f_ASAP7_75t_L g480 ( .A(n_472), .Y(n_480) );
OR2x2_ASAP7_75t_L g492 ( .A(n_472), .B(n_493), .Y(n_492) );
INVx2_ASAP7_75t_L g506 ( .A(n_472), .Y(n_506) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
AOI22xp33_ASAP7_75t_L g998 ( .A1(n_475), .A2(n_482), .B1(n_999), .B2(n_1000), .Y(n_998) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_475), .A2(n_482), .B1(n_1070), .B2(n_1071), .Y(n_1069) );
AOI22xp33_ASAP7_75t_SL g1140 ( .A1(n_475), .A2(n_482), .B1(n_1130), .B2(n_1141), .Y(n_1140) );
AOI22xp33_ASAP7_75t_SL g1232 ( .A1(n_475), .A2(n_482), .B1(n_1225), .B2(n_1233), .Y(n_1232) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_475), .A2(n_482), .B1(n_1435), .B2(n_1436), .Y(n_1434) );
AOI22xp33_ASAP7_75t_L g1516 ( .A1(n_475), .A2(n_482), .B1(n_1517), .B2(n_1518), .Y(n_1516) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_479), .Y(n_475) );
AND2x4_ASAP7_75t_L g482 ( .A(n_476), .B(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g769 ( .A(n_476), .B(n_479), .Y(n_769) );
A2O1A1Ixp33_ASAP7_75t_L g1428 ( .A1(n_476), .A2(n_1429), .B(n_1431), .C(n_1434), .Y(n_1428) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx3_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g486 ( .A(n_478), .Y(n_486) );
BUFx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g522 ( .A(n_480), .B(n_523), .Y(n_522) );
INVx2_ASAP7_75t_L g612 ( .A(n_480), .Y(n_612) );
NAND2x1p5_ASAP7_75t_L g632 ( .A(n_480), .B(n_484), .Y(n_632) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_482), .Y(n_770) );
AOI22xp33_ASAP7_75t_SL g848 ( .A1(n_482), .A2(n_830), .B1(n_849), .B2(n_850), .Y(n_848) );
BUFx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
CKINVDCx8_ASAP7_75t_R g772 ( .A(n_485), .Y(n_772) );
CKINVDCx8_ASAP7_75t_R g828 ( .A(n_485), .Y(n_828) );
OAI31xp33_ASAP7_75t_L g1427 ( .A1(n_485), .A2(n_1428), .A3(n_1437), .B(n_1439), .Y(n_1427) );
INVx1_ASAP7_75t_L g491 ( .A(n_486), .Y(n_491) );
OR2x6_ASAP7_75t_L g496 ( .A(n_486), .B(n_497), .Y(n_496) );
OR2x4_ASAP7_75t_L g501 ( .A(n_486), .B(n_492), .Y(n_501) );
NAND3x1_ASAP7_75t_L g527 ( .A(n_486), .B(n_528), .C(n_530), .Y(n_527) );
AND2x4_ASAP7_75t_L g579 ( .A(n_486), .B(n_580), .Y(n_579) );
NAND2x1p5_ASAP7_75t_L g605 ( .A(n_486), .B(n_530), .Y(n_605) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx3_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
BUFx2_ASAP7_75t_L g774 ( .A(n_490), .Y(n_774) );
INVx2_ASAP7_75t_SL g1067 ( .A(n_490), .Y(n_1067) );
BUFx2_ASAP7_75t_L g1438 ( .A(n_490), .Y(n_1438) );
OR2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g502 ( .A(n_491), .B(n_503), .Y(n_502) );
INVx2_ASAP7_75t_L g584 ( .A(n_492), .Y(n_584) );
BUFx3_ASAP7_75t_L g696 ( .A(n_492), .Y(n_696) );
BUFx3_ASAP7_75t_L g894 ( .A(n_492), .Y(n_894) );
BUFx4f_ASAP7_75t_L g1026 ( .A(n_492), .Y(n_1026) );
INVx1_ASAP7_75t_L g516 ( .A(n_493), .Y(n_516) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVxp67_ASAP7_75t_L g505 ( .A(n_494), .Y(n_505) );
INVx2_ASAP7_75t_L g926 ( .A(n_495), .Y(n_926) );
AOI22xp33_ASAP7_75t_L g1593 ( .A1(n_495), .A2(n_502), .B1(n_1594), .B2(n_1595), .Y(n_1593) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g776 ( .A(n_496), .Y(n_776) );
INVx1_ASAP7_75t_L g834 ( .A(n_496), .Y(n_834) );
BUFx3_ASAP7_75t_L g1074 ( .A(n_496), .Y(n_1074) );
BUFx3_ASAP7_75t_L g799 ( .A(n_497), .Y(n_799) );
INVx1_ASAP7_75t_L g901 ( .A(n_497), .Y(n_901) );
BUFx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g623 ( .A(n_498), .Y(n_623) );
INVx2_ASAP7_75t_L g930 ( .A(n_500), .Y(n_930) );
AOI22xp33_ASAP7_75t_L g1601 ( .A1(n_500), .A2(n_1067), .B1(n_1602), .B2(n_1603), .Y(n_1601) );
INVx2_ASAP7_75t_SL g500 ( .A(n_501), .Y(n_500) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_501), .Y(n_762) );
INVx2_ASAP7_75t_SL g843 ( .A(n_501), .Y(n_843) );
INVx1_ASAP7_75t_L g996 ( .A(n_501), .Y(n_996) );
INVx1_ASAP7_75t_L g1937 ( .A(n_501), .Y(n_1937) );
INVx1_ASAP7_75t_L g763 ( .A(n_502), .Y(n_763) );
INVx1_ASAP7_75t_L g826 ( .A(n_502), .Y(n_826) );
INVx2_ASAP7_75t_L g844 ( .A(n_502), .Y(n_844) );
INVxp67_ASAP7_75t_L g925 ( .A(n_502), .Y(n_925) );
INVx1_ASAP7_75t_L g1073 ( .A(n_502), .Y(n_1073) );
BUFx6f_ASAP7_75t_L g519 ( .A(n_503), .Y(n_519) );
INVx1_ASAP7_75t_L g709 ( .A(n_503), .Y(n_709) );
BUFx6f_ASAP7_75t_L g898 ( .A(n_503), .Y(n_898) );
INVx2_ASAP7_75t_L g992 ( .A(n_503), .Y(n_992) );
INVx2_ASAP7_75t_L g1921 ( .A(n_503), .Y(n_1921) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
BUFx8_ASAP7_75t_L g592 ( .A(n_504), .Y(n_592) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_504), .Y(n_703) );
INVx2_ASAP7_75t_L g797 ( .A(n_504), .Y(n_797) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g515 ( .A(n_506), .B(n_516), .Y(n_515) );
AOI33xp33_ASAP7_75t_L g507 ( .A1(n_508), .A2(n_512), .A3(n_518), .B1(n_524), .B2(n_525), .B3(n_531), .Y(n_507) );
NAND3xp33_ASAP7_75t_L g943 ( .A(n_508), .B(n_944), .C(n_947), .Y(n_943) );
BUFx3_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
AOI33xp33_ASAP7_75t_L g594 ( .A1(n_509), .A2(n_595), .A3(n_599), .B1(n_601), .B2(n_603), .B3(n_606), .Y(n_594) );
AOI33xp33_ASAP7_75t_L g1338 ( .A1(n_509), .A2(n_603), .A3(n_1339), .B1(n_1340), .B2(n_1341), .B3(n_1345), .Y(n_1338) );
NAND3xp33_ASAP7_75t_L g1443 ( .A(n_509), .B(n_1444), .C(n_1445), .Y(n_1443) );
INVx1_ASAP7_75t_L g685 ( .A(n_510), .Y(n_685) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g541 ( .A(n_511), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g1279 ( .A(n_511), .B(n_626), .Y(n_1279) );
BUFx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
INVx1_ASAP7_75t_L g1582 ( .A(n_514), .Y(n_1582) );
BUFx3_ASAP7_75t_L g514 ( .A(n_515), .Y(n_514) );
INVx8_ASAP7_75t_L g533 ( .A(n_515), .Y(n_533) );
BUFx3_ASAP7_75t_L g598 ( .A(n_515), .Y(n_598) );
NAND2x1p5_ASAP7_75t_L g636 ( .A(n_515), .B(n_579), .Y(n_636) );
HB1xp67_ASAP7_75t_L g1305 ( .A(n_515), .Y(n_1305) );
INVx1_ASAP7_75t_L g985 ( .A(n_519), .Y(n_985) );
INVx1_ASAP7_75t_L g1510 ( .A(n_519), .Y(n_1510) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx2_ASAP7_75t_R g600 ( .A(n_521), .Y(n_600) );
INVx1_ASAP7_75t_L g953 ( .A(n_521), .Y(n_953) );
INVx5_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
BUFx12f_ASAP7_75t_L g602 ( .A(n_522), .Y(n_602) );
BUFx3_ASAP7_75t_L g1308 ( .A(n_522), .Y(n_1308) );
BUFx3_ASAP7_75t_L g1344 ( .A(n_522), .Y(n_1344) );
INVx1_ASAP7_75t_L g617 ( .A(n_523), .Y(n_617) );
BUFx2_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g904 ( .A(n_526), .Y(n_904) );
BUFx2_ASAP7_75t_L g1925 ( .A(n_526), .Y(n_1925) );
INVx3_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx3_ASAP7_75t_L g713 ( .A(n_527), .Y(n_713) );
OAI33xp33_ASAP7_75t_L g1505 ( .A1(n_527), .A2(n_782), .A3(n_1506), .B1(n_1508), .B2(n_1509), .B3(n_1511), .Y(n_1505) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g578 ( .A(n_529), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g1254 ( .A(n_529), .B(n_642), .Y(n_1254) );
AOI22xp33_ASAP7_75t_L g1431 ( .A1(n_532), .A2(n_703), .B1(n_1432), .B2(n_1433), .Y(n_1431) );
INVx8_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g607 ( .A(n_533), .Y(n_607) );
CKINVDCx5p33_ASAP7_75t_R g1299 ( .A(n_533), .Y(n_1299) );
INVx2_ASAP7_75t_L g1334 ( .A(n_533), .Y(n_1334) );
HB1xp67_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
AOI33xp33_ASAP7_75t_L g536 ( .A1(n_537), .A2(n_543), .A3(n_550), .B1(n_559), .B2(n_563), .B3(n_567), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
OAI33xp33_ASAP7_75t_L g721 ( .A1(n_538), .A2(n_722), .A3(n_730), .B1(n_738), .B2(n_740), .B3(n_741), .Y(n_721) );
OAI33xp33_ASAP7_75t_L g804 ( .A1(n_538), .A2(n_740), .A3(n_805), .B1(n_809), .B2(n_810), .B3(n_814), .Y(n_804) );
OAI33xp33_ASAP7_75t_L g1208 ( .A1(n_538), .A2(n_889), .A3(n_1209), .B1(n_1212), .B2(n_1216), .B3(n_1218), .Y(n_1208) );
OAI33xp33_ASAP7_75t_L g1490 ( .A1(n_538), .A2(n_889), .A3(n_1491), .B1(n_1496), .B2(n_1499), .B3(n_1502), .Y(n_1490) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g866 ( .A(n_540), .Y(n_866) );
INVx2_ASAP7_75t_L g1048 ( .A(n_540), .Y(n_1048) );
INVx1_ASAP7_75t_L g1169 ( .A(n_540), .Y(n_1169) );
INVx1_ASAP7_75t_L g1269 ( .A(n_540), .Y(n_1269) );
AND2x4_ASAP7_75t_L g540 ( .A(n_541), .B(n_542), .Y(n_540) );
OR2x6_ASAP7_75t_L g604 ( .A(n_541), .B(n_605), .Y(n_604) );
INVx1_ASAP7_75t_L g1326 ( .A(n_541), .Y(n_1326) );
INVx1_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
INVx2_ASAP7_75t_L g1275 ( .A(n_545), .Y(n_1275) );
INVx2_ASAP7_75t_L g1560 ( .A(n_545), .Y(n_1560) );
INVx2_ASAP7_75t_SL g1563 ( .A(n_545), .Y(n_1563) );
INVx1_ASAP7_75t_L g1571 ( .A(n_545), .Y(n_1571) );
INVx1_ASAP7_75t_SL g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
BUFx3_ASAP7_75t_L g935 ( .A(n_548), .Y(n_935) );
BUFx3_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_549), .Y(n_569) );
BUFx3_ASAP7_75t_L g681 ( .A(n_549), .Y(n_681) );
INVx2_ASAP7_75t_L g1256 ( .A(n_549), .Y(n_1256) );
BUFx3_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g649 ( .A(n_553), .B(n_642), .Y(n_649) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_553), .B(n_642), .Y(n_1290) );
INVx2_ASAP7_75t_L g1368 ( .A(n_553), .Y(n_1368) );
INVx1_ASAP7_75t_L g1557 ( .A(n_553), .Y(n_1557) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
AOI221xp5_ASAP7_75t_L g1564 ( .A1(n_556), .A2(n_1373), .B1(n_1413), .B2(n_1552), .C(n_1565), .Y(n_1564) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g562 ( .A(n_558), .Y(n_562) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx2_ASAP7_75t_L g740 ( .A(n_563), .Y(n_740) );
CKINVDCx5p33_ASAP7_75t_R g889 ( .A(n_563), .Y(n_889) );
NAND3xp33_ASAP7_75t_L g938 ( .A(n_563), .B(n_939), .C(n_942), .Y(n_938) );
AND2x4_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
INVx1_ASAP7_75t_SL g655 ( .A(n_564), .Y(n_655) );
OAI21xp33_ASAP7_75t_L g1377 ( .A1(n_564), .A2(n_877), .B(n_1378), .Y(n_1377) );
INVx4_ASAP7_75t_L g1401 ( .A(n_564), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1479 ( .A1(n_564), .A2(n_673), .B1(n_877), .B2(n_1480), .C(n_1481), .Y(n_1479) );
NAND2xp5_ASAP7_75t_L g1914 ( .A(n_564), .B(n_565), .Y(n_1914) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
AND2x4_ASAP7_75t_L g641 ( .A(n_569), .B(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_569), .Y(n_658) );
INVx1_ASAP7_75t_L g1464 ( .A(n_569), .Y(n_1464) );
AND3x1_ASAP7_75t_L g571 ( .A(n_572), .B(n_618), .C(n_638), .Y(n_571) );
NOR3xp33_ASAP7_75t_L g572 ( .A(n_573), .B(n_581), .C(n_593), .Y(n_572) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OAI211xp5_ASAP7_75t_SL g1576 ( .A1(n_574), .A2(n_691), .B(n_1577), .C(n_1583), .Y(n_1576) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g1350 ( .A1(n_575), .A2(n_1351), .B1(n_1352), .B2(n_1353), .C(n_1354), .Y(n_1350) );
AOI221xp5_ASAP7_75t_L g1456 ( .A1(n_575), .A2(n_1351), .B1(n_1353), .B2(n_1457), .C(n_1458), .Y(n_1456) );
AND2x4_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
AND2x2_ASAP7_75t_L g610 ( .A(n_577), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_L g614 ( .A(n_577), .B(n_615), .Y(n_614) );
AND2x4_ASAP7_75t_SL g1351 ( .A(n_577), .B(n_611), .Y(n_1351) );
AND2x4_ASAP7_75t_SL g1353 ( .A(n_577), .B(n_615), .Y(n_1353) );
AND2x4_ASAP7_75t_L g577 ( .A(n_578), .B(n_579), .Y(n_577) );
OR2x2_ASAP7_75t_L g624 ( .A(n_578), .B(n_625), .Y(n_624) );
AND2x6_ASAP7_75t_L g1294 ( .A(n_579), .B(n_611), .Y(n_1294) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_579), .B(n_617), .Y(n_1296) );
INVx1_ASAP7_75t_L g1302 ( .A(n_579), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1539 ( .A(n_582), .B(n_1540), .Y(n_1539) );
OR2x6_ASAP7_75t_L g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx2_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g716 ( .A(n_584), .Y(n_716) );
INVxp67_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g1544 ( .A(n_586), .B(n_1423), .Y(n_1544) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx1_ASAP7_75t_L g591 ( .A(n_587), .Y(n_591) );
OR2x2_ASAP7_75t_L g621 ( .A(n_587), .B(n_622), .Y(n_621) );
OR2x2_ASAP7_75t_L g630 ( .A(n_587), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g1313 ( .A(n_588), .Y(n_1313) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_590), .B(n_1348), .Y(n_1347) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_590), .B(n_1447), .Y(n_1446) );
AND2x4_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
AND2x4_ASAP7_75t_L g1333 ( .A(n_591), .B(n_1334), .Y(n_1333) );
INVx3_ASAP7_75t_L g952 ( .A(n_592), .Y(n_952) );
INVx2_ASAP7_75t_SL g1107 ( .A(n_592), .Y(n_1107) );
INVx3_ASAP7_75t_L g1161 ( .A(n_592), .Y(n_1161) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_608), .Y(n_593) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
BUFx3_ASAP7_75t_L g948 ( .A(n_598), .Y(n_948) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_602), .A2(n_1300), .B1(n_1410), .B2(n_1430), .Y(n_1429) );
NAND3xp33_ASAP7_75t_L g1452 ( .A(n_603), .B(n_1453), .C(n_1454), .Y(n_1452) );
INVx1_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
OAI33xp33_ASAP7_75t_L g981 ( .A1(n_604), .A2(n_782), .A3(n_982), .B1(n_984), .B2(n_987), .B3(n_991), .Y(n_981) );
OAI33xp33_ASAP7_75t_L g1095 ( .A1(n_604), .A2(n_1096), .A3(n_1097), .B1(n_1101), .B2(n_1105), .B3(n_1109), .Y(n_1095) );
INVx3_ASAP7_75t_L g1317 ( .A(n_605), .Y(n_1317) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B1(n_613), .B2(n_614), .Y(n_608) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_619), .A2(n_627), .B(n_628), .Y(n_618) );
INVx8_ASAP7_75t_L g619 ( .A(n_620), .Y(n_619) );
AND2x4_ASAP7_75t_L g620 ( .A(n_621), .B(n_624), .Y(n_620) );
INVx1_ASAP7_75t_L g1336 ( .A(n_621), .Y(n_1336) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
BUFx6f_ASAP7_75t_L g706 ( .A(n_623), .Y(n_706) );
INVx1_ASAP7_75t_L g1250 ( .A(n_624), .Y(n_1250) );
INVx1_ASAP7_75t_L g668 ( .A(n_626), .Y(n_668) );
HB1xp67_ASAP7_75t_L g1375 ( .A(n_626), .Y(n_1375) );
AND2x4_ASAP7_75t_L g629 ( .A(n_630), .B(n_633), .Y(n_629) );
INVx2_ASAP7_75t_L g1331 ( .A(n_630), .Y(n_1331) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_631), .Y(n_699) );
INVx3_ASAP7_75t_L g719 ( .A(n_631), .Y(n_719) );
INVx4_ASAP7_75t_L g766 ( .A(n_631), .Y(n_766) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
BUFx3_ASAP7_75t_L g787 ( .A(n_632), .Y(n_787) );
BUFx2_ASAP7_75t_L g990 ( .A(n_632), .Y(n_990) );
INVx1_ASAP7_75t_L g1633 ( .A(n_634), .Y(n_1633) );
OR2x2_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
OR2x6_ASAP7_75t_L g1386 ( .A(n_636), .B(n_637), .Y(n_1386) );
OAI21xp5_ASAP7_75t_SL g638 ( .A1(n_639), .A2(n_660), .B(n_682), .Y(n_638) );
INVx3_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx2_ASAP7_75t_L g1365 ( .A(n_642), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1573 ( .A(n_642), .B(n_1255), .Y(n_1573) );
AOI22xp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B1(n_647), .B2(n_648), .Y(n_643) );
INVx1_ASAP7_75t_L g1618 ( .A(n_645), .Y(n_1618) );
BUFx6f_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
AND2x4_ASAP7_75t_L g1286 ( .A(n_646), .B(n_1287), .Y(n_1286) );
BUFx6f_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g1621 ( .A(n_649), .Y(n_1621) );
AOI21xp5_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_656), .B(n_659), .Y(n_650) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
BUFx2_ASAP7_75t_L g934 ( .A(n_653), .Y(n_934) );
A2O1A1Ixp33_ASAP7_75t_SL g1409 ( .A1(n_657), .A2(n_1375), .B(n_1410), .C(n_1411), .Y(n_1409) );
AOI211xp5_ASAP7_75t_SL g1629 ( .A1(n_659), .A2(n_1575), .B(n_1598), .C(n_1630), .Y(n_1629) );
INVx2_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx4_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
BUFx3_ASAP7_75t_L g1575 ( .A(n_664), .Y(n_1575) );
INVx2_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
INVx2_ASAP7_75t_L g1631 ( .A(n_666), .Y(n_1631) );
NOR2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
INVx1_ASAP7_75t_L g1413 ( .A(n_667), .Y(n_1413) );
INVx1_ASAP7_75t_L g1477 ( .A(n_668), .Y(n_1477) );
OAI211xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_671), .B(n_675), .C(n_680), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g1124 ( .A1(n_671), .A2(n_880), .B1(n_1099), .B2(n_1111), .Y(n_1124) );
INVx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g1063 ( .A(n_672), .Y(n_1063) );
INVx2_ASAP7_75t_L g1217 ( .A(n_672), .Y(n_1217) );
INVx1_ASAP7_75t_L g1524 ( .A(n_672), .Y(n_1524) );
INVx4_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
BUFx4f_ASAP7_75t_L g854 ( .A(n_673), .Y(n_854) );
BUFx4f_ASAP7_75t_L g882 ( .A(n_673), .Y(n_882) );
BUFx4f_ASAP7_75t_L g1009 ( .A(n_673), .Y(n_1009) );
BUFx4f_ASAP7_75t_L g1056 ( .A(n_673), .Y(n_1056) );
BUFx6f_ASAP7_75t_L g1215 ( .A(n_673), .Y(n_1215) );
OR2x6_ASAP7_75t_L g1276 ( .A(n_673), .B(n_1277), .Y(n_1276) );
BUFx6f_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
BUFx3_ASAP7_75t_L g737 ( .A(n_674), .Y(n_737) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g941 ( .A(n_677), .Y(n_941) );
INVx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g1359 ( .A1(n_679), .A2(n_1217), .B1(n_1360), .B2(n_1361), .C(n_1362), .Y(n_1359) );
INVx1_ASAP7_75t_L g1406 ( .A(n_679), .Y(n_1406) );
OAI221xp5_ASAP7_75t_L g1465 ( .A1(n_679), .A2(n_1217), .B1(n_1466), .B2(n_1467), .C(n_1468), .Y(n_1465) );
INVx2_ASAP7_75t_L g1558 ( .A(n_679), .Y(n_1558) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g1615 ( .A1(n_683), .A2(n_1616), .B(n_1629), .Y(n_1615) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
BUFx2_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI31xp33_ASAP7_75t_L g1355 ( .A1(n_685), .A2(n_1356), .A3(n_1363), .B(n_1376), .Y(n_1355) );
HB1xp67_ASAP7_75t_L g1393 ( .A(n_685), .Y(n_1393) );
OAI31xp33_ASAP7_75t_L g1461 ( .A1(n_685), .A2(n_1462), .A3(n_1469), .B(n_1478), .Y(n_1461) );
INVx1_ASAP7_75t_L g835 ( .A(n_686), .Y(n_835) );
XOR2x2_ASAP7_75t_L g686 ( .A(n_687), .B(n_778), .Y(n_686) );
AND3x1_ASAP7_75t_L g688 ( .A(n_689), .B(n_742), .C(n_760), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_721), .Y(n_689) );
OAI33xp33_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_694), .A3(n_700), .B1(n_707), .B2(n_712), .B3(n_714), .Y(n_690) );
OAI33xp33_ASAP7_75t_L g1150 ( .A1(n_691), .A2(n_1042), .A3(n_1151), .B1(n_1154), .B2(n_1159), .B3(n_1163), .Y(n_1150) );
OAI33xp33_ASAP7_75t_L g1962 ( .A1(n_691), .A2(n_1042), .A3(n_1963), .B1(n_1966), .B2(n_1969), .B3(n_1972), .Y(n_1962) );
BUFx4f_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
BUFx8_ASAP7_75t_L g782 ( .A(n_692), .Y(n_782) );
BUFx4f_ASAP7_75t_L g1022 ( .A(n_692), .Y(n_1022) );
BUFx2_ASAP7_75t_L g1096 ( .A(n_692), .Y(n_1096) );
BUFx2_ASAP7_75t_L g1323 ( .A(n_693), .Y(n_1323) );
OAI22xp33_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_696), .B1(n_697), .B2(n_698), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g722 ( .A1(n_695), .A2(n_717), .B1(n_723), .B2(n_727), .Y(n_722) );
OAI22xp33_ASAP7_75t_L g783 ( .A1(n_696), .A2(n_784), .B1(n_785), .B2(n_786), .Y(n_783) );
OAI22xp33_ASAP7_75t_L g800 ( .A1(n_696), .A2(n_801), .B1(n_802), .B2(n_803), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g1109 ( .A1(n_696), .A2(n_1110), .B1(n_1111), .B2(n_1112), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1315 ( .A1(n_696), .A2(n_1267), .B1(n_1273), .B2(n_1316), .C(n_1317), .Y(n_1315) );
OAI22xp33_ASAP7_75t_L g1650 ( .A1(n_696), .A2(n_1165), .B1(n_1651), .B2(n_1652), .Y(n_1650) );
OAI22xp5_ASAP7_75t_L g738 ( .A1(n_697), .A2(n_720), .B1(n_731), .B2(n_739), .Y(n_738) );
HB1xp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g1040 ( .A(n_699), .Y(n_1040) );
OAI22xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_704), .B2(n_705), .Y(n_700) );
OAI22xp5_ASAP7_75t_L g730 ( .A1(n_701), .A2(n_708), .B1(n_731), .B2(n_735), .Y(n_730) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx5_ASAP7_75t_L g791 ( .A(n_703), .Y(n_791) );
INVx3_ASAP7_75t_L g1033 ( .A(n_703), .Y(n_1033) );
INVx2_ASAP7_75t_SL g1343 ( .A(n_703), .Y(n_1343) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_704), .A2(n_710), .B1(n_725), .B2(n_727), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g788 ( .A1(n_705), .A2(n_789), .B1(n_790), .B2(n_792), .Y(n_788) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_705), .A2(n_972), .B1(n_980), .B2(n_992), .Y(n_991) );
OAI22xp5_ASAP7_75t_L g1202 ( .A1(n_705), .A2(n_790), .B1(n_1203), .B2(n_1204), .Y(n_1202) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_705), .A2(n_897), .B1(n_1319), .B2(n_1320), .Y(n_1318) );
OAI221xp5_ASAP7_75t_L g1416 ( .A1(n_705), .A2(n_1417), .B1(n_1418), .B2(n_1419), .C(n_1420), .Y(n_1416) );
OAI221xp5_ASAP7_75t_L g1421 ( .A1(n_705), .A2(n_1404), .B1(n_1422), .B2(n_1424), .C(n_1425), .Y(n_1421) );
OAI22xp5_ASAP7_75t_L g1508 ( .A1(n_705), .A2(n_1422), .B1(n_1497), .B2(n_1503), .Y(n_1508) );
OAI221xp5_ASAP7_75t_L g1605 ( .A1(n_705), .A2(n_1037), .B1(n_1606), .B2(n_1607), .C(n_1608), .Y(n_1605) );
CKINVDCx8_ASAP7_75t_R g705 ( .A(n_706), .Y(n_705) );
INVx3_ASAP7_75t_L g711 ( .A(n_706), .Y(n_711) );
INVx3_ASAP7_75t_L g986 ( .A(n_706), .Y(n_986) );
INVx1_ASAP7_75t_L g1104 ( .A(n_706), .Y(n_1104) );
INVx3_ASAP7_75t_L g1922 ( .A(n_706), .Y(n_1922) );
OAI22xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_710), .B2(n_711), .Y(n_707) );
OAI22xp5_ASAP7_75t_L g1199 ( .A1(n_709), .A2(n_899), .B1(n_1200), .B2(n_1201), .Y(n_1199) );
OAI22xp5_ASAP7_75t_L g1043 ( .A1(n_711), .A2(n_1044), .B1(n_1045), .B2(n_1046), .Y(n_1043) );
OAI22xp5_ASAP7_75t_L g1159 ( .A1(n_711), .A2(n_1160), .B1(n_1161), .B2(n_1162), .Y(n_1159) );
OAI22xp5_ASAP7_75t_L g1969 ( .A1(n_711), .A2(n_1031), .B1(n_1970), .B2(n_1971), .Y(n_1969) );
OAI33xp33_ASAP7_75t_L g781 ( .A1(n_712), .A2(n_782), .A3(n_783), .B1(n_788), .B2(n_793), .B3(n_800), .Y(n_781) );
OAI33xp33_ASAP7_75t_L g1193 ( .A1(n_712), .A2(n_782), .A3(n_1194), .B1(n_1199), .B2(n_1202), .B3(n_1205), .Y(n_1193) );
OAI33xp33_ASAP7_75t_L g1642 ( .A1(n_712), .A2(n_1021), .A3(n_1643), .B1(n_1647), .B2(n_1650), .B3(n_1653), .Y(n_1642) );
CKINVDCx5p33_ASAP7_75t_R g712 ( .A(n_713), .Y(n_712) );
NAND3xp33_ASAP7_75t_L g949 ( .A(n_713), .B(n_950), .C(n_954), .Y(n_949) );
INVx2_ASAP7_75t_L g1042 ( .A(n_713), .Y(n_1042) );
INVx2_ASAP7_75t_L g1426 ( .A(n_713), .Y(n_1426) );
NAND3xp33_ASAP7_75t_L g1583 ( .A(n_713), .B(n_1584), .C(n_1585), .Y(n_1583) );
OAI22xp33_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_717), .B1(n_718), .B2(n_720), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g1097 ( .A1(n_715), .A2(n_1098), .B1(n_1099), .B2(n_1100), .Y(n_1097) );
BUFx4f_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_716), .A2(n_966), .B1(n_974), .B2(n_983), .Y(n_982) );
OAI22xp33_ASAP7_75t_L g987 ( .A1(n_716), .A2(n_967), .B1(n_976), .B2(n_988), .Y(n_987) );
OAI22xp5_ASAP7_75t_L g1647 ( .A1(n_716), .A2(n_1165), .B1(n_1648), .B2(n_1649), .Y(n_1647) );
INVx2_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx2_ASAP7_75t_L g847 ( .A(n_719), .Y(n_847) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
BUFx6f_ASAP7_75t_L g807 ( .A(n_726), .Y(n_807) );
INVx4_ASAP7_75t_L g1381 ( .A(n_726), .Y(n_1381) );
OAI22xp5_ASAP7_75t_L g814 ( .A1(n_727), .A2(n_792), .B1(n_798), .B2(n_815), .Y(n_814) );
OAI22xp33_ASAP7_75t_L g1168 ( .A1(n_727), .A2(n_815), .B1(n_1152), .B2(n_1164), .Y(n_1168) );
OAI22xp5_ASAP7_75t_L g1660 ( .A1(n_727), .A2(n_869), .B1(n_1646), .B2(n_1655), .Y(n_1660) );
OAI22xp33_ASAP7_75t_L g1976 ( .A1(n_727), .A2(n_815), .B1(n_1964), .B2(n_1973), .Y(n_1976) );
INVx6_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx5_ASAP7_75t_L g887 ( .A(n_728), .Y(n_887) );
BUFx6f_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g808 ( .A(n_729), .Y(n_808) );
INVx2_ASAP7_75t_L g872 ( .A(n_729), .Y(n_872) );
INVx2_ASAP7_75t_L g969 ( .A(n_729), .Y(n_969) );
INVx2_ASAP7_75t_SL g1053 ( .A(n_729), .Y(n_1053) );
INVx4_ASAP7_75t_L g1119 ( .A(n_729), .Y(n_1119) );
INVx2_ASAP7_75t_L g1472 ( .A(n_729), .Y(n_1472) );
INVx1_ASAP7_75t_L g1984 ( .A(n_729), .Y(n_1984) );
OAI22xp5_ASAP7_75t_L g809 ( .A1(n_731), .A2(n_735), .B1(n_789), .B2(n_794), .Y(n_809) );
OAI22xp5_ASAP7_75t_L g1216 ( .A1(n_731), .A2(n_1198), .B1(n_1207), .B2(n_1217), .Y(n_1216) );
INVx4_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx2_ASAP7_75t_L g1362 ( .A(n_733), .Y(n_1362) );
INVx2_ASAP7_75t_L g1468 ( .A(n_733), .Y(n_1468) );
INVx2_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
BUFx2_ASAP7_75t_L g813 ( .A(n_734), .Y(n_813) );
BUFx3_ASAP7_75t_L g877 ( .A(n_734), .Y(n_877) );
BUFx2_ASAP7_75t_L g1116 ( .A(n_734), .Y(n_1116) );
INVx1_ASAP7_75t_L g1214 ( .A(n_734), .Y(n_1214) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_735), .A2(n_880), .B1(n_971), .B2(n_972), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g1171 ( .A1(n_735), .A2(n_1055), .B1(n_1153), .B2(n_1166), .Y(n_1171) );
OAI22xp5_ASAP7_75t_L g1499 ( .A1(n_735), .A2(n_1213), .B1(n_1500), .B2(n_1501), .Y(n_1499) );
OAI211xp5_ASAP7_75t_L g1567 ( .A1(n_735), .A2(n_1568), .B(n_1569), .C(n_1570), .Y(n_1567) );
OAI22xp5_ASAP7_75t_L g1658 ( .A1(n_735), .A2(n_880), .B1(n_1644), .B2(n_1654), .Y(n_1658) );
OAI22xp5_ASAP7_75t_L g1977 ( .A1(n_735), .A2(n_1967), .B1(n_1970), .B2(n_1978), .Y(n_1977) );
OAI22xp33_ASAP7_75t_L g1980 ( .A1(n_735), .A2(n_1965), .B1(n_1974), .B2(n_1981), .Y(n_1980) );
INVx5_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
INVx2_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_SL g739 ( .A(n_737), .Y(n_739) );
BUFx3_ASAP7_75t_L g747 ( .A(n_737), .Y(n_747) );
OR2x2_ASAP7_75t_L g1257 ( .A(n_737), .B(n_1254), .Y(n_1257) );
NAND2xp5_ASAP7_75t_L g1371 ( .A(n_737), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_737), .B(n_1475), .Y(n_1474) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_739), .A2(n_785), .B1(n_802), .B2(n_811), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g1659 ( .A1(n_739), .A2(n_811), .B1(n_1649), .B2(n_1652), .Y(n_1659) );
OAI33xp33_ASAP7_75t_L g1047 ( .A1(n_740), .A2(n_1048), .A3(n_1049), .B1(n_1054), .B2(n_1057), .B3(n_1058), .Y(n_1047) );
OAI33xp33_ASAP7_75t_L g1167 ( .A1(n_740), .A2(n_1168), .A3(n_1169), .B1(n_1170), .B2(n_1171), .B3(n_1172), .Y(n_1167) );
OAI33xp33_ASAP7_75t_L g1656 ( .A1(n_740), .A2(n_1269), .A3(n_1657), .B1(n_1658), .B2(n_1659), .B3(n_1660), .Y(n_1656) );
OAI33xp33_ASAP7_75t_L g1975 ( .A1(n_740), .A2(n_1169), .A3(n_1976), .B1(n_1977), .B2(n_1980), .B3(n_1982), .Y(n_1975) );
OAI31xp33_ASAP7_75t_L g742 ( .A1(n_743), .A2(n_745), .A3(n_754), .B(n_759), .Y(n_742) );
BUFx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g1223 ( .A(n_747), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g1622 ( .A1(n_747), .A2(n_1623), .B(n_1624), .C(n_1625), .Y(n_1622) );
OAI211xp5_ASAP7_75t_SL g1626 ( .A1(n_747), .A2(n_1610), .B(n_1627), .C(n_1628), .Y(n_1626) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_751), .B1(n_752), .B2(n_753), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g856 ( .A1(n_750), .A2(n_752), .B1(n_849), .B2(n_857), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g1224 ( .A1(n_750), .A2(n_752), .B1(n_1225), .B2(n_1226), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1525 ( .A1(n_750), .A2(n_1517), .B1(n_1526), .B2(n_1528), .Y(n_1525) );
AOI22xp33_ASAP7_75t_L g1671 ( .A1(n_750), .A2(n_1526), .B1(n_1665), .B2(n_1672), .Y(n_1671) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_751), .A2(n_768), .B1(n_770), .B2(n_771), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_752), .A2(n_1086), .B1(n_1178), .B2(n_1189), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1997 ( .A1(n_752), .A2(n_1086), .B1(n_1990), .B2(n_1998), .Y(n_1997) );
BUFx6f_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
BUFx2_ASAP7_75t_L g859 ( .A(n_756), .Y(n_859) );
INVx1_ASAP7_75t_L g1080 ( .A(n_756), .Y(n_1080) );
HB1xp67_ASAP7_75t_L g1942 ( .A(n_756), .Y(n_1942) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g860 ( .A(n_758), .Y(n_860) );
INVx1_ASAP7_75t_L g1015 ( .A(n_758), .Y(n_1015) );
OAI31xp33_ASAP7_75t_L g1219 ( .A1(n_759), .A2(n_1220), .A3(n_1221), .B(n_1227), .Y(n_1219) );
OAI31xp33_ASAP7_75t_L g1521 ( .A1(n_759), .A2(n_1522), .A3(n_1523), .B(n_1529), .Y(n_1521) );
OAI31xp33_ASAP7_75t_L g1668 ( .A1(n_759), .A2(n_1669), .A3(n_1670), .B(n_1673), .Y(n_1668) );
OAI31xp33_ASAP7_75t_SL g1938 ( .A1(n_759), .A2(n_1939), .A3(n_1941), .B(n_1944), .Y(n_1938) );
OAI31xp33_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_764), .A3(n_773), .B(n_777), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g905 ( .A1(n_765), .A2(n_871), .B1(n_883), .B2(n_892), .Y(n_905) );
INVx2_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
INVx1_ASAP7_75t_L g895 ( .A(n_766), .Y(n_895) );
INVx1_ASAP7_75t_L g983 ( .A(n_766), .Y(n_983) );
INVx2_ASAP7_75t_L g1316 ( .A(n_766), .Y(n_1316) );
INVx1_ASAP7_75t_L g1512 ( .A(n_766), .Y(n_1512) );
AOI22xp33_ASAP7_75t_L g928 ( .A1(n_768), .A2(n_770), .B1(n_917), .B2(n_918), .Y(n_928) );
AOI22xp33_ASAP7_75t_L g1177 ( .A1(n_768), .A2(n_770), .B1(n_1178), .B2(n_1179), .Y(n_1177) );
AOI22xp33_ASAP7_75t_L g1989 ( .A1(n_768), .A2(n_770), .B1(n_1990), .B2(n_1991), .Y(n_1989) );
BUFx3_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
BUFx3_ASAP7_75t_L g830 ( .A(n_769), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_770), .A2(n_820), .B1(n_830), .B2(n_831), .Y(n_829) );
AOI222xp33_ASAP7_75t_L g1596 ( .A1(n_770), .A2(n_830), .B1(n_1597), .B2(n_1598), .C1(n_1599), .C2(n_1600), .Y(n_1596) );
AOI22xp33_ASAP7_75t_L g1664 ( .A1(n_770), .A2(n_830), .B1(n_1665), .B2(n_1666), .Y(n_1664) );
AOI22xp33_ASAP7_75t_L g1932 ( .A1(n_770), .A2(n_830), .B1(n_1933), .B2(n_1934), .Y(n_1932) );
INVx1_ASAP7_75t_L g775 ( .A(n_776), .Y(n_775) );
OAI31xp33_ASAP7_75t_L g824 ( .A1(n_777), .A2(n_825), .A3(n_827), .B(n_832), .Y(n_824) );
OAI31xp33_ASAP7_75t_SL g1064 ( .A1(n_777), .A2(n_1065), .A3(n_1068), .B(n_1072), .Y(n_1064) );
OAI31xp33_ASAP7_75t_L g1929 ( .A1(n_777), .A2(n_1930), .A3(n_1931), .B(n_1935), .Y(n_1929) );
AND3x1_ASAP7_75t_L g779 ( .A(n_780), .B(n_816), .C(n_824), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g780 ( .A(n_781), .B(n_804), .Y(n_780) );
OAI33xp33_ASAP7_75t_L g890 ( .A1(n_782), .A2(n_891), .A3(n_896), .B1(n_902), .B2(n_903), .B3(n_905), .Y(n_890) );
OAI22xp33_ASAP7_75t_L g805 ( .A1(n_784), .A2(n_801), .B1(n_806), .B2(n_808), .Y(n_805) );
HB1xp67_ASAP7_75t_L g786 ( .A(n_787), .Y(n_786) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_787), .Y(n_803) );
BUFx6f_ASAP7_75t_L g1028 ( .A(n_787), .Y(n_1028) );
INVx2_ASAP7_75t_L g1139 ( .A(n_787), .Y(n_1139) );
OAI22xp5_ASAP7_75t_L g1653 ( .A1(n_790), .A2(n_799), .B1(n_1654), .B2(n_1655), .Y(n_1653) );
BUFx3_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_791), .A2(n_878), .B1(n_888), .B2(n_899), .Y(n_902) );
INVx8_ASAP7_75t_L g1157 ( .A(n_791), .Y(n_1157) );
OAI22xp5_ASAP7_75t_L g793 ( .A1(n_794), .A2(n_795), .B1(n_798), .B2(n_799), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g1037 ( .A(n_796), .Y(n_1037) );
INVx1_ASAP7_75t_L g796 ( .A(n_797), .Y(n_796) );
BUFx2_ASAP7_75t_L g946 ( .A(n_797), .Y(n_946) );
INVx3_ASAP7_75t_L g1423 ( .A(n_797), .Y(n_1423) );
OAI22xp5_ASAP7_75t_L g1154 ( .A1(n_799), .A2(n_1155), .B1(n_1156), .B2(n_1158), .Y(n_1154) );
OAI22xp5_ASAP7_75t_L g1966 ( .A1(n_799), .A2(n_1156), .B1(n_1967), .B2(n_1968), .Y(n_1966) );
INVx2_ASAP7_75t_L g806 ( .A(n_807), .Y(n_806) );
INVx2_ASAP7_75t_L g815 ( .A(n_807), .Y(n_815) );
INVx3_ASAP7_75t_L g979 ( .A(n_807), .Y(n_979) );
INVx2_ASAP7_75t_SL g1050 ( .A(n_807), .Y(n_1050) );
OAI22xp33_ASAP7_75t_L g1657 ( .A1(n_808), .A2(n_885), .B1(n_1648), .B2(n_1651), .Y(n_1657) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx4_ASAP7_75t_L g880 ( .A(n_812), .Y(n_880) );
INVx2_ASAP7_75t_L g975 ( .A(n_812), .Y(n_975) );
INVx2_ASAP7_75t_L g1055 ( .A(n_812), .Y(n_1055) );
INVx4_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
OAI31xp33_ASAP7_75t_L g816 ( .A1(n_817), .A2(n_818), .A3(n_822), .B(n_823), .Y(n_816) );
OAI31xp33_ASAP7_75t_L g852 ( .A1(n_823), .A2(n_853), .A3(n_858), .B(n_861), .Y(n_852) );
OAI31xp33_ASAP7_75t_L g1075 ( .A1(n_823), .A2(n_1076), .A3(n_1078), .B(n_1084), .Y(n_1075) );
OAI31xp33_ASAP7_75t_L g1182 ( .A1(n_823), .A2(n_1183), .A3(n_1184), .B(n_1185), .Y(n_1182) );
OAI31xp33_ASAP7_75t_SL g1993 ( .A1(n_823), .A2(n_1994), .A3(n_1995), .B(n_1996), .Y(n_1993) );
NAND4xp25_ASAP7_75t_L g1592 ( .A(n_828), .B(n_1593), .C(n_1596), .D(n_1601), .Y(n_1592) );
INVx1_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
XOR2xp5_ASAP7_75t_L g836 ( .A(n_837), .B(n_960), .Y(n_836) );
OAI22xp5_ASAP7_75t_L g837 ( .A1(n_838), .A2(n_906), .B1(n_958), .B2(n_959), .Y(n_837) );
INVx1_ASAP7_75t_L g958 ( .A(n_838), .Y(n_958) );
NAND3xp33_ASAP7_75t_L g839 ( .A(n_840), .B(n_852), .C(n_862), .Y(n_839) );
INVx2_ASAP7_75t_SL g842 ( .A(n_843), .Y(n_842) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_847), .Y(n_846) );
OAI211xp5_ASAP7_75t_L g1321 ( .A1(n_847), .A2(n_1272), .B(n_1322), .C(n_1324), .Y(n_1321) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_854), .A2(n_874), .B1(n_875), .B2(n_878), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g973 ( .A1(n_854), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
OAI22xp5_ASAP7_75t_L g1115 ( .A1(n_854), .A2(n_1102), .B1(n_1106), .B2(n_1116), .Y(n_1115) );
INVx1_ASAP7_75t_L g1187 ( .A(n_854), .Y(n_1187) );
OAI22xp5_ASAP7_75t_L g1496 ( .A1(n_854), .A2(n_975), .B1(n_1497), .B2(n_1498), .Y(n_1496) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_863), .B(n_890), .Y(n_862) );
OAI33xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_867), .A3(n_873), .B1(n_879), .B2(n_884), .B3(n_889), .Y(n_863) );
OAI33xp33_ASAP7_75t_L g964 ( .A1(n_864), .A2(n_889), .A3(n_965), .B1(n_970), .B2(n_973), .B3(n_977), .Y(n_964) );
INVx1_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx2_ASAP7_75t_SL g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_SL g937 ( .A(n_866), .Y(n_937) );
OAI22xp33_ASAP7_75t_L g867 ( .A1(n_868), .A2(n_869), .B1(n_871), .B2(n_872), .Y(n_867) );
OAI22xp33_ASAP7_75t_L g891 ( .A1(n_868), .A2(n_881), .B1(n_892), .B2(n_895), .Y(n_891) );
BUFx3_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
BUFx6f_ASAP7_75t_L g1118 ( .A(n_870), .Y(n_1118) );
INVx2_ASAP7_75t_SL g1211 ( .A(n_870), .Y(n_1211) );
BUFx3_ASAP7_75t_L g1266 ( .A(n_870), .Y(n_1266) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_872), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_977) );
OAI22xp33_ASAP7_75t_L g1218 ( .A1(n_872), .A2(n_1201), .B1(n_1204), .B2(n_1210), .Y(n_1218) );
OAI22xp5_ASAP7_75t_L g896 ( .A1(n_874), .A2(n_886), .B1(n_897), .B2(n_899), .Y(n_896) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_875), .A2(n_1027), .B1(n_1046), .B2(n_1051), .Y(n_1057) );
INVx3_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
OAI22xp5_ASAP7_75t_L g1170 ( .A1(n_877), .A2(n_1056), .B1(n_1155), .B2(n_1160), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1981 ( .A(n_877), .Y(n_1981) );
OAI22xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_881), .B1(n_882), .B2(n_883), .Y(n_879) );
OAI221xp5_ASAP7_75t_L g1271 ( .A1(n_882), .A2(n_1213), .B1(n_1272), .B2(n_1273), .C(n_1274), .Y(n_1271) );
OAI211xp5_ASAP7_75t_SL g1398 ( .A1(n_882), .A2(n_1399), .B(n_1400), .C(n_1402), .Y(n_1398) );
OAI211xp5_ASAP7_75t_SL g1403 ( .A1(n_882), .A2(n_1404), .B(n_1405), .C(n_1407), .Y(n_1403) );
OAI22xp5_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_886), .B1(n_887), .B2(n_888), .Y(n_884) );
OAI22xp33_ASAP7_75t_L g965 ( .A1(n_885), .A2(n_966), .B1(n_967), .B2(n_968), .Y(n_965) );
OAI22xp5_ASAP7_75t_L g1120 ( .A1(n_885), .A2(n_1103), .B1(n_1108), .B2(n_1121), .Y(n_1120) );
OAI22xp33_ASAP7_75t_L g1172 ( .A1(n_887), .A2(n_1059), .B1(n_1158), .B2(n_1162), .Y(n_1172) );
OAI22xp33_ASAP7_75t_L g1209 ( .A1(n_887), .A2(n_1195), .B1(n_1206), .B2(n_1210), .Y(n_1209) );
OAI22xp5_ASAP7_75t_L g1502 ( .A1(n_887), .A2(n_1210), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
OAI21xp5_ASAP7_75t_L g1270 ( .A1(n_889), .A2(n_1271), .B(n_1276), .Y(n_1270) );
OAI22xp33_ASAP7_75t_L g1151 ( .A1(n_892), .A2(n_1028), .B1(n_1152), .B2(n_1153), .Y(n_1151) );
OAI22xp33_ASAP7_75t_L g1163 ( .A1(n_892), .A2(n_1164), .B1(n_1165), .B2(n_1166), .Y(n_1163) );
OAI22xp33_ASAP7_75t_L g1205 ( .A1(n_892), .A2(n_1176), .B1(n_1206), .B2(n_1207), .Y(n_1205) );
OAI22xp33_ASAP7_75t_L g1963 ( .A1(n_892), .A2(n_1028), .B1(n_1964), .B2(n_1965), .Y(n_1963) );
OAI22xp33_ASAP7_75t_L g1972 ( .A1(n_892), .A2(n_1028), .B1(n_1973), .B2(n_1974), .Y(n_1972) );
INVx2_ASAP7_75t_L g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
INVx1_ASAP7_75t_L g1197 ( .A(n_894), .Y(n_1197) );
INVx2_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
INVx2_ASAP7_75t_SL g1417 ( .A(n_898), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1509 ( .A1(n_899), .A2(n_1498), .B1(n_1504), .B2(n_1510), .Y(n_1509) );
OAI221xp5_ASAP7_75t_L g1577 ( .A1(n_899), .A2(n_992), .B1(n_1578), .B2(n_1579), .C(n_1580), .Y(n_1577) );
OAI22xp33_ASAP7_75t_SL g1643 ( .A1(n_899), .A2(n_1644), .B1(n_1645), .B2(n_1646), .Y(n_1643) );
INVx3_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
BUFx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g1035 ( .A(n_901), .Y(n_1035) );
INVx1_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx2_ASAP7_75t_L g959 ( .A(n_906), .Y(n_959) );
INVx1_ASAP7_75t_L g956 ( .A(n_907), .Y(n_956) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_908), .B(n_923), .C(n_931), .Y(n_907) );
OAI21xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_919), .B(n_922), .Y(n_908) );
INVx2_ASAP7_75t_L g1943 ( .A(n_912), .Y(n_1943) );
INVx2_ASAP7_75t_L g912 ( .A(n_913), .Y(n_912) );
OAI31xp33_ASAP7_75t_SL g1003 ( .A1(n_922), .A2(n_1004), .A3(n_1008), .B(n_1014), .Y(n_1003) );
OAI31xp33_ASAP7_75t_L g1125 ( .A1(n_922), .A2(n_1126), .A3(n_1127), .B(n_1132), .Y(n_1125) );
AND4x1_ASAP7_75t_L g931 ( .A(n_932), .B(n_938), .C(n_943), .D(n_949), .Y(n_931) );
NAND3xp33_ASAP7_75t_L g932 ( .A(n_933), .B(n_936), .C(n_937), .Y(n_932) );
HB1xp67_ASAP7_75t_L g940 ( .A(n_941), .Y(n_940) );
INVx2_ASAP7_75t_L g1261 ( .A(n_941), .Y(n_1261) );
INVx2_ASAP7_75t_L g945 ( .A(n_946), .Y(n_945) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_946), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1101) );
OAI221xp5_ASAP7_75t_L g1609 ( .A1(n_946), .A2(n_986), .B1(n_1610), .B2(n_1611), .C(n_1612), .Y(n_1609) );
INVx1_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_961), .A2(n_1016), .B1(n_1017), .B2(n_1089), .Y(n_960) );
INVx2_ASAP7_75t_SL g1089 ( .A(n_961), .Y(n_1089) );
NAND3xp33_ASAP7_75t_L g962 ( .A(n_963), .B(n_993), .C(n_1003), .Y(n_962) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_964), .B(n_981), .Y(n_963) );
OAI22xp5_ASAP7_75t_L g1264 ( .A1(n_968), .A2(n_1265), .B1(n_1266), .B2(n_1267), .Y(n_1264) );
BUFx6f_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
OAI22xp5_ASAP7_75t_L g984 ( .A1(n_971), .A2(n_978), .B1(n_985), .B2(n_986), .Y(n_984) );
HB1xp67_ASAP7_75t_L g1231 ( .A(n_983), .Y(n_1231) );
OAI22xp5_ASAP7_75t_L g1105 ( .A1(n_986), .A2(n_1106), .B1(n_1107), .B2(n_1108), .Y(n_1105) );
OAI22xp5_ASAP7_75t_L g1926 ( .A1(n_986), .A2(n_1906), .B1(n_1917), .B2(n_1927), .Y(n_1926) );
INVx1_ASAP7_75t_L g988 ( .A(n_989), .Y(n_988) );
INVx1_ASAP7_75t_L g1100 ( .A(n_989), .Y(n_1100) );
INVxp67_ASAP7_75t_L g1988 ( .A(n_989), .Y(n_1988) );
INVx1_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1113 ( .A(n_990), .Y(n_1113) );
OAI31xp33_ASAP7_75t_L g993 ( .A1(n_994), .A2(n_997), .A3(n_1001), .B(n_1002), .Y(n_993) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
OAI31xp33_ASAP7_75t_SL g1133 ( .A1(n_1002), .A2(n_1134), .A3(n_1135), .B(n_1137), .Y(n_1133) );
INVx1_ASAP7_75t_L g1005 ( .A(n_1006), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
INVx2_ASAP7_75t_L g1010 ( .A(n_1011), .Y(n_1010) );
INVx2_ASAP7_75t_L g1128 ( .A(n_1011), .Y(n_1128) );
INVx2_ASAP7_75t_SL g1016 ( .A(n_1017), .Y(n_1016) );
NAND3xp33_ASAP7_75t_L g1018 ( .A(n_1019), .B(n_1064), .C(n_1075), .Y(n_1018) );
NOR2xp33_ASAP7_75t_SL g1019 ( .A(n_1020), .B(n_1047), .Y(n_1019) );
OAI33xp33_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1023), .A3(n_1029), .B1(n_1036), .B2(n_1042), .B3(n_1043), .Y(n_1020) );
OAI22xp33_ASAP7_75t_L g1415 ( .A1(n_1021), .A2(n_1416), .B1(n_1421), .B2(n_1426), .Y(n_1415) );
OAI22xp5_ASAP7_75t_L g1604 ( .A1(n_1021), .A2(n_1042), .B1(n_1605), .B2(n_1609), .Y(n_1604) );
OAI33xp33_ASAP7_75t_L g1918 ( .A1(n_1021), .A2(n_1919), .A3(n_1920), .B1(n_1923), .B2(n_1924), .B3(n_1926), .Y(n_1918) );
BUFx3_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
OAI22xp33_ASAP7_75t_L g1023 ( .A1(n_1024), .A2(n_1025), .B1(n_1027), .B2(n_1028), .Y(n_1023) );
OAI22xp5_ASAP7_75t_L g1049 ( .A1(n_1024), .A2(n_1045), .B1(n_1050), .B2(n_1051), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g1025 ( .A(n_1026), .Y(n_1025) );
HB1xp67_ASAP7_75t_L g1044 ( .A(n_1026), .Y(n_1044) );
INVx1_ASAP7_75t_L g1928 ( .A(n_1026), .Y(n_1928) );
OAI22xp5_ASAP7_75t_L g1923 ( .A1(n_1028), .A2(n_1510), .B1(n_1902), .B2(n_1911), .Y(n_1923) );
OAI22xp33_ASAP7_75t_SL g1029 ( .A1(n_1030), .A2(n_1031), .B1(n_1034), .B2(n_1035), .Y(n_1029) );
OAI22xp5_ASAP7_75t_L g1054 ( .A1(n_1030), .A2(n_1038), .B1(n_1055), .B2(n_1056), .Y(n_1054) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_1032), .A2(n_1285), .B1(n_1288), .B2(n_1305), .Y(n_1304) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
OAI22xp33_ASAP7_75t_L g1058 ( .A1(n_1034), .A2(n_1041), .B1(n_1059), .B2(n_1063), .Y(n_1058) );
OAI22xp5_ASAP7_75t_L g1036 ( .A1(n_1037), .A2(n_1038), .B1(n_1039), .B2(n_1041), .Y(n_1036) );
OAI22xp33_ASAP7_75t_L g1919 ( .A1(n_1039), .A2(n_1044), .B1(n_1905), .B2(n_1916), .Y(n_1919) );
INVx2_ASAP7_75t_SL g1039 ( .A(n_1040), .Y(n_1039) );
OAI33xp33_ASAP7_75t_L g1114 ( .A1(n_1048), .A2(n_1115), .A3(n_1117), .B1(n_1120), .B2(n_1122), .B3(n_1124), .Y(n_1114) );
OAI33xp33_ASAP7_75t_L g1899 ( .A1(n_1048), .A2(n_1900), .A3(n_1904), .B1(n_1909), .B2(n_1912), .B3(n_1915), .Y(n_1899) );
INVx1_ASAP7_75t_L g1051 ( .A(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
OAI22xp33_ASAP7_75t_L g1491 ( .A1(n_1053), .A2(n_1492), .B1(n_1493), .B2(n_1495), .Y(n_1491) );
OAI22xp5_ASAP7_75t_L g1982 ( .A1(n_1059), .A2(n_1968), .B1(n_1971), .B2(n_1983), .Y(n_1982) );
INVx1_ASAP7_75t_L g1059 ( .A(n_1060), .Y(n_1059) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1136 ( .A(n_1067), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1085 ( .A1(n_1070), .A2(n_1086), .B1(n_1087), .B2(n_1088), .Y(n_1085) );
INVx1_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_SL g1082 ( .A(n_1083), .Y(n_1082) );
AOI22xp33_ASAP7_75t_L g1945 ( .A1(n_1086), .A2(n_1526), .B1(n_1933), .B2(n_1946), .Y(n_1945) );
INVx1_ASAP7_75t_L g1142 ( .A(n_1090), .Y(n_1142) );
HB1xp67_ASAP7_75t_L g1090 ( .A(n_1091), .Y(n_1090) );
XNOR2xp5_ASAP7_75t_L g1091 ( .A(n_1092), .B(n_1093), .Y(n_1091) );
AND3x1_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1125), .C(n_1133), .Y(n_1093) );
NOR2xp33_ASAP7_75t_SL g1094 ( .A(n_1095), .B(n_1114), .Y(n_1094) );
OAI22xp33_ASAP7_75t_L g1117 ( .A1(n_1098), .A2(n_1110), .B1(n_1118), .B2(n_1119), .Y(n_1117) );
INVxp67_ASAP7_75t_SL g1112 ( .A(n_1113), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g1176 ( .A(n_1113), .Y(n_1176) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1113), .Y(n_1507) );
OAI22xp5_ASAP7_75t_L g1900 ( .A1(n_1116), .A2(n_1901), .B1(n_1902), .B2(n_1903), .Y(n_1900) );
OAI22xp5_ASAP7_75t_L g1915 ( .A1(n_1116), .A2(n_1907), .B1(n_1916), .B2(n_1917), .Y(n_1915) );
OAI22xp5_ASAP7_75t_L g1379 ( .A1(n_1119), .A2(n_1380), .B1(n_1381), .B2(n_1382), .Y(n_1379) );
INVx2_ASAP7_75t_L g1908 ( .A(n_1119), .Y(n_1908) );
INVx2_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
INVx1_ASAP7_75t_L g1138 ( .A(n_1139), .Y(n_1138) );
INVx2_ASAP7_75t_L g1165 ( .A(n_1139), .Y(n_1165) );
INVx1_ASAP7_75t_L g1143 ( .A(n_1144), .Y(n_1143) );
AOI22xp5_ASAP7_75t_L g1144 ( .A1(n_1145), .A2(n_1146), .B1(n_1190), .B2(n_1235), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1146), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_1147), .Y(n_1146) );
AND3x1_ASAP7_75t_L g1148 ( .A(n_1149), .B(n_1173), .C(n_1182), .Y(n_1148) );
NOR2xp33_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1167), .Y(n_1149) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
INVx1_ASAP7_75t_L g1645 ( .A(n_1157), .Y(n_1645) );
OAI22xp33_ASAP7_75t_L g1194 ( .A1(n_1165), .A2(n_1195), .B1(n_1196), .B2(n_1198), .Y(n_1194) );
HB1xp67_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1235 ( .A(n_1190), .Y(n_1235) );
NAND3xp33_ASAP7_75t_L g1191 ( .A(n_1192), .B(n_1219), .C(n_1228), .Y(n_1191) );
NOR2xp33_ASAP7_75t_L g1192 ( .A(n_1193), .B(n_1208), .Y(n_1192) );
OAI22xp33_ASAP7_75t_L g1506 ( .A1(n_1196), .A2(n_1492), .B1(n_1500), .B2(n_1507), .Y(n_1506) );
OAI22xp33_ASAP7_75t_L g1511 ( .A1(n_1196), .A2(n_1495), .B1(n_1501), .B2(n_1512), .Y(n_1511) );
INVx2_ASAP7_75t_L g1196 ( .A(n_1197), .Y(n_1196) );
OAI22xp5_ASAP7_75t_SL g1212 ( .A1(n_1200), .A2(n_1203), .B1(n_1213), .B2(n_1215), .Y(n_1212) );
OAI22xp5_ASAP7_75t_L g1904 ( .A1(n_1210), .A2(n_1905), .B1(n_1906), .B2(n_1907), .Y(n_1904) );
OAI22xp33_ASAP7_75t_L g1909 ( .A1(n_1210), .A2(n_1215), .B1(n_1910), .B2(n_1911), .Y(n_1909) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
INVx2_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
HB1xp67_ASAP7_75t_L g1903 ( .A(n_1215), .Y(n_1903) );
INVx1_ASAP7_75t_L g1222 ( .A(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1237 ( .A(n_1238), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1239), .Y(n_1238) );
XNOR2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1484), .Y(n_1239) );
INVx3_ASAP7_75t_SL g1240 ( .A(n_1241), .Y(n_1240) );
BUFx3_ASAP7_75t_L g1241 ( .A(n_1242), .Y(n_1241) );
OA22x2_ASAP7_75t_L g1242 ( .A1(n_1243), .A2(n_1244), .B1(n_1388), .B2(n_1483), .Y(n_1242) );
INVx1_ASAP7_75t_L g1243 ( .A(n_1244), .Y(n_1243) );
XOR2xp5_ASAP7_75t_L g1244 ( .A(n_1245), .B(n_1327), .Y(n_1244) );
XNOR2x1_ASAP7_75t_L g1245 ( .A(n_1246), .B(n_1247), .Y(n_1245) );
NAND4xp75_ASAP7_75t_L g1247 ( .A(n_1248), .B(n_1258), .C(n_1284), .D(n_1291), .Y(n_1247) );
INVx1_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
INVx1_ASAP7_75t_L g1251 ( .A(n_1252), .Y(n_1251) );
AND2x4_ASAP7_75t_L g1252 ( .A(n_1253), .B(n_1255), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
INVx3_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1256), .Y(n_1408) );
AOI211x1_ASAP7_75t_L g1258 ( .A1(n_1259), .A2(n_1268), .B(n_1270), .C(n_1280), .Y(n_1258) );
INVx2_ASAP7_75t_L g1260 ( .A(n_1261), .Y(n_1260) );
BUFx2_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
AOI221xp5_ASAP7_75t_L g1366 ( .A1(n_1263), .A2(n_1348), .B1(n_1354), .B2(n_1367), .C(n_1369), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g1470 ( .A1(n_1263), .A2(n_1367), .B1(n_1447), .B2(n_1458), .C(n_1471), .Y(n_1470) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NAND2x2_ASAP7_75t_L g1281 ( .A(n_1278), .B(n_1282), .Y(n_1281) );
INVx2_ASAP7_75t_L g1278 ( .A(n_1279), .Y(n_1278) );
INVx2_ASAP7_75t_SL g1282 ( .A(n_1283), .Y(n_1282) );
AOI22xp5_ASAP7_75t_L g1284 ( .A1(n_1285), .A2(n_1286), .B1(n_1288), .B2(n_1289), .Y(n_1284) );
INVx3_ASAP7_75t_L g1540 ( .A(n_1286), .Y(n_1540) );
AND2x4_ASAP7_75t_L g1289 ( .A(n_1287), .B(n_1290), .Y(n_1289) );
INVx2_ASAP7_75t_L g1545 ( .A(n_1289), .Y(n_1545) );
OAI31xp67_ASAP7_75t_L g1291 ( .A1(n_1292), .A2(n_1303), .A3(n_1314), .B(n_1325), .Y(n_1291) );
INVx4_ASAP7_75t_L g1293 ( .A(n_1294), .Y(n_1293) );
INVx2_ASAP7_75t_L g1295 ( .A(n_1296), .Y(n_1295) );
A2O1A1Ixp33_ASAP7_75t_L g1297 ( .A1(n_1298), .A2(n_1299), .B(n_1300), .C(n_1301), .Y(n_1297) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
AOI21xp33_ASAP7_75t_L g1303 ( .A1(n_1304), .A2(n_1306), .B(n_1311), .Y(n_1303) );
AOI22xp33_ASAP7_75t_L g1306 ( .A1(n_1307), .A2(n_1308), .B1(n_1309), .B2(n_1310), .Y(n_1306) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
HB1xp67_ASAP7_75t_L g1312 ( .A(n_1313), .Y(n_1312) );
OAI21xp5_ASAP7_75t_SL g1314 ( .A1(n_1315), .A2(n_1318), .B(n_1321), .Y(n_1314) );
AOI31xp33_ASAP7_75t_L g1553 ( .A1(n_1325), .A2(n_1554), .A3(n_1567), .B(n_1572), .Y(n_1553) );
BUFx2_ASAP7_75t_L g1325 ( .A(n_1326), .Y(n_1325) );
XNOR2x1_ASAP7_75t_L g1327 ( .A(n_1328), .B(n_1387), .Y(n_1327) );
OR2x2_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1349), .Y(n_1328) );
NAND3xp33_ASAP7_75t_L g1329 ( .A(n_1330), .B(n_1338), .C(n_1347), .Y(n_1329) );
AOI222xp33_ASAP7_75t_L g1330 ( .A1(n_1331), .A2(n_1332), .B1(n_1333), .B2(n_1335), .C1(n_1336), .C2(n_1337), .Y(n_1330) );
AOI222xp33_ASAP7_75t_L g1448 ( .A1(n_1331), .A2(n_1333), .B1(n_1336), .B2(n_1449), .C1(n_1450), .C2(n_1451), .Y(n_1448) );
AOI22xp5_ASAP7_75t_L g1550 ( .A1(n_1331), .A2(n_1336), .B1(n_1551), .B2(n_1552), .Y(n_1550) );
INVx2_ASAP7_75t_L g1342 ( .A(n_1343), .Y(n_1342) );
NAND3xp33_ASAP7_75t_SL g1349 ( .A(n_1350), .B(n_1355), .C(n_1383), .Y(n_1349) );
INVx1_ASAP7_75t_L g1548 ( .A(n_1351), .Y(n_1548) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1353), .Y(n_1549) );
INVx1_ASAP7_75t_L g1357 ( .A(n_1358), .Y(n_1357) );
OAI21xp33_ASAP7_75t_L g1363 ( .A1(n_1364), .A2(n_1366), .B(n_1370), .Y(n_1363) );
OAI21xp5_ASAP7_75t_SL g1469 ( .A1(n_1364), .A2(n_1470), .B(n_1473), .Y(n_1469) );
INVxp67_ASAP7_75t_L g1364 ( .A(n_1365), .Y(n_1364) );
OAI21xp5_ASAP7_75t_L g1395 ( .A1(n_1365), .A2(n_1396), .B(n_1397), .Y(n_1395) );
INVx2_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1373), .Y(n_1414) );
AOI22xp5_ASAP7_75t_L g1475 ( .A1(n_1373), .A2(n_1449), .B1(n_1457), .B2(n_1476), .Y(n_1475) );
INVx1_ASAP7_75t_L g1373 ( .A(n_1374), .Y(n_1373) );
INVx1_ASAP7_75t_L g1566 ( .A(n_1375), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1384), .B(n_1385), .Y(n_1383) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1385), .B(n_1460), .Y(n_1459) );
INVx5_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
INVx3_ASAP7_75t_L g1536 ( .A(n_1386), .Y(n_1536) );
XNOR2xp5_ASAP7_75t_L g1388 ( .A(n_1389), .B(n_1440), .Y(n_1388) );
XOR2xp5_ASAP7_75t_L g1483 ( .A(n_1389), .B(n_1440), .Y(n_1483) );
XNOR2x1_ASAP7_75t_L g1389 ( .A(n_1390), .B(n_1391), .Y(n_1389) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1427), .Y(n_1391) );
AOI21xp5_ASAP7_75t_L g1392 ( .A1(n_1393), .A2(n_1394), .B(n_1415), .Y(n_1392) );
NAND4xp25_ASAP7_75t_L g1394 ( .A(n_1395), .B(n_1398), .C(n_1403), .D(n_1409), .Y(n_1394) );
INVx1_ASAP7_75t_L g1412 ( .A(n_1413), .Y(n_1412) );
INVx2_ASAP7_75t_L g1422 ( .A(n_1423), .Y(n_1422) );
XNOR2x1_ASAP7_75t_L g1440 ( .A(n_1441), .B(n_1482), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1455), .Y(n_1441) );
NAND4xp25_ASAP7_75t_SL g1442 ( .A(n_1443), .B(n_1446), .C(n_1448), .D(n_1452), .Y(n_1442) );
NAND3xp33_ASAP7_75t_SL g1455 ( .A(n_1456), .B(n_1459), .C(n_1461), .Y(n_1455) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1979 ( .A(n_1468), .Y(n_1979) );
AO22x2_ASAP7_75t_L g1484 ( .A1(n_1485), .A2(n_1486), .B1(n_1636), .B2(n_1637), .Y(n_1484) );
INVx1_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
AO22x2_ASAP7_75t_L g1486 ( .A1(n_1487), .A2(n_1530), .B1(n_1531), .B2(n_1635), .Y(n_1486) );
INVx1_ASAP7_75t_L g1635 ( .A(n_1487), .Y(n_1635) );
NAND3xp33_ASAP7_75t_L g1488 ( .A(n_1489), .B(n_1513), .C(n_1521), .Y(n_1488) );
NOR2xp33_ASAP7_75t_L g1489 ( .A(n_1490), .B(n_1505), .Y(n_1489) );
INVx1_ASAP7_75t_L g1493 ( .A(n_1494), .Y(n_1493) );
OAI31xp33_ASAP7_75t_L g1513 ( .A1(n_1514), .A2(n_1515), .A3(n_1519), .B(n_1520), .Y(n_1513) );
OAI31xp33_ASAP7_75t_L g1661 ( .A1(n_1520), .A2(n_1662), .A3(n_1663), .B(n_1667), .Y(n_1661) );
OAI31xp33_ASAP7_75t_L g1985 ( .A1(n_1520), .A2(n_1986), .A3(n_1987), .B(n_1992), .Y(n_1985) );
INVx2_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
INVx2_ASAP7_75t_L g1530 ( .A(n_1531), .Y(n_1530) );
XOR2x2_ASAP7_75t_L g1531 ( .A(n_1532), .B(n_1589), .Y(n_1531) );
INVx1_ASAP7_75t_L g1587 ( .A(n_1533), .Y(n_1587) );
NAND3xp33_ASAP7_75t_L g1533 ( .A(n_1534), .B(n_1537), .C(n_1546), .Y(n_1533) );
NAND2xp5_ASAP7_75t_L g1534 ( .A(n_1535), .B(n_1536), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_1535), .A2(n_1573), .B1(n_1574), .B2(n_1575), .Y(n_1572) );
AOI22xp33_ASAP7_75t_L g1537 ( .A1(n_1538), .A2(n_1539), .B1(n_1541), .B2(n_1542), .Y(n_1537) );
NAND2x1_ASAP7_75t_L g1542 ( .A(n_1543), .B(n_1545), .Y(n_1542) );
INVx2_ASAP7_75t_SL g1543 ( .A(n_1544), .Y(n_1543) );
NOR3xp33_ASAP7_75t_SL g1546 ( .A(n_1547), .B(n_1553), .C(n_1576), .Y(n_1546) );
NAND2xp5_ASAP7_75t_L g1562 ( .A(n_1551), .B(n_1563), .Y(n_1562) );
AOI21xp5_ASAP7_75t_L g1554 ( .A1(n_1555), .A2(n_1559), .B(n_1561), .Y(n_1554) );
INVx2_ASAP7_75t_SL g1556 ( .A(n_1557), .Y(n_1556) );
AOI21xp5_ASAP7_75t_L g1561 ( .A1(n_1562), .A2(n_1564), .B(n_1566), .Y(n_1561) );
INVx2_ASAP7_75t_L g1619 ( .A(n_1573), .Y(n_1619) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1590 ( .A(n_1591), .Y(n_1590) );
NAND2xp5_ASAP7_75t_L g1632 ( .A(n_1599), .B(n_1633), .Y(n_1632) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1600), .Y(n_1614) );
INVx1_ASAP7_75t_L g1613 ( .A(n_1614), .Y(n_1613) );
NOR2xp33_ASAP7_75t_L g1616 ( .A(n_1617), .B(n_1620), .Y(n_1616) );
INVx1_ASAP7_75t_L g1636 ( .A(n_1637), .Y(n_1636) );
INVx1_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
INVx1_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
NAND3xp33_ASAP7_75t_L g1640 ( .A(n_1641), .B(n_1661), .C(n_1668), .Y(n_1640) );
NOR2xp33_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1656), .Y(n_1641) );
OAI221xp5_ASAP7_75t_L g1674 ( .A1(n_1675), .A2(n_1893), .B1(n_1896), .B2(n_1947), .C(n_1953), .Y(n_1674) );
AOI21xp5_ASAP7_75t_L g1675 ( .A1(n_1676), .A2(n_1817), .B(n_1865), .Y(n_1675) );
NAND5xp2_ASAP7_75t_L g1676 ( .A(n_1677), .B(n_1739), .C(n_1780), .D(n_1795), .E(n_1810), .Y(n_1676) );
AOI211xp5_ASAP7_75t_SL g1677 ( .A1(n_1678), .A2(n_1703), .B(n_1721), .C(n_1732), .Y(n_1677) );
AND2x2_ASAP7_75t_L g1678 ( .A(n_1679), .B(n_1694), .Y(n_1678) );
OR2x2_ASAP7_75t_L g1802 ( .A(n_1679), .B(n_1704), .Y(n_1802) );
A2O1A1Ixp33_ASAP7_75t_SL g1810 ( .A1(n_1679), .A2(n_1794), .B(n_1811), .C(n_1814), .Y(n_1810) );
INVx2_ASAP7_75t_L g1815 ( .A(n_1679), .Y(n_1815) );
NAND2xp5_ASAP7_75t_SL g1821 ( .A(n_1679), .B(n_1753), .Y(n_1821) );
NAND2xp5_ASAP7_75t_L g1837 ( .A(n_1679), .B(n_1838), .Y(n_1837) );
INVx2_ASAP7_75t_L g1679 ( .A(n_1680), .Y(n_1679) );
INVx3_ASAP7_75t_L g1731 ( .A(n_1680), .Y(n_1731) );
NOR2xp33_ASAP7_75t_L g1755 ( .A(n_1680), .B(n_1707), .Y(n_1755) );
NOR2xp33_ASAP7_75t_L g1759 ( .A(n_1680), .B(n_1760), .Y(n_1759) );
AND2x2_ASAP7_75t_L g1763 ( .A(n_1680), .B(n_1707), .Y(n_1763) );
NAND2xp5_ASAP7_75t_L g1831 ( .A(n_1680), .B(n_1782), .Y(n_1831) );
AND2x2_ASAP7_75t_L g1858 ( .A(n_1680), .B(n_1722), .Y(n_1858) );
AND2x2_ASAP7_75t_L g1680 ( .A(n_1681), .B(n_1689), .Y(n_1680) );
AND2x4_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1684), .Y(n_1682) );
AND2x6_ASAP7_75t_L g1687 ( .A(n_1683), .B(n_1688), .Y(n_1687) );
AND2x6_ASAP7_75t_L g1690 ( .A(n_1683), .B(n_1691), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1683), .B(n_1693), .Y(n_1692) );
AND2x2_ASAP7_75t_L g1701 ( .A(n_1683), .B(n_1693), .Y(n_1701) );
AND2x2_ASAP7_75t_L g1709 ( .A(n_1683), .B(n_1693), .Y(n_1709) );
AND2x2_ASAP7_75t_L g1684 ( .A(n_1685), .B(n_1686), .Y(n_1684) );
INVx2_ASAP7_75t_L g1895 ( .A(n_1690), .Y(n_1895) );
OAI21xp5_ASAP7_75t_L g2000 ( .A1(n_1691), .A2(n_2001), .B(n_2002), .Y(n_2000) );
INVx1_ASAP7_75t_L g1694 ( .A(n_1695), .Y(n_1694) );
OR2x2_ASAP7_75t_L g1741 ( .A(n_1695), .B(n_1722), .Y(n_1741) );
AOI21xp33_ASAP7_75t_L g1867 ( .A1(n_1695), .A2(n_1802), .B(n_1805), .Y(n_1867) );
OR2x2_ASAP7_75t_L g1695 ( .A(n_1696), .B(n_1699), .Y(n_1695) );
INVx1_ASAP7_75t_L g1730 ( .A(n_1696), .Y(n_1730) );
INVx1_ASAP7_75t_L g1765 ( .A(n_1696), .Y(n_1765) );
INVx1_ASAP7_75t_L g1782 ( .A(n_1696), .Y(n_1782) );
AND2x2_ASAP7_75t_L g1826 ( .A(n_1696), .B(n_1699), .Y(n_1826) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1698), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1738 ( .A(n_1699), .B(n_1730), .Y(n_1738) );
NAND2xp5_ASAP7_75t_L g1772 ( .A(n_1699), .B(n_1723), .Y(n_1772) );
AND2x2_ASAP7_75t_L g1794 ( .A(n_1699), .B(n_1722), .Y(n_1794) );
NAND2xp5_ASAP7_75t_L g1885 ( .A(n_1699), .B(n_1815), .Y(n_1885) );
AND2x2_ASAP7_75t_L g1699 ( .A(n_1700), .B(n_1702), .Y(n_1699) );
AND2x4_ASAP7_75t_L g1750 ( .A(n_1700), .B(n_1702), .Y(n_1750) );
NAND2xp5_ASAP7_75t_L g1703 ( .A(n_1704), .B(n_1718), .Y(n_1703) );
INVx1_ASAP7_75t_L g1704 ( .A(n_1705), .Y(n_1704) );
AND2x2_ASAP7_75t_L g1727 ( .A(n_1705), .B(n_1728), .Y(n_1727) );
AND2x2_ASAP7_75t_L g1705 ( .A(n_1706), .B(n_1711), .Y(n_1705) );
OR2x2_ASAP7_75t_L g1786 ( .A(n_1706), .B(n_1733), .Y(n_1786) );
AND2x2_ASAP7_75t_L g1798 ( .A(n_1706), .B(n_1799), .Y(n_1798) );
AND2x2_ASAP7_75t_L g1813 ( .A(n_1706), .B(n_1753), .Y(n_1813) );
AND2x2_ASAP7_75t_L g1816 ( .A(n_1706), .B(n_1774), .Y(n_1816) );
OR2x2_ASAP7_75t_L g1820 ( .A(n_1706), .B(n_1821), .Y(n_1820) );
AOI321xp33_ASAP7_75t_L g1850 ( .A1(n_1706), .A2(n_1851), .A3(n_1852), .B1(n_1853), .B2(n_1855), .C(n_1856), .Y(n_1850) );
AND2x2_ASAP7_75t_L g1876 ( .A(n_1706), .B(n_1781), .Y(n_1876) );
AND2x2_ASAP7_75t_L g1881 ( .A(n_1706), .B(n_1882), .Y(n_1881) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_1707), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1719 ( .A(n_1707), .B(n_1720), .Y(n_1719) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1707), .B(n_1778), .Y(n_1777) );
AND2x2_ASAP7_75t_L g1838 ( .A(n_1707), .B(n_1711), .Y(n_1838) );
OR2x2_ASAP7_75t_L g1844 ( .A(n_1707), .B(n_1779), .Y(n_1844) );
NAND2xp5_ASAP7_75t_L g1854 ( .A(n_1707), .B(n_1799), .Y(n_1854) );
AND2x2_ASAP7_75t_L g1707 ( .A(n_1708), .B(n_1710), .Y(n_1707) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1708), .B(n_1710), .Y(n_1744) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1711), .Y(n_1760) );
NAND2xp5_ASAP7_75t_L g1874 ( .A(n_1711), .B(n_1815), .Y(n_1874) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1715), .Y(n_1711) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1712), .Y(n_1735) );
INVx1_ASAP7_75t_L g1799 ( .A(n_1712), .Y(n_1799) );
NAND2xp5_ASAP7_75t_L g1712 ( .A(n_1713), .B(n_1714), .Y(n_1712) );
INVx1_ASAP7_75t_L g1720 ( .A(n_1715), .Y(n_1720) );
AND2x2_ASAP7_75t_L g1734 ( .A(n_1715), .B(n_1735), .Y(n_1734) );
OR2x2_ASAP7_75t_L g1754 ( .A(n_1715), .B(n_1735), .Y(n_1754) );
INVx1_ASAP7_75t_L g1779 ( .A(n_1715), .Y(n_1779) );
NAND2xp5_ASAP7_75t_L g1715 ( .A(n_1716), .B(n_1717), .Y(n_1715) );
CKINVDCx14_ASAP7_75t_R g1718 ( .A(n_1719), .Y(n_1718) );
A2O1A1Ixp33_ASAP7_75t_L g1866 ( .A1(n_1719), .A2(n_1809), .B(n_1851), .C(n_1867), .Y(n_1866) );
AND2x2_ASAP7_75t_L g1774 ( .A(n_1720), .B(n_1735), .Y(n_1774) );
NOR2xp33_ASAP7_75t_L g1721 ( .A(n_1722), .B(n_1726), .Y(n_1721) );
INVx3_ASAP7_75t_L g1722 ( .A(n_1723), .Y(n_1722) );
AND2x2_ASAP7_75t_L g1757 ( .A(n_1723), .B(n_1758), .Y(n_1757) );
NOR2xp33_ASAP7_75t_L g1789 ( .A(n_1723), .B(n_1764), .Y(n_1789) );
INVx3_ASAP7_75t_L g1809 ( .A(n_1723), .Y(n_1809) );
AND2x2_ASAP7_75t_L g1839 ( .A(n_1723), .B(n_1782), .Y(n_1839) );
OR2x2_ASAP7_75t_L g1841 ( .A(n_1723), .B(n_1738), .Y(n_1841) );
AND2x2_ASAP7_75t_L g1849 ( .A(n_1723), .B(n_1764), .Y(n_1849) );
AND2x2_ASAP7_75t_L g1855 ( .A(n_1723), .B(n_1737), .Y(n_1855) );
AND2x2_ASAP7_75t_L g1880 ( .A(n_1723), .B(n_1826), .Y(n_1880) );
AND2x4_ASAP7_75t_SL g1723 ( .A(n_1724), .B(n_1725), .Y(n_1723) );
INVxp67_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
AOI221xp5_ASAP7_75t_L g1818 ( .A1(n_1727), .A2(n_1738), .B1(n_1794), .B2(n_1819), .C(n_1824), .Y(n_1818) );
OAI21xp33_ASAP7_75t_L g1770 ( .A1(n_1728), .A2(n_1771), .B(n_1773), .Y(n_1770) );
INVx1_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
NAND2xp5_ASAP7_75t_L g1729 ( .A(n_1730), .B(n_1731), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1749 ( .A(n_1730), .B(n_1750), .Y(n_1749) );
NAND2xp5_ASAP7_75t_L g1736 ( .A(n_1731), .B(n_1737), .Y(n_1736) );
INVx1_ASAP7_75t_L g1746 ( .A(n_1731), .Y(n_1746) );
NOR2xp33_ASAP7_75t_L g1781 ( .A(n_1731), .B(n_1754), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1731), .B(n_1734), .Y(n_1791) );
O2A1O1Ixp33_ASAP7_75t_L g1890 ( .A1(n_1731), .A2(n_1741), .B(n_1891), .C(n_1892), .Y(n_1890) );
NOR2xp33_ASAP7_75t_L g1732 ( .A(n_1733), .B(n_1736), .Y(n_1732) );
OR2x2_ASAP7_75t_L g1870 ( .A(n_1733), .B(n_1744), .Y(n_1870) );
INVx1_ASAP7_75t_L g1733 ( .A(n_1734), .Y(n_1733) );
NAND2xp5_ASAP7_75t_L g1745 ( .A(n_1734), .B(n_1746), .Y(n_1745) );
AND2x2_ASAP7_75t_L g1828 ( .A(n_1734), .B(n_1755), .Y(n_1828) );
NAND3xp33_ASAP7_75t_L g1832 ( .A(n_1734), .B(n_1758), .C(n_1833), .Y(n_1832) );
AND2x2_ASAP7_75t_L g1887 ( .A(n_1734), .B(n_1763), .Y(n_1887) );
INVx1_ASAP7_75t_L g1882 ( .A(n_1735), .Y(n_1882) );
NOR2xp33_ASAP7_75t_L g1775 ( .A(n_1736), .B(n_1776), .Y(n_1775) );
INVx1_ASAP7_75t_L g1801 ( .A(n_1736), .Y(n_1801) );
AND2x2_ASAP7_75t_L g1851 ( .A(n_1737), .B(n_1746), .Y(n_1851) );
INVx2_ASAP7_75t_SL g1737 ( .A(n_1738), .Y(n_1737) );
AOI211xp5_ASAP7_75t_L g1739 ( .A1(n_1740), .A2(n_1742), .B(n_1747), .C(n_1775), .Y(n_1739) );
INVx1_ASAP7_75t_L g1740 ( .A(n_1741), .Y(n_1740) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
OR2x2_ASAP7_75t_L g1743 ( .A(n_1744), .B(n_1745), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1744), .B(n_1774), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1806 ( .A(n_1744), .B(n_1753), .Y(n_1806) );
AOI32xp33_ASAP7_75t_L g1857 ( .A1(n_1744), .A2(n_1789), .A3(n_1858), .B1(n_1859), .B2(n_1861), .Y(n_1857) );
OAI211xp5_ASAP7_75t_L g1856 ( .A1(n_1745), .A2(n_1848), .B(n_1857), .C(n_1862), .Y(n_1856) );
AND2x2_ASAP7_75t_L g1833 ( .A(n_1746), .B(n_1834), .Y(n_1833) );
AND2x2_ASAP7_75t_L g1861 ( .A(n_1746), .B(n_1774), .Y(n_1861) );
OAI211xp5_ASAP7_75t_SL g1747 ( .A1(n_1748), .A2(n_1751), .B(n_1756), .C(n_1770), .Y(n_1747) );
INVx1_ASAP7_75t_L g1748 ( .A(n_1749), .Y(n_1748) );
AOI221xp5_ASAP7_75t_L g1875 ( .A1(n_1749), .A2(n_1814), .B1(n_1855), .B2(n_1876), .C(n_1877), .Y(n_1875) );
INVx2_ASAP7_75t_L g1758 ( .A(n_1750), .Y(n_1758) );
CKINVDCx6p67_ASAP7_75t_R g1808 ( .A(n_1750), .Y(n_1808) );
NAND2xp5_ASAP7_75t_L g1829 ( .A(n_1750), .B(n_1830), .Y(n_1829) );
INVx1_ASAP7_75t_L g1751 ( .A(n_1752), .Y(n_1751) );
AND2x2_ASAP7_75t_L g1752 ( .A(n_1753), .B(n_1755), .Y(n_1752) );
NAND2xp5_ASAP7_75t_L g1762 ( .A(n_1753), .B(n_1763), .Y(n_1762) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
AND2x2_ASAP7_75t_L g1823 ( .A(n_1755), .B(n_1774), .Y(n_1823) );
INVx1_ASAP7_75t_L g1878 ( .A(n_1755), .Y(n_1878) );
AOI221xp5_ASAP7_75t_L g1756 ( .A1(n_1757), .A2(n_1759), .B1(n_1761), .B2(n_1764), .C(n_1766), .Y(n_1756) );
OAI22xp5_ASAP7_75t_L g1783 ( .A1(n_1757), .A2(n_1758), .B1(n_1784), .B2(n_1786), .Y(n_1783) );
INVx1_ASAP7_75t_L g1845 ( .A(n_1757), .Y(n_1845) );
OAI22xp5_ASAP7_75t_L g1819 ( .A1(n_1758), .A2(n_1807), .B1(n_1820), .B2(n_1822), .Y(n_1819) );
INVx1_ASAP7_75t_L g1892 ( .A(n_1759), .Y(n_1892) );
OAI22xp5_ASAP7_75t_L g1787 ( .A1(n_1760), .A2(n_1788), .B1(n_1790), .B2(n_1792), .Y(n_1787) );
NAND2xp5_ASAP7_75t_L g1859 ( .A(n_1760), .B(n_1860), .Y(n_1859) );
INVx1_ASAP7_75t_L g1761 ( .A(n_1762), .Y(n_1761) );
NAND2xp5_ASAP7_75t_L g1785 ( .A(n_1762), .B(n_1782), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1793 ( .A(n_1764), .B(n_1794), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1764), .B(n_1887), .Y(n_1886) );
INVx1_ASAP7_75t_L g1764 ( .A(n_1765), .Y(n_1764) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1767), .Y(n_1766) );
INVx1_ASAP7_75t_L g1864 ( .A(n_1767), .Y(n_1864) );
AND2x2_ASAP7_75t_L g1767 ( .A(n_1768), .B(n_1769), .Y(n_1767) );
O2A1O1Ixp33_ASAP7_75t_L g1888 ( .A1(n_1771), .A2(n_1828), .B(n_1889), .C(n_1890), .Y(n_1888) );
INVx1_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
INVx1_ASAP7_75t_L g1891 ( .A(n_1773), .Y(n_1891) );
INVx1_ASAP7_75t_L g1860 ( .A(n_1774), .Y(n_1860) );
NAND2xp5_ASAP7_75t_L g1811 ( .A(n_1776), .B(n_1812), .Y(n_1811) );
INVx1_ASAP7_75t_L g1776 ( .A(n_1777), .Y(n_1776) );
A2O1A1Ixp33_ASAP7_75t_L g1883 ( .A1(n_1777), .A2(n_1852), .B(n_1884), .C(n_1886), .Y(n_1883) );
INVx1_ASAP7_75t_L g1778 ( .A(n_1779), .Y(n_1778) );
O2A1O1Ixp33_ASAP7_75t_L g1780 ( .A1(n_1781), .A2(n_1782), .B(n_1783), .C(n_1787), .Y(n_1780) );
NAND2xp5_ASAP7_75t_L g1804 ( .A(n_1781), .B(n_1782), .Y(n_1804) );
INVx1_ASAP7_75t_L g1834 ( .A(n_1782), .Y(n_1834) );
INVxp67_ASAP7_75t_L g1784 ( .A(n_1785), .Y(n_1784) );
NOR2xp33_ASAP7_75t_L g1847 ( .A(n_1786), .B(n_1848), .Y(n_1847) );
INVx1_ASAP7_75t_L g1788 ( .A(n_1789), .Y(n_1788) );
INVx1_ASAP7_75t_L g1790 ( .A(n_1791), .Y(n_1790) );
AOI21xp33_ASAP7_75t_L g1872 ( .A1(n_1792), .A2(n_1873), .B(n_1874), .Y(n_1872) );
INVx1_ASAP7_75t_L g1792 ( .A(n_1793), .Y(n_1792) );
AOI221xp5_ASAP7_75t_L g1868 ( .A1(n_1794), .A2(n_1830), .B1(n_1869), .B2(n_1871), .C(n_1872), .Y(n_1868) );
OAI21xp33_ASAP7_75t_L g1795 ( .A1(n_1796), .A2(n_1803), .B(n_1809), .Y(n_1795) );
OAI21xp33_ASAP7_75t_L g1796 ( .A1(n_1797), .A2(n_1800), .B(n_1802), .Y(n_1796) );
NOR2xp33_ASAP7_75t_L g1830 ( .A(n_1797), .B(n_1831), .Y(n_1830) );
INVx1_ASAP7_75t_L g1797 ( .A(n_1798), .Y(n_1797) );
INVxp67_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
AOI21xp33_ASAP7_75t_SL g1803 ( .A1(n_1804), .A2(n_1805), .B(n_1807), .Y(n_1803) );
INVx1_ASAP7_75t_L g1889 ( .A(n_1804), .Y(n_1889) );
CKINVDCx5p33_ASAP7_75t_R g1805 ( .A(n_1806), .Y(n_1805) );
CKINVDCx6p67_ASAP7_75t_R g1807 ( .A(n_1808), .Y(n_1807) );
INVx2_ASAP7_75t_L g1852 ( .A(n_1809), .Y(n_1852) );
OAI221xp5_ASAP7_75t_L g1840 ( .A1(n_1812), .A2(n_1841), .B1(n_1842), .B2(n_1845), .C(n_1846), .Y(n_1840) );
INVx1_ASAP7_75t_L g1812 ( .A(n_1813), .Y(n_1812) );
AND2x2_ASAP7_75t_L g1814 ( .A(n_1815), .B(n_1816), .Y(n_1814) );
NOR2xp33_ASAP7_75t_L g1843 ( .A(n_1815), .B(n_1844), .Y(n_1843) );
NAND3xp33_ASAP7_75t_L g1817 ( .A(n_1818), .B(n_1835), .C(n_1850), .Y(n_1817) );
AOI211xp5_ASAP7_75t_L g1877 ( .A1(n_1821), .A2(n_1878), .B(n_1879), .C(n_1881), .Y(n_1877) );
INVx1_ASAP7_75t_L g1822 ( .A(n_1823), .Y(n_1822) );
OAI211xp5_ASAP7_75t_L g1824 ( .A1(n_1825), .A2(n_1827), .B(n_1829), .C(n_1832), .Y(n_1824) );
CKINVDCx14_ASAP7_75t_R g1825 ( .A(n_1826), .Y(n_1825) );
INVx1_ASAP7_75t_L g1827 ( .A(n_1828), .Y(n_1827) );
O2A1O1Ixp33_ASAP7_75t_L g1835 ( .A1(n_1828), .A2(n_1836), .B(n_1839), .C(n_1840), .Y(n_1835) );
INVx1_ASAP7_75t_L g1836 ( .A(n_1837), .Y(n_1836) );
INVx1_ASAP7_75t_L g1873 ( .A(n_1838), .Y(n_1873) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1841), .Y(n_1871) );
INVx1_ASAP7_75t_L g1842 ( .A(n_1843), .Y(n_1842) );
INVxp67_ASAP7_75t_SL g1846 ( .A(n_1847), .Y(n_1846) );
INVx1_ASAP7_75t_L g1848 ( .A(n_1849), .Y(n_1848) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1854), .Y(n_1853) );
INVx1_ASAP7_75t_L g1862 ( .A(n_1863), .Y(n_1862) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1864), .Y(n_1863) );
NAND5xp2_ASAP7_75t_SL g1865 ( .A(n_1866), .B(n_1868), .C(n_1875), .D(n_1883), .E(n_1888), .Y(n_1865) );
INVx1_ASAP7_75t_L g1869 ( .A(n_1870), .Y(n_1869) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1880), .Y(n_1879) );
INVx1_ASAP7_75t_L g1884 ( .A(n_1885), .Y(n_1884) );
CKINVDCx20_ASAP7_75t_R g1893 ( .A(n_1894), .Y(n_1893) );
CKINVDCx20_ASAP7_75t_R g1894 ( .A(n_1895), .Y(n_1894) );
NAND3xp33_ASAP7_75t_L g1897 ( .A(n_1898), .B(n_1929), .C(n_1938), .Y(n_1897) );
NOR2xp33_ASAP7_75t_L g1898 ( .A(n_1899), .B(n_1918), .Y(n_1898) );
OAI22xp5_ASAP7_75t_L g1920 ( .A1(n_1901), .A2(n_1910), .B1(n_1921), .B2(n_1922), .Y(n_1920) );
INVx2_ASAP7_75t_L g1907 ( .A(n_1908), .Y(n_1907) );
INVx2_ASAP7_75t_L g1912 ( .A(n_1913), .Y(n_1912) );
INVx1_ASAP7_75t_L g1913 ( .A(n_1914), .Y(n_1913) );
INVx1_ASAP7_75t_L g1924 ( .A(n_1925), .Y(n_1924) );
INVx2_ASAP7_75t_L g1927 ( .A(n_1928), .Y(n_1927) );
INVx1_ASAP7_75t_L g1936 ( .A(n_1937), .Y(n_1936) );
CKINVDCx20_ASAP7_75t_R g1947 ( .A(n_1948), .Y(n_1947) );
CKINVDCx20_ASAP7_75t_R g1948 ( .A(n_1949), .Y(n_1948) );
INVx3_ASAP7_75t_L g1949 ( .A(n_1950), .Y(n_1949) );
BUFx3_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
HB1xp67_ASAP7_75t_L g1954 ( .A(n_1955), .Y(n_1954) );
BUFx3_ASAP7_75t_L g1955 ( .A(n_1956), .Y(n_1955) );
INVxp33_ASAP7_75t_L g1957 ( .A(n_1958), .Y(n_1957) );
INVx1_ASAP7_75t_L g1959 ( .A(n_1960), .Y(n_1959) );
AND3x1_ASAP7_75t_L g1960 ( .A(n_1961), .B(n_1985), .C(n_1993), .Y(n_1960) );
NOR2xp33_ASAP7_75t_L g1961 ( .A(n_1962), .B(n_1975), .Y(n_1961) );
INVx1_ASAP7_75t_L g1978 ( .A(n_1979), .Y(n_1978) );
BUFx3_ASAP7_75t_L g1983 ( .A(n_1984), .Y(n_1983) );
HB1xp67_ASAP7_75t_L g1999 ( .A(n_2000), .Y(n_1999) );
INVx1_ASAP7_75t_L g2002 ( .A(n_2003), .Y(n_2002) );
endmodule