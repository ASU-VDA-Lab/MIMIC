module fake_netlist_1_10075_n_664 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_664);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_664;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_243;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_409;
wire n_315;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_440;
wire n_106;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_25), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_32), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_7), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_8), .Y(n_92) );
INVx2_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_79), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_4), .Y(n_95) );
INVx2_ASAP7_75t_L g96 ( .A(n_11), .Y(n_96) );
CKINVDCx5p33_ASAP7_75t_R g97 ( .A(n_76), .Y(n_97) );
CKINVDCx5p33_ASAP7_75t_R g98 ( .A(n_35), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_85), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_18), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_63), .Y(n_101) );
NAND2xp5_ASAP7_75t_L g102 ( .A(n_19), .B(n_64), .Y(n_102) );
INVx2_ASAP7_75t_SL g103 ( .A(n_7), .Y(n_103) );
INVxp67_ASAP7_75t_SL g104 ( .A(n_61), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_26), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_21), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_50), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_55), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_59), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_48), .Y(n_111) );
INVxp67_ASAP7_75t_L g112 ( .A(n_18), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_57), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_51), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_39), .Y(n_115) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_60), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_72), .Y(n_118) );
INVxp33_ASAP7_75t_L g119 ( .A(n_15), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_66), .Y(n_120) );
INVx2_ASAP7_75t_SL g121 ( .A(n_49), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_5), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_80), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_86), .Y(n_124) );
INVx2_ASAP7_75t_L g125 ( .A(n_30), .Y(n_125) );
INVxp67_ASAP7_75t_SL g126 ( .A(n_15), .Y(n_126) );
CKINVDCx14_ASAP7_75t_R g127 ( .A(n_1), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_58), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_52), .Y(n_129) );
OAI21x1_ASAP7_75t_L g130 ( .A1(n_93), .A2(n_40), .B(n_87), .Y(n_130) );
INVx4_ASAP7_75t_L g131 ( .A(n_115), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g132 ( .A(n_103), .B(n_0), .Y(n_132) );
BUFx12f_ASAP7_75t_L g133 ( .A(n_89), .Y(n_133) );
INVxp67_ASAP7_75t_L g134 ( .A(n_108), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_119), .B(n_0), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_93), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_96), .Y(n_137) );
INVx4_ASAP7_75t_L g138 ( .A(n_115), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_125), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_125), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_90), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_127), .B(n_96), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_90), .Y(n_144) );
INVx3_ASAP7_75t_L g145 ( .A(n_94), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_94), .Y(n_146) );
AND2x4_ASAP7_75t_L g147 ( .A(n_121), .B(n_1), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_121), .B(n_2), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_99), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_103), .Y(n_151) );
INVx1_ASAP7_75t_L g152 ( .A(n_101), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_101), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_106), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_106), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_116), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_107), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_130), .Y(n_158) );
AND2x6_ASAP7_75t_L g159 ( .A(n_147), .B(n_107), .Y(n_159) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_130), .Y(n_160) );
INVxp67_ASAP7_75t_L g161 ( .A(n_143), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_130), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_142), .Y(n_163) );
INVx4_ASAP7_75t_L g164 ( .A(n_147), .Y(n_164) );
INVx4_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
INVx2_ASAP7_75t_SL g166 ( .A(n_144), .Y(n_166) );
AND2x6_ASAP7_75t_SL g167 ( .A(n_132), .B(n_91), .Y(n_167) );
INVx2_ASAP7_75t_L g168 ( .A(n_142), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_147), .Y(n_169) );
OR2x2_ASAP7_75t_L g170 ( .A(n_131), .B(n_112), .Y(n_170) );
AND2x2_ASAP7_75t_L g171 ( .A(n_143), .B(n_91), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_143), .B(n_95), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_144), .B(n_111), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_142), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_131), .B(n_111), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_142), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_147), .B(n_114), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_136), .Y(n_178) );
INVx3_ASAP7_75t_L g179 ( .A(n_142), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_131), .B(n_114), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
BUFx2_ASAP7_75t_L g182 ( .A(n_131), .Y(n_182) );
BUFx3_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_145), .Y(n_184) );
OR2x6_ASAP7_75t_L g185 ( .A(n_131), .B(n_95), .Y(n_185) );
BUFx8_ASAP7_75t_SL g186 ( .A(n_156), .Y(n_186) );
INVx4_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_146), .B(n_117), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_145), .Y(n_189) );
HB1xp67_ASAP7_75t_L g190 ( .A(n_138), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_138), .B(n_97), .Y(n_191) );
INVx2_ASAP7_75t_L g192 ( .A(n_187), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_185), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_182), .B(n_138), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_187), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_183), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_190), .B(n_134), .Y(n_197) );
INVx1_ASAP7_75t_L g198 ( .A(n_179), .Y(n_198) );
CKINVDCx20_ASAP7_75t_R g199 ( .A(n_186), .Y(n_199) );
CKINVDCx5p33_ASAP7_75t_R g200 ( .A(n_185), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_183), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_179), .Y(n_202) );
AOI22xp33_ASAP7_75t_L g203 ( .A1(n_159), .A2(n_135), .B1(n_138), .B2(n_148), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_185), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_160), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_182), .B(n_138), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_183), .B(n_134), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_170), .B(n_151), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_185), .A2(n_135), .B1(n_148), .B2(n_154), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_190), .B(n_151), .Y(n_210) );
AND2x2_ASAP7_75t_L g211 ( .A(n_161), .B(n_135), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_187), .Y(n_212) );
INVxp67_ASAP7_75t_L g213 ( .A(n_170), .Y(n_213) );
NAND3xp33_ASAP7_75t_SL g214 ( .A(n_161), .B(n_122), .C(n_105), .Y(n_214) );
NOR2xp67_ASAP7_75t_L g215 ( .A(n_164), .B(n_145), .Y(n_215) );
INVx1_ASAP7_75t_SL g216 ( .A(n_185), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_187), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_179), .Y(n_218) );
INVx1_ASAP7_75t_L g219 ( .A(n_179), .Y(n_219) );
INVx2_ASAP7_75t_SL g220 ( .A(n_164), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_168), .Y(n_221) );
HB1xp67_ASAP7_75t_L g222 ( .A(n_171), .Y(n_222) );
INVx5_ASAP7_75t_L g223 ( .A(n_159), .Y(n_223) );
NAND2xp33_ASAP7_75t_L g224 ( .A(n_159), .B(n_146), .Y(n_224) );
AO22x1_ASAP7_75t_L g225 ( .A1(n_159), .A2(n_177), .B1(n_158), .B2(n_162), .Y(n_225) );
HB1xp67_ASAP7_75t_L g226 ( .A(n_171), .Y(n_226) );
AND2x4_ASAP7_75t_L g227 ( .A(n_172), .B(n_149), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_168), .Y(n_228) );
BUFx3_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_172), .B(n_149), .Y(n_230) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_166), .B(n_133), .Y(n_231) );
INVx3_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_175), .B(n_152), .Y(n_233) );
OR2x6_ASAP7_75t_L g234 ( .A(n_164), .B(n_165), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_165), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_228), .Y(n_236) );
OAI33xp33_ASAP7_75t_L g237 ( .A1(n_210), .A2(n_188), .A3(n_173), .B1(n_132), .B2(n_153), .B3(n_154), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_213), .B(n_180), .Y(n_238) );
BUFx12f_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_221), .Y(n_240) );
INVx5_ASAP7_75t_L g241 ( .A(n_234), .Y(n_241) );
AND2x2_ASAP7_75t_L g242 ( .A(n_211), .B(n_165), .Y(n_242) );
BUFx6f_ASAP7_75t_L g243 ( .A(n_229), .Y(n_243) );
INVx8_ASAP7_75t_L g244 ( .A(n_234), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_SL g245 ( .A1(n_208), .A2(n_162), .B(n_158), .C(n_169), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_197), .B(n_159), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_227), .B(n_159), .Y(n_247) );
AND2x2_ASAP7_75t_SL g248 ( .A(n_193), .B(n_165), .Y(n_248) );
OAI22xp33_ASAP7_75t_L g249 ( .A1(n_200), .A2(n_188), .B1(n_173), .B2(n_169), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_222), .Y(n_250) );
AOI22xp33_ASAP7_75t_L g251 ( .A1(n_193), .A2(n_159), .B1(n_177), .B2(n_169), .Y(n_251) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_225), .A2(n_158), .B(n_162), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_226), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_227), .B(n_177), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_228), .Y(n_255) );
NOR2xp33_ASAP7_75t_L g256 ( .A(n_211), .B(n_191), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_225), .A2(n_169), .B(n_166), .Y(n_257) );
INVx2_ASAP7_75t_L g258 ( .A(n_221), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_223), .Y(n_259) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_229), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_227), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_227), .B(n_177), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_192), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_230), .B(n_177), .Y(n_264) );
CKINVDCx20_ASAP7_75t_R g265 ( .A(n_199), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_234), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_192), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_230), .B(n_166), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_195), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_195), .Y(n_270) );
INVx4_ASAP7_75t_L g271 ( .A(n_204), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_212), .Y(n_272) );
OR2x2_ASAP7_75t_SL g273 ( .A(n_214), .B(n_167), .Y(n_273) );
INVx5_ASAP7_75t_L g274 ( .A(n_234), .Y(n_274) );
INVx6_ASAP7_75t_L g275 ( .A(n_223), .Y(n_275) );
AOI21xp33_ASAP7_75t_L g276 ( .A1(n_216), .A2(n_133), .B(n_184), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_207), .B(n_167), .Y(n_277) );
INVx2_ASAP7_75t_L g278 ( .A(n_212), .Y(n_278) );
OAI22xp5_ASAP7_75t_L g279 ( .A1(n_204), .A2(n_189), .B1(n_184), .B2(n_163), .Y(n_279) );
AOI22xp33_ASAP7_75t_L g280 ( .A1(n_277), .A2(n_230), .B1(n_201), .B2(n_196), .Y(n_280) );
OA21x2_ASAP7_75t_L g281 ( .A1(n_252), .A2(n_157), .B(n_150), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_258), .Y(n_282) );
OAI21x1_ASAP7_75t_L g283 ( .A1(n_257), .A2(n_150), .B(n_157), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_258), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_236), .Y(n_285) );
NOR2xp33_ASAP7_75t_SL g286 ( .A(n_244), .B(n_229), .Y(n_286) );
OAI21x1_ASAP7_75t_L g287 ( .A1(n_240), .A2(n_150), .B(n_157), .Y(n_287) );
INVx1_ASAP7_75t_SL g288 ( .A(n_241), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_244), .B(n_196), .Y(n_289) );
OA21x2_ASAP7_75t_L g290 ( .A1(n_240), .A2(n_117), .B(n_129), .Y(n_290) );
AOI22xp33_ASAP7_75t_L g291 ( .A1(n_250), .A2(n_230), .B1(n_201), .B2(n_177), .Y(n_291) );
AO31x2_ASAP7_75t_L g292 ( .A1(n_236), .A2(n_139), .A3(n_136), .B(n_141), .Y(n_292) );
OAI22xp33_ASAP7_75t_L g293 ( .A1(n_244), .A2(n_209), .B1(n_234), .B2(n_233), .Y(n_293) );
OAI21x1_ASAP7_75t_L g294 ( .A1(n_255), .A2(n_124), .B(n_120), .Y(n_294) );
INVxp67_ASAP7_75t_L g295 ( .A(n_242), .Y(n_295) );
OAI21x1_ASAP7_75t_L g296 ( .A1(n_255), .A2(n_124), .B(n_120), .Y(n_296) );
INVx2_ASAP7_75t_L g297 ( .A(n_263), .Y(n_297) );
AOI22xp33_ASAP7_75t_L g298 ( .A1(n_253), .A2(n_177), .B1(n_203), .B2(n_209), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_263), .Y(n_299) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_266), .A2(n_128), .B(n_123), .Y(n_300) );
BUFx2_ASAP7_75t_SL g301 ( .A(n_241), .Y(n_301) );
O2A1O1Ixp33_ASAP7_75t_SL g302 ( .A1(n_245), .A2(n_102), .B(n_231), .C(n_219), .Y(n_302) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_244), .A2(n_223), .B1(n_215), .B2(n_133), .Y(n_303) );
AOI22x1_ASAP7_75t_L g304 ( .A1(n_269), .A2(n_160), .B1(n_205), .B2(n_178), .Y(n_304) );
A2O1A1Ixp33_ASAP7_75t_L g305 ( .A1(n_256), .A2(n_215), .B(n_224), .C(n_232), .Y(n_305) );
INVx3_ASAP7_75t_SL g306 ( .A(n_241), .Y(n_306) );
AOI21x1_ASAP7_75t_L g307 ( .A1(n_246), .A2(n_141), .B(n_136), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_269), .Y(n_308) );
OAI21x1_ASAP7_75t_L g309 ( .A1(n_266), .A2(n_279), .B(n_278), .Y(n_309) );
OAI21x1_ASAP7_75t_L g310 ( .A1(n_266), .A2(n_128), .B(n_123), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_242), .B(n_177), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_232), .Y(n_312) );
OR2x2_ASAP7_75t_SL g313 ( .A(n_273), .B(n_100), .Y(n_313) );
OA21x2_ASAP7_75t_L g314 ( .A1(n_267), .A2(n_129), .B(n_155), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_278), .A2(n_198), .B(n_202), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_282), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_295), .B(n_261), .Y(n_317) );
AOI22xp33_ASAP7_75t_L g318 ( .A1(n_293), .A2(n_237), .B1(n_248), .B2(n_268), .Y(n_318) );
OR2x2_ASAP7_75t_L g319 ( .A(n_282), .B(n_238), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_284), .B(n_248), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_306), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g323 ( .A1(n_284), .A2(n_249), .B1(n_271), .B2(n_241), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_285), .Y(n_325) );
AOI21xp5_ASAP7_75t_L g326 ( .A1(n_302), .A2(n_205), .B(n_160), .Y(n_326) );
AND2x4_ASAP7_75t_L g327 ( .A(n_289), .B(n_241), .Y(n_327) );
OAI22xp33_ASAP7_75t_L g328 ( .A1(n_286), .A2(n_274), .B1(n_239), .B2(n_271), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_298), .A2(n_239), .B1(n_274), .B2(n_276), .Y(n_329) );
OAI21xp5_ASAP7_75t_L g330 ( .A1(n_287), .A2(n_267), .B(n_270), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_285), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_297), .Y(n_332) );
NAND2x1p5_ASAP7_75t_L g333 ( .A(n_288), .B(n_274), .Y(n_333) );
OA21x2_ASAP7_75t_L g334 ( .A1(n_309), .A2(n_141), .B(n_139), .Y(n_334) );
OAI22xp33_ASAP7_75t_L g335 ( .A1(n_286), .A2(n_274), .B1(n_271), .B2(n_265), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_295), .B(n_274), .Y(n_336) );
AOI22xp33_ASAP7_75t_L g337 ( .A1(n_280), .A2(n_254), .B1(n_247), .B2(n_262), .Y(n_337) );
AO21x2_ASAP7_75t_L g338 ( .A1(n_309), .A2(n_139), .B(n_153), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_297), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_312), .B(n_270), .Y(n_340) );
OAI21x1_ASAP7_75t_L g341 ( .A1(n_304), .A2(n_272), .B(n_202), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_312), .A2(n_264), .B1(n_206), .B2(n_194), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_297), .B(n_299), .Y(n_343) );
OA21x2_ASAP7_75t_L g344 ( .A1(n_283), .A2(n_155), .B(n_152), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_291), .A2(n_251), .B1(n_92), .B2(n_126), .C(n_100), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_316), .B(n_299), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_332), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_322), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_316), .B(n_299), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_320), .B(n_340), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_320), .B(n_308), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_327), .B(n_288), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_318), .A2(n_301), .B1(n_306), .B2(n_289), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_340), .B(n_308), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_332), .Y(n_356) );
INVx3_ASAP7_75t_L g357 ( .A(n_321), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_324), .B(n_308), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_324), .B(n_281), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_325), .B(n_281), .Y(n_360) );
INVxp67_ASAP7_75t_SL g361 ( .A(n_343), .Y(n_361) );
BUFx2_ASAP7_75t_L g362 ( .A(n_333), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_325), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_319), .B(n_292), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_331), .B(n_339), .Y(n_365) );
OR2x2_ASAP7_75t_L g366 ( .A(n_319), .B(n_292), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_331), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_339), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_332), .B(n_290), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_317), .B(n_281), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_327), .B(n_290), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_321), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_338), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_338), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_348), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_347), .Y(n_376) );
INVxp67_ASAP7_75t_SL g377 ( .A(n_367), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_338), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_348), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_364), .Y(n_380) );
OAI22xp5_ASAP7_75t_SL g381 ( .A1(n_354), .A2(n_265), .B1(n_313), .B2(n_273), .Y(n_381) );
INVxp67_ASAP7_75t_L g382 ( .A(n_365), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_364), .B(n_313), .Y(n_383) );
NAND3xp33_ASAP7_75t_L g384 ( .A(n_373), .B(n_137), .C(n_140), .Y(n_384) );
OAI321xp33_ASAP7_75t_L g385 ( .A1(n_367), .A2(n_335), .A3(n_328), .B1(n_345), .B2(n_323), .C(n_329), .Y(n_385) );
NAND3xp33_ASAP7_75t_SL g386 ( .A(n_366), .B(n_109), .C(n_333), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_347), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_350), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_347), .Y(n_389) );
AND2x4_ASAP7_75t_L g390 ( .A(n_371), .B(n_327), .Y(n_390) );
AND2x4_ASAP7_75t_L g391 ( .A(n_371), .B(n_327), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_366), .B(n_323), .Y(n_392) );
AOI22xp5_ASAP7_75t_L g393 ( .A1(n_353), .A2(n_336), .B1(n_337), .B2(n_301), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_356), .Y(n_394) );
NOR3xp33_ASAP7_75t_L g395 ( .A(n_355), .B(n_109), .C(n_140), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g396 ( .A(n_351), .B(n_104), .Y(n_396) );
INVx3_ASAP7_75t_SL g397 ( .A(n_353), .Y(n_397) );
NOR3xp33_ASAP7_75t_SL g398 ( .A(n_355), .B(n_303), .C(n_110), .Y(n_398) );
INVx2_ASAP7_75t_L g399 ( .A(n_356), .Y(n_399) );
INVx2_ASAP7_75t_SL g400 ( .A(n_372), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_356), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_350), .Y(n_402) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_137), .B1(n_113), .B2(n_342), .C(n_305), .Y(n_403) );
AND2x4_ASAP7_75t_SL g404 ( .A(n_353), .B(n_321), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_365), .B(n_334), .Y(n_405) );
OAI221xp5_ASAP7_75t_L g406 ( .A1(n_374), .A2(n_333), .B1(n_306), .B2(n_330), .C(n_289), .Y(n_406) );
AOI221xp5_ASAP7_75t_L g407 ( .A1(n_374), .A2(n_330), .B1(n_178), .B2(n_311), .C(n_163), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_363), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_363), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_382), .B(n_352), .Y(n_410) );
INVx1_ASAP7_75t_SL g411 ( .A(n_397), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_380), .B(n_368), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_378), .B(n_352), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_383), .B(n_368), .Y(n_414) );
AND2x2_ASAP7_75t_L g415 ( .A(n_378), .B(n_369), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_381), .B(n_362), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_383), .B(n_361), .Y(n_417) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_375), .B(n_369), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_376), .Y(n_419) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_375), .Y(n_421) );
OR2x2_ASAP7_75t_L g422 ( .A(n_377), .B(n_362), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_390), .Y(n_423) );
OR2x2_ASAP7_75t_L g424 ( .A(n_390), .B(n_346), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_405), .B(n_359), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_379), .B(n_346), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_387), .Y(n_427) );
AND3x2_ASAP7_75t_L g428 ( .A(n_395), .B(n_353), .C(n_358), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_405), .B(n_359), .Y(n_429) );
NAND4xp25_ASAP7_75t_SL g430 ( .A(n_392), .B(n_349), .C(n_358), .D(n_360), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_390), .B(n_372), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_387), .Y(n_432) );
AND2x2_ASAP7_75t_L g433 ( .A(n_391), .B(n_372), .Y(n_433) );
AND2x2_ASAP7_75t_L g434 ( .A(n_391), .B(n_360), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_400), .B(n_357), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_391), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_397), .B(n_349), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_396), .B(n_357), .Y(n_438) );
AND2x2_ASAP7_75t_L g439 ( .A(n_402), .B(n_357), .Y(n_439) );
NOR2x1_ASAP7_75t_L g440 ( .A(n_386), .B(n_357), .Y(n_440) );
NAND4xp25_ASAP7_75t_L g441 ( .A(n_393), .B(n_370), .C(n_311), .D(n_326), .Y(n_441) );
INVx3_ASAP7_75t_SL g442 ( .A(n_404), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_400), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_379), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_402), .B(n_370), .Y(n_445) );
NOR2xp67_ASAP7_75t_SL g446 ( .A(n_406), .B(n_321), .Y(n_446) );
NAND3xp33_ASAP7_75t_L g447 ( .A(n_398), .B(n_290), .C(n_178), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_389), .Y(n_448) );
OR2x2_ASAP7_75t_L g449 ( .A(n_408), .B(n_292), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_388), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_388), .B(n_292), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_389), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_394), .Y(n_453) );
NOR2x1_ASAP7_75t_L g454 ( .A(n_384), .B(n_321), .Y(n_454) );
OAI21xp33_ASAP7_75t_L g455 ( .A1(n_392), .A2(n_178), .B(n_300), .Y(n_455) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_394), .Y(n_456) );
NAND3xp33_ASAP7_75t_L g457 ( .A(n_403), .B(n_290), .C(n_178), .Y(n_457) );
NAND2x1_ASAP7_75t_L g458 ( .A(n_408), .B(n_409), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_409), .B(n_292), .Y(n_459) );
AND2x4_ASAP7_75t_SL g460 ( .A(n_399), .B(n_321), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_425), .B(n_399), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_458), .Y(n_462) );
AND4x1_ASAP7_75t_L g463 ( .A(n_446), .B(n_407), .C(n_3), .D(n_4), .Y(n_463) );
OR2x2_ASAP7_75t_L g464 ( .A(n_424), .B(n_401), .Y(n_464) );
AND2x2_ASAP7_75t_L g465 ( .A(n_413), .B(n_404), .Y(n_465) );
OAI31xp33_ASAP7_75t_L g466 ( .A1(n_416), .A2(n_401), .A3(n_385), .B(n_5), .Y(n_466) );
NAND3xp33_ASAP7_75t_L g467 ( .A(n_438), .B(n_314), .C(n_178), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_413), .B(n_334), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_425), .B(n_334), .Y(n_469) );
OAI21xp33_ASAP7_75t_SL g470 ( .A1(n_411), .A2(n_310), .B(n_300), .Y(n_470) );
BUFx2_ASAP7_75t_L g471 ( .A(n_442), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_420), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_429), .B(n_334), .Y(n_473) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_437), .Y(n_474) );
AO211x2_ASAP7_75t_L g475 ( .A1(n_447), .A2(n_2), .B(n_3), .C(n_6), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_429), .B(n_292), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_415), .B(n_6), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_420), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_415), .B(n_8), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_412), .B(n_9), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_410), .B(n_314), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_414), .B(n_417), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_421), .B(n_314), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_444), .B(n_314), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_434), .B(n_9), .Y(n_485) );
OAI211xp5_ASAP7_75t_L g486 ( .A1(n_416), .A2(n_310), .B(n_294), .C(n_296), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_450), .B(n_10), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_443), .B(n_10), .Y(n_489) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_442), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_434), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_422), .Y(n_492) );
OR2x2_ASAP7_75t_L g493 ( .A(n_445), .B(n_11), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_426), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_419), .Y(n_495) );
OR2x2_ASAP7_75t_L g496 ( .A(n_418), .B(n_13), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_423), .B(n_13), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_428), .B(n_14), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_428), .B(n_14), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_451), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_459), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_431), .B(n_16), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_439), .B(n_16), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_439), .B(n_17), .Y(n_504) );
OR2x6_ASAP7_75t_L g505 ( .A(n_440), .B(n_289), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_419), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_427), .B(n_281), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_427), .B(n_344), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_432), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_432), .B(n_344), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_448), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_448), .B(n_344), .Y(n_512) );
OAI22xp5_ASAP7_75t_L g513 ( .A1(n_454), .A2(n_289), .B1(n_344), .B2(n_307), .Y(n_513) );
AND2x2_ASAP7_75t_L g514 ( .A(n_433), .B(n_17), .Y(n_514) );
OR2x2_ASAP7_75t_L g515 ( .A(n_423), .B(n_294), .Y(n_515) );
OR2x2_ASAP7_75t_L g516 ( .A(n_423), .B(n_296), .Y(n_516) );
NOR2xp33_ASAP7_75t_L g517 ( .A(n_436), .B(n_20), .Y(n_517) );
NAND4xp25_ASAP7_75t_L g518 ( .A(n_441), .B(n_198), .C(n_219), .D(n_176), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_452), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_452), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_500), .B(n_436), .Y(n_521) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_488), .B(n_436), .Y(n_522) );
INVx2_ASAP7_75t_SL g523 ( .A(n_490), .Y(n_523) );
INVx2_ASAP7_75t_L g524 ( .A(n_478), .Y(n_524) );
HB1xp67_ASAP7_75t_L g525 ( .A(n_474), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_471), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_461), .B(n_449), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_501), .B(n_453), .Y(n_528) );
OAI22xp5_ASAP7_75t_L g529 ( .A1(n_505), .A2(n_435), .B1(n_455), .B2(n_457), .Y(n_529) );
OAI22xp5_ASAP7_75t_L g530 ( .A1(n_505), .A2(n_435), .B1(n_460), .B2(n_453), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g531 ( .A1(n_505), .A2(n_490), .B1(n_498), .B2(n_499), .Y(n_531) );
INVx1_ASAP7_75t_SL g532 ( .A(n_490), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_470), .A2(n_430), .B(n_460), .Y(n_533) );
OAI22xp33_ASAP7_75t_L g534 ( .A1(n_518), .A2(n_497), .B1(n_467), .B2(n_493), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_494), .B(n_456), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_491), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_465), .B(n_456), .Y(n_537) );
OAI22xp33_ASAP7_75t_L g538 ( .A1(n_518), .A2(n_456), .B1(n_160), .B2(n_307), .Y(n_538) );
AOI21xp33_ASAP7_75t_L g539 ( .A1(n_466), .A2(n_456), .B(n_118), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_492), .B(n_287), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_482), .B(n_341), .Y(n_541) );
NOR3x1_ASAP7_75t_L g542 ( .A(n_480), .B(n_283), .C(n_315), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_461), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_477), .B(n_315), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_472), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_479), .B(n_341), .Y(n_546) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_513), .A2(n_304), .B(n_205), .Y(n_547) );
INVx1_ASAP7_75t_SL g548 ( .A(n_464), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_495), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_462), .B(n_22), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_506), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_509), .Y(n_552) );
OAI21xp5_ASAP7_75t_L g553 ( .A1(n_466), .A2(n_98), .B(n_272), .Y(n_553) );
BUFx2_ASAP7_75t_L g554 ( .A(n_502), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g555 ( .A1(n_476), .A2(n_160), .B1(n_260), .B2(n_243), .Y(n_555) );
BUFx2_ASAP7_75t_L g556 ( .A(n_514), .Y(n_556) );
INVx2_ASAP7_75t_SL g557 ( .A(n_485), .Y(n_557) );
AND2x2_ASAP7_75t_L g558 ( .A(n_468), .B(n_23), .Y(n_558) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_489), .A2(n_160), .B1(n_174), .B2(n_176), .C(n_189), .Y(n_559) );
NAND2xp33_ASAP7_75t_SL g560 ( .A(n_513), .B(n_260), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_511), .B(n_519), .Y(n_561) );
A2O1A1Ixp33_ASAP7_75t_L g562 ( .A1(n_517), .A2(n_259), .B(n_260), .C(n_243), .Y(n_562) );
AOI21xp33_ASAP7_75t_L g563 ( .A1(n_496), .A2(n_24), .B(n_27), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_481), .B(n_28), .Y(n_564) );
OAI21xp33_ASAP7_75t_SL g565 ( .A1(n_469), .A2(n_29), .B(n_31), .Y(n_565) );
OAI221xp5_ASAP7_75t_L g566 ( .A1(n_463), .A2(n_218), .B1(n_259), .B2(n_174), .C(n_243), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_520), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_487), .Y(n_568) );
AOI221xp5_ASAP7_75t_L g569 ( .A1(n_503), .A2(n_168), .B1(n_181), .B2(n_218), .C(n_205), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_469), .B(n_33), .Y(n_570) );
INVx2_ASAP7_75t_SL g571 ( .A(n_504), .Y(n_571) );
OAI21xp33_ASAP7_75t_L g572 ( .A1(n_473), .A2(n_205), .B(n_181), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_475), .A2(n_260), .B1(n_243), .B2(n_275), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_525), .B(n_473), .Y(n_574) );
A2O1A1Ixp33_ASAP7_75t_L g575 ( .A1(n_526), .A2(n_486), .B(n_515), .C(n_516), .Y(n_575) );
INVx2_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
OAI21xp33_ASAP7_75t_L g577 ( .A1(n_522), .A2(n_484), .B(n_483), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_543), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g579 ( .A(n_526), .B(n_512), .Y(n_579) );
AOI21xp33_ASAP7_75t_SL g580 ( .A1(n_534), .A2(n_512), .B(n_510), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_551), .Y(n_581) );
O2A1O1Ixp33_ASAP7_75t_L g582 ( .A1(n_565), .A2(n_510), .B(n_508), .C(n_507), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_552), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_548), .B(n_508), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_568), .B(n_507), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_536), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_524), .Y(n_587) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_560), .A2(n_181), .B(n_223), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_527), .B(n_34), .Y(n_589) );
AOI22xp33_ASAP7_75t_SL g590 ( .A1(n_554), .A2(n_260), .B1(n_243), .B2(n_275), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_541), .B(n_36), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_549), .Y(n_592) );
OAI211xp5_ASAP7_75t_L g593 ( .A1(n_533), .A2(n_223), .B(n_232), .C(n_41), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_521), .B(n_37), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_528), .Y(n_595) );
AOI32xp33_ASAP7_75t_L g596 ( .A1(n_534), .A2(n_232), .A3(n_42), .B1(n_43), .B2(n_44), .Y(n_596) );
INVxp67_ASAP7_75t_L g597 ( .A(n_571), .Y(n_597) );
AOI22xp33_ASAP7_75t_SL g598 ( .A1(n_556), .A2(n_275), .B1(n_223), .B2(n_46), .Y(n_598) );
OAI21xp33_ASAP7_75t_L g599 ( .A1(n_522), .A2(n_38), .B(n_45), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_561), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_567), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_545), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_535), .B(n_47), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_540), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_523), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_557), .B(n_53), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_546), .B(n_54), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_537), .B(n_56), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_532), .Y(n_609) );
AND2x2_ASAP7_75t_L g610 ( .A(n_609), .B(n_531), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_595), .Y(n_611) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_582), .A2(n_530), .B(n_529), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_580), .B(n_544), .Y(n_613) );
NOR3xp33_ASAP7_75t_L g614 ( .A(n_596), .B(n_539), .C(n_553), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_601), .Y(n_615) );
INVx1_ASAP7_75t_L g616 ( .A(n_578), .Y(n_616) );
OAI21xp5_ASAP7_75t_L g617 ( .A1(n_582), .A2(n_533), .B(n_538), .Y(n_617) );
OAI221xp5_ASAP7_75t_L g618 ( .A1(n_575), .A2(n_560), .B1(n_566), .B2(n_573), .C(n_563), .Y(n_618) );
BUFx2_ASAP7_75t_L g619 ( .A(n_576), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_597), .A2(n_559), .B1(n_555), .B2(n_538), .C(n_569), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_600), .B(n_542), .Y(n_621) );
BUFx3_ASAP7_75t_L g622 ( .A(n_605), .Y(n_622) );
OAI21xp5_ASAP7_75t_L g623 ( .A1(n_593), .A2(n_547), .B(n_562), .Y(n_623) );
AOI22xp5_ASAP7_75t_L g624 ( .A1(n_597), .A2(n_558), .B1(n_570), .B2(n_550), .Y(n_624) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_593), .B(n_547), .C(n_562), .D(n_564), .Y(n_625) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_604), .B(n_572), .Y(n_626) );
NOR2xp33_ASAP7_75t_SL g627 ( .A(n_599), .B(n_275), .Y(n_627) );
OA22x2_ASAP7_75t_L g628 ( .A1(n_574), .A2(n_62), .B1(n_65), .B2(n_67), .Y(n_628) );
INVx1_ASAP7_75t_SL g629 ( .A(n_585), .Y(n_629) );
AOI22xp33_ASAP7_75t_L g630 ( .A1(n_577), .A2(n_235), .B1(n_220), .B2(n_70), .Y(n_630) );
AOI22x1_ASAP7_75t_L g631 ( .A1(n_588), .A2(n_68), .B1(n_69), .B2(n_71), .Y(n_631) );
NOR3xp33_ASAP7_75t_SL g632 ( .A(n_617), .B(n_606), .C(n_591), .Y(n_632) );
NAND4xp25_ASAP7_75t_L g633 ( .A(n_614), .B(n_598), .C(n_590), .D(n_588), .Y(n_633) );
NOR3xp33_ASAP7_75t_L g634 ( .A(n_612), .B(n_598), .C(n_607), .Y(n_634) );
INVxp33_ASAP7_75t_L g635 ( .A(n_610), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_613), .A2(n_579), .B1(n_586), .B2(n_581), .C(n_583), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_622), .A2(n_584), .B1(n_590), .B2(n_587), .Y(n_637) );
AOI211xp5_ASAP7_75t_L g638 ( .A1(n_614), .A2(n_589), .B(n_608), .C(n_594), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_621), .B(n_602), .Y(n_639) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_611), .Y(n_640) );
NOR3xp33_ASAP7_75t_SL g641 ( .A(n_618), .B(n_603), .C(n_75), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_621), .A2(n_592), .B1(n_235), .B2(n_220), .Y(n_642) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_623), .A2(n_73), .B(n_77), .Y(n_643) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_622), .A2(n_78), .B1(n_81), .B2(n_82), .Y(n_644) );
NAND3x1_ASAP7_75t_L g645 ( .A(n_634), .B(n_620), .C(n_624), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_633), .B(n_625), .C(n_626), .Y(n_646) );
AND2x2_ASAP7_75t_L g647 ( .A(n_635), .B(n_629), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_636), .B(n_616), .Y(n_648) );
NOR3xp33_ASAP7_75t_L g649 ( .A(n_637), .B(n_615), .C(n_619), .Y(n_649) );
AND2x4_ASAP7_75t_L g650 ( .A(n_639), .B(n_630), .Y(n_650) );
NOR2xp67_ASAP7_75t_L g651 ( .A(n_642), .B(n_630), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g652 ( .A1(n_646), .A2(n_640), .B(n_643), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_645), .A2(n_651), .B1(n_647), .B2(n_649), .Y(n_653) );
OR4x2_ASAP7_75t_L g654 ( .A(n_650), .B(n_632), .C(n_638), .D(n_641), .Y(n_654) );
OAI211xp5_ASAP7_75t_SL g655 ( .A1(n_648), .A2(n_644), .B(n_628), .C(n_627), .Y(n_655) );
INVx2_ASAP7_75t_SL g656 ( .A(n_654), .Y(n_656) );
XNOR2xp5_ASAP7_75t_L g657 ( .A(n_653), .B(n_628), .Y(n_657) );
XNOR2xp5_ASAP7_75t_L g658 ( .A(n_652), .B(n_631), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_656), .Y(n_659) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_658), .A2(n_655), .B(n_217), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_659), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_661), .A2(n_657), .B1(n_660), .B2(n_217), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_662), .Y(n_663) );
AOI22xp33_ASAP7_75t_SL g664 ( .A1(n_663), .A2(n_83), .B1(n_84), .B2(n_88), .Y(n_664) );
endmodule