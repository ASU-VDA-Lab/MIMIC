module fake_ariane_2523_n_2284 (n_8, n_24, n_7, n_22, n_43, n_1, n_49, n_6, n_13, n_20, n_27, n_48, n_29, n_17, n_4, n_41, n_50, n_38, n_2, n_47, n_18, n_32, n_28, n_37, n_9, n_51, n_45, n_11, n_34, n_26, n_3, n_46, n_14, n_0, n_52, n_36, n_33, n_44, n_19, n_30, n_39, n_40, n_31, n_42, n_16, n_5, n_12, n_15, n_53, n_21, n_23, n_35, n_10, n_54, n_25, n_2284);

input n_8;
input n_24;
input n_7;
input n_22;
input n_43;
input n_1;
input n_49;
input n_6;
input n_13;
input n_20;
input n_27;
input n_48;
input n_29;
input n_17;
input n_4;
input n_41;
input n_50;
input n_38;
input n_2;
input n_47;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_51;
input n_45;
input n_11;
input n_34;
input n_26;
input n_3;
input n_46;
input n_14;
input n_0;
input n_52;
input n_36;
input n_33;
input n_44;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_42;
input n_16;
input n_5;
input n_12;
input n_15;
input n_53;
input n_21;
input n_23;
input n_35;
input n_10;
input n_54;
input n_25;

output n_2284;

wire n_913;
wire n_1681;
wire n_2163;
wire n_1486;
wire n_1507;
wire n_1938;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_2131;
wire n_423;
wire n_1383;
wire n_2182;
wire n_603;
wire n_373;
wire n_2135;
wire n_1250;
wire n_2030;
wire n_1169;
wire n_789;
wire n_850;
wire n_1916;
wire n_610;
wire n_245;
wire n_1713;
wire n_96;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_2002;
wire n_1463;
wire n_2243;
wire n_1238;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_2013;
wire n_1566;
wire n_189;
wire n_717;
wire n_72;
wire n_2006;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_57;
wire n_1706;
wire n_2207;
wire n_117;
wire n_524;
wire n_1214;
wire n_634;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_2042;
wire n_2123;
wire n_1853;
wire n_764;
wire n_1503;
wire n_2238;
wire n_462;
wire n_1196;
wire n_1181;
wire n_1999;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_137;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_2084;
wire n_568;
wire n_2278;
wire n_1088;
wire n_77;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_2248;
wire n_813;
wire n_419;
wire n_1985;
wire n_146;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1909;
wire n_2156;
wire n_1184;
wire n_1961;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1979;
wire n_1277;
wire n_2107;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_2221;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1974;
wire n_1736;
wire n_1018;
wire n_2200;
wire n_69;
wire n_259;
wire n_953;
wire n_1364;
wire n_143;
wire n_1888;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_1944;
wire n_331;
wire n_559;
wire n_2233;
wire n_267;
wire n_495;
wire n_1988;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_1936;
wire n_2149;
wire n_2277;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_2078;
wire n_1145;
wire n_971;
wire n_2201;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_2232;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_2227;
wire n_1539;
wire n_884;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_2192;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_93;
wire n_859;
wire n_1765;
wire n_108;
wire n_1889;
wire n_587;
wire n_1977;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_2060;
wire n_1850;
wire n_238;
wire n_365;
wire n_2004;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_136;
wire n_192;
wire n_661;
wire n_2098;
wire n_1751;
wire n_300;
wire n_533;
wire n_1917;
wire n_104;
wire n_1924;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_2045;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_2061;
wire n_2094;
wire n_1354;
wire n_1790;
wire n_149;
wire n_1213;
wire n_237;
wire n_2043;
wire n_780;
wire n_1918;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1949;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_2077;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1947;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_2038;
wire n_2263;
wire n_2116;
wire n_2271;
wire n_2145;
wire n_1838;
wire n_1594;
wire n_680;
wire n_1935;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_2281;
wire n_1432;
wire n_94;
wire n_2245;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_65;
wire n_123;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_2216;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_135;
wire n_947;
wire n_2134;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_102;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_78;
wire n_2166;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_2185;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_2015;
wire n_1972;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_2202;
wire n_2072;
wire n_306;
wire n_92;
wire n_203;
wire n_436;
wire n_150;
wire n_324;
wire n_2087;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_111;
wire n_274;
wire n_967;
wire n_1083;
wire n_2161;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_2155;
wire n_615;
wire n_1139;
wire n_76;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_159;
wire n_2172;
wire n_892;
wire n_1880;
wire n_959;
wire n_2257;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_2219;
wire n_1855;
wire n_2100;
wire n_144;
wire n_990;
wire n_1623;
wire n_1903;
wire n_867;
wire n_2147;
wire n_1226;
wire n_2224;
wire n_944;
wire n_749;
wire n_1932;
wire n_1780;
wire n_1970;
wire n_1920;
wire n_2083;
wire n_815;
wire n_542;
wire n_2167;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_2273;
wire n_1433;
wire n_1911;
wire n_1825;
wire n_1908;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_2066;
wire n_964;
wire n_1627;
wire n_2220;
wire n_382;
wire n_489;
wire n_80;
wire n_2274;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_1914;
wire n_155;
wire n_2253;
wire n_934;
wire n_2213;
wire n_1447;
wire n_1220;
wire n_356;
wire n_2019;
wire n_698;
wire n_2130;
wire n_1674;
wire n_2021;
wire n_2025;
wire n_2160;
wire n_1992;
wire n_124;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_2142;
wire n_1633;
wire n_404;
wire n_172;
wire n_1913;
wire n_2069;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_2261;
wire n_1455;
wire n_299;
wire n_836;
wire n_2223;
wire n_1279;
wire n_2144;
wire n_564;
wire n_133;
wire n_66;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_2262;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_2120;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_2041;
wire n_2113;
wire n_1933;
wire n_1651;
wire n_85;
wire n_130;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_2168;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_138;
wire n_162;
wire n_264;
wire n_441;
wire n_1951;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_73;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_2132;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_1943;
wire n_194;
wire n_1802;
wire n_2178;
wire n_2112;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_145;
wire n_2146;
wire n_1868;
wire n_59;
wire n_1501;
wire n_2241;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_2099;
wire n_487;
wire n_1518;
wire n_1456;
wire n_90;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2129;
wire n_855;
wire n_158;
wire n_808;
wire n_1365;
wire n_553;
wire n_2059;
wire n_1439;
wire n_814;
wire n_578;
wire n_2074;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_2122;
wire n_120;
wire n_320;
wire n_1414;
wire n_1134;
wire n_2067;
wire n_1484;
wire n_1901;
wire n_647;
wire n_2055;
wire n_2027;
wire n_1423;
wire n_2117;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_1939;
wire n_2242;
wire n_1906;
wire n_529;
wire n_1899;
wire n_2195;
wire n_502;
wire n_2194;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_2159;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_2267;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_2102;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_2023;
wire n_1278;
wire n_707;
wire n_129;
wire n_126;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_2075;
wire n_1945;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_2031;
wire n_2118;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_2225;
wire n_986;
wire n_1104;
wire n_1963;
wire n_729;
wire n_887;
wire n_2057;
wire n_2218;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_2125;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_2184;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_2254;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_2033;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_2217;
wire n_221;
wire n_321;
wire n_86;
wire n_2226;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_2214;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_2256;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_2190;
wire n_1478;
wire n_1883;
wire n_1969;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_84;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1927;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_70;
wire n_343;
wire n_1222;
wire n_1844;
wire n_2283;
wire n_582;
wire n_1957;
wire n_1953;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_1919;
wire n_534;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_2266;
wire n_560;
wire n_890;
wire n_842;
wire n_148;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1907;
wire n_1793;
wire n_61;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1975;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_2119;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1990;
wire n_1372;
wire n_476;
wire n_832;
wire n_55;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_2008;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_2127;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_2211;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_2071;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_2082;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_2140;
wire n_873;
wire n_1301;
wire n_1748;
wire n_2157;
wire n_1966;
wire n_1243;
wire n_2171;
wire n_1400;
wire n_342;
wire n_2035;
wire n_1466;
wire n_1527;
wire n_1513;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_2128;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1993;
wire n_1545;
wire n_134;
wire n_1257;
wire n_1480;
wire n_1954;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_157;
wire n_2137;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_2265;
wire n_687;
wire n_797;
wire n_2026;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_2106;
wire n_97;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_2272;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_2091;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_1929;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_295;
wire n_1658;
wire n_190;
wire n_2249;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_64;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1997;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1733;
wire n_1856;
wire n_2016;
wire n_1524;
wire n_1118;
wire n_943;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_71;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1984;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_1971;
wire n_586;
wire n_1324;
wire n_1429;
wire n_2064;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_2022;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_1987;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_87;
wire n_714;
wire n_2170;
wire n_790;
wire n_2244;
wire n_2143;
wire n_354;
wire n_140;
wire n_725;
wire n_1577;
wire n_151;
wire n_1448;
wire n_2198;
wire n_1009;
wire n_230;
wire n_1133;
wire n_154;
wire n_883;
wire n_142;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_2279;
wire n_594;
wire n_2222;
wire n_1995;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_2076;
wire n_2133;
wire n_2203;
wire n_833;
wire n_1426;
wire n_2250;
wire n_2247;
wire n_2230;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_75;
wire n_2001;
wire n_1047;
wire n_95;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_2158;
wire n_152;
wire n_169;
wire n_106;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_2173;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_2070;
wire n_2136;
wire n_426;
wire n_433;
wire n_398;
wire n_62;
wire n_210;
wire n_1090;
wire n_1367;
wire n_2044;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_128;
wire n_224;
wire n_82;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_2020;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1976;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_1958;
wire n_467;
wire n_2177;
wire n_1511;
wire n_1422;
wire n_1965;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_81;
wire n_538;
wire n_1517;
wire n_2036;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_2003;
wire n_2210;
wire n_1307;
wire n_1128;
wire n_2053;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_141;
wire n_846;
wire n_1398;
wire n_1921;
wire n_1356;
wire n_1341;
wire n_2234;
wire n_1504;
wire n_1955;
wire n_2110;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_56;
wire n_60;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_89;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_1948;
wire n_74;
wire n_810;
wire n_1290;
wire n_181;
wire n_1959;
wire n_617;
wire n_543;
wire n_1362;
wire n_2121;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_1960;
wire n_2068;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1968;
wire n_107;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_2196;
wire n_1038;
wire n_1978;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_1940;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_58;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_2007;
wire n_526;
wire n_1994;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_125;
wire n_1973;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_161;
wire n_1814;
wire n_532;
wire n_2154;
wire n_2236;
wire n_1789;
wire n_763;
wire n_1986;
wire n_2174;
wire n_99;
wire n_540;
wire n_216;
wire n_692;
wire n_2054;
wire n_1857;
wire n_984;
wire n_1687;
wire n_2073;
wire n_223;
wire n_2150;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_2046;
wire n_1816;
wire n_1910;
wire n_1756;
wire n_1606;
wire n_2189;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_2093;
wire n_2018;
wire n_1772;
wire n_67;
wire n_1014;
wire n_724;
wire n_2204;
wire n_1427;
wire n_1481;
wire n_2040;
wire n_493;
wire n_1311;
wire n_2199;
wire n_1956;
wire n_1589;
wire n_114;
wire n_2151;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_2231;
wire n_697;
wire n_622;
wire n_1626;
wire n_1962;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_2114;
wire n_1175;
wire n_132;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2180;
wire n_580;
wire n_1579;
wire n_494;
wire n_2181;
wire n_434;
wire n_2014;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_2276;
wire n_1805;
wire n_2282;
wire n_981;
wire n_2141;
wire n_1110;
wire n_1758;
wire n_2270;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_2251;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_2010;
wire n_1054;
wire n_508;
wire n_118;
wire n_121;
wire n_1679;
wire n_2126;
wire n_1952;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_116;
wire n_653;
wire n_1445;
wire n_1317;
wire n_2050;
wire n_2197;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_160;
wire n_119;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_1980;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_1998;
wire n_2165;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_2169;
wire n_341;
wire n_1270;
wire n_109;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_2028;
wire n_919;
wire n_1663;
wire n_2092;
wire n_2175;
wire n_1625;
wire n_2086;
wire n_1926;
wire n_318;
wire n_1458;
wire n_244;
wire n_103;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_2176;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_139;
wire n_1922;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_2138;
wire n_2065;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_1930;
wire n_765;
wire n_1809;
wire n_1904;
wire n_1843;
wire n_122;
wire n_2000;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_2096;
wire n_2186;
wire n_1530;
wire n_2215;
wire n_631;
wire n_399;
wire n_1170;
wire n_2258;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1937;
wire n_2012;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_2039;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_2212;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_2268;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_2252;
wire n_2111;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_153;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_2024;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_2103;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_115;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_2062;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_2153;
wire n_1510;
wire n_2139;
wire n_1099;
wire n_839;
wire n_79;
wire n_1754;
wire n_759;
wire n_567;
wire n_91;
wire n_240;
wire n_369;
wire n_1727;
wire n_2235;
wire n_1991;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_2260;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_1902;
wire n_997;
wire n_635;
wire n_2206;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_2034;
wire n_1845;
wire n_1934;
wire n_2101;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_2104;
wire n_1265;
wire n_1576;
wire n_2105;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_2088;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_88;
wire n_2005;
wire n_2048;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_2108;
wire n_1039;
wire n_2246;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_2191;
wire n_1497;
wire n_1866;
wire n_2056;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1941;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_1915;
wire n_723;
wire n_1393;
wire n_2240;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_2085;
wire n_1686;
wire n_1964;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_2188;
wire n_1982;
wire n_2097;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_2193;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1983;
wire n_1041;
wire n_2115;
wire n_993;
wire n_1862;
wire n_948;
wire n_2017;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1923;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_1946;
wire n_2148;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_2051;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_68;
wire n_1896;
wire n_2164;
wire n_1732;
wire n_415;
wire n_1967;
wire n_2179;
wire n_63;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_2052;
wire n_537;
wire n_1063;
wire n_991;
wire n_2183;
wire n_2205;
wire n_83;
wire n_2275;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1799;
wire n_1707;
wire n_2080;
wire n_2058;
wire n_1126;
wire n_2029;
wire n_195;
wire n_1846;
wire n_1912;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_110;
wire n_304;
wire n_1639;
wire n_583;
wire n_2209;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_1928;
wire n_98;
wire n_946;
wire n_757;
wire n_2047;
wire n_375;
wire n_113;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_2269;
wire n_472;
wire n_937;
wire n_1474;
wire n_2081;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_156;
wire n_174;
wire n_275;
wire n_100;
wire n_1794;
wire n_1375;
wire n_147;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_2229;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_105;
wire n_1051;
wire n_719;
wire n_131;
wire n_1102;
wire n_263;
wire n_360;
wire n_2255;
wire n_1129;
wire n_1252;
wire n_2239;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_101;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1905;
wire n_1569;
wire n_289;
wire n_112;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_2063;
wire n_177;
wire n_1925;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_2079;
wire n_1228;
wire n_2152;
wire n_1931;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_2259;
wire n_849;
wire n_2095;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_1989;
wire n_447;
wire n_1421;
wire n_2208;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_2228;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_1981;
wire n_2037;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_127;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_2089;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g55 ( 
.A(n_8),
.Y(n_55)
);

CKINVDCx5p33_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx5p33_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

CKINVDCx5p33_ASAP7_75t_R g59 ( 
.A(n_12),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g60 ( 
.A(n_14),
.Y(n_60)
);

CKINVDCx5p33_ASAP7_75t_R g61 ( 
.A(n_25),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

CKINVDCx5p33_ASAP7_75t_R g63 ( 
.A(n_22),
.Y(n_63)
);

CKINVDCx5p33_ASAP7_75t_R g64 ( 
.A(n_33),
.Y(n_64)
);

CKINVDCx5p33_ASAP7_75t_R g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_24),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g70 ( 
.A(n_41),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_44),
.Y(n_73)
);

CKINVDCx5p33_ASAP7_75t_R g74 ( 
.A(n_39),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_40),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_32),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_25),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_23),
.Y(n_79)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_17),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_36),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_4),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g83 ( 
.A(n_9),
.Y(n_83)
);

BUFx8_ASAP7_75t_SL g84 ( 
.A(n_22),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_44),
.Y(n_85)
);

CKINVDCx5p33_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_50),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_40),
.Y(n_88)
);

CKINVDCx5p33_ASAP7_75t_R g89 ( 
.A(n_5),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_6),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_6),
.Y(n_91)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_52),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_9),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_47),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_20),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_21),
.Y(n_98)
);

CKINVDCx5p33_ASAP7_75t_R g99 ( 
.A(n_45),
.Y(n_99)
);

CKINVDCx5p33_ASAP7_75t_R g100 ( 
.A(n_3),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_14),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_19),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_20),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_8),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_10),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_12),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_37),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_68),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_62),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_68),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_68),
.Y(n_116)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_66),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_71),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_60),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_71),
.Y(n_121)
);

CKINVDCx5p33_ASAP7_75t_R g122 ( 
.A(n_84),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_60),
.Y(n_123)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_87),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_87),
.Y(n_125)
);

INVxp67_ASAP7_75t_SL g126 ( 
.A(n_58),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_94),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_94),
.Y(n_128)
);

AND2x4_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_66),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_92),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_111),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_111),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_115),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_114),
.A2(n_69),
.B1(n_95),
.B2(n_107),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_69),
.B1(n_112),
.B2(n_123),
.Y(n_144)
);

AND2x4_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_66),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_119),
.A2(n_123),
.B1(n_114),
.B2(n_112),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_126),
.A2(n_95),
.B1(n_97),
.B2(n_107),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

CKINVDCx5p33_ASAP7_75t_R g149 ( 
.A(n_119),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_117),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_117),
.Y(n_153)
);

AND2x6_ASAP7_75t_L g154 ( 
.A(n_124),
.B(n_66),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_117),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_125),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_125),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_110),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_127),
.Y(n_160)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_150),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_146),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_92),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_141),
.B(n_127),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_141),
.B(n_127),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_128),
.B1(n_92),
.B2(n_126),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_147),
.A2(n_128),
.B1(n_97),
.B2(n_65),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_150),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_150),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_157),
.B(n_128),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_150),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_110),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_150),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_150),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_132),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_158),
.B(n_153),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_157),
.B(n_131),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_142),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_142),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_146),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_157),
.B(n_131),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_132),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_132),
.Y(n_197)
);

AND2x4_ASAP7_75t_L g198 ( 
.A(n_131),
.B(n_97),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_110),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_147),
.A2(n_143),
.B1(n_144),
.B2(n_158),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_153),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_134),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_155),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_151),
.B(n_113),
.Y(n_204)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_142),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g206 ( 
.A(n_155),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

NAND2xp33_ASAP7_75t_SL g208 ( 
.A(n_131),
.B(n_59),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_134),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g210 ( 
.A(n_155),
.Y(n_210)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_153),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_151),
.B(n_113),
.Y(n_212)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_131),
.B(n_113),
.Y(n_213)
);

INVx3_ASAP7_75t_L g214 ( 
.A(n_153),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_142),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_134),
.Y(n_217)
);

INVx3_ASAP7_75t_L g218 ( 
.A(n_153),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_135),
.Y(n_219)
);

OAI21x1_ASAP7_75t_L g220 ( 
.A1(n_130),
.A2(n_120),
.B(n_118),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_142),
.B(n_72),
.Y(n_221)
);

AND2x4_ASAP7_75t_L g222 ( 
.A(n_129),
.B(n_58),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_135),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_142),
.B(n_72),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_142),
.Y(n_225)
);

AND2x4_ASAP7_75t_L g226 ( 
.A(n_129),
.B(n_67),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_151),
.B(n_152),
.Y(n_227)
);

AND2x6_ASAP7_75t_L g228 ( 
.A(n_129),
.B(n_67),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_129),
.B(n_145),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_142),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_227),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_166),
.A2(n_144),
.B1(n_143),
.B2(n_129),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_227),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_166),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_220),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_227),
.Y(n_236)
);

INVx4_ASAP7_75t_L g237 ( 
.A(n_173),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_182),
.B(n_139),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_220),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_178),
.B(n_129),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_187),
.Y(n_241)
);

AND2x2_ASAP7_75t_SL g242 ( 
.A(n_166),
.B(n_129),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_195),
.Y(n_243)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_229),
.Y(n_244)
);

INVx2_ASAP7_75t_SL g245 ( 
.A(n_182),
.Y(n_245)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_178),
.B(n_129),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

INVx3_ASAP7_75t_L g248 ( 
.A(n_195),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_178),
.B(n_151),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_187),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_195),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_220),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_203),
.B(n_210),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_178),
.B(n_152),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

AOI22xp33_ASAP7_75t_L g256 ( 
.A1(n_200),
.A2(n_144),
.B1(n_145),
.B2(n_154),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

CKINVDCx6p67_ASAP7_75t_R g258 ( 
.A(n_228),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_189),
.B(n_145),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_203),
.B(n_139),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_187),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_189),
.B(n_152),
.Y(n_262)
);

INVx6_ASAP7_75t_L g263 ( 
.A(n_195),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_187),
.Y(n_264)
);

AND2x4_ASAP7_75t_L g265 ( 
.A(n_229),
.B(n_145),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_192),
.Y(n_266)
);

CKINVDCx11_ASAP7_75t_R g267 ( 
.A(n_163),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

AND2x4_ASAP7_75t_L g269 ( 
.A(n_229),
.B(n_145),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_192),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_182),
.B(n_139),
.Y(n_271)
);

AND2x6_ASAP7_75t_L g272 ( 
.A(n_198),
.B(n_145),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_195),
.Y(n_273)
);

AND2x6_ASAP7_75t_L g274 ( 
.A(n_198),
.B(n_145),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_220),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_192),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_189),
.B(n_152),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_203),
.B(n_139),
.Y(n_278)
);

AND2x6_ASAP7_75t_L g279 ( 
.A(n_198),
.B(n_145),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_210),
.B(n_139),
.Y(n_280)
);

AND2x6_ASAP7_75t_L g281 ( 
.A(n_198),
.B(n_160),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_192),
.Y(n_282)
);

INVx4_ASAP7_75t_L g283 ( 
.A(n_173),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_189),
.B(n_194),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_200),
.B(n_140),
.Y(n_285)
);

AND2x4_ASAP7_75t_L g286 ( 
.A(n_229),
.B(n_156),
.Y(n_286)
);

OR2x6_ASAP7_75t_L g287 ( 
.A(n_200),
.B(n_140),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_195),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_210),
.B(n_140),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_171),
.A2(n_154),
.B1(n_160),
.B2(n_156),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_196),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_196),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_196),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_182),
.Y(n_294)
);

AND2x6_ASAP7_75t_L g295 ( 
.A(n_198),
.B(n_160),
.Y(n_295)
);

INVx2_ASAP7_75t_SL g296 ( 
.A(n_182),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_194),
.B(n_213),
.Y(n_297)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_195),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_194),
.B(n_140),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_171),
.A2(n_154),
.B1(n_160),
.B2(n_156),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g301 ( 
.A1(n_171),
.A2(n_154),
.B1(n_140),
.B2(n_156),
.Y(n_301)
);

AND2x6_ASAP7_75t_L g302 ( 
.A(n_198),
.B(n_135),
.Y(n_302)
);

BUFx4f_ASAP7_75t_L g303 ( 
.A(n_228),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_L g304 ( 
.A1(n_208),
.A2(n_154),
.B1(n_84),
.B2(n_142),
.Y(n_304)
);

BUFx10_ASAP7_75t_L g305 ( 
.A(n_198),
.Y(n_305)
);

NAND2xp33_ASAP7_75t_L g306 ( 
.A(n_195),
.B(n_154),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_196),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_194),
.B(n_146),
.Y(n_308)
);

INVx4_ASAP7_75t_L g309 ( 
.A(n_173),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_193),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_206),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_206),
.B(n_172),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_202),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_202),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g315 ( 
.A(n_213),
.B(n_159),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_163),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_202),
.Y(n_317)
);

BUFx4f_ASAP7_75t_L g318 ( 
.A(n_228),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_202),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_207),
.Y(n_320)
);

INVx4_ASAP7_75t_L g321 ( 
.A(n_173),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_207),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_207),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_207),
.Y(n_324)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_195),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g326 ( 
.A(n_213),
.B(n_159),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_206),
.B(n_149),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g328 ( 
.A(n_172),
.Y(n_328)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_213),
.B(n_159),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_206),
.B(n_59),
.Y(n_330)
);

AND2x6_ASAP7_75t_L g331 ( 
.A(n_198),
.B(n_172),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_209),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_209),
.Y(n_333)
);

AND2x4_ASAP7_75t_L g334 ( 
.A(n_206),
.B(n_154),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_208),
.B(n_149),
.Y(n_335)
);

BUFx6f_ASAP7_75t_SL g336 ( 
.A(n_228),
.Y(n_336)
);

INVx5_ASAP7_75t_L g337 ( 
.A(n_173),
.Y(n_337)
);

INVx2_ASAP7_75t_L g338 ( 
.A(n_209),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_209),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_217),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_228),
.A2(n_154),
.B1(n_142),
.B2(n_77),
.Y(n_341)
);

OR2x6_ASAP7_75t_L g342 ( 
.A(n_222),
.B(n_116),
.Y(n_342)
);

BUFx4f_ASAP7_75t_L g343 ( 
.A(n_228),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_217),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_217),
.Y(n_345)
);

INVx4_ASAP7_75t_L g346 ( 
.A(n_173),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_199),
.B(n_135),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_217),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_222),
.B(n_61),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_223),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_193),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_201),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_193),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g354 ( 
.A(n_299),
.B(n_201),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_253),
.B(n_222),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g356 ( 
.A(n_242),
.B(n_201),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_276),
.Y(n_357)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_276),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_327),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_276),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_312),
.A2(n_228),
.B1(n_188),
.B2(n_226),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_242),
.B(n_245),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_331),
.A2(n_228),
.B1(n_188),
.B2(n_226),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_241),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

INVx2_ASAP7_75t_SL g366 ( 
.A(n_305),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_231),
.B(n_222),
.Y(n_367)
);

NAND2xp33_ASAP7_75t_L g368 ( 
.A(n_331),
.B(n_173),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_242),
.B(n_201),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_231),
.B(n_222),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_233),
.B(n_222),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_241),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_292),
.Y(n_373)
);

OAI21xp33_ASAP7_75t_L g374 ( 
.A1(n_260),
.A2(n_278),
.B(n_284),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_233),
.B(n_222),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_292),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_245),
.B(n_201),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_250),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_250),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_261),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_236),
.B(n_222),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_236),
.B(n_297),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_331),
.A2(n_285),
.B1(n_287),
.B2(n_234),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_296),
.B(n_201),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_240),
.B(n_226),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_285),
.B(n_188),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_261),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_264),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_240),
.B(n_226),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_246),
.B(n_226),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_L g392 ( 
.A(n_335),
.B(n_226),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_296),
.A2(n_218),
.B1(n_214),
.B2(n_211),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_331),
.A2(n_228),
.B1(n_226),
.B2(n_212),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_294),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_246),
.B(n_259),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_259),
.B(n_226),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_294),
.B(n_280),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_264),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_305),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_289),
.B(n_201),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_249),
.B(n_199),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_266),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_254),
.B(n_199),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_315),
.B(n_169),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_315),
.B(n_169),
.Y(n_406)
);

A2O1A1Ixp33_ASAP7_75t_L g407 ( 
.A1(n_262),
.A2(n_212),
.B(n_169),
.C(n_170),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_326),
.B(n_170),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_305),
.B(n_201),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_326),
.B(n_170),
.Y(n_410)
);

NOR2xp67_ASAP7_75t_L g411 ( 
.A(n_266),
.B(n_211),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_329),
.B(n_165),
.Y(n_412)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_331),
.A2(n_228),
.B1(n_221),
.B2(n_224),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_329),
.B(n_165),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_314),
.Y(n_415)
);

INVxp67_ASAP7_75t_L g416 ( 
.A(n_308),
.Y(n_416)
);

INVx2_ASAP7_75t_SL g417 ( 
.A(n_305),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_314),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_277),
.B(n_165),
.Y(n_419)
);

NAND2xp33_ASAP7_75t_L g420 ( 
.A(n_331),
.B(n_173),
.Y(n_420)
);

A2O1A1Ixp33_ASAP7_75t_L g421 ( 
.A1(n_256),
.A2(n_212),
.B(n_223),
.C(n_219),
.Y(n_421)
);

INVx2_ASAP7_75t_SL g422 ( 
.A(n_303),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_286),
.B(n_165),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_286),
.B(n_168),
.Y(n_424)
);

INVx8_ASAP7_75t_L g425 ( 
.A(n_281),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_270),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_323),
.Y(n_427)
);

AND2x6_ASAP7_75t_SL g428 ( 
.A(n_287),
.B(n_77),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_331),
.A2(n_228),
.B1(n_223),
.B2(n_197),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_301),
.B(n_201),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_303),
.B(n_201),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_308),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_303),
.B(n_201),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_286),
.B(n_168),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_286),
.B(n_168),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_SL g436 ( 
.A(n_287),
.B(n_228),
.Y(n_436)
);

BUFx6f_ASAP7_75t_L g437 ( 
.A(n_243),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_303),
.B(n_201),
.Y(n_438)
);

INVxp33_ASAP7_75t_L g439 ( 
.A(n_267),
.Y(n_439)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_232),
.B(n_223),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_244),
.B(n_168),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_331),
.B(n_181),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g443 ( 
.A1(n_287),
.A2(n_228),
.B1(n_197),
.B2(n_219),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_265),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_R g445 ( 
.A(n_336),
.B(n_181),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_270),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_310),
.B(n_351),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_323),
.Y(n_448)
);

BUFx6f_ASAP7_75t_L g449 ( 
.A(n_243),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_282),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_318),
.B(n_211),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_287),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_282),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_244),
.B(n_181),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_318),
.B(n_343),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g456 ( 
.A(n_265),
.B(n_183),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_244),
.B(n_181),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_323),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_265),
.B(n_185),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_311),
.B(n_185),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g461 ( 
.A(n_318),
.B(n_211),
.Y(n_461)
);

INVx4_ASAP7_75t_L g462 ( 
.A(n_258),
.Y(n_462)
);

NAND2xp33_ASAP7_75t_L g463 ( 
.A(n_243),
.B(n_173),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_291),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_291),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_265),
.B(n_185),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_293),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_269),
.B(n_185),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_269),
.B(n_176),
.Y(n_469)
);

AND2x4_ASAP7_75t_L g470 ( 
.A(n_269),
.B(n_228),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_293),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_269),
.B(n_183),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_359),
.B(n_272),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_444),
.B(n_470),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_353),
.B(n_272),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_357),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_425),
.Y(n_478)
);

INVx1_ASAP7_75t_SL g479 ( 
.A(n_447),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_382),
.B(n_272),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_416),
.B(n_272),
.Y(n_481)
);

NOR2xp67_ASAP7_75t_L g482 ( 
.A(n_432),
.B(n_395),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_364),
.Y(n_483)
);

AOI22xp33_ASAP7_75t_L g484 ( 
.A1(n_392),
.A2(n_274),
.B1(n_272),
.B2(n_279),
.Y(n_484)
);

OR2x4_ASAP7_75t_L g485 ( 
.A(n_441),
.B(n_459),
.Y(n_485)
);

INVx2_ASAP7_75t_SL g486 ( 
.A(n_425),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g487 ( 
.A(n_456),
.B(n_342),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_444),
.Y(n_488)
);

INVx2_ASAP7_75t_SL g489 ( 
.A(n_425),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_470),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_342),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_372),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_372),
.Y(n_493)
);

INVx3_ASAP7_75t_SL g494 ( 
.A(n_470),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_472),
.B(n_272),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_357),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_378),
.Y(n_497)
);

AND2x2_ASAP7_75t_L g498 ( 
.A(n_472),
.B(n_342),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

BUFx3_ASAP7_75t_L g500 ( 
.A(n_470),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_437),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_405),
.B(n_272),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_428),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_406),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_429),
.B(n_243),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_408),
.B(n_410),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_396),
.B(n_342),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_429),
.B(n_243),
.Y(n_508)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_466),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_358),
.Y(n_510)
);

BUFx3_ASAP7_75t_L g511 ( 
.A(n_437),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_387),
.A2(n_295),
.B1(n_281),
.B2(n_302),
.Y(n_512)
);

INVx2_ASAP7_75t_SL g513 ( 
.A(n_445),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_378),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_379),
.Y(n_515)
);

BUFx8_ASAP7_75t_L g516 ( 
.A(n_440),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_379),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_398),
.B(n_330),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_394),
.A2(n_316),
.B1(n_290),
.B2(n_300),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_355),
.B(n_402),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_380),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_358),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_404),
.B(n_440),
.Y(n_523)
);

BUFx3_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_367),
.B(n_272),
.Y(n_525)
);

BUFx2_ASAP7_75t_L g526 ( 
.A(n_442),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_380),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_370),
.B(n_274),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_SL g529 ( 
.A1(n_394),
.A2(n_290),
.B1(n_300),
.B2(n_304),
.Y(n_529)
);

INVx3_ASAP7_75t_SL g530 ( 
.A(n_452),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_428),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_371),
.B(n_274),
.Y(n_532)
);

OAI21xp33_ASAP7_75t_L g533 ( 
.A1(n_374),
.A2(n_342),
.B(n_349),
.Y(n_533)
);

NOR2xp67_ASAP7_75t_L g534 ( 
.A(n_384),
.B(n_238),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_437),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_374),
.B(n_243),
.Y(n_536)
);

AND2x4_ASAP7_75t_L g537 ( 
.A(n_462),
.B(n_334),
.Y(n_537)
);

INVx5_ASAP7_75t_L g538 ( 
.A(n_437),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_388),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_388),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_SL g541 ( 
.A(n_443),
.B(n_268),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_L g542 ( 
.A1(n_361),
.A2(n_318),
.B1(n_343),
.B2(n_258),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_389),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g544 ( 
.A(n_375),
.B(n_274),
.Y(n_544)
);

OR2x6_ASAP7_75t_L g545 ( 
.A(n_462),
.B(n_334),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_381),
.B(n_274),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_468),
.B(n_271),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_389),
.B(n_399),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_471),
.B(n_399),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_403),
.B(n_274),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_360),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_403),
.B(n_274),
.Y(n_552)
);

AOI221xp5_ASAP7_75t_SL g553 ( 
.A1(n_421),
.A2(n_347),
.B1(n_350),
.B2(n_340),
.C(n_322),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_426),
.B(n_471),
.Y(n_554)
);

INVx4_ASAP7_75t_L g555 ( 
.A(n_462),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_366),
.Y(n_556)
);

NAND2x1p5_ASAP7_75t_L g557 ( 
.A(n_366),
.B(n_334),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_L g558 ( 
.A(n_426),
.B(n_274),
.Y(n_558)
);

INVx5_ASAP7_75t_L g559 ( 
.A(n_449),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_446),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_446),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_360),
.Y(n_562)
);

INVx4_ASAP7_75t_L g563 ( 
.A(n_449),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_L g564 ( 
.A(n_450),
.B(n_279),
.Y(n_564)
);

HB1xp67_ASAP7_75t_L g565 ( 
.A(n_423),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_365),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_443),
.B(n_268),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_365),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_450),
.B(n_279),
.Y(n_569)
);

AO22x1_ASAP7_75t_L g570 ( 
.A1(n_439),
.A2(n_295),
.B1(n_281),
.B2(n_302),
.Y(n_570)
);

INVx4_ASAP7_75t_L g571 ( 
.A(n_449),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_384),
.B(n_436),
.Y(n_572)
);

AND3x1_ASAP7_75t_SL g573 ( 
.A(n_453),
.B(n_101),
.C(n_90),
.Y(n_573)
);

INVx5_ASAP7_75t_L g574 ( 
.A(n_449),
.Y(n_574)
);

AO22x1_ASAP7_75t_L g575 ( 
.A1(n_452),
.A2(n_295),
.B1(n_281),
.B2(n_302),
.Y(n_575)
);

AND3x2_ASAP7_75t_SL g576 ( 
.A(n_368),
.B(n_333),
.C(n_324),
.Y(n_576)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_362),
.A2(n_295),
.B1(n_281),
.B2(n_302),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_453),
.Y(n_578)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_368),
.A2(n_295),
.B1(n_281),
.B2(n_302),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_373),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_463),
.A2(n_283),
.B(n_237),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

NAND2x1p5_ASAP7_75t_L g583 ( 
.A(n_400),
.B(n_334),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_449),
.B(n_268),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_397),
.B(n_324),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_361),
.B(n_413),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_373),
.Y(n_587)
);

OAI21xp5_ASAP7_75t_L g588 ( 
.A1(n_407),
.A2(n_313),
.B(n_307),
.Y(n_588)
);

OR2x2_ASAP7_75t_L g589 ( 
.A(n_386),
.B(n_324),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_376),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_422),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g592 ( 
.A(n_469),
.B(n_333),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_467),
.B(n_279),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_467),
.B(n_279),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_464),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_465),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_465),
.Y(n_597)
);

AND2x2_ASAP7_75t_L g598 ( 
.A(n_390),
.B(n_333),
.Y(n_598)
);

BUFx2_ASAP7_75t_L g599 ( 
.A(n_391),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_376),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_383),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_412),
.B(n_279),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_383),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_L g604 ( 
.A(n_400),
.B(n_281),
.Y(n_604)
);

OR2x6_ASAP7_75t_L g605 ( 
.A(n_356),
.B(n_338),
.Y(n_605)
);

OAI22xp5_ASAP7_75t_L g606 ( 
.A1(n_363),
.A2(n_343),
.B1(n_350),
.B2(n_340),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_415),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_415),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_418),
.Y(n_609)
);

INVx4_ASAP7_75t_L g610 ( 
.A(n_417),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_414),
.B(n_279),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_424),
.B(n_279),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_434),
.B(n_281),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_417),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_363),
.A2(n_336),
.B1(n_295),
.B2(n_302),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_435),
.A2(n_343),
.B1(n_419),
.B2(n_454),
.Y(n_616)
);

INVx2_ASAP7_75t_SL g617 ( 
.A(n_422),
.Y(n_617)
);

NOR2x1_ASAP7_75t_R g618 ( 
.A(n_369),
.B(n_61),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_418),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_457),
.B(n_338),
.Y(n_620)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_420),
.A2(n_295),
.B1(n_302),
.B2(n_336),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_R g622 ( 
.A(n_420),
.B(n_336),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_427),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_427),
.B(n_338),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_455),
.B(n_344),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_523),
.B(n_460),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_520),
.B(n_448),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_506),
.B(n_448),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_476),
.B(n_458),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_622),
.B(n_615),
.Y(n_630)
);

NAND2xp33_ASAP7_75t_SL g631 ( 
.A(n_622),
.B(n_529),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_599),
.B(n_458),
.Y(n_632)
);

NAND2xp33_ASAP7_75t_SL g633 ( 
.A(n_606),
.B(n_268),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_599),
.B(n_344),
.Y(n_634)
);

NAND2xp33_ASAP7_75t_SL g635 ( 
.A(n_519),
.B(n_268),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_SL g636 ( 
.A(n_548),
.B(n_268),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_SL g637 ( 
.A(n_549),
.B(n_237),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_482),
.B(n_344),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_504),
.B(n_348),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_592),
.B(n_547),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_480),
.B(n_348),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_SL g642 ( 
.A(n_512),
.B(n_348),
.Y(n_642)
);

AND2x4_ASAP7_75t_L g643 ( 
.A(n_500),
.B(n_411),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_485),
.B(n_63),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_479),
.B(n_307),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_509),
.B(n_411),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_SL g647 ( 
.A(n_589),
.B(n_313),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_589),
.B(n_317),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_473),
.B(n_317),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_585),
.B(n_319),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_585),
.B(n_319),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_598),
.B(n_320),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_SL g653 ( 
.A(n_494),
.B(n_237),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_598),
.B(n_320),
.Y(n_654)
);

NAND2xp33_ASAP7_75t_SL g655 ( 
.A(n_494),
.B(n_237),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_556),
.B(n_322),
.Y(n_656)
);

NAND2xp5_ASAP7_75t_L g657 ( 
.A(n_565),
.B(n_332),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_556),
.B(n_332),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_579),
.B(n_339),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_SL g660 ( 
.A(n_538),
.B(n_339),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_538),
.B(n_345),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_538),
.B(n_345),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_538),
.B(n_337),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_475),
.B(n_295),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_483),
.B(n_492),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_SL g666 ( 
.A(n_554),
.B(n_283),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_538),
.B(n_337),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_559),
.B(n_337),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_SL g669 ( 
.A(n_484),
.B(n_283),
.Y(n_669)
);

AND2x4_ASAP7_75t_L g670 ( 
.A(n_500),
.B(n_409),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_559),
.B(n_337),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_SL g672 ( 
.A(n_559),
.B(n_337),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_493),
.B(n_183),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_SL g674 ( 
.A(n_559),
.B(n_337),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_530),
.B(n_204),
.Y(n_675)
);

NAND2xp33_ASAP7_75t_SL g676 ( 
.A(n_530),
.B(n_283),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_559),
.B(n_401),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_574),
.B(n_309),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_SL g679 ( 
.A(n_574),
.B(n_309),
.Y(n_679)
);

NAND2xp33_ASAP7_75t_SL g680 ( 
.A(n_487),
.B(n_309),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_574),
.B(n_309),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_574),
.B(n_321),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_574),
.B(n_321),
.Y(n_683)
);

NAND2xp33_ASAP7_75t_SL g684 ( 
.A(n_501),
.B(n_535),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_502),
.B(n_321),
.Y(n_685)
);

AND2x4_ASAP7_75t_L g686 ( 
.A(n_474),
.B(n_302),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_537),
.B(n_321),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_SL g688 ( 
.A(n_501),
.B(n_346),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_537),
.B(n_346),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_537),
.B(n_346),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_577),
.B(n_346),
.Y(n_691)
);

AND3x1_ASAP7_75t_L g692 ( 
.A(n_518),
.B(n_101),
.C(n_90),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_534),
.B(n_354),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_SL g694 ( 
.A(n_507),
.B(n_377),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_497),
.B(n_197),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_SL g696 ( 
.A(n_501),
.B(n_463),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_507),
.B(n_385),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_526),
.B(n_248),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_526),
.B(n_248),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_620),
.B(n_248),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_613),
.B(n_248),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_602),
.B(n_251),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_611),
.B(n_251),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_SL g704 ( 
.A(n_501),
.B(n_431),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_550),
.B(n_552),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_474),
.B(n_251),
.Y(n_706)
);

NAND2xp33_ASAP7_75t_SL g707 ( 
.A(n_501),
.B(n_433),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_514),
.B(n_219),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_558),
.B(n_564),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_569),
.B(n_251),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_593),
.B(n_255),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_515),
.B(n_204),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_517),
.B(n_204),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_521),
.B(n_228),
.Y(n_714)
);

NAND2xp33_ASAP7_75t_SL g715 ( 
.A(n_535),
.B(n_542),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_527),
.B(n_63),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_594),
.B(n_255),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_539),
.B(n_64),
.Y(n_718)
);

NAND2xp5_ASAP7_75t_SL g719 ( 
.A(n_610),
.B(n_255),
.Y(n_719)
);

NAND2xp33_ASAP7_75t_SL g720 ( 
.A(n_535),
.B(n_438),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_610),
.B(n_255),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_474),
.B(n_257),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_610),
.B(n_503),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_540),
.B(n_64),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_604),
.B(n_341),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_543),
.B(n_65),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_560),
.B(n_70),
.Y(n_727)
);

NAND2xp33_ASAP7_75t_SL g728 ( 
.A(n_487),
.B(n_451),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_503),
.B(n_257),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_531),
.B(n_257),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_SL g731 ( 
.A(n_491),
.B(n_461),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_561),
.B(n_70),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_490),
.B(n_73),
.Y(n_733)
);

NAND2xp33_ASAP7_75t_SL g734 ( 
.A(n_491),
.B(n_257),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_SL g735 ( 
.A(n_498),
.B(n_273),
.Y(n_735)
);

NAND2xp33_ASAP7_75t_SL g736 ( 
.A(n_498),
.B(n_273),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_531),
.B(n_273),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_SL g738 ( 
.A(n_495),
.B(n_273),
.Y(n_738)
);

NAND2xp33_ASAP7_75t_SL g739 ( 
.A(n_555),
.B(n_288),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_525),
.B(n_288),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_528),
.B(n_288),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_532),
.B(n_288),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_544),
.B(n_298),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_490),
.B(n_298),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_546),
.B(n_298),
.Y(n_745)
);

NAND2xp33_ASAP7_75t_SL g746 ( 
.A(n_535),
.B(n_298),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_612),
.B(n_325),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_621),
.B(n_325),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_513),
.B(n_325),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_513),
.B(n_325),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_SL g751 ( 
.A(n_618),
.B(n_73),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_578),
.B(n_74),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_582),
.B(n_74),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_481),
.B(n_352),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_617),
.B(n_352),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_617),
.B(n_352),
.Y(n_756)
);

NAND2xp33_ASAP7_75t_SL g757 ( 
.A(n_555),
.B(n_352),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_555),
.B(n_535),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_591),
.B(n_393),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_SL g760 ( 
.A(n_499),
.B(n_82),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_591),
.B(n_235),
.Y(n_761)
);

NAND2xp33_ASAP7_75t_SL g762 ( 
.A(n_499),
.B(n_82),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_595),
.B(n_103),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_596),
.B(n_597),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_SL g765 ( 
.A(n_499),
.B(n_103),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_591),
.B(n_235),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_SL g767 ( 
.A(n_499),
.B(n_104),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_SL g768 ( 
.A(n_533),
.B(n_235),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_545),
.B(n_430),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_614),
.B(n_239),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_SL g771 ( 
.A(n_614),
.B(n_239),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_SL g772 ( 
.A(n_499),
.B(n_104),
.Y(n_772)
);

NAND2xp33_ASAP7_75t_SL g773 ( 
.A(n_478),
.B(n_106),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_SL g774 ( 
.A(n_478),
.B(n_106),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_616),
.B(n_239),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_557),
.B(n_247),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_557),
.B(n_583),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_583),
.B(n_247),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_516),
.B(n_247),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_SL g780 ( 
.A(n_516),
.B(n_252),
.Y(n_780)
);

NAND2xp33_ASAP7_75t_SL g781 ( 
.A(n_486),
.B(n_108),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_SL g782 ( 
.A(n_516),
.B(n_252),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_485),
.B(n_108),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_488),
.B(n_176),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_SL g785 ( 
.A(n_563),
.B(n_252),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_SL g786 ( 
.A(n_486),
.B(n_275),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_489),
.B(n_275),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_489),
.B(n_275),
.Y(n_788)
);

NAND2xp33_ASAP7_75t_SL g789 ( 
.A(n_563),
.B(n_176),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_L g790 ( 
.A(n_600),
.B(n_603),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_511),
.B(n_221),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_609),
.B(n_136),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_590),
.B(n_55),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_790),
.Y(n_794)
);

BUFx12f_ASAP7_75t_L g795 ( 
.A(n_675),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_665),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_764),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_692),
.A2(n_586),
.B1(n_572),
.B2(n_573),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_769),
.Y(n_799)
);

BUFx8_ASAP7_75t_L g800 ( 
.A(n_733),
.Y(n_800)
);

BUFx6f_ASAP7_75t_L g801 ( 
.A(n_706),
.Y(n_801)
);

AND2x2_ASAP7_75t_L g802 ( 
.A(n_769),
.B(n_624),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_768),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_629),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_744),
.B(n_624),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_645),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_640),
.B(n_619),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_SL g808 ( 
.A1(n_644),
.A2(n_109),
.B1(n_102),
.B2(n_105),
.Y(n_808)
);

AND3x1_ASAP7_75t_SL g809 ( 
.A(n_751),
.B(n_105),
.C(n_102),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_744),
.B(n_624),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_626),
.B(n_477),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_631),
.B(n_563),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_657),
.B(n_477),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_793),
.B(n_496),
.Y(n_814)
);

AND2x2_ASAP7_75t_L g815 ( 
.A(n_744),
.B(n_624),
.Y(n_815)
);

NAND2x1p5_ASAP7_75t_L g816 ( 
.A(n_779),
.B(n_572),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_712),
.B(n_496),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_761),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_635),
.A2(n_586),
.B(n_604),
.C(n_567),
.Y(n_819)
);

INVx2_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

NAND2x1p5_ASAP7_75t_L g821 ( 
.A(n_780),
.B(n_541),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_766),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_627),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_706),
.Y(n_824)
);

CKINVDCx5p33_ASAP7_75t_R g825 ( 
.A(n_783),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_713),
.B(n_510),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_631),
.B(n_571),
.Y(n_827)
);

BUFx3_ASAP7_75t_L g828 ( 
.A(n_706),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_635),
.A2(n_570),
.B1(n_545),
.B2(n_575),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_723),
.B(n_56),
.Y(n_830)
);

BUFx6f_ASAP7_75t_L g831 ( 
.A(n_722),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_643),
.B(n_571),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_673),
.B(n_510),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_722),
.B(n_605),
.Y(n_834)
);

AND3x1_ASAP7_75t_SL g835 ( 
.A(n_773),
.B(n_109),
.C(n_1),
.Y(n_835)
);

AND3x1_ASAP7_75t_SL g836 ( 
.A(n_774),
.B(n_0),
.C(n_1),
.Y(n_836)
);

INVx3_ASAP7_75t_L g837 ( 
.A(n_722),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_716),
.B(n_522),
.Y(n_838)
);

INVx2_ASAP7_75t_SL g839 ( 
.A(n_758),
.Y(n_839)
);

NAND3xp33_ASAP7_75t_SL g840 ( 
.A(n_718),
.B(n_88),
.C(n_57),
.Y(n_840)
);

INVx5_ASAP7_75t_L g841 ( 
.A(n_643),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_782),
.Y(n_842)
);

AND2x2_ASAP7_75t_L g843 ( 
.A(n_650),
.B(n_605),
.Y(n_843)
);

OAI22xp5_ASAP7_75t_L g844 ( 
.A1(n_725),
.A2(n_686),
.B1(n_726),
.B2(n_724),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_651),
.B(n_605),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_727),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_705),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_633),
.A2(n_541),
.B(n_567),
.C(n_588),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_732),
.B(n_522),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_652),
.B(n_605),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_643),
.B(n_571),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_785),
.Y(n_852)
);

BUFx2_ASAP7_75t_L g853 ( 
.A(n_785),
.Y(n_853)
);

BUFx6f_ASAP7_75t_L g854 ( 
.A(n_686),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_654),
.B(n_590),
.Y(n_855)
);

AOI221xp5_ASAP7_75t_L g856 ( 
.A1(n_752),
.A2(n_96),
.B1(n_76),
.B2(n_75),
.C(n_98),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_753),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_670),
.B(n_551),
.Y(n_858)
);

NAND2x1p5_ASAP7_75t_L g859 ( 
.A(n_642),
.B(n_505),
.Y(n_859)
);

INVx2_ASAP7_75t_L g860 ( 
.A(n_709),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_SL g861 ( 
.A1(n_763),
.A2(n_100),
.B1(n_80),
.B2(n_81),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_781),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_630),
.A2(n_545),
.B1(n_623),
.B2(n_608),
.Y(n_863)
);

OAI21xp5_ASAP7_75t_L g864 ( 
.A1(n_759),
.A2(n_536),
.B(n_553),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_670),
.B(n_725),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_639),
.B(n_551),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_632),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_647),
.B(n_562),
.Y(n_868)
);

CKINVDCx6p67_ASAP7_75t_R g869 ( 
.A(n_729),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_686),
.B(n_576),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_641),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_792),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_670),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_695),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_648),
.B(n_562),
.Y(n_875)
);

INVx3_ASAP7_75t_L g876 ( 
.A(n_664),
.Y(n_876)
);

AND2x2_ASAP7_75t_SL g877 ( 
.A(n_633),
.B(n_576),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_708),
.B(n_784),
.Y(n_878)
);

BUFx6f_ASAP7_75t_L g879 ( 
.A(n_663),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_694),
.B(n_566),
.Y(n_880)
);

INVxp67_ASAP7_75t_L g881 ( 
.A(n_638),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_697),
.B(n_566),
.Y(n_882)
);

AOI22xp5_ASAP7_75t_L g883 ( 
.A1(n_728),
.A2(n_545),
.B1(n_508),
.B2(n_505),
.Y(n_883)
);

INVx4_ASAP7_75t_L g884 ( 
.A(n_684),
.Y(n_884)
);

INVx5_ASAP7_75t_L g885 ( 
.A(n_684),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_702),
.Y(n_886)
);

AOI22xp33_ASAP7_75t_L g887 ( 
.A1(n_630),
.A2(n_601),
.B1(n_623),
.B2(n_608),
.Y(n_887)
);

OAI22xp5_ASAP7_75t_L g888 ( 
.A1(n_659),
.A2(n_508),
.B1(n_625),
.B2(n_536),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_634),
.B(n_568),
.Y(n_889)
);

INVx2_ASAP7_75t_L g890 ( 
.A(n_703),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_L g891 ( 
.A(n_646),
.B(n_568),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_740),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_776),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_730),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_777),
.B(n_580),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_693),
.A2(n_580),
.B1(n_607),
.B2(n_601),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_778),
.Y(n_897)
);

BUFx3_ASAP7_75t_L g898 ( 
.A(n_714),
.Y(n_898)
);

AND2x2_ASAP7_75t_L g899 ( 
.A(n_698),
.B(n_587),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_760),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_775),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_699),
.B(n_587),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_731),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_770),
.B(n_511),
.Y(n_904)
);

AOI21xp33_ASAP7_75t_L g905 ( 
.A1(n_791),
.A2(n_607),
.B(n_224),
.Y(n_905)
);

AND2x2_ASAP7_75t_SL g906 ( 
.A(n_734),
.B(n_306),
.Y(n_906)
);

BUFx8_ASAP7_75t_L g907 ( 
.A(n_762),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_715),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_649),
.B(n_524),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_656),
.B(n_136),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_735),
.B(n_524),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_658),
.B(n_136),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_771),
.B(n_584),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_737),
.B(n_136),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_636),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_736),
.B(n_625),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_676),
.B(n_584),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_636),
.Y(n_918)
);

HB1xp67_ASAP7_75t_L g919 ( 
.A(n_747),
.Y(n_919)
);

BUFx3_ASAP7_75t_L g920 ( 
.A(n_696),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_741),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_742),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_700),
.B(n_138),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_715),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_L g925 ( 
.A(n_749),
.B(n_138),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_765),
.A2(n_221),
.B1(n_224),
.B2(n_154),
.Y(n_926)
);

AND2x2_ASAP7_75t_SL g927 ( 
.A(n_680),
.B(n_116),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_787),
.Y(n_928)
);

AND2x2_ASAP7_75t_L g929 ( 
.A(n_701),
.B(n_159),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_788),
.Y(n_930)
);

AND2x2_ASAP7_75t_L g931 ( 
.A(n_743),
.B(n_159),
.Y(n_931)
);

BUFx2_ASAP7_75t_SL g932 ( 
.A(n_677),
.Y(n_932)
);

NAND2x1p5_ASAP7_75t_L g933 ( 
.A(n_748),
.B(n_581),
.Y(n_933)
);

INVx1_ASAP7_75t_SL g934 ( 
.A(n_767),
.Y(n_934)
);

AOI22xp5_ASAP7_75t_L g935 ( 
.A1(n_772),
.A2(n_91),
.B1(n_79),
.B2(n_99),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_745),
.B(n_159),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_754),
.B(n_130),
.Y(n_937)
);

INVx1_ASAP7_75t_L g938 ( 
.A(n_696),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_710),
.B(n_130),
.Y(n_939)
);

A2O1A1Ixp33_ASAP7_75t_SL g940 ( 
.A1(n_637),
.A2(n_130),
.B(n_138),
.C(n_148),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_750),
.B(n_138),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_789),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_687),
.B(n_133),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_711),
.Y(n_944)
);

NAND2x1p5_ASAP7_75t_L g945 ( 
.A(n_691),
.B(n_211),
.Y(n_945)
);

INVx4_ASAP7_75t_L g946 ( 
.A(n_746),
.Y(n_946)
);

INVx5_ASAP7_75t_SL g947 ( 
.A(n_927),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_901),
.Y(n_948)
);

BUFx4f_ASAP7_75t_L g949 ( 
.A(n_927),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_798),
.A2(n_756),
.B(n_755),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_901),
.Y(n_951)
);

OAI21x1_ASAP7_75t_SL g952 ( 
.A1(n_946),
.A2(n_746),
.B(n_757),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_924),
.Y(n_953)
);

INVx6_ASAP7_75t_L g954 ( 
.A(n_841),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_938),
.Y(n_955)
);

INVx2_ASAP7_75t_SL g956 ( 
.A(n_885),
.Y(n_956)
);

AND2x2_ASAP7_75t_L g957 ( 
.A(n_796),
.B(n_116),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_853),
.Y(n_958)
);

AOI21x1_ASAP7_75t_L g959 ( 
.A1(n_917),
.A2(n_660),
.B(n_661),
.Y(n_959)
);

AND2x2_ASAP7_75t_L g960 ( 
.A(n_796),
.B(n_118),
.Y(n_960)
);

OAI21x1_ASAP7_75t_L g961 ( 
.A1(n_933),
.A2(n_685),
.B(n_717),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_924),
.Y(n_962)
);

AO21x2_ASAP7_75t_L g963 ( 
.A1(n_864),
.A2(n_721),
.B(n_719),
.Y(n_963)
);

OAI21x1_ASAP7_75t_L g964 ( 
.A1(n_933),
.A2(n_683),
.B(n_678),
.Y(n_964)
);

INVx1_ASAP7_75t_SL g965 ( 
.A(n_846),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_885),
.Y(n_966)
);

BUFx12f_ASAP7_75t_L g967 ( 
.A(n_800),
.Y(n_967)
);

OR2x6_ASAP7_75t_L g968 ( 
.A(n_908),
.B(n_689),
.Y(n_968)
);

OAI21x1_ASAP7_75t_L g969 ( 
.A1(n_933),
.A2(n_679),
.B(n_681),
.Y(n_969)
);

AND2x2_ASAP7_75t_L g970 ( 
.A(n_877),
.B(n_118),
.Y(n_970)
);

OAI21x1_ASAP7_75t_L g971 ( 
.A1(n_938),
.A2(n_682),
.B(n_671),
.Y(n_971)
);

BUFx12f_ASAP7_75t_L g972 ( 
.A(n_800),
.Y(n_972)
);

BUFx12f_ASAP7_75t_L g973 ( 
.A(n_800),
.Y(n_973)
);

AOI21x1_ASAP7_75t_L g974 ( 
.A1(n_844),
.A2(n_662),
.B(n_674),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_846),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_920),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_820),
.Y(n_977)
);

INVxp33_ASAP7_75t_L g978 ( 
.A(n_806),
.Y(n_978)
);

BUFx6f_ASAP7_75t_L g979 ( 
.A(n_885),
.Y(n_979)
);

OAI21x1_ASAP7_75t_L g980 ( 
.A1(n_859),
.A2(n_667),
.B(n_668),
.Y(n_980)
);

AND2x4_ASAP7_75t_L g981 ( 
.A(n_885),
.B(n_690),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_859),
.A2(n_672),
.B(n_130),
.Y(n_982)
);

AO21x2_ASAP7_75t_L g983 ( 
.A1(n_803),
.A2(n_120),
.B(n_121),
.Y(n_983)
);

OAI21x1_ASAP7_75t_L g984 ( 
.A1(n_859),
.A2(n_130),
.B(n_148),
.Y(n_984)
);

OAI21x1_ASAP7_75t_L g985 ( 
.A1(n_888),
.A2(n_133),
.B(n_148),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_893),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_885),
.B(n_920),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_885),
.Y(n_988)
);

OAI21x1_ASAP7_75t_L g989 ( 
.A1(n_915),
.A2(n_133),
.B(n_148),
.Y(n_989)
);

INVx6_ASAP7_75t_SL g990 ( 
.A(n_904),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_915),
.A2(n_133),
.B(n_148),
.Y(n_991)
);

BUFx2_ASAP7_75t_L g992 ( 
.A(n_853),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_884),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_893),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_884),
.Y(n_995)
);

BUFx12f_ASAP7_75t_L g996 ( 
.A(n_857),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_797),
.B(n_120),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_918),
.Y(n_998)
);

INVx6_ASAP7_75t_L g999 ( 
.A(n_841),
.Y(n_999)
);

OAI21x1_ASAP7_75t_SL g1000 ( 
.A1(n_946),
.A2(n_739),
.B(n_666),
.Y(n_1000)
);

INVx2_ASAP7_75t_SL g1001 ( 
.A(n_841),
.Y(n_1001)
);

OAI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_798),
.A2(n_637),
.B(n_666),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_918),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_897),
.Y(n_1004)
);

BUFx2_ASAP7_75t_SL g1005 ( 
.A(n_884),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_797),
.Y(n_1006)
);

AND2x4_ASAP7_75t_L g1007 ( 
.A(n_908),
.B(n_133),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_897),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_820),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_852),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_823),
.Y(n_1011)
);

BUFx10_ASAP7_75t_L g1012 ( 
.A(n_927),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_852),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_794),
.Y(n_1014)
);

AND2x2_ASAP7_75t_L g1015 ( 
.A(n_877),
.B(n_865),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_877),
.A2(n_688),
.B(n_653),
.Y(n_1016)
);

OAI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_848),
.A2(n_704),
.B(n_720),
.Y(n_1017)
);

AND2x4_ASAP7_75t_L g1018 ( 
.A(n_799),
.B(n_137),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_946),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_816),
.A2(n_137),
.B(n_786),
.Y(n_1020)
);

BUFx6f_ASAP7_75t_L g1021 ( 
.A(n_841),
.Y(n_1021)
);

INVx5_ASAP7_75t_L g1022 ( 
.A(n_870),
.Y(n_1022)
);

BUFx2_ASAP7_75t_SL g1023 ( 
.A(n_841),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_794),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_803),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_SL g1026 ( 
.A(n_903),
.B(n_738),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_841),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_812),
.A2(n_121),
.B(n_137),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_847),
.Y(n_1029)
);

BUFx12f_ASAP7_75t_L g1030 ( 
.A(n_857),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_823),
.Y(n_1031)
);

AOI22x1_ASAP7_75t_L g1032 ( 
.A1(n_942),
.A2(n_89),
.B1(n_85),
.B2(n_86),
.Y(n_1032)
);

OAI21x1_ASAP7_75t_L g1033 ( 
.A1(n_816),
.A2(n_137),
.B(n_121),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_847),
.Y(n_1034)
);

INVx1_ASAP7_75t_SL g1035 ( 
.A(n_795),
.Y(n_1035)
);

INVx1_ASAP7_75t_SL g1036 ( 
.A(n_795),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_867),
.Y(n_1037)
);

NAND2x1p5_ASAP7_75t_L g1038 ( 
.A(n_916),
.B(n_688),
.Y(n_1038)
);

BUFx6f_ASAP7_75t_L g1039 ( 
.A(n_801),
.Y(n_1039)
);

BUFx2_ASAP7_75t_L g1040 ( 
.A(n_913),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_860),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_799),
.B(n_669),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_816),
.A2(n_137),
.B(n_190),
.Y(n_1043)
);

HB1xp67_ASAP7_75t_L g1044 ( 
.A(n_860),
.Y(n_1044)
);

BUFx3_ASAP7_75t_L g1045 ( 
.A(n_870),
.Y(n_1045)
);

INVx2_ASAP7_75t_SL g1046 ( 
.A(n_867),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_804),
.Y(n_1047)
);

BUFx12f_ASAP7_75t_L g1048 ( 
.A(n_825),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_802),
.B(n_142),
.Y(n_1049)
);

INVx6_ASAP7_75t_L g1050 ( 
.A(n_907),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_945),
.A2(n_205),
.B(n_190),
.Y(n_1051)
);

INVx6_ASAP7_75t_L g1052 ( 
.A(n_907),
.Y(n_1052)
);

AO21x2_ASAP7_75t_L g1053 ( 
.A1(n_905),
.A2(n_191),
.B(n_190),
.Y(n_1053)
);

AO21x2_ASAP7_75t_L g1054 ( 
.A1(n_895),
.A2(n_191),
.B(n_190),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_804),
.Y(n_1055)
);

BUFx12f_ASAP7_75t_L g1056 ( 
.A(n_825),
.Y(n_1056)
);

BUFx3_ASAP7_75t_L g1057 ( 
.A(n_870),
.Y(n_1057)
);

AO21x2_ASAP7_75t_L g1058 ( 
.A1(n_891),
.A2(n_191),
.B(n_190),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_818),
.Y(n_1059)
);

BUFx2_ASAP7_75t_SL g1060 ( 
.A(n_870),
.Y(n_1060)
);

CKINVDCx20_ASAP7_75t_R g1061 ( 
.A(n_862),
.Y(n_1061)
);

BUFx2_ASAP7_75t_R g1062 ( 
.A(n_903),
.Y(n_1062)
);

OAI21x1_ASAP7_75t_SL g1063 ( 
.A1(n_839),
.A2(n_878),
.B(n_829),
.Y(n_1063)
);

INVx3_ASAP7_75t_L g1064 ( 
.A(n_913),
.Y(n_1064)
);

BUFx10_ASAP7_75t_L g1065 ( 
.A(n_942),
.Y(n_1065)
);

INVx3_ASAP7_75t_L g1066 ( 
.A(n_913),
.Y(n_1066)
);

AO21x2_ASAP7_75t_L g1067 ( 
.A1(n_818),
.A2(n_191),
.B(n_205),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_822),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_874),
.B(n_83),
.Y(n_1069)
);

INVx3_ASAP7_75t_SL g1070 ( 
.A(n_842),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_822),
.Y(n_1071)
);

AOI22xp5_ASAP7_75t_L g1072 ( 
.A1(n_808),
.A2(n_669),
.B1(n_707),
.B2(n_704),
.Y(n_1072)
);

OAI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_935),
.A2(n_720),
.B(n_707),
.Y(n_1073)
);

BUFx3_ASAP7_75t_L g1074 ( 
.A(n_870),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_801),
.Y(n_1075)
);

INVx2_ASAP7_75t_SL g1076 ( 
.A(n_839),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1006),
.B(n_865),
.Y(n_1077)
);

BUFx12f_ASAP7_75t_L g1078 ( 
.A(n_967),
.Y(n_1078)
);

INVx2_ASAP7_75t_SL g1079 ( 
.A(n_1076),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_948),
.Y(n_1080)
);

CKINVDCx11_ASAP7_75t_R g1081 ( 
.A(n_1061),
.Y(n_1081)
);

CKINVDCx6p67_ASAP7_75t_R g1082 ( 
.A(n_967),
.Y(n_1082)
);

INVx6_ASAP7_75t_L g1083 ( 
.A(n_972),
.Y(n_1083)
);

CKINVDCx11_ASAP7_75t_R g1084 ( 
.A(n_972),
.Y(n_1084)
);

AOI22xp33_ASAP7_75t_L g1085 ( 
.A1(n_949),
.A2(n_870),
.B1(n_898),
.B2(n_814),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_SL g1086 ( 
.A1(n_1060),
.A2(n_870),
.B1(n_907),
.B2(n_842),
.Y(n_1086)
);

BUFx4f_ASAP7_75t_SL g1087 ( 
.A(n_973),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_1009),
.Y(n_1088)
);

BUFx10_ASAP7_75t_L g1089 ( 
.A(n_1050),
.Y(n_1089)
);

AOI22xp33_ASAP7_75t_L g1090 ( 
.A1(n_949),
.A2(n_898),
.B1(n_858),
.B2(n_882),
.Y(n_1090)
);

INVx1_ASAP7_75t_SL g1091 ( 
.A(n_1070),
.Y(n_1091)
);

INVx2_ASAP7_75t_L g1092 ( 
.A(n_1009),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_966),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_949),
.A2(n_858),
.B1(n_882),
.B2(n_880),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1009),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_1070),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_958),
.Y(n_1097)
);

AOI22xp33_ASAP7_75t_L g1098 ( 
.A1(n_949),
.A2(n_880),
.B1(n_845),
.B2(n_850),
.Y(n_1098)
);

AOI22xp33_ASAP7_75t_L g1099 ( 
.A1(n_1045),
.A2(n_845),
.B1(n_843),
.B2(n_850),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1014),
.B(n_874),
.Y(n_1100)
);

AOI22xp33_ASAP7_75t_SL g1101 ( 
.A1(n_1060),
.A2(n_900),
.B1(n_873),
.B2(n_932),
.Y(n_1101)
);

INVx4_ASAP7_75t_L g1102 ( 
.A(n_987),
.Y(n_1102)
);

AOI22xp33_ASAP7_75t_SL g1103 ( 
.A1(n_1045),
.A2(n_873),
.B1(n_932),
.B2(n_934),
.Y(n_1103)
);

CKINVDCx16_ASAP7_75t_R g1104 ( 
.A(n_973),
.Y(n_1104)
);

INVx1_ASAP7_75t_L g1105 ( 
.A(n_948),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_1011),
.Y(n_1106)
);

BUFx12f_ASAP7_75t_L g1107 ( 
.A(n_996),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_966),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_1072),
.A2(n_819),
.B1(n_869),
.B2(n_894),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_996),
.Y(n_1110)
);

AOI22xp33_ASAP7_75t_L g1111 ( 
.A1(n_1045),
.A2(n_843),
.B1(n_855),
.B2(n_802),
.Y(n_1111)
);

BUFx2_ASAP7_75t_L g1112 ( 
.A(n_958),
.Y(n_1112)
);

BUFx3_ASAP7_75t_L g1113 ( 
.A(n_1050),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_SL g1114 ( 
.A(n_1030),
.Y(n_1114)
);

OAI22xp33_ASAP7_75t_L g1115 ( 
.A1(n_1072),
.A2(n_883),
.B1(n_821),
.B2(n_869),
.Y(n_1115)
);

BUFx12f_ASAP7_75t_L g1116 ( 
.A(n_1030),
.Y(n_1116)
);

INVx6_ASAP7_75t_L g1117 ( 
.A(n_1022),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1011),
.Y(n_1118)
);

INVx2_ASAP7_75t_L g1119 ( 
.A(n_1011),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1031),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_1031),
.Y(n_1121)
);

CKINVDCx11_ASAP7_75t_R g1122 ( 
.A(n_1048),
.Y(n_1122)
);

AND2x2_ASAP7_75t_L g1123 ( 
.A(n_1064),
.B(n_824),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_1048),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_1070),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_951),
.Y(n_1126)
);

AOI22xp33_ASAP7_75t_SL g1127 ( 
.A1(n_1057),
.A2(n_830),
.B1(n_821),
.B2(n_834),
.Y(n_1127)
);

CKINVDCx11_ASAP7_75t_R g1128 ( 
.A(n_1056),
.Y(n_1128)
);

AOI22xp33_ASAP7_75t_L g1129 ( 
.A1(n_1057),
.A2(n_855),
.B1(n_876),
.B2(n_863),
.Y(n_1129)
);

CKINVDCx11_ASAP7_75t_R g1130 ( 
.A(n_1056),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1031),
.Y(n_1131)
);

BUFx12f_ASAP7_75t_L g1132 ( 
.A(n_1050),
.Y(n_1132)
);

CKINVDCx11_ASAP7_75t_R g1133 ( 
.A(n_965),
.Y(n_1133)
);

OAI22xp5_ASAP7_75t_L g1134 ( 
.A1(n_947),
.A2(n_975),
.B1(n_1002),
.B2(n_968),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_951),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1025),
.Y(n_1136)
);

AOI22xp33_ASAP7_75t_SL g1137 ( 
.A1(n_1057),
.A2(n_821),
.B1(n_834),
.B2(n_906),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_966),
.Y(n_1138)
);

OAI22xp5_ASAP7_75t_L g1139 ( 
.A1(n_947),
.A2(n_968),
.B1(n_1073),
.B2(n_1017),
.Y(n_1139)
);

OAI22xp5_ASAP7_75t_L g1140 ( 
.A1(n_947),
.A2(n_827),
.B1(n_926),
.B2(n_824),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1025),
.Y(n_1141)
);

AOI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1074),
.A2(n_876),
.B1(n_872),
.B2(n_849),
.Y(n_1142)
);

INVx3_ASAP7_75t_L g1143 ( 
.A(n_966),
.Y(n_1143)
);

OAI22xp5_ASAP7_75t_L g1144 ( 
.A1(n_947),
.A2(n_837),
.B1(n_824),
.B2(n_828),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_1055),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_1035),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_1074),
.A2(n_876),
.B1(n_872),
.B2(n_838),
.Y(n_1147)
);

INVx2_ASAP7_75t_SL g1148 ( 
.A(n_1076),
.Y(n_1148)
);

INVx3_ASAP7_75t_L g1149 ( 
.A(n_966),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_1022),
.Y(n_1150)
);

INVx1_ASAP7_75t_SL g1151 ( 
.A(n_1036),
.Y(n_1151)
);

AOI22xp33_ASAP7_75t_L g1152 ( 
.A1(n_1074),
.A2(n_889),
.B1(n_840),
.B2(n_902),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1014),
.B(n_944),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_992),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_987),
.Y(n_1155)
);

INVx6_ASAP7_75t_L g1156 ( 
.A(n_1022),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_986),
.Y(n_1157)
);

OAI21xp5_ASAP7_75t_SL g1158 ( 
.A1(n_992),
.A2(n_836),
.B(n_835),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_986),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_1055),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_1022),
.A2(n_889),
.B1(n_902),
.B2(n_899),
.Y(n_1161)
);

AOI22xp33_ASAP7_75t_L g1162 ( 
.A1(n_1022),
.A2(n_899),
.B1(n_909),
.B2(n_887),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_994),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1064),
.B(n_837),
.Y(n_1164)
);

INVx6_ASAP7_75t_L g1165 ( 
.A(n_1022),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_1050),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_947),
.A2(n_837),
.B1(n_828),
.B2(n_831),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1063),
.A2(n_906),
.B1(n_815),
.B2(n_810),
.Y(n_1168)
);

AOI22xp33_ASAP7_75t_SL g1169 ( 
.A1(n_1063),
.A2(n_906),
.B1(n_815),
.B2(n_810),
.Y(n_1169)
);

AOI22xp33_ASAP7_75t_SL g1170 ( 
.A1(n_970),
.A2(n_805),
.B1(n_854),
.B2(n_861),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1055),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_994),
.Y(n_1172)
);

AOI22xp33_ASAP7_75t_L g1173 ( 
.A1(n_970),
.A2(n_909),
.B1(n_871),
.B2(n_892),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1024),
.B(n_944),
.Y(n_1174)
);

INVx1_ASAP7_75t_L g1175 ( 
.A(n_1004),
.Y(n_1175)
);

AOI22xp33_ASAP7_75t_L g1176 ( 
.A1(n_957),
.A2(n_871),
.B1(n_892),
.B2(n_886),
.Y(n_1176)
);

INVx1_ASAP7_75t_SL g1177 ( 
.A(n_1062),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_1052),
.Y(n_1178)
);

BUFx8_ASAP7_75t_L g1179 ( 
.A(n_1019),
.Y(n_1179)
);

OAI21xp5_ASAP7_75t_SL g1180 ( 
.A1(n_1016),
.A2(n_856),
.B(n_809),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_987),
.Y(n_1181)
);

AND2x2_ASAP7_75t_L g1182 ( 
.A(n_1064),
.B(n_805),
.Y(n_1182)
);

INVx6_ASAP7_75t_L g1183 ( 
.A(n_1052),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1004),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_SL g1185 ( 
.A1(n_1052),
.A2(n_854),
.B1(n_831),
.B2(n_801),
.Y(n_1185)
);

AOI22xp33_ASAP7_75t_L g1186 ( 
.A1(n_957),
.A2(n_921),
.B1(n_922),
.B2(n_890),
.Y(n_1186)
);

INVx1_ASAP7_75t_L g1187 ( 
.A(n_1008),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_SL g1188 ( 
.A1(n_1012),
.A2(n_854),
.B1(n_801),
.B2(n_831),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_960),
.A2(n_1015),
.B1(n_1029),
.B2(n_1041),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1012),
.A2(n_854),
.B1(n_801),
.B2(n_831),
.Y(n_1190)
);

AOI22xp5_ASAP7_75t_L g1191 ( 
.A1(n_960),
.A2(n_881),
.B1(n_854),
.B2(n_807),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_1052),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1015),
.A2(n_922),
.B1(n_886),
.B2(n_890),
.Y(n_1193)
);

AO22x1_ASAP7_75t_L g1194 ( 
.A1(n_987),
.A2(n_904),
.B1(n_928),
.B2(n_930),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_1008),
.Y(n_1195)
);

AOI22xp33_ASAP7_75t_L g1196 ( 
.A1(n_1029),
.A2(n_921),
.B1(n_904),
.B2(n_896),
.Y(n_1196)
);

INVx1_ASAP7_75t_SL g1197 ( 
.A(n_976),
.Y(n_1197)
);

AOI21xp5_ASAP7_75t_L g1198 ( 
.A1(n_1109),
.A2(n_952),
.B(n_1000),
.Y(n_1198)
);

HB1xp67_ASAP7_75t_L g1199 ( 
.A(n_1097),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_L g1200 ( 
.A(n_1079),
.B(n_953),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1158),
.A2(n_1032),
.B(n_1069),
.Y(n_1201)
);

OAI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1158),
.A2(n_1032),
.B(n_1059),
.Y(n_1202)
);

INVx4_ASAP7_75t_SL g1203 ( 
.A(n_1117),
.Y(n_1203)
);

OAI21xp5_ASAP7_75t_L g1204 ( 
.A1(n_1180),
.A2(n_1068),
.B(n_1059),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1142),
.A2(n_1003),
.B(n_998),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_L g1206 ( 
.A1(n_1152),
.A2(n_983),
.B1(n_1041),
.B2(n_1034),
.Y(n_1206)
);

NAND2xp5_ASAP7_75t_L g1207 ( 
.A(n_1079),
.B(n_953),
.Y(n_1207)
);

HB1xp67_ASAP7_75t_L g1208 ( 
.A(n_1097),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1102),
.Y(n_1209)
);

OA21x2_ASAP7_75t_L g1210 ( 
.A1(n_1147),
.A2(n_1003),
.B(n_998),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_1080),
.Y(n_1211)
);

OA21x2_ASAP7_75t_L g1212 ( 
.A1(n_1153),
.A2(n_1003),
.B(n_998),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1080),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1105),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1088),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_1105),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1126),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1112),
.Y(n_1218)
);

OR2x6_ASAP7_75t_L g1219 ( 
.A(n_1194),
.B(n_1023),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1180),
.A2(n_988),
.B(n_950),
.C(n_976),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1148),
.B(n_962),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1126),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1135),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1115),
.A2(n_952),
.B(n_1000),
.Y(n_1224)
);

AOI221xp5_ASAP7_75t_L g1225 ( 
.A1(n_1139),
.A2(n_1024),
.B1(n_978),
.B2(n_1034),
.C(n_997),
.Y(n_1225)
);

AOI22xp33_ASAP7_75t_SL g1226 ( 
.A1(n_1134),
.A2(n_1012),
.B1(n_976),
.B2(n_1023),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1140),
.A2(n_1026),
.B(n_911),
.Y(n_1227)
);

AOI22xp5_ASAP7_75t_L g1228 ( 
.A1(n_1170),
.A2(n_1012),
.B1(n_1049),
.B2(n_968),
.Y(n_1228)
);

A2O1A1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1086),
.A2(n_988),
.B(n_976),
.C(n_956),
.Y(n_1229)
);

NAND2xp5_ASAP7_75t_SL g1230 ( 
.A(n_1148),
.B(n_1019),
.Y(n_1230)
);

INVx2_ASAP7_75t_L g1231 ( 
.A(n_1088),
.Y(n_1231)
);

AOI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1194),
.A2(n_1071),
.B(n_1068),
.Y(n_1232)
);

A2O1A1Ixp33_ASAP7_75t_L g1233 ( 
.A1(n_1085),
.A2(n_988),
.B(n_956),
.C(n_1040),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_L g1234 ( 
.A(n_1112),
.B(n_962),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1102),
.B(n_1064),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1144),
.A2(n_1038),
.B(n_993),
.Y(n_1236)
);

BUFx5_ASAP7_75t_L g1237 ( 
.A(n_1132),
.Y(n_1237)
);

OAI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1168),
.A2(n_1071),
.B(n_1038),
.Y(n_1238)
);

INVx2_ASAP7_75t_L g1239 ( 
.A(n_1092),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1093),
.A2(n_974),
.B(n_969),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_1102),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1135),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_1136),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1136),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_SL g1245 ( 
.A(n_1154),
.B(n_1019),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1185),
.A2(n_1038),
.B(n_993),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1141),
.Y(n_1247)
);

AND2x4_ASAP7_75t_L g1248 ( 
.A(n_1155),
.B(n_1066),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1185),
.A2(n_993),
.B(n_940),
.Y(n_1249)
);

OAI211xp5_ASAP7_75t_L g1250 ( 
.A1(n_1154),
.A2(n_1013),
.B(n_955),
.C(n_1040),
.Y(n_1250)
);

OAI21x1_ASAP7_75t_L g1251 ( 
.A1(n_1093),
.A2(n_974),
.B(n_969),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1092),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1095),
.Y(n_1253)
);

OA21x2_ASAP7_75t_L g1254 ( 
.A1(n_1174),
.A2(n_1013),
.B(n_955),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1077),
.B(n_955),
.Y(n_1255)
);

A2O1A1Ixp33_ASAP7_75t_L g1256 ( 
.A1(n_1169),
.A2(n_1191),
.B(n_1103),
.C(n_1137),
.Y(n_1256)
);

AOI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1167),
.A2(n_993),
.B(n_655),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_1095),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1106),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1182),
.B(n_1066),
.Y(n_1260)
);

CKINVDCx11_ASAP7_75t_R g1261 ( 
.A(n_1081),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_1084),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1141),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1077),
.B(n_1066),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_1182),
.B(n_1066),
.Y(n_1265)
);

AOI221xp5_ASAP7_75t_L g1266 ( 
.A1(n_1189),
.A2(n_1100),
.B1(n_1173),
.B2(n_1195),
.C(n_1187),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1157),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1197),
.A2(n_995),
.B(n_968),
.Y(n_1268)
);

AOI21xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1104),
.A2(n_968),
.B(n_995),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1157),
.B(n_1044),
.Y(n_1270)
);

OAI21x1_ASAP7_75t_L g1271 ( 
.A1(n_1093),
.A2(n_964),
.B(n_961),
.Y(n_1271)
);

INVx4_ASAP7_75t_L g1272 ( 
.A(n_1083),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1159),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1197),
.A2(n_995),
.B(n_1019),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1108),
.A2(n_964),
.B(n_961),
.Y(n_1275)
);

OA21x2_ASAP7_75t_L g1276 ( 
.A1(n_1106),
.A2(n_1047),
.B(n_977),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1159),
.B(n_1010),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1129),
.A2(n_1196),
.B1(n_1098),
.B2(n_1162),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1163),
.Y(n_1279)
);

AOI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1163),
.A2(n_959),
.B(n_1028),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1155),
.B(n_1010),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_SL g1282 ( 
.A(n_1091),
.B(n_1019),
.Y(n_1282)
);

AND2x2_ASAP7_75t_L g1283 ( 
.A(n_1155),
.B(n_1010),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1172),
.Y(n_1284)
);

NAND2xp5_ASAP7_75t_L g1285 ( 
.A(n_1172),
.B(n_1010),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1175),
.B(n_1037),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1175),
.B(n_1037),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1184),
.B(n_1046),
.Y(n_1288)
);

OA21x2_ASAP7_75t_L g1289 ( 
.A1(n_1118),
.A2(n_1047),
.B(n_977),
.Y(n_1289)
);

OAI21xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1096),
.A2(n_995),
.B(n_1001),
.Y(n_1290)
);

OAI221xp5_ASAP7_75t_L g1291 ( 
.A1(n_1127),
.A2(n_1046),
.B1(n_811),
.B2(n_919),
.C(n_813),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1101),
.A2(n_1019),
.B(n_1001),
.Y(n_1292)
);

AO21x2_ASAP7_75t_L g1293 ( 
.A1(n_1191),
.A2(n_983),
.B(n_1058),
.Y(n_1293)
);

AOI221xp5_ASAP7_75t_L g1294 ( 
.A1(n_1184),
.A2(n_930),
.B1(n_928),
.B2(n_1018),
.C(n_1049),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1187),
.Y(n_1295)
);

OA21x2_ASAP7_75t_L g1296 ( 
.A1(n_1118),
.A2(n_971),
.B(n_1020),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1181),
.B(n_1042),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1195),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1151),
.B(n_1007),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_SL g1300 ( 
.A(n_1181),
.B(n_966),
.Y(n_1300)
);

OR2x2_ASAP7_75t_L g1301 ( 
.A(n_1181),
.B(n_1042),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1108),
.A2(n_832),
.B(n_851),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1123),
.B(n_1007),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1099),
.A2(n_983),
.B1(n_990),
.B2(n_1049),
.Y(n_1304)
);

NOR2xp33_ASAP7_75t_L g1305 ( 
.A(n_1125),
.B(n_1065),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1123),
.B(n_1007),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1164),
.B(n_1042),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1119),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1108),
.A2(n_980),
.B(n_971),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1078),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1119),
.Y(n_1311)
);

INVx2_ASAP7_75t_L g1312 ( 
.A(n_1120),
.Y(n_1312)
);

OA21x2_ASAP7_75t_L g1313 ( 
.A1(n_1120),
.A2(n_1020),
.B(n_991),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1121),
.Y(n_1314)
);

BUFx2_ASAP7_75t_SL g1315 ( 
.A(n_1125),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1164),
.Y(n_1316)
);

CKINVDCx6p67_ASAP7_75t_R g1317 ( 
.A(n_1078),
.Y(n_1317)
);

AND2x2_ASAP7_75t_L g1318 ( 
.A(n_1138),
.B(n_1143),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1138),
.A2(n_980),
.B(n_991),
.Y(n_1319)
);

AOI21xp5_ASAP7_75t_L g1320 ( 
.A1(n_1138),
.A2(n_981),
.B(n_1042),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1121),
.Y(n_1321)
);

OAI22xp5_ASAP7_75t_L g1322 ( 
.A1(n_1178),
.A2(n_1005),
.B1(n_1007),
.B2(n_981),
.Y(n_1322)
);

INVx2_ASAP7_75t_L g1323 ( 
.A(n_1131),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1188),
.B(n_979),
.Y(n_1324)
);

OA21x2_ASAP7_75t_L g1325 ( 
.A1(n_1131),
.A2(n_989),
.B(n_985),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1143),
.A2(n_981),
.B(n_1042),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1193),
.B(n_1039),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1186),
.A2(n_959),
.B(n_1033),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1145),
.Y(n_1329)
);

A2O1A1Ixp33_ASAP7_75t_L g1330 ( 
.A1(n_1090),
.A2(n_979),
.B(n_1027),
.C(n_981),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1145),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1176),
.B(n_1039),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1160),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1160),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1094),
.A2(n_1111),
.B1(n_1161),
.B2(n_990),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1143),
.A2(n_979),
.B(n_963),
.Y(n_1336)
);

INVx2_ASAP7_75t_L g1337 ( 
.A(n_1171),
.Y(n_1337)
);

OAI21xp33_ASAP7_75t_L g1338 ( 
.A1(n_1204),
.A2(n_1146),
.B(n_1149),
.Y(n_1338)
);

AOI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1278),
.A2(n_1122),
.B1(n_1128),
.B2(n_1130),
.Y(n_1339)
);

AND2x2_ASAP7_75t_L g1340 ( 
.A(n_1260),
.B(n_1104),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1211),
.Y(n_1341)
);

AOI211xp5_ASAP7_75t_L g1342 ( 
.A1(n_1256),
.A2(n_1177),
.B(n_1146),
.C(n_1192),
.Y(n_1342)
);

AND2x2_ASAP7_75t_L g1343 ( 
.A(n_1260),
.B(n_1113),
.Y(n_1343)
);

OAI22xp33_ASAP7_75t_L g1344 ( 
.A1(n_1228),
.A2(n_1165),
.B1(n_1156),
.B2(n_1150),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1199),
.Y(n_1345)
);

NAND2xp5_ASAP7_75t_L g1346 ( 
.A(n_1208),
.B(n_1149),
.Y(n_1346)
);

OAI21xp5_ASAP7_75t_L g1347 ( 
.A1(n_1256),
.A2(n_1190),
.B(n_1033),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1220),
.A2(n_1183),
.B1(n_1005),
.B2(n_1083),
.Y(n_1348)
);

AOI222xp33_ASAP7_75t_L g1349 ( 
.A1(n_1201),
.A2(n_1110),
.B1(n_1107),
.B2(n_1116),
.C1(n_1124),
.C2(n_1087),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1220),
.A2(n_979),
.B(n_1149),
.Y(n_1350)
);

OAI221xp5_ASAP7_75t_L g1351 ( 
.A1(n_1202),
.A2(n_1083),
.B1(n_1171),
.B2(n_1183),
.C(n_1113),
.Y(n_1351)
);

AOI222xp33_ASAP7_75t_L g1352 ( 
.A1(n_1225),
.A2(n_1107),
.B1(n_1110),
.B2(n_1124),
.C1(n_1116),
.C2(n_1114),
.Y(n_1352)
);

INVx2_ASAP7_75t_SL g1353 ( 
.A(n_1310),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1206),
.A2(n_990),
.B1(n_1049),
.B2(n_831),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1218),
.B(n_1192),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1265),
.B(n_1082),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1264),
.B(n_1039),
.Y(n_1357)
);

OAI211xp5_ASAP7_75t_L g1358 ( 
.A1(n_1290),
.A2(n_1133),
.B(n_914),
.C(n_923),
.Y(n_1358)
);

INVx3_ASAP7_75t_L g1359 ( 
.A(n_1272),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1261),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1265),
.B(n_1082),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1213),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1335),
.A2(n_990),
.B1(n_1083),
.B2(n_1183),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1304),
.A2(n_1183),
.B1(n_1165),
.B2(n_1156),
.Y(n_1364)
);

OAI22xp33_ASAP7_75t_L g1365 ( 
.A1(n_1219),
.A2(n_1165),
.B1(n_1156),
.B2(n_1150),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1214),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1205),
.A2(n_1117),
.B1(n_1150),
.B2(n_1165),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1216),
.Y(n_1368)
);

AOI221xp5_ASAP7_75t_L g1369 ( 
.A1(n_1266),
.A2(n_1291),
.B1(n_1238),
.B2(n_1250),
.C(n_1294),
.Y(n_1369)
);

CKINVDCx6p67_ASAP7_75t_R g1370 ( 
.A(n_1261),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1227),
.A2(n_1132),
.B1(n_1156),
.B2(n_1150),
.Y(n_1371)
);

AOI221xp5_ASAP7_75t_L g1372 ( 
.A1(n_1255),
.A2(n_1018),
.B1(n_817),
.B2(n_826),
.C(n_833),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1316),
.B(n_1089),
.Y(n_1373)
);

INVx3_ASAP7_75t_L g1374 ( 
.A(n_1272),
.Y(n_1374)
);

HB1xp67_ASAP7_75t_L g1375 ( 
.A(n_1234),
.Y(n_1375)
);

OR2x2_ASAP7_75t_L g1376 ( 
.A(n_1264),
.B(n_1039),
.Y(n_1376)
);

NOR2xp33_ASAP7_75t_L g1377 ( 
.A(n_1315),
.B(n_1065),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1310),
.Y(n_1378)
);

O2A1O1Ixp33_ASAP7_75t_L g1379 ( 
.A1(n_1229),
.A2(n_868),
.B(n_875),
.C(n_912),
.Y(n_1379)
);

OAI211xp5_ASAP7_75t_L g1380 ( 
.A1(n_1198),
.A2(n_910),
.B(n_925),
.C(n_941),
.Y(n_1380)
);

AOI22xp33_ASAP7_75t_L g1381 ( 
.A1(n_1205),
.A2(n_1117),
.B1(n_963),
.B2(n_979),
.Y(n_1381)
);

NAND3xp33_ASAP7_75t_L g1382 ( 
.A(n_1200),
.B(n_1039),
.C(n_1075),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1307),
.B(n_1089),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1217),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1205),
.A2(n_1117),
.B1(n_963),
.B2(n_979),
.Y(n_1385)
);

NAND3xp33_ASAP7_75t_L g1386 ( 
.A(n_1207),
.B(n_1039),
.C(n_1075),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1222),
.Y(n_1387)
);

AOI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1332),
.A2(n_954),
.B1(n_999),
.B2(n_1027),
.Y(n_1388)
);

AND2x4_ASAP7_75t_L g1389 ( 
.A(n_1203),
.B(n_1021),
.Y(n_1389)
);

BUFx2_ASAP7_75t_L g1390 ( 
.A(n_1262),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_SL g1391 ( 
.A1(n_1210),
.A2(n_954),
.B1(n_999),
.B2(n_1021),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1286),
.B(n_1075),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1276),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1210),
.A2(n_954),
.B1(n_999),
.B2(n_866),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1223),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1276),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1210),
.A2(n_954),
.B1(n_999),
.B2(n_1018),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1276),
.Y(n_1398)
);

AOI22xp33_ASAP7_75t_L g1399 ( 
.A1(n_1293),
.A2(n_1018),
.B1(n_1058),
.B2(n_1054),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1242),
.Y(n_1400)
);

NOR2xp67_ASAP7_75t_L g1401 ( 
.A(n_1262),
.B(n_1021),
.Y(n_1401)
);

AOI22xp33_ASAP7_75t_SL g1402 ( 
.A1(n_1219),
.A2(n_1021),
.B1(n_1065),
.B2(n_1089),
.Y(n_1402)
);

CKINVDCx11_ASAP7_75t_R g1403 ( 
.A(n_1317),
.Y(n_1403)
);

AOI211x1_ASAP7_75t_L g1404 ( 
.A1(n_1224),
.A2(n_1028),
.B(n_931),
.C(n_936),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1293),
.A2(n_1058),
.B1(n_1054),
.B2(n_1021),
.Y(n_1405)
);

AOI22xp33_ASAP7_75t_L g1406 ( 
.A1(n_1293),
.A2(n_1054),
.B1(n_1021),
.B2(n_929),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1287),
.B(n_1075),
.Y(n_1407)
);

OAI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1236),
.A2(n_1229),
.B(n_1269),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1307),
.B(n_1166),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1243),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_SL g1411 ( 
.A(n_1246),
.B(n_1065),
.Y(n_1411)
);

A2O1A1Ixp33_ASAP7_75t_L g1412 ( 
.A1(n_1233),
.A2(n_1075),
.B(n_985),
.C(n_93),
.Y(n_1412)
);

AOI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1327),
.A2(n_1075),
.B(n_929),
.Y(n_1413)
);

AOI22xp33_ASAP7_75t_SL g1414 ( 
.A1(n_1219),
.A2(n_1166),
.B1(n_1179),
.B2(n_879),
.Y(n_1414)
);

AND2x2_ASAP7_75t_L g1415 ( 
.A(n_1297),
.B(n_1166),
.Y(n_1415)
);

AO31x2_ASAP7_75t_L g1416 ( 
.A1(n_1233),
.A2(n_943),
.A3(n_1067),
.B(n_1053),
.Y(n_1416)
);

OAI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1226),
.A2(n_879),
.B1(n_945),
.B2(n_931),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1244),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1221),
.Y(n_1419)
);

BUFx12f_ASAP7_75t_L g1420 ( 
.A(n_1272),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1328),
.A2(n_936),
.B1(n_1067),
.B2(n_1053),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1324),
.A2(n_879),
.B(n_1043),
.C(n_937),
.Y(n_1422)
);

HB1xp67_ASAP7_75t_L g1423 ( 
.A(n_1277),
.Y(n_1423)
);

AOI222xp33_ASAP7_75t_L g1424 ( 
.A1(n_1324),
.A2(n_154),
.B1(n_937),
.B2(n_939),
.C1(n_7),
.C2(n_10),
.Y(n_1424)
);

CKINVDCx5p33_ASAP7_75t_R g1425 ( 
.A(n_1317),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1219),
.A2(n_1067),
.B1(n_1053),
.B2(n_939),
.Y(n_1426)
);

OAI211xp5_ASAP7_75t_L g1427 ( 
.A1(n_1268),
.A2(n_0),
.B(n_2),
.C(n_5),
.Y(n_1427)
);

NOR2x1_ASAP7_75t_R g1428 ( 
.A(n_1237),
.B(n_1179),
.Y(n_1428)
);

AOI221xp5_ASAP7_75t_L g1429 ( 
.A1(n_1270),
.A2(n_879),
.B1(n_11),
.B2(n_13),
.C(n_15),
.Y(n_1429)
);

OAI211xp5_ASAP7_75t_L g1430 ( 
.A1(n_1245),
.A2(n_7),
.B(n_11),
.C(n_13),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1247),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1232),
.A2(n_989),
.B(n_1043),
.Y(n_1432)
);

INVx4_ASAP7_75t_L g1433 ( 
.A(n_1237),
.Y(n_1433)
);

BUFx12f_ASAP7_75t_L g1434 ( 
.A(n_1235),
.Y(n_1434)
);

AND2x2_ASAP7_75t_L g1435 ( 
.A(n_1297),
.B(n_1235),
.Y(n_1435)
);

INVx3_ASAP7_75t_L g1436 ( 
.A(n_1235),
.Y(n_1436)
);

NAND2x1p5_ASAP7_75t_L g1437 ( 
.A(n_1282),
.B(n_879),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1288),
.B(n_1179),
.Y(n_1438)
);

OAI33xp33_ASAP7_75t_L g1439 ( 
.A1(n_1285),
.A2(n_1298),
.A3(n_1284),
.B1(n_1295),
.B2(n_1273),
.B3(n_1279),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1299),
.A2(n_154),
.B1(n_1179),
.B2(n_945),
.Y(n_1440)
);

NAND3xp33_ASAP7_75t_L g1441 ( 
.A(n_1245),
.B(n_191),
.C(n_205),
.Y(n_1441)
);

AOI22xp33_ASAP7_75t_L g1442 ( 
.A1(n_1308),
.A2(n_154),
.B1(n_982),
.B2(n_984),
.Y(n_1442)
);

AOI22xp33_ASAP7_75t_L g1443 ( 
.A1(n_1321),
.A2(n_1334),
.B1(n_1333),
.B2(n_1331),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1329),
.A2(n_154),
.B1(n_982),
.B2(n_984),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1301),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1263),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1254),
.A2(n_154),
.B1(n_1051),
.B2(n_263),
.Y(n_1447)
);

OAI211xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1282),
.A2(n_16),
.B(n_18),
.C(n_21),
.Y(n_1448)
);

AOI22xp33_ASAP7_75t_L g1449 ( 
.A1(n_1254),
.A2(n_154),
.B1(n_1051),
.B2(n_263),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1254),
.A2(n_154),
.B1(n_263),
.B2(n_230),
.Y(n_1450)
);

AOI211xp5_ASAP7_75t_L g1451 ( 
.A1(n_1330),
.A2(n_18),
.B(n_23),
.C(n_24),
.Y(n_1451)
);

OAI22xp5_ASAP7_75t_SL g1452 ( 
.A1(n_1305),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_1452)
);

OR2x2_ASAP7_75t_L g1453 ( 
.A(n_1303),
.B(n_26),
.Y(n_1453)
);

AOI221xp5_ASAP7_75t_L g1454 ( 
.A1(n_1267),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.C(n_31),
.Y(n_1454)
);

INVx3_ASAP7_75t_L g1455 ( 
.A(n_1248),
.Y(n_1455)
);

OAI22xp5_ASAP7_75t_SL g1456 ( 
.A1(n_1301),
.A2(n_31),
.B1(n_32),
.B2(n_34),
.Y(n_1456)
);

OA21x2_ASAP7_75t_L g1457 ( 
.A1(n_1336),
.A2(n_205),
.B(n_230),
.Y(n_1457)
);

HB1xp67_ASAP7_75t_L g1458 ( 
.A(n_1212),
.Y(n_1458)
);

AND2x4_ASAP7_75t_L g1459 ( 
.A(n_1203),
.B(n_34),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1240),
.A2(n_205),
.B(n_230),
.Y(n_1460)
);

BUFx6f_ASAP7_75t_L g1461 ( 
.A(n_1240),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1248),
.B(n_35),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1251),
.A2(n_215),
.B(n_230),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1212),
.B(n_35),
.Y(n_1464)
);

OAI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1330),
.A2(n_36),
.B1(n_37),
.B2(n_38),
.Y(n_1465)
);

OR2x6_ASAP7_75t_L g1466 ( 
.A(n_1292),
.B(n_1320),
.Y(n_1466)
);

AOI221xp5_ASAP7_75t_L g1467 ( 
.A1(n_1215),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.C(n_45),
.Y(n_1467)
);

OAI211xp5_ASAP7_75t_L g1468 ( 
.A1(n_1230),
.A2(n_42),
.B(n_46),
.C(n_230),
.Y(n_1468)
);

AOI22xp33_ASAP7_75t_L g1469 ( 
.A1(n_1212),
.A2(n_263),
.B1(n_216),
.B2(n_215),
.Y(n_1469)
);

OAI221xp5_ASAP7_75t_L g1470 ( 
.A1(n_1326),
.A2(n_1337),
.B1(n_1253),
.B2(n_1323),
.C(n_1239),
.Y(n_1470)
);

INVx4_ASAP7_75t_L g1471 ( 
.A(n_1237),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1215),
.A2(n_263),
.B1(n_216),
.B2(n_215),
.Y(n_1472)
);

AOI21xp5_ASAP7_75t_L g1473 ( 
.A1(n_1257),
.A2(n_215),
.B(n_216),
.Y(n_1473)
);

AOI22xp33_ASAP7_75t_L g1474 ( 
.A1(n_1231),
.A2(n_216),
.B1(n_215),
.B2(n_46),
.Y(n_1474)
);

AOI22xp5_ASAP7_75t_L g1475 ( 
.A1(n_1322),
.A2(n_216),
.B1(n_179),
.B2(n_162),
.Y(n_1475)
);

NAND2xp5_ASAP7_75t_L g1476 ( 
.A(n_1318),
.B(n_49),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1302),
.A2(n_1230),
.B(n_1249),
.Y(n_1477)
);

AOI211xp5_ASAP7_75t_L g1478 ( 
.A1(n_1300),
.A2(n_179),
.B(n_162),
.C(n_164),
.Y(n_1478)
);

AOI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1231),
.A2(n_225),
.B1(n_162),
.B2(n_164),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1337),
.Y(n_1480)
);

AOI21xp5_ASAP7_75t_L g1481 ( 
.A1(n_1300),
.A2(n_179),
.B(n_162),
.Y(n_1481)
);

INVx4_ASAP7_75t_L g1482 ( 
.A(n_1237),
.Y(n_1482)
);

AOI22xp33_ASAP7_75t_L g1483 ( 
.A1(n_1239),
.A2(n_1252),
.B1(n_1323),
.B2(n_1314),
.Y(n_1483)
);

OAI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1252),
.A2(n_1259),
.B1(n_1253),
.B2(n_1314),
.C(n_1258),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_L g1485 ( 
.A1(n_1258),
.A2(n_225),
.B1(n_162),
.B2(n_164),
.Y(n_1485)
);

INVx1_ASAP7_75t_SL g1486 ( 
.A(n_1370),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1393),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1393),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1466),
.B(n_1436),
.Y(n_1489)
);

AND2x4_ASAP7_75t_L g1490 ( 
.A(n_1466),
.B(n_1203),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1464),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1341),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1362),
.Y(n_1493)
);

BUFx3_ASAP7_75t_L g1494 ( 
.A(n_1360),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1466),
.B(n_1318),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1366),
.Y(n_1496)
);

AND2x4_ASAP7_75t_SL g1497 ( 
.A(n_1459),
.B(n_1248),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1368),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1384),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1461),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1369),
.A2(n_1306),
.B1(n_1274),
.B2(n_1209),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1436),
.B(n_1209),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1396),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1387),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1455),
.B(n_1209),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1395),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1396),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1455),
.B(n_1435),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1400),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1340),
.B(n_1241),
.Y(n_1510)
);

AND2x2_ASAP7_75t_L g1511 ( 
.A(n_1356),
.B(n_1241),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1361),
.B(n_1241),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1373),
.B(n_1281),
.Y(n_1513)
);

INVxp67_ASAP7_75t_SL g1514 ( 
.A(n_1458),
.Y(n_1514)
);

NAND2x1_ASAP7_75t_L g1515 ( 
.A(n_1359),
.B(n_1281),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1398),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1375),
.B(n_1419),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1345),
.B(n_1283),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1423),
.B(n_1283),
.Y(n_1519)
);

BUFx2_ASAP7_75t_L g1520 ( 
.A(n_1477),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1346),
.B(n_1343),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1410),
.Y(n_1522)
);

AOI21xp5_ASAP7_75t_SL g1523 ( 
.A1(n_1459),
.A2(n_1296),
.B(n_1203),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1357),
.B(n_1271),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1418),
.B(n_1311),
.Y(n_1525)
);

INVx2_ASAP7_75t_SL g1526 ( 
.A(n_1461),
.Y(n_1526)
);

AO31x2_ASAP7_75t_L g1527 ( 
.A1(n_1398),
.A2(n_1311),
.A3(n_1259),
.B(n_1312),
.Y(n_1527)
);

OR2x2_ASAP7_75t_L g1528 ( 
.A(n_1431),
.B(n_1312),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1446),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1480),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1443),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1461),
.Y(n_1532)
);

BUFx3_ASAP7_75t_L g1533 ( 
.A(n_1360),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1443),
.Y(n_1534)
);

CKINVDCx5p33_ASAP7_75t_R g1535 ( 
.A(n_1403),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1390),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1359),
.B(n_1275),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1374),
.B(n_1275),
.Y(n_1538)
);

INVxp67_ASAP7_75t_SL g1539 ( 
.A(n_1342),
.Y(n_1539)
);

AOI22xp33_ASAP7_75t_L g1540 ( 
.A1(n_1339),
.A2(n_1289),
.B1(n_1296),
.B2(n_1251),
.Y(n_1540)
);

HB1xp67_ASAP7_75t_L g1541 ( 
.A(n_1461),
.Y(n_1541)
);

BUFx3_ASAP7_75t_L g1542 ( 
.A(n_1420),
.Y(n_1542)
);

NOR2x1_ASAP7_75t_L g1543 ( 
.A(n_1408),
.B(n_1296),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1392),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1407),
.B(n_1309),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1374),
.B(n_1383),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1376),
.B(n_1271),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1355),
.B(n_1309),
.Y(n_1548)
);

BUFx3_ASAP7_75t_L g1549 ( 
.A(n_1420),
.Y(n_1549)
);

AND2x2_ASAP7_75t_L g1550 ( 
.A(n_1409),
.B(n_1319),
.Y(n_1550)
);

AND2x2_ASAP7_75t_L g1551 ( 
.A(n_1338),
.B(n_1319),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1437),
.B(n_1313),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1457),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1457),
.Y(n_1554)
);

AND2x4_ASAP7_75t_L g1555 ( 
.A(n_1389),
.B(n_1401),
.Y(n_1555)
);

INVx4_ASAP7_75t_L g1556 ( 
.A(n_1425),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1453),
.B(n_1289),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1378),
.Y(n_1558)
);

INVx2_ASAP7_75t_L g1559 ( 
.A(n_1457),
.Y(n_1559)
);

HB1xp67_ASAP7_75t_L g1560 ( 
.A(n_1382),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1386),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1437),
.B(n_1313),
.Y(n_1562)
);

INVx2_ASAP7_75t_SL g1563 ( 
.A(n_1434),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1462),
.B(n_1289),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1470),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1421),
.B(n_1280),
.Y(n_1566)
);

AND2x2_ASAP7_75t_L g1567 ( 
.A(n_1434),
.B(n_1313),
.Y(n_1567)
);

INVx2_ASAP7_75t_L g1568 ( 
.A(n_1484),
.Y(n_1568)
);

OAI22xp33_ASAP7_75t_SL g1569 ( 
.A1(n_1465),
.A2(n_1237),
.B1(n_1325),
.B2(n_167),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1463),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1415),
.B(n_1237),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1389),
.B(n_1237),
.Y(n_1572)
);

BUFx3_ASAP7_75t_L g1573 ( 
.A(n_1378),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1421),
.B(n_1325),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1402),
.B(n_1325),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1378),
.B(n_225),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1438),
.B(n_179),
.Y(n_1577)
);

AND2x2_ASAP7_75t_L g1578 ( 
.A(n_1378),
.B(n_225),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1372),
.B(n_179),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1379),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1353),
.B(n_225),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1339),
.A2(n_174),
.B1(n_164),
.B2(n_167),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1483),
.Y(n_1583)
);

INVx3_ASAP7_75t_L g1584 ( 
.A(n_1433),
.Y(n_1584)
);

INVx1_ASAP7_75t_L g1585 ( 
.A(n_1483),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1414),
.B(n_1433),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1422),
.B(n_164),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1347),
.A2(n_175),
.B1(n_167),
.B2(n_184),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1367),
.B(n_225),
.Y(n_1589)
);

INVx2_ASAP7_75t_SL g1590 ( 
.A(n_1471),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1471),
.B(n_167),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1476),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1388),
.Y(n_1593)
);

BUFx6f_ASAP7_75t_L g1594 ( 
.A(n_1460),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1371),
.Y(n_1595)
);

INVx2_ASAP7_75t_L g1596 ( 
.A(n_1463),
.Y(n_1596)
);

AO21x2_ASAP7_75t_L g1597 ( 
.A1(n_1427),
.A2(n_167),
.B(n_184),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1351),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1381),
.B(n_225),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1381),
.B(n_225),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1385),
.B(n_225),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1411),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1411),
.Y(n_1603)
);

AO31x2_ASAP7_75t_L g1604 ( 
.A1(n_1422),
.A2(n_184),
.A3(n_175),
.B(n_174),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1463),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1527),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1522),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1522),
.Y(n_1608)
);

OA21x2_ASAP7_75t_L g1609 ( 
.A1(n_1520),
.A2(n_1385),
.B(n_1394),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1527),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1494),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_1535),
.Y(n_1612)
);

HB1xp67_ASAP7_75t_L g1613 ( 
.A(n_1492),
.Y(n_1613)
);

AOI211xp5_ASAP7_75t_L g1614 ( 
.A1(n_1520),
.A2(n_1452),
.B(n_1358),
.C(n_1456),
.Y(n_1614)
);

INVx5_ASAP7_75t_SL g1615 ( 
.A(n_1597),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1527),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1527),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1451),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1492),
.Y(n_1619)
);

AOI221xp5_ASAP7_75t_L g1620 ( 
.A1(n_1580),
.A2(n_1439),
.B1(n_1429),
.B2(n_1445),
.C(n_1454),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1495),
.B(n_1377),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_SL g1622 ( 
.A1(n_1539),
.A2(n_1574),
.B1(n_1566),
.B2(n_1531),
.Y(n_1622)
);

AND2x4_ASAP7_75t_L g1623 ( 
.A(n_1490),
.B(n_1482),
.Y(n_1623)
);

OAI21x1_ASAP7_75t_L g1624 ( 
.A1(n_1543),
.A2(n_1394),
.B(n_1350),
.Y(n_1624)
);

AOI21x1_ASAP7_75t_L g1625 ( 
.A1(n_1541),
.A2(n_1348),
.B(n_1473),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1539),
.A2(n_1467),
.B(n_1430),
.C(n_1448),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1493),
.Y(n_1627)
);

BUFx2_ASAP7_75t_SL g1628 ( 
.A(n_1556),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1501),
.A2(n_1412),
.B(n_1365),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1491),
.B(n_1352),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1493),
.Y(n_1631)
);

AND2x4_ASAP7_75t_L g1632 ( 
.A(n_1490),
.B(n_1482),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1496),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1495),
.B(n_1377),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1491),
.B(n_1517),
.Y(n_1635)
);

NAND4xp25_ASAP7_75t_L g1636 ( 
.A(n_1536),
.B(n_1349),
.C(n_1424),
.D(n_1404),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1517),
.B(n_1363),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1363),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1496),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1566),
.B(n_1416),
.Y(n_1640)
);

AOI221xp5_ASAP7_75t_L g1641 ( 
.A1(n_1531),
.A2(n_1406),
.B1(n_1413),
.B2(n_1397),
.C(n_1468),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1498),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1498),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1527),
.Y(n_1644)
);

OAI21x1_ASAP7_75t_L g1645 ( 
.A1(n_1543),
.A2(n_1397),
.B(n_1406),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1527),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1499),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1592),
.B(n_1474),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1499),
.Y(n_1649)
);

BUFx3_ASAP7_75t_L g1650 ( 
.A(n_1494),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1527),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1495),
.B(n_1391),
.Y(n_1652)
);

OAI22xp33_ASAP7_75t_L g1653 ( 
.A1(n_1574),
.A2(n_1417),
.B1(n_1344),
.B2(n_1475),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1504),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1487),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1487),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1487),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1504),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1536),
.B(n_1474),
.Y(n_1659)
);

AOI211xp5_ASAP7_75t_L g1660 ( 
.A1(n_1501),
.A2(n_1412),
.B(n_1380),
.C(n_1478),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1506),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1506),
.Y(n_1662)
);

INVx2_ASAP7_75t_SL g1663 ( 
.A(n_1494),
.Y(n_1663)
);

OAI22xp5_ASAP7_75t_L g1664 ( 
.A1(n_1588),
.A2(n_1364),
.B1(n_1426),
.B2(n_1354),
.Y(n_1664)
);

AND2x4_ASAP7_75t_L g1665 ( 
.A(n_1490),
.B(n_1416),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1509),
.Y(n_1666)
);

NOR2xp33_ASAP7_75t_L g1667 ( 
.A(n_1486),
.B(n_1428),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1509),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1529),
.Y(n_1669)
);

AOI211xp5_ASAP7_75t_L g1670 ( 
.A1(n_1569),
.A2(n_1441),
.B(n_1432),
.C(n_1416),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1602),
.B(n_1364),
.Y(n_1671)
);

OAI21x1_ASAP7_75t_L g1672 ( 
.A1(n_1500),
.A2(n_1405),
.B(n_1399),
.Y(n_1672)
);

AO21x2_ASAP7_75t_L g1673 ( 
.A1(n_1514),
.A2(n_1481),
.B(n_1416),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1529),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1602),
.B(n_1426),
.Y(n_1675)
);

AND2x4_ASAP7_75t_L g1676 ( 
.A(n_1490),
.B(n_1354),
.Y(n_1676)
);

OAI21xp33_ASAP7_75t_L g1677 ( 
.A1(n_1561),
.A2(n_1440),
.B(n_1405),
.Y(n_1677)
);

OAI21x1_ASAP7_75t_L g1678 ( 
.A1(n_1500),
.A2(n_1399),
.B(n_1469),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1489),
.B(n_1440),
.Y(n_1679)
);

AND2x4_ASAP7_75t_SL g1680 ( 
.A(n_1556),
.B(n_1447),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1603),
.B(n_1469),
.Y(n_1681)
);

AND2x2_ASAP7_75t_L g1682 ( 
.A(n_1489),
.B(n_1447),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1561),
.Y(n_1683)
);

AO21x2_ASAP7_75t_L g1684 ( 
.A1(n_1514),
.A2(n_1450),
.B(n_1449),
.Y(n_1684)
);

AND2x2_ASAP7_75t_L g1685 ( 
.A(n_1489),
.B(n_1449),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1486),
.B(n_1450),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1488),
.Y(n_1687)
);

OAI21x1_ASAP7_75t_L g1688 ( 
.A1(n_1500),
.A2(n_1442),
.B(n_1444),
.Y(n_1688)
);

OAI21x1_ASAP7_75t_L g1689 ( 
.A1(n_1500),
.A2(n_1442),
.B(n_1444),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1528),
.Y(n_1690)
);

NOR2xp67_ASAP7_75t_L g1691 ( 
.A(n_1556),
.B(n_1485),
.Y(n_1691)
);

AOI21xp5_ASAP7_75t_L g1692 ( 
.A1(n_1523),
.A2(n_1485),
.B(n_1479),
.Y(n_1692)
);

INVx2_ASAP7_75t_L g1693 ( 
.A(n_1488),
.Y(n_1693)
);

AOI22xp33_ASAP7_75t_L g1694 ( 
.A1(n_1534),
.A2(n_1479),
.B1(n_1472),
.B2(n_174),
.Y(n_1694)
);

OA21x2_ASAP7_75t_L g1695 ( 
.A1(n_1534),
.A2(n_1585),
.B(n_1583),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1488),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1533),
.Y(n_1697)
);

INVx4_ASAP7_75t_R g1698 ( 
.A(n_1533),
.Y(n_1698)
);

OA21x2_ASAP7_75t_L g1699 ( 
.A1(n_1583),
.A2(n_1472),
.B(n_184),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1528),
.Y(n_1700)
);

OAI21x1_ASAP7_75t_L g1701 ( 
.A1(n_1523),
.A2(n_184),
.B(n_174),
.Y(n_1701)
);

NAND4xp25_ASAP7_75t_L g1702 ( 
.A(n_1533),
.B(n_211),
.C(n_218),
.D(n_214),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1558),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1508),
.B(n_225),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_SL g1705 ( 
.A1(n_1569),
.A2(n_225),
.B1(n_173),
.B2(n_180),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1557),
.A2(n_174),
.B(n_175),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1503),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1525),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1603),
.B(n_225),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1525),
.Y(n_1710)
);

HB1xp67_ASAP7_75t_L g1711 ( 
.A(n_1611),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1613),
.Y(n_1712)
);

INVx2_ASAP7_75t_L g1713 ( 
.A(n_1606),
.Y(n_1713)
);

AOI221xp5_ASAP7_75t_L g1714 ( 
.A1(n_1622),
.A2(n_1585),
.B1(n_1540),
.B2(n_1565),
.C(n_1560),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1611),
.B(n_1586),
.Y(n_1715)
);

BUFx3_ASAP7_75t_L g1716 ( 
.A(n_1612),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1639),
.Y(n_1717)
);

OAI31xp33_ASAP7_75t_L g1718 ( 
.A1(n_1626),
.A2(n_1565),
.A3(n_1598),
.B(n_1589),
.Y(n_1718)
);

OR2x6_ASAP7_75t_SL g1719 ( 
.A(n_1630),
.B(n_1595),
.Y(n_1719)
);

INVx1_ASAP7_75t_L g1720 ( 
.A(n_1627),
.Y(n_1720)
);

AOI31xp33_ASAP7_75t_L g1721 ( 
.A1(n_1614),
.A2(n_1563),
.A3(n_1586),
.B(n_1560),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1697),
.B(n_1650),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1606),
.Y(n_1723)
);

INVx1_ASAP7_75t_L g1724 ( 
.A(n_1627),
.Y(n_1724)
);

BUFx2_ASAP7_75t_L g1725 ( 
.A(n_1650),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1697),
.B(n_1508),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1621),
.B(n_1573),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1631),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1621),
.B(n_1573),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_L g1730 ( 
.A(n_1612),
.B(n_1556),
.Y(n_1730)
);

INVx4_ASAP7_75t_L g1731 ( 
.A(n_1663),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1631),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1683),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1634),
.B(n_1663),
.Y(n_1734)
);

AND2x4_ASAP7_75t_SL g1735 ( 
.A(n_1623),
.B(n_1558),
.Y(n_1735)
);

INVx3_ASAP7_75t_L g1736 ( 
.A(n_1673),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1634),
.B(n_1573),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1607),
.B(n_1619),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1633),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1633),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1623),
.B(n_1558),
.Y(n_1741)
);

AND2x4_ASAP7_75t_L g1742 ( 
.A(n_1623),
.B(n_1526),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1642),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1642),
.Y(n_1744)
);

INVx4_ASAP7_75t_L g1745 ( 
.A(n_1703),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1632),
.B(n_1558),
.Y(n_1746)
);

NOR2xp67_ASAP7_75t_L g1747 ( 
.A(n_1652),
.B(n_1584),
.Y(n_1747)
);

AND2x4_ASAP7_75t_L g1748 ( 
.A(n_1632),
.B(n_1526),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1610),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1632),
.B(n_1558),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1704),
.B(n_1558),
.Y(n_1751)
);

AO21x2_ASAP7_75t_L g1752 ( 
.A1(n_1640),
.A2(n_1532),
.B(n_1541),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1660),
.A2(n_1595),
.B1(n_1563),
.B2(n_1593),
.Y(n_1753)
);

NOR2xp33_ASAP7_75t_L g1754 ( 
.A(n_1618),
.B(n_1542),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1610),
.Y(n_1755)
);

INVx4_ASAP7_75t_L g1756 ( 
.A(n_1703),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1635),
.B(n_1690),
.Y(n_1757)
);

INVx2_ASAP7_75t_L g1758 ( 
.A(n_1616),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1673),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1704),
.B(n_1558),
.Y(n_1760)
);

INVx4_ASAP7_75t_L g1761 ( 
.A(n_1703),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1652),
.B(n_1563),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1686),
.Y(n_1763)
);

NAND3xp33_ASAP7_75t_L g1764 ( 
.A(n_1620),
.B(n_1532),
.C(n_1582),
.Y(n_1764)
);

AOI221xp5_ASAP7_75t_L g1765 ( 
.A1(n_1675),
.A2(n_1575),
.B1(n_1568),
.B2(n_1557),
.C(n_1551),
.Y(n_1765)
);

AOI22xp33_ASAP7_75t_L g1766 ( 
.A1(n_1695),
.A2(n_1568),
.B1(n_1598),
.B2(n_1597),
.Y(n_1766)
);

OR2x2_ASAP7_75t_L g1767 ( 
.A(n_1700),
.B(n_1544),
.Y(n_1767)
);

INVx2_ASAP7_75t_L g1768 ( 
.A(n_1616),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1617),
.Y(n_1769)
);

AND2x2_ASAP7_75t_L g1770 ( 
.A(n_1628),
.B(n_1542),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1654),
.Y(n_1771)
);

AND2x2_ASAP7_75t_L g1772 ( 
.A(n_1628),
.B(n_1542),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1607),
.B(n_1643),
.Y(n_1773)
);

OR2x2_ASAP7_75t_L g1774 ( 
.A(n_1700),
.B(n_1544),
.Y(n_1774)
);

BUFx2_ASAP7_75t_L g1775 ( 
.A(n_1647),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1629),
.B(n_1555),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1681),
.B(n_1564),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1667),
.B(n_1549),
.Y(n_1778)
);

OAI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1692),
.A2(n_1564),
.B1(n_1568),
.B2(n_1589),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1654),
.Y(n_1780)
);

NAND3xp33_ASAP7_75t_SL g1781 ( 
.A(n_1670),
.B(n_1575),
.C(n_1551),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1649),
.B(n_1530),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1658),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1625),
.B(n_1549),
.Y(n_1784)
);

AND2x2_ASAP7_75t_L g1785 ( 
.A(n_1625),
.B(n_1549),
.Y(n_1785)
);

AOI22xp33_ASAP7_75t_SL g1786 ( 
.A1(n_1695),
.A2(n_1567),
.B1(n_1551),
.B2(n_1589),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1608),
.B(n_1497),
.Y(n_1787)
);

AOI22xp33_ASAP7_75t_SL g1788 ( 
.A1(n_1695),
.A2(n_1567),
.B1(n_1597),
.B2(n_1562),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1679),
.B(n_1497),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1679),
.B(n_1497),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1679),
.B(n_1546),
.Y(n_1791)
);

AOI33xp33_ASAP7_75t_L g1792 ( 
.A1(n_1653),
.A2(n_1593),
.A3(n_1567),
.B1(n_1562),
.B2(n_1552),
.B3(n_1532),
.Y(n_1792)
);

BUFx2_ASAP7_75t_L g1793 ( 
.A(n_1668),
.Y(n_1793)
);

HB1xp67_ASAP7_75t_L g1794 ( 
.A(n_1659),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1658),
.Y(n_1795)
);

NAND3xp33_ASAP7_75t_L g1796 ( 
.A(n_1636),
.B(n_1579),
.C(n_1587),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1661),
.Y(n_1797)
);

INVx2_ASAP7_75t_L g1798 ( 
.A(n_1617),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1648),
.B(n_1546),
.Y(n_1799)
);

OR2x2_ASAP7_75t_L g1800 ( 
.A(n_1796),
.B(n_1669),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1791),
.B(n_1691),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1775),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1775),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1791),
.B(n_1550),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1736),
.Y(n_1805)
);

NAND2xp5_ASAP7_75t_L g1806 ( 
.A(n_1799),
.B(n_1677),
.Y(n_1806)
);

OR2x2_ASAP7_75t_L g1807 ( 
.A(n_1796),
.B(n_1661),
.Y(n_1807)
);

AND2x2_ASAP7_75t_L g1808 ( 
.A(n_1727),
.B(n_1550),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1736),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1727),
.B(n_1550),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1793),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1733),
.B(n_1662),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1793),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1720),
.Y(n_1814)
);

HB1xp67_ASAP7_75t_L g1815 ( 
.A(n_1711),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1729),
.B(n_1584),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1736),
.Y(n_1817)
);

AND2x4_ASAP7_75t_L g1818 ( 
.A(n_1789),
.B(n_1676),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1789),
.B(n_1676),
.Y(n_1819)
);

BUFx2_ASAP7_75t_L g1820 ( 
.A(n_1778),
.Y(n_1820)
);

OR2x2_ASAP7_75t_L g1821 ( 
.A(n_1757),
.B(n_1662),
.Y(n_1821)
);

AND2x4_ASAP7_75t_L g1822 ( 
.A(n_1790),
.B(n_1676),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1715),
.B(n_1682),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1715),
.B(n_1682),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1720),
.Y(n_1825)
);

NOR2x1_ASAP7_75t_L g1826 ( 
.A(n_1721),
.B(n_1637),
.Y(n_1826)
);

AND2x4_ASAP7_75t_SL g1827 ( 
.A(n_1790),
.B(n_1698),
.Y(n_1827)
);

AND2x4_ASAP7_75t_L g1828 ( 
.A(n_1734),
.B(n_1722),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1763),
.B(n_1685),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1724),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1757),
.B(n_1666),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1763),
.B(n_1685),
.Y(n_1832)
);

NOR4xp25_ASAP7_75t_SL g1833 ( 
.A(n_1714),
.B(n_1641),
.C(n_1674),
.D(n_1666),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1721),
.B(n_1714),
.C(n_1753),
.Y(n_1834)
);

AND2x4_ASAP7_75t_SL g1835 ( 
.A(n_1734),
.B(n_1572),
.Y(n_1835)
);

AND2x2_ASAP7_75t_SL g1836 ( 
.A(n_1784),
.B(n_1785),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1762),
.Y(n_1837)
);

AND2x4_ASAP7_75t_L g1838 ( 
.A(n_1722),
.B(n_1674),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1725),
.B(n_1671),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1736),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1759),
.Y(n_1841)
);

INVx3_ASAP7_75t_L g1842 ( 
.A(n_1759),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1724),
.Y(n_1843)
);

OR2x2_ASAP7_75t_L g1844 ( 
.A(n_1767),
.B(n_1708),
.Y(n_1844)
);

INVx2_ASAP7_75t_L g1845 ( 
.A(n_1759),
.Y(n_1845)
);

INVx1_ASAP7_75t_SL g1846 ( 
.A(n_1716),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1786),
.B(n_1665),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1716),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1728),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1725),
.B(n_1638),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1728),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1729),
.B(n_1584),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1726),
.B(n_1708),
.Y(n_1853)
);

NAND2xp5_ASAP7_75t_L g1854 ( 
.A(n_1753),
.B(n_1762),
.Y(n_1854)
);

HB1xp67_ASAP7_75t_L g1855 ( 
.A(n_1726),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1732),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1737),
.B(n_1584),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1737),
.B(n_1590),
.Y(n_1858)
);

NAND2xp67_ASAP7_75t_L g1859 ( 
.A(n_1778),
.B(n_1680),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1732),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1735),
.B(n_1590),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1716),
.Y(n_1862)
);

INVx1_ASAP7_75t_SL g1863 ( 
.A(n_1719),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1735),
.B(n_1590),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1767),
.B(n_1710),
.Y(n_1865)
);

AND2x2_ASAP7_75t_L g1866 ( 
.A(n_1735),
.B(n_1521),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1739),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1741),
.B(n_1521),
.Y(n_1868)
);

HB1xp67_ASAP7_75t_L g1869 ( 
.A(n_1747),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1741),
.B(n_1521),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1739),
.Y(n_1871)
);

INVx2_ASAP7_75t_L g1872 ( 
.A(n_1759),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1746),
.B(n_1502),
.Y(n_1873)
);

AND2x2_ASAP7_75t_L g1874 ( 
.A(n_1746),
.B(n_1502),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1719),
.Y(n_1875)
);

OR2x6_ASAP7_75t_L g1876 ( 
.A(n_1794),
.B(n_1624),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1774),
.B(n_1710),
.Y(n_1877)
);

AND2x4_ASAP7_75t_L g1878 ( 
.A(n_1731),
.B(n_1680),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1750),
.B(n_1505),
.Y(n_1879)
);

AND2x4_ASAP7_75t_L g1880 ( 
.A(n_1731),
.B(n_1624),
.Y(n_1880)
);

NOR2xp33_ASAP7_75t_R g1881 ( 
.A(n_1730),
.B(n_1581),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1740),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_SL g1883 ( 
.A(n_1833),
.B(n_1792),
.C(n_1718),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1815),
.Y(n_1884)
);

AOI22xp5_ASAP7_75t_L g1885 ( 
.A1(n_1834),
.A2(n_1781),
.B1(n_1786),
.B2(n_1765),
.Y(n_1885)
);

INVx1_ASAP7_75t_SL g1886 ( 
.A(n_1820),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1820),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1827),
.B(n_1770),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1827),
.B(n_1770),
.Y(n_1889)
);

NOR4xp25_ASAP7_75t_L g1890 ( 
.A(n_1863),
.B(n_1781),
.C(n_1765),
.D(n_1764),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1837),
.B(n_1712),
.Y(n_1891)
);

AND4x1_ASAP7_75t_L g1892 ( 
.A(n_1826),
.B(n_1754),
.C(n_1718),
.D(n_1764),
.Y(n_1892)
);

INVx1_ASAP7_75t_SL g1893 ( 
.A(n_1875),
.Y(n_1893)
);

OAI22xp5_ASAP7_75t_SL g1894 ( 
.A1(n_1854),
.A2(n_1788),
.B1(n_1766),
.B2(n_1717),
.Y(n_1894)
);

OR2x2_ASAP7_75t_L g1895 ( 
.A(n_1807),
.B(n_1823),
.Y(n_1895)
);

NOR2xp33_ASAP7_75t_R g1896 ( 
.A(n_1846),
.B(n_1772),
.Y(n_1896)
);

AND2x4_ASAP7_75t_SL g1897 ( 
.A(n_1828),
.B(n_1772),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1855),
.Y(n_1898)
);

NAND4xp75_ASAP7_75t_L g1899 ( 
.A(n_1836),
.B(n_1784),
.C(n_1785),
.D(n_1747),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1828),
.B(n_1787),
.Y(n_1900)
);

OR2x2_ASAP7_75t_L g1901 ( 
.A(n_1807),
.B(n_1712),
.Y(n_1901)
);

OR2x2_ASAP7_75t_L g1902 ( 
.A(n_1824),
.B(n_1717),
.Y(n_1902)
);

NAND4xp75_ASAP7_75t_L g1903 ( 
.A(n_1836),
.B(n_1776),
.C(n_1609),
.D(n_1750),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1805),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1828),
.B(n_1787),
.Y(n_1905)
);

OR2x2_ASAP7_75t_L g1906 ( 
.A(n_1800),
.B(n_1738),
.Y(n_1906)
);

AND2x2_ASAP7_75t_L g1907 ( 
.A(n_1878),
.B(n_1742),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1878),
.B(n_1742),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1805),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1809),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1809),
.Y(n_1911)
);

HB1xp67_ASAP7_75t_L g1912 ( 
.A(n_1801),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1878),
.B(n_1742),
.Y(n_1913)
);

AND2x2_ASAP7_75t_L g1914 ( 
.A(n_1868),
.B(n_1870),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1868),
.B(n_1742),
.Y(n_1915)
);

NAND3xp33_ASAP7_75t_L g1916 ( 
.A(n_1847),
.B(n_1788),
.C(n_1731),
.Y(n_1916)
);

AND2x2_ASAP7_75t_L g1917 ( 
.A(n_1870),
.B(n_1748),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1817),
.Y(n_1918)
);

AOI22xp5_ASAP7_75t_L g1919 ( 
.A1(n_1876),
.A2(n_1779),
.B1(n_1777),
.B2(n_1609),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1817),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1840),
.Y(n_1921)
);

XOR2x2_ASAP7_75t_L g1922 ( 
.A(n_1829),
.B(n_1609),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1866),
.B(n_1748),
.Y(n_1923)
);

NOR2xp33_ASAP7_75t_L g1924 ( 
.A(n_1848),
.B(n_1731),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1840),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1853),
.B(n_1777),
.Y(n_1926)
);

INVx2_ASAP7_75t_SL g1927 ( 
.A(n_1818),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1853),
.B(n_1751),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1866),
.B(n_1748),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1876),
.Y(n_1930)
);

XNOR2x2_ASAP7_75t_L g1931 ( 
.A(n_1862),
.B(n_1645),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1853),
.B(n_1751),
.Y(n_1932)
);

NOR2xp33_ASAP7_75t_L g1933 ( 
.A(n_1832),
.B(n_1748),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1838),
.B(n_1760),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1876),
.Y(n_1935)
);

HB1xp67_ASAP7_75t_L g1936 ( 
.A(n_1801),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1876),
.Y(n_1937)
);

OAI21xp5_ASAP7_75t_L g1938 ( 
.A1(n_1806),
.A2(n_1645),
.B(n_1640),
.Y(n_1938)
);

INVx2_ASAP7_75t_SL g1939 ( 
.A(n_1818),
.Y(n_1939)
);

AOI22xp5_ASAP7_75t_L g1940 ( 
.A1(n_1818),
.A2(n_1664),
.B1(n_1615),
.B2(n_1684),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1841),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1841),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1816),
.B(n_1760),
.Y(n_1943)
);

INVx2_ASAP7_75t_L g1944 ( 
.A(n_1819),
.Y(n_1944)
);

NOR4xp75_ASAP7_75t_L g1945 ( 
.A(n_1839),
.B(n_1738),
.C(n_1773),
.D(n_1782),
.Y(n_1945)
);

XNOR2xp5_ASAP7_75t_L g1946 ( 
.A(n_1859),
.B(n_1702),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1845),
.Y(n_1947)
);

XNOR2xp5_ASAP7_75t_L g1948 ( 
.A(n_1859),
.B(n_1705),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1838),
.B(n_1773),
.Y(n_1949)
);

INVx2_ASAP7_75t_L g1950 ( 
.A(n_1819),
.Y(n_1950)
);

INVx2_ASAP7_75t_L g1951 ( 
.A(n_1819),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1816),
.B(n_1740),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1838),
.B(n_1743),
.Y(n_1953)
);

XNOR2x1_ASAP7_75t_L g1954 ( 
.A(n_1800),
.B(n_1672),
.Y(n_1954)
);

NOR2xp33_ASAP7_75t_L g1955 ( 
.A(n_1850),
.B(n_1774),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1845),
.Y(n_1956)
);

OR2x2_ASAP7_75t_L g1957 ( 
.A(n_1821),
.B(n_1782),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1852),
.B(n_1743),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1931),
.Y(n_1959)
);

INVx1_ASAP7_75t_L g1960 ( 
.A(n_1887),
.Y(n_1960)
);

NAND2x1_ASAP7_75t_L g1961 ( 
.A(n_1927),
.B(n_1880),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_L g1962 ( 
.A(n_1914),
.B(n_1822),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1914),
.B(n_1890),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1915),
.B(n_1858),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1887),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1906),
.B(n_1811),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_SL g1967 ( 
.A(n_1892),
.B(n_1880),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1915),
.B(n_1858),
.Y(n_1968)
);

AOI22xp5_ASAP7_75t_L g1969 ( 
.A1(n_1883),
.A2(n_1822),
.B1(n_1880),
.B2(n_1804),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1906),
.B(n_1811),
.Y(n_1970)
);

AND2x2_ASAP7_75t_L g1971 ( 
.A(n_1917),
.B(n_1822),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1886),
.B(n_1802),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1917),
.B(n_1852),
.Y(n_1973)
);

OAI21xp5_ASAP7_75t_SL g1974 ( 
.A1(n_1885),
.A2(n_1869),
.B(n_1857),
.Y(n_1974)
);

OAI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1919),
.A2(n_1842),
.B1(n_1865),
.B2(n_1877),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_L g1976 ( 
.A(n_1955),
.B(n_1803),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1952),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_L g1978 ( 
.A(n_1912),
.B(n_1813),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1900),
.B(n_1857),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1952),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1900),
.B(n_1905),
.Y(n_1981)
);

INVx2_ASAP7_75t_SL g1982 ( 
.A(n_1897),
.Y(n_1982)
);

AND2x2_ASAP7_75t_L g1983 ( 
.A(n_1905),
.B(n_1835),
.Y(n_1983)
);

AND2x2_ASAP7_75t_L g1984 ( 
.A(n_1927),
.B(n_1835),
.Y(n_1984)
);

OR2x2_ASAP7_75t_L g1985 ( 
.A(n_1895),
.B(n_1813),
.Y(n_1985)
);

INVxp33_ASAP7_75t_L g1986 ( 
.A(n_1896),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1936),
.B(n_1821),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1939),
.B(n_1923),
.Y(n_1988)
);

AND2x2_ASAP7_75t_L g1989 ( 
.A(n_1939),
.B(n_1804),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1923),
.B(n_1808),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1958),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1958),
.Y(n_1992)
);

INVx1_ASAP7_75t_L g1993 ( 
.A(n_1904),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1944),
.B(n_1831),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1896),
.Y(n_1995)
);

NOR2xp33_ASAP7_75t_L g1996 ( 
.A(n_1897),
.B(n_1831),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1931),
.Y(n_1997)
);

AOI221xp5_ASAP7_75t_L g1998 ( 
.A1(n_1894),
.A2(n_1872),
.B1(n_1882),
.B2(n_1814),
.C(n_1867),
.Y(n_1998)
);

NAND2x1p5_ASAP7_75t_L g1999 ( 
.A(n_1893),
.B(n_1842),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1944),
.B(n_1881),
.Y(n_2000)
);

AOI22xp5_ASAP7_75t_L g2001 ( 
.A1(n_1922),
.A2(n_1673),
.B1(n_1872),
.B2(n_1808),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1929),
.B(n_1810),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1909),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_L g2004 ( 
.A(n_1950),
.B(n_1844),
.Y(n_2004)
);

NOR2xp33_ASAP7_75t_L g2005 ( 
.A(n_1888),
.B(n_1812),
.Y(n_2005)
);

AOI32xp33_ASAP7_75t_L g2006 ( 
.A1(n_1954),
.A2(n_1810),
.A3(n_1842),
.B1(n_1814),
.B2(n_1825),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1950),
.B(n_1844),
.Y(n_2007)
);

NOR2xp33_ASAP7_75t_L g2008 ( 
.A(n_1888),
.B(n_1812),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1951),
.B(n_1865),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1929),
.B(n_1861),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1907),
.B(n_1861),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1916),
.B(n_1895),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1901),
.B(n_1877),
.Y(n_2013)
);

OAI22xp5_ASAP7_75t_L g2014 ( 
.A1(n_1903),
.A2(n_1879),
.B1(n_1874),
.B2(n_1873),
.Y(n_2014)
);

INVx2_ASAP7_75t_SL g2015 ( 
.A(n_1907),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1908),
.B(n_1864),
.Y(n_2016)
);

OAI21xp33_ASAP7_75t_L g2017 ( 
.A1(n_1969),
.A2(n_1933),
.B(n_1946),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1981),
.Y(n_2018)
);

OAI22xp5_ASAP7_75t_L g2019 ( 
.A1(n_1959),
.A2(n_1899),
.B1(n_1901),
.B2(n_1948),
.Y(n_2019)
);

INVx2_ASAP7_75t_SL g2020 ( 
.A(n_1971),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1989),
.Y(n_2021)
);

XNOR2xp5_ASAP7_75t_L g2022 ( 
.A(n_1971),
.B(n_1922),
.Y(n_2022)
);

OAI22xp5_ASAP7_75t_SL g2023 ( 
.A1(n_1963),
.A2(n_1951),
.B1(n_1946),
.B2(n_1884),
.Y(n_2023)
);

XNOR2xp5_ASAP7_75t_L g2024 ( 
.A(n_2014),
.B(n_1945),
.Y(n_2024)
);

AOI22xp33_ASAP7_75t_L g2025 ( 
.A1(n_1959),
.A2(n_1954),
.B1(n_1938),
.B2(n_1930),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1989),
.Y(n_2026)
);

NAND3xp33_ASAP7_75t_L g2027 ( 
.A(n_1998),
.B(n_1924),
.C(n_1898),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1981),
.Y(n_2028)
);

OR4x1_ASAP7_75t_L g2029 ( 
.A(n_1982),
.B(n_1918),
.C(n_1956),
.D(n_1910),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_2013),
.Y(n_2030)
);

INVx1_ASAP7_75t_SL g2031 ( 
.A(n_1997),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_2013),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1997),
.A2(n_1930),
.B1(n_1935),
.B2(n_1937),
.Y(n_2033)
);

NAND3xp33_ASAP7_75t_L g2034 ( 
.A(n_1967),
.B(n_1937),
.C(n_1935),
.Y(n_2034)
);

AOI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_2001),
.A2(n_1940),
.B1(n_1899),
.B2(n_1948),
.Y(n_2035)
);

INVx2_ASAP7_75t_SL g2036 ( 
.A(n_1988),
.Y(n_2036)
);

INVxp67_ASAP7_75t_L g2037 ( 
.A(n_1988),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_L g2038 ( 
.A(n_2012),
.B(n_1926),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1990),
.Y(n_2039)
);

AOI22xp5_ASAP7_75t_L g2040 ( 
.A1(n_1975),
.A2(n_1943),
.B1(n_1908),
.B2(n_1913),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1999),
.Y(n_2041)
);

AOI21xp33_ASAP7_75t_SL g2042 ( 
.A1(n_1967),
.A2(n_1902),
.B(n_1889),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1990),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_2002),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_2012),
.A2(n_1949),
.B(n_1891),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2002),
.Y(n_2046)
);

A2O1A1Ixp33_ASAP7_75t_L g2047 ( 
.A1(n_2006),
.A2(n_1957),
.B(n_1920),
.C(n_1947),
.Y(n_2047)
);

AOI221xp5_ASAP7_75t_L g2048 ( 
.A1(n_1974),
.A2(n_1925),
.B1(n_1911),
.B2(n_1942),
.C(n_1941),
.Y(n_2048)
);

AOI22xp33_ASAP7_75t_L g2049 ( 
.A1(n_1999),
.A2(n_1615),
.B1(n_1758),
.B2(n_1798),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_1985),
.A2(n_1957),
.B1(n_1902),
.B2(n_1921),
.Y(n_2050)
);

INVx1_ASAP7_75t_L g2051 ( 
.A(n_1985),
.Y(n_2051)
);

O2A1O1Ixp33_ASAP7_75t_L g2052 ( 
.A1(n_1995),
.A2(n_1986),
.B(n_1960),
.C(n_1965),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1977),
.Y(n_2053)
);

A2O1A1Ixp33_ASAP7_75t_L g2054 ( 
.A1(n_1986),
.A2(n_1672),
.B(n_1843),
.C(n_1825),
.Y(n_2054)
);

XOR2x2_ASAP7_75t_L g2055 ( 
.A(n_1961),
.B(n_1889),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1980),
.Y(n_2056)
);

NAND3xp33_ASAP7_75t_L g2057 ( 
.A(n_2005),
.B(n_1913),
.C(n_1953),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1991),
.Y(n_2058)
);

AOI22xp33_ASAP7_75t_L g2059 ( 
.A1(n_1993),
.A2(n_1615),
.B1(n_1798),
.B2(n_1769),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1992),
.Y(n_2060)
);

AND2x4_ASAP7_75t_L g2061 ( 
.A(n_2015),
.B(n_1943),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_L g2062 ( 
.A(n_1962),
.B(n_1928),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1994),
.Y(n_2063)
);

AOI22xp5_ASAP7_75t_L g2064 ( 
.A1(n_2010),
.A2(n_1932),
.B1(n_1934),
.B2(n_1752),
.Y(n_2064)
);

INVx1_ASAP7_75t_L g2065 ( 
.A(n_2004),
.Y(n_2065)
);

AO32x1_ASAP7_75t_L g2066 ( 
.A1(n_2019),
.A2(n_1982),
.A3(n_2015),
.B1(n_1984),
.B2(n_2016),
.Y(n_2066)
);

AOI211x1_ASAP7_75t_L g2067 ( 
.A1(n_2019),
.A2(n_1968),
.B(n_1964),
.C(n_1987),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_2061),
.B(n_1979),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_2028),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_2061),
.Y(n_2070)
);

OAI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2038),
.A2(n_1976),
.B1(n_1966),
.B2(n_1970),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2018),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_2036),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2020),
.B(n_1964),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2039),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2043),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_2055),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2037),
.B(n_1968),
.Y(n_2078)
);

NOR2xp33_ASAP7_75t_L g2079 ( 
.A(n_2042),
.B(n_1979),
.Y(n_2079)
);

OAI221xp5_ASAP7_75t_L g2080 ( 
.A1(n_2031),
.A2(n_2007),
.B1(n_2009),
.B2(n_1970),
.C(n_1966),
.Y(n_2080)
);

NAND2xp33_ASAP7_75t_SL g2081 ( 
.A(n_2038),
.B(n_2011),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2025),
.A2(n_1615),
.B1(n_1713),
.B2(n_1723),
.Y(n_2082)
);

OAI21xp5_ASAP7_75t_L g2083 ( 
.A1(n_2045),
.A2(n_1978),
.B(n_1972),
.Y(n_2083)
);

OR2x2_ASAP7_75t_L g2084 ( 
.A(n_2044),
.B(n_1973),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_2045),
.B(n_1973),
.Y(n_2085)
);

INVx1_ASAP7_75t_SL g2086 ( 
.A(n_2046),
.Y(n_2086)
);

OAI221xp5_ASAP7_75t_L g2087 ( 
.A1(n_2031),
.A2(n_2003),
.B1(n_2008),
.B2(n_2000),
.C(n_1996),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2030),
.Y(n_2088)
);

AOI21xp33_ASAP7_75t_L g2089 ( 
.A1(n_2052),
.A2(n_1867),
.B(n_1843),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_SL g2090 ( 
.A(n_2057),
.B(n_2017),
.Y(n_2090)
);

OAI221xp5_ASAP7_75t_L g2091 ( 
.A1(n_2022),
.A2(n_2016),
.B1(n_2011),
.B2(n_2010),
.C(n_1830),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2032),
.Y(n_2092)
);

INVx1_ASAP7_75t_L g2093 ( 
.A(n_2021),
.Y(n_2093)
);

INVx2_ASAP7_75t_L g2094 ( 
.A(n_2029),
.Y(n_2094)
);

AOI21xp33_ASAP7_75t_L g2095 ( 
.A1(n_2052),
.A2(n_1882),
.B(n_1830),
.Y(n_2095)
);

INVxp67_ASAP7_75t_SL g2096 ( 
.A(n_2051),
.Y(n_2096)
);

BUFx2_ASAP7_75t_L g2097 ( 
.A(n_2026),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2062),
.B(n_1984),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_L g2099 ( 
.A(n_2041),
.B(n_1983),
.Y(n_2099)
);

BUFx3_ASAP7_75t_L g2100 ( 
.A(n_2063),
.Y(n_2100)
);

OAI21xp33_ASAP7_75t_L g2101 ( 
.A1(n_2040),
.A2(n_1983),
.B(n_1864),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_2034),
.Y(n_2102)
);

OAI21xp33_ASAP7_75t_SL g2103 ( 
.A1(n_2048),
.A2(n_1745),
.B(n_1756),
.Y(n_2103)
);

AOI22xp5_ASAP7_75t_L g2104 ( 
.A1(n_2023),
.A2(n_2035),
.B1(n_2033),
.B2(n_2024),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_2065),
.Y(n_2105)
);

AOI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_2064),
.A2(n_1752),
.B1(n_1526),
.B2(n_1849),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_2053),
.Y(n_2107)
);

OAI21xp33_ASAP7_75t_L g2108 ( 
.A1(n_2027),
.A2(n_2047),
.B(n_2054),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_2050),
.B(n_2048),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_2060),
.Y(n_2110)
);

OAI22xp5_ASAP7_75t_L g2111 ( 
.A1(n_2049),
.A2(n_1856),
.B1(n_1851),
.B2(n_1860),
.Y(n_2111)
);

NAND2xp5_ASAP7_75t_L g2112 ( 
.A(n_2056),
.B(n_1871),
.Y(n_2112)
);

AOI22xp5_ASAP7_75t_L g2113 ( 
.A1(n_2102),
.A2(n_2059),
.B1(n_2058),
.B2(n_1752),
.Y(n_2113)
);

AOI211xp5_ASAP7_75t_L g2114 ( 
.A1(n_2108),
.A2(n_2071),
.B(n_2109),
.C(n_2083),
.Y(n_2114)
);

HB1xp67_ASAP7_75t_L g2115 ( 
.A(n_2084),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2070),
.B(n_1873),
.Y(n_2116)
);

XOR2x2_ASAP7_75t_L g2117 ( 
.A(n_2104),
.B(n_1752),
.Y(n_2117)
);

OAI32xp33_ASAP7_75t_L g2118 ( 
.A1(n_2085),
.A2(n_1761),
.A3(n_1756),
.B1(n_1745),
.B2(n_1797),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_2074),
.Y(n_2119)
);

OAI31xp33_ASAP7_75t_L g2120 ( 
.A1(n_2080),
.A2(n_1665),
.A3(n_1744),
.B(n_1771),
.Y(n_2120)
);

INVx1_ASAP7_75t_SL g2121 ( 
.A(n_2081),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2097),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_2066),
.Y(n_2123)
);

INVxp67_ASAP7_75t_L g2124 ( 
.A(n_2079),
.Y(n_2124)
);

INVxp67_ASAP7_75t_L g2125 ( 
.A(n_2068),
.Y(n_2125)
);

AOI221xp5_ASAP7_75t_L g2126 ( 
.A1(n_2071),
.A2(n_1744),
.B1(n_1771),
.B2(n_1780),
.C(n_1797),
.Y(n_2126)
);

INVx1_ASAP7_75t_L g2127 ( 
.A(n_2066),
.Y(n_2127)
);

OAI21xp33_ASAP7_75t_L g2128 ( 
.A1(n_2090),
.A2(n_1879),
.B(n_1874),
.Y(n_2128)
);

AOI22xp5_ASAP7_75t_L g2129 ( 
.A1(n_2077),
.A2(n_1795),
.B1(n_1783),
.B2(n_1780),
.Y(n_2129)
);

OAI22xp5_ASAP7_75t_L g2130 ( 
.A1(n_2067),
.A2(n_1783),
.B1(n_1795),
.B2(n_1761),
.Y(n_2130)
);

AO21x1_ASAP7_75t_L g2131 ( 
.A1(n_2083),
.A2(n_1745),
.B(n_1756),
.Y(n_2131)
);

AOI21xp5_ASAP7_75t_L g2132 ( 
.A1(n_2066),
.A2(n_1745),
.B(n_1756),
.Y(n_2132)
);

OAI21xp33_ASAP7_75t_SL g2133 ( 
.A1(n_2089),
.A2(n_1761),
.B(n_1769),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2096),
.B(n_1761),
.Y(n_2134)
);

OAI21xp33_ASAP7_75t_L g2135 ( 
.A1(n_2101),
.A2(n_1665),
.B(n_1709),
.Y(n_2135)
);

NOR2xp33_ASAP7_75t_L g2136 ( 
.A(n_2098),
.B(n_1655),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_2078),
.Y(n_2137)
);

OR2x2_ASAP7_75t_L g2138 ( 
.A(n_2086),
.B(n_2072),
.Y(n_2138)
);

AND2x2_ASAP7_75t_L g2139 ( 
.A(n_2069),
.B(n_1519),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2100),
.Y(n_2140)
);

NAND2xp5_ASAP7_75t_SL g2141 ( 
.A(n_2094),
.B(n_1655),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2088),
.Y(n_2142)
);

BUFx3_ASAP7_75t_L g2143 ( 
.A(n_2073),
.Y(n_2143)
);

AOI31xp33_ASAP7_75t_L g2144 ( 
.A1(n_2099),
.A2(n_1581),
.A3(n_1572),
.B(n_1578),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2092),
.B(n_1656),
.Y(n_2145)
);

OAI221xp5_ASAP7_75t_L g2146 ( 
.A1(n_2106),
.A2(n_1798),
.B1(n_1769),
.B2(n_1768),
.C(n_1758),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_L g2147 ( 
.A(n_2091),
.B(n_2103),
.Y(n_2147)
);

INVx2_ASAP7_75t_L g2148 ( 
.A(n_2116),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2115),
.Y(n_2149)
);

AND2x2_ASAP7_75t_L g2150 ( 
.A(n_2125),
.B(n_2075),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_2128),
.B(n_2107),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2138),
.Y(n_2152)
);

NOR3x1_ASAP7_75t_L g2153 ( 
.A(n_2123),
.B(n_2087),
.C(n_2076),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_2122),
.Y(n_2154)
);

NAND3xp33_ASAP7_75t_L g2155 ( 
.A(n_2114),
.B(n_2093),
.C(n_2110),
.Y(n_2155)
);

INVxp67_ASAP7_75t_L g2156 ( 
.A(n_2134),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_L g2157 ( 
.A(n_2121),
.B(n_2136),
.Y(n_2157)
);

INVxp33_ASAP7_75t_SL g2158 ( 
.A(n_2147),
.Y(n_2158)
);

INVx1_ASAP7_75t_SL g2159 ( 
.A(n_2143),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_SL g2160 ( 
.A(n_2127),
.B(n_2089),
.Y(n_2160)
);

AOI211xp5_ASAP7_75t_L g2161 ( 
.A1(n_2124),
.A2(n_2095),
.B(n_2111),
.C(n_2105),
.Y(n_2161)
);

NAND2xp5_ASAP7_75t_L g2162 ( 
.A(n_2140),
.B(n_2112),
.Y(n_2162)
);

NOR2xp33_ASAP7_75t_L g2163 ( 
.A(n_2134),
.B(n_2133),
.Y(n_2163)
);

INVx1_ASAP7_75t_L g2164 ( 
.A(n_2139),
.Y(n_2164)
);

CKINVDCx5p33_ASAP7_75t_R g2165 ( 
.A(n_2137),
.Y(n_2165)
);

NOR2xp33_ASAP7_75t_L g2166 ( 
.A(n_2119),
.B(n_2095),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_2145),
.Y(n_2167)
);

AND4x1_ASAP7_75t_L g2168 ( 
.A(n_2129),
.B(n_2082),
.C(n_2112),
.D(n_2111),
.Y(n_2168)
);

NAND2xp5_ASAP7_75t_SL g2169 ( 
.A(n_2132),
.B(n_1713),
.Y(n_2169)
);

O2A1O1Ixp5_ASAP7_75t_SL g2170 ( 
.A1(n_2142),
.A2(n_1723),
.B(n_1758),
.C(n_1755),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2145),
.Y(n_2171)
);

NOR2xp33_ASAP7_75t_SL g2172 ( 
.A(n_2132),
.B(n_1576),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2144),
.B(n_1678),
.Y(n_2173)
);

OA21x2_ASAP7_75t_L g2174 ( 
.A1(n_2160),
.A2(n_2113),
.B(n_2131),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_2148),
.Y(n_2175)
);

NOR2xp33_ASAP7_75t_L g2176 ( 
.A(n_2158),
.B(n_2141),
.Y(n_2176)
);

AOI211xp5_ASAP7_75t_L g2177 ( 
.A1(n_2160),
.A2(n_2155),
.B(n_2166),
.C(n_2149),
.Y(n_2177)
);

OAI221xp5_ASAP7_75t_L g2178 ( 
.A1(n_2166),
.A2(n_2117),
.B1(n_2120),
.B2(n_2146),
.C(n_2135),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_SL g2179 ( 
.A(n_2159),
.B(n_2130),
.Y(n_2179)
);

O2A1O1Ixp33_ASAP7_75t_SL g2180 ( 
.A1(n_2157),
.A2(n_2118),
.B(n_2126),
.C(n_2146),
.Y(n_2180)
);

AOI222xp33_ASAP7_75t_L g2181 ( 
.A1(n_2169),
.A2(n_2126),
.B1(n_1768),
.B2(n_1755),
.C1(n_1749),
.C2(n_1723),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2150),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2152),
.B(n_2164),
.Y(n_2183)
);

NOR4xp25_ASAP7_75t_L g2184 ( 
.A(n_2151),
.B(n_1768),
.C(n_1755),
.D(n_1749),
.Y(n_2184)
);

NAND3xp33_ASAP7_75t_L g2185 ( 
.A(n_2161),
.B(n_1749),
.C(n_1713),
.Y(n_2185)
);

A2O1A1Ixp33_ASAP7_75t_L g2186 ( 
.A1(n_2167),
.A2(n_1707),
.B(n_1656),
.C(n_1696),
.Y(n_2186)
);

OAI211xp5_ASAP7_75t_L g2187 ( 
.A1(n_2162),
.A2(n_1515),
.B(n_1706),
.C(n_1537),
.Y(n_2187)
);

AOI221xp5_ASAP7_75t_SL g2188 ( 
.A1(n_2156),
.A2(n_2163),
.B1(n_2154),
.B2(n_2169),
.C(n_2171),
.Y(n_2188)
);

AOI221xp5_ASAP7_75t_L g2189 ( 
.A1(n_2173),
.A2(n_2163),
.B1(n_2165),
.B2(n_2172),
.C(n_2153),
.Y(n_2189)
);

NAND4xp25_ASAP7_75t_L g2190 ( 
.A(n_2168),
.B(n_1576),
.C(n_1578),
.D(n_1577),
.Y(n_2190)
);

NOR2x1_ASAP7_75t_L g2191 ( 
.A(n_2170),
.B(n_1515),
.Y(n_2191)
);

AOI21xp5_ASAP7_75t_L g2192 ( 
.A1(n_2160),
.A2(n_1707),
.B(n_1696),
.Y(n_2192)
);

OAI221xp5_ASAP7_75t_L g2193 ( 
.A1(n_2160),
.A2(n_1693),
.B1(n_1687),
.B2(n_1657),
.C(n_1646),
.Y(n_2193)
);

AOI22xp33_ASAP7_75t_L g2194 ( 
.A1(n_2160),
.A2(n_1651),
.B1(n_1644),
.B2(n_1646),
.Y(n_2194)
);

INVxp67_ASAP7_75t_SL g2195 ( 
.A(n_2177),
.Y(n_2195)
);

AOI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2176),
.A2(n_1657),
.B1(n_1693),
.B2(n_1687),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_2183),
.Y(n_2197)
);

INVxp67_ASAP7_75t_L g2198 ( 
.A(n_2182),
.Y(n_2198)
);

INVx2_ASAP7_75t_L g2199 ( 
.A(n_2175),
.Y(n_2199)
);

A2O1A1Ixp33_ASAP7_75t_SL g2200 ( 
.A1(n_2178),
.A2(n_1538),
.B(n_1537),
.C(n_1644),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_2174),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2174),
.Y(n_2202)
);

INVx1_ASAP7_75t_L g2203 ( 
.A(n_2185),
.Y(n_2203)
);

AOI221xp5_ASAP7_75t_L g2204 ( 
.A1(n_2184),
.A2(n_2192),
.B1(n_2193),
.B2(n_2189),
.C(n_2180),
.Y(n_2204)
);

INVxp67_ASAP7_75t_SL g2205 ( 
.A(n_2179),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_2191),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2187),
.A2(n_1548),
.B1(n_1545),
.B2(n_1538),
.Y(n_2207)
);

NOR4xp25_ASAP7_75t_L g2208 ( 
.A(n_2188),
.B(n_1651),
.C(n_1503),
.D(n_1516),
.Y(n_2208)
);

AOI22xp5_ASAP7_75t_L g2209 ( 
.A1(n_2181),
.A2(n_1516),
.B1(n_1503),
.B2(n_1507),
.Y(n_2209)
);

INVxp67_ASAP7_75t_L g2210 ( 
.A(n_2190),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2194),
.A2(n_2186),
.B1(n_1548),
.B2(n_1545),
.Y(n_2211)
);

O2A1O1Ixp33_ASAP7_75t_L g2212 ( 
.A1(n_2177),
.A2(n_1516),
.B(n_1507),
.C(n_1587),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2183),
.Y(n_2213)
);

OAI22xp5_ASAP7_75t_L g2214 ( 
.A1(n_2177),
.A2(n_1507),
.B1(n_1577),
.B2(n_1518),
.Y(n_2214)
);

OAI22xp5_ASAP7_75t_L g2215 ( 
.A1(n_2177),
.A2(n_1518),
.B1(n_1524),
.B2(n_1547),
.Y(n_2215)
);

A2O1A1Ixp33_ASAP7_75t_L g2216 ( 
.A1(n_2201),
.A2(n_1678),
.B(n_1701),
.C(n_1547),
.Y(n_2216)
);

AOI311xp33_ASAP7_75t_L g2217 ( 
.A1(n_2195),
.A2(n_1530),
.A3(n_1579),
.B(n_1505),
.C(n_1519),
.Y(n_2217)
);

AOI222xp33_ASAP7_75t_L g2218 ( 
.A1(n_2202),
.A2(n_1599),
.B1(n_1601),
.B2(n_1600),
.C1(n_1562),
.C2(n_1552),
.Y(n_2218)
);

NAND2xp5_ASAP7_75t_L g2219 ( 
.A(n_2205),
.B(n_1684),
.Y(n_2219)
);

OAI211xp5_ASAP7_75t_SL g2220 ( 
.A1(n_2204),
.A2(n_1570),
.B(n_1596),
.C(n_1605),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_2199),
.Y(n_2221)
);

NAND4xp25_ASAP7_75t_L g2222 ( 
.A(n_2197),
.B(n_1572),
.C(n_1555),
.D(n_1694),
.Y(n_2222)
);

OAI211xp5_ASAP7_75t_L g2223 ( 
.A1(n_2206),
.A2(n_1701),
.B(n_1571),
.C(n_1547),
.Y(n_2223)
);

OAI22xp5_ASAP7_75t_L g2224 ( 
.A1(n_2198),
.A2(n_1524),
.B1(n_1572),
.B2(n_1519),
.Y(n_2224)
);

OAI22xp33_ASAP7_75t_L g2225 ( 
.A1(n_2203),
.A2(n_1559),
.B1(n_1553),
.B2(n_1554),
.Y(n_2225)
);

AOI221xp5_ASAP7_75t_SL g2226 ( 
.A1(n_2213),
.A2(n_1524),
.B1(n_1510),
.B2(n_1512),
.C(n_1511),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2208),
.B(n_1684),
.Y(n_2227)
);

O2A1O1Ixp33_ASAP7_75t_L g2228 ( 
.A1(n_2210),
.A2(n_1597),
.B(n_1552),
.C(n_1596),
.Y(n_2228)
);

AOI322xp5_ASAP7_75t_L g2229 ( 
.A1(n_2209),
.A2(n_1599),
.A3(n_1600),
.B1(n_1601),
.B2(n_1553),
.C1(n_1554),
.C2(n_1559),
.Y(n_2229)
);

NAND4xp25_ASAP7_75t_L g2230 ( 
.A(n_2200),
.B(n_1555),
.C(n_1591),
.D(n_1571),
.Y(n_2230)
);

OAI21x1_ASAP7_75t_SL g2231 ( 
.A1(n_2212),
.A2(n_2214),
.B(n_2215),
.Y(n_2231)
);

AOI22xp33_ASAP7_75t_L g2232 ( 
.A1(n_2211),
.A2(n_1554),
.B1(n_1559),
.B2(n_1553),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2221),
.B(n_2208),
.Y(n_2233)
);

NAND3xp33_ASAP7_75t_L g2234 ( 
.A(n_2219),
.B(n_2196),
.C(n_2207),
.Y(n_2234)
);

AOI221xp5_ASAP7_75t_L g2235 ( 
.A1(n_2220),
.A2(n_1570),
.B1(n_1596),
.B2(n_1605),
.C(n_1600),
.Y(n_2235)
);

OAI221xp5_ASAP7_75t_L g2236 ( 
.A1(n_2232),
.A2(n_1605),
.B1(n_1570),
.B2(n_1594),
.C(n_1699),
.Y(n_2236)
);

AOI221xp5_ASAP7_75t_L g2237 ( 
.A1(n_2227),
.A2(n_1601),
.B1(n_1599),
.B2(n_1594),
.C(n_1591),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_2231),
.Y(n_2238)
);

AOI211xp5_ASAP7_75t_L g2239 ( 
.A1(n_2222),
.A2(n_1555),
.B(n_1689),
.C(n_1688),
.Y(n_2239)
);

AOI221xp5_ASAP7_75t_SL g2240 ( 
.A1(n_2230),
.A2(n_1512),
.B1(n_1511),
.B2(n_1510),
.C(n_1513),
.Y(n_2240)
);

NOR2xp33_ASAP7_75t_L g2241 ( 
.A(n_2228),
.B(n_1689),
.Y(n_2241)
);

OAI211xp5_ASAP7_75t_SL g2242 ( 
.A1(n_2223),
.A2(n_214),
.B(n_218),
.C(n_211),
.Y(n_2242)
);

AOI22xp5_ASAP7_75t_L g2243 ( 
.A1(n_2234),
.A2(n_2225),
.B1(n_2226),
.B2(n_2218),
.Y(n_2243)
);

OAI221xp5_ASAP7_75t_L g2244 ( 
.A1(n_2238),
.A2(n_2233),
.B1(n_2242),
.B2(n_2241),
.C(n_2239),
.Y(n_2244)
);

NOR2xp33_ASAP7_75t_L g2245 ( 
.A(n_2235),
.B(n_2224),
.Y(n_2245)
);

INVx1_ASAP7_75t_L g2246 ( 
.A(n_2237),
.Y(n_2246)
);

NOR2x1_ASAP7_75t_L g2247 ( 
.A(n_2236),
.B(n_2216),
.Y(n_2247)
);

OAI22xp5_ASAP7_75t_L g2248 ( 
.A1(n_2240),
.A2(n_2217),
.B1(n_2229),
.B2(n_1591),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2238),
.B(n_1688),
.Y(n_2249)
);

OR3x1_ASAP7_75t_L g2250 ( 
.A(n_2238),
.B(n_1591),
.C(n_1513),
.Y(n_2250)
);

AOI22xp5_ASAP7_75t_L g2251 ( 
.A1(n_2234),
.A2(n_1594),
.B1(n_1699),
.B2(n_1604),
.Y(n_2251)
);

OA21x2_ASAP7_75t_L g2252 ( 
.A1(n_2244),
.A2(n_175),
.B(n_1699),
.Y(n_2252)
);

NAND4xp75_ASAP7_75t_L g2253 ( 
.A(n_2247),
.B(n_175),
.C(n_1604),
.D(n_1594),
.Y(n_2253)
);

NOR2xp67_ASAP7_75t_SL g2254 ( 
.A(n_2246),
.B(n_211),
.Y(n_2254)
);

NAND5xp2_ASAP7_75t_L g2255 ( 
.A(n_2243),
.B(n_1604),
.C(n_1594),
.D(n_218),
.E(n_214),
.Y(n_2255)
);

NAND4xp25_ASAP7_75t_SL g2256 ( 
.A(n_2249),
.B(n_1594),
.C(n_1604),
.D(n_218),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_2250),
.B(n_1594),
.Y(n_2257)
);

XNOR2x1_ASAP7_75t_L g2258 ( 
.A(n_2248),
.B(n_218),
.Y(n_2258)
);

INVx2_ASAP7_75t_L g2259 ( 
.A(n_2245),
.Y(n_2259)
);

INVx1_ASAP7_75t_L g2260 ( 
.A(n_2251),
.Y(n_2260)
);

AOI21xp5_ASAP7_75t_L g2261 ( 
.A1(n_2259),
.A2(n_218),
.B(n_214),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_2257),
.Y(n_2262)
);

INVx2_ASAP7_75t_L g2263 ( 
.A(n_2252),
.Y(n_2263)
);

NOR4xp25_ASAP7_75t_L g2264 ( 
.A(n_2260),
.B(n_2256),
.C(n_2258),
.D(n_2254),
.Y(n_2264)
);

INVx1_ASAP7_75t_SL g2265 ( 
.A(n_2253),
.Y(n_2265)
);

NAND3xp33_ASAP7_75t_SL g2266 ( 
.A(n_2255),
.B(n_1604),
.C(n_218),
.Y(n_2266)
);

OAI221xp5_ASAP7_75t_L g2267 ( 
.A1(n_2252),
.A2(n_214),
.B1(n_173),
.B2(n_180),
.C(n_177),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_2257),
.Y(n_2268)
);

XOR2x1_ASAP7_75t_L g2269 ( 
.A(n_2263),
.B(n_2268),
.Y(n_2269)
);

NAND2xp5_ASAP7_75t_L g2270 ( 
.A(n_2262),
.B(n_1604),
.Y(n_2270)
);

INVx3_ASAP7_75t_L g2271 ( 
.A(n_2265),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_2267),
.Y(n_2272)
);

OAI22xp5_ASAP7_75t_SL g2273 ( 
.A1(n_2271),
.A2(n_2264),
.B1(n_2266),
.B2(n_2261),
.Y(n_2273)
);

OAI22xp5_ASAP7_75t_L g2274 ( 
.A1(n_2272),
.A2(n_214),
.B1(n_173),
.B2(n_180),
.Y(n_2274)
);

OAI22xp5_ASAP7_75t_L g2275 ( 
.A1(n_2273),
.A2(n_2270),
.B1(n_2269),
.B2(n_214),
.Y(n_2275)
);

OAI211xp5_ASAP7_75t_SL g2276 ( 
.A1(n_2275),
.A2(n_2274),
.B(n_177),
.C(n_186),
.Y(n_2276)
);

AOI31xp33_ASAP7_75t_L g2277 ( 
.A1(n_2276),
.A2(n_1604),
.A3(n_180),
.B(n_177),
.Y(n_2277)
);

AOI22xp5_ASAP7_75t_L g2278 ( 
.A1(n_2277),
.A2(n_180),
.B1(n_177),
.B2(n_161),
.Y(n_2278)
);

OAI221xp5_ASAP7_75t_L g2279 ( 
.A1(n_2278),
.A2(n_161),
.B1(n_177),
.B2(n_186),
.C(n_180),
.Y(n_2279)
);

AOI22xp5_ASAP7_75t_L g2280 ( 
.A1(n_2279),
.A2(n_180),
.B1(n_177),
.B2(n_161),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2280),
.Y(n_2281)
);

OR2x6_ASAP7_75t_L g2282 ( 
.A(n_2281),
.B(n_161),
.Y(n_2282)
);

OAI22xp5_ASAP7_75t_SL g2283 ( 
.A1(n_2282),
.A2(n_180),
.B1(n_177),
.B2(n_161),
.Y(n_2283)
);

AOI22xp5_ASAP7_75t_L g2284 ( 
.A1(n_2283),
.A2(n_161),
.B1(n_177),
.B2(n_186),
.Y(n_2284)
);


endmodule