module fake_jpeg_21291_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx11_ASAP7_75t_SL g19 ( 
.A(n_12),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_9),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_18),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_39),
.B(n_40),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_9),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_26),
.B(n_0),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_48),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_26),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_26),
.Y(n_44)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_39),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_0),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_54),
.B(n_56),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_36),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_36),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_63),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_39),
.B(n_32),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_67),
.Y(n_73)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_68),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_64),
.A2(n_48),
.B1(n_45),
.B2(n_41),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_69),
.A2(n_20),
.B1(n_37),
.B2(n_52),
.Y(n_109)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_70),
.Y(n_100)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_71),
.A2(n_78),
.B1(n_80),
.B2(n_92),
.Y(n_113)
);

BUFx16f_ASAP7_75t_L g74 ( 
.A(n_53),
.Y(n_74)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_51),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_75),
.B(n_53),
.Y(n_120)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_76),
.Y(n_121)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_48),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_83),
.B(n_88),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g84 ( 
.A(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_84),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

CKINVDCx9p33_ASAP7_75t_R g87 ( 
.A(n_57),
.Y(n_87)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_87),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_57),
.B(n_41),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_55),
.A2(n_22),
.B1(n_27),
.B2(n_28),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_29),
.B(n_19),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_68),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_51),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_50),
.A2(n_27),
.B1(n_22),
.B2(n_20),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_98),
.B1(n_43),
.B2(n_44),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_46),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_95),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_58),
.B(n_46),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_49),
.B(n_44),
.Y(n_98)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_94),
.B(n_43),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_99),
.A2(n_66),
.B(n_21),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_83),
.B(n_43),
.C(n_44),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_98),
.C(n_77),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

OAI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_79),
.A2(n_45),
.B1(n_20),
.B2(n_22),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_104),
.A2(n_111),
.B1(n_123),
.B2(n_124),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_69),
.B(n_88),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_109),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_79),
.A2(n_37),
.B1(n_50),
.B2(n_38),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_58),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_114),
.B(n_115),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_58),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_117),
.A2(n_30),
.B1(n_29),
.B2(n_28),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_81),
.B(n_96),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_118),
.B(n_77),
.Y(n_149)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_97),
.Y(n_119)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_120),
.Y(n_154)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_125),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_91),
.A2(n_50),
.B1(n_27),
.B2(n_38),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_66),
.B1(n_67),
.B2(n_32),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_98),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_128),
.B(n_146),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_130),
.B(n_112),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_102),
.A2(n_71),
.B1(n_127),
.B2(n_100),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_134),
.A2(n_137),
.B(n_150),
.Y(n_165)
);

INVx3_ASAP7_75t_SL g138 ( 
.A(n_126),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_142),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_99),
.A2(n_82),
.B1(n_80),
.B2(n_78),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_140),
.A2(n_150),
.B(n_125),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_118),
.B(n_86),
.Y(n_141)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_107),
.B(n_106),
.Y(n_142)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_116),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_145),
.Y(n_181)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_113),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_144),
.Y(n_182)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_121),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_101),
.B(n_110),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_100),
.B(n_76),
.Y(n_147)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_147),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_127),
.B(n_77),
.Y(n_148)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_148),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_149),
.B(n_151),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_115),
.A2(n_2),
.B(n_3),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_17),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_109),
.A2(n_33),
.B1(n_23),
.B2(n_92),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_152),
.A2(n_124),
.B1(n_123),
.B2(n_111),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_102),
.B(n_74),
.Y(n_153)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_153),
.Y(n_175)
);

AND2x6_ASAP7_75t_L g155 ( 
.A(n_99),
.B(n_31),
.Y(n_155)
);

NAND2xp33_ASAP7_75t_R g162 ( 
.A(n_155),
.B(n_105),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_159),
.A2(n_160),
.B1(n_164),
.B2(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_135),
.A2(n_114),
.B1(n_103),
.B2(n_117),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_155),
.B(n_105),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_161),
.B(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_162),
.A2(n_165),
.B1(n_31),
.B2(n_34),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_122),
.B1(n_119),
.B2(n_108),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_108),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_176),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_167),
.B(n_185),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_174),
.B(n_179),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_129),
.A2(n_131),
.B1(n_132),
.B2(n_152),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_131),
.A2(n_23),
.B(n_33),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_129),
.A2(n_112),
.B1(n_121),
.B2(n_116),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_177),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_132),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_178),
.B(n_180),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_140),
.A2(n_21),
.B(n_35),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_146),
.B(n_24),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_144),
.A2(n_128),
.B1(n_149),
.B2(n_154),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_139),
.B(n_24),
.Y(n_184)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_184),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_130),
.B(n_31),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_134),
.A2(n_21),
.B(n_35),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_186),
.A2(n_73),
.B(n_35),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_137),
.A2(n_24),
.B1(n_25),
.B2(n_21),
.Y(n_187)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_187),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_188),
.B(n_156),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_140),
.B(n_74),
.C(n_47),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_140),
.C(n_156),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_190),
.B(n_185),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_167),
.B(n_156),
.C(n_138),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_47),
.C(n_53),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_195),
.A2(n_188),
.B1(n_183),
.B2(n_186),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_206),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_158),
.B(n_145),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_199),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_181),
.Y(n_201)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_201),
.Y(n_234)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_177),
.Y(n_202)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_202),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_208),
.B(n_215),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_138),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_176),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_85),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g237 ( 
.A(n_207),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_175),
.B(n_169),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_184),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_210),
.B(n_212),
.Y(n_221)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_166),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_213),
.B(n_214),
.Y(n_228)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g215 ( 
.A(n_164),
.B(n_34),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_72),
.A3(n_73),
.B1(n_34),
.B2(n_25),
.Y(n_217)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_161),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_219),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_168),
.B(n_72),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_195),
.A2(n_157),
.B(n_172),
.Y(n_222)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_222),
.A2(n_215),
.B(n_196),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_229),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_193),
.A2(n_179),
.B(n_174),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_224),
.B(n_226),
.Y(n_261)
);

AND2x4_ASAP7_75t_SL g227 ( 
.A(n_193),
.B(n_189),
.Y(n_227)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_227),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_211),
.B(n_170),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_191),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_231),
.B(n_236),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_211),
.B(n_170),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g255 ( 
.A(n_232),
.B(n_198),
.Y(n_255)
);

NAND3xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_180),
.C(n_10),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g249 ( 
.A(n_233),
.B(n_8),
.C(n_15),
.Y(n_249)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_157),
.B(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_216),
.A2(n_160),
.B1(n_178),
.B2(n_187),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_239),
.A2(n_206),
.B1(n_205),
.B2(n_196),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_200),
.A2(n_159),
.B1(n_182),
.B2(n_11),
.Y(n_241)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_241),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_200),
.A2(n_10),
.B1(n_16),
.B2(n_15),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_201),
.B(n_9),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_243),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_244),
.B(n_194),
.C(n_190),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_2),
.Y(n_245)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_245),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_249),
.B(n_230),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_254),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_225),
.A2(n_208),
.B1(n_205),
.B2(n_192),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_251),
.A2(n_259),
.B1(n_265),
.B2(n_224),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_252),
.A2(n_235),
.B1(n_227),
.B2(n_240),
.Y(n_271)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_229),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_255),
.B(n_257),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_232),
.B(n_214),
.C(n_213),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_258),
.B(n_264),
.C(n_227),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_220),
.A2(n_210),
.B1(n_192),
.B2(n_198),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_227),
.B(n_202),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_221),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_244),
.B(n_191),
.C(n_47),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_220),
.A2(n_8),
.B1(n_16),
.B2(n_14),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_234),
.Y(n_266)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_266),
.Y(n_276)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_270),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_262),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_260),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_281),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_256),
.Y(n_286)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_280),
.Y(n_295)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_222),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_236),
.Y(n_297)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_258),
.B(n_221),
.C(n_238),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_247),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_283),
.B(n_237),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_261),
.A2(n_231),
.B1(n_239),
.B2(n_228),
.Y(n_284)
);

OAI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_284),
.A2(n_260),
.B1(n_263),
.B2(n_246),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_296),
.B1(n_283),
.B2(n_276),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_288),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_280),
.B(n_245),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_287),
.B(n_294),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_256),
.Y(n_288)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_284),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_297),
.Y(n_305)
);

AOI321xp33_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_228),
.A3(n_267),
.B1(n_254),
.B2(n_225),
.C(n_255),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_291),
.A2(n_237),
.B(n_12),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_277),
.B(n_264),
.C(n_251),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_299),
.B(n_7),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_292),
.A2(n_295),
.B1(n_270),
.B2(n_290),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_308),
.B1(n_311),
.B2(n_307),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_278),
.C(n_282),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_302),
.B(n_306),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_303),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_293),
.A2(n_282),
.B1(n_268),
.B2(n_238),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_304),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_312),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_298),
.A2(n_7),
.B1(n_16),
.B2(n_14),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_6),
.B(n_14),
.Y(n_309)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_309),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_299),
.B(n_6),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_311),
.B(n_5),
.Y(n_315)
);

OR2x2_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_5),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_313),
.B(n_315),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_305),
.B(n_12),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_319),
.B(n_321),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_13),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_314),
.B(n_310),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_322),
.B(n_323),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_316),
.B(n_304),
.Y(n_323)
);

INVx11_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_324),
.A2(n_326),
.B(n_328),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_312),
.C(n_302),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g328 ( 
.A1(n_318),
.A2(n_300),
.B(n_13),
.Y(n_328)
);

XNOR2x1_ASAP7_75t_L g329 ( 
.A(n_327),
.B(n_300),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_329),
.Y(n_332)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_332),
.A2(n_331),
.A3(n_318),
.B1(n_330),
.B2(n_325),
.C1(n_317),
.C2(n_4),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_333),
.Y(n_334)
);

AOI322xp5_ASAP7_75t_L g335 ( 
.A1(n_334),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_47),
.C1(n_325),
.C2(n_331),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_3),
.B1(n_4),
.B2(n_47),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_47),
.Y(n_338)
);


endmodule