module fake_netlist_6_4595_n_1004 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_209, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_210, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_211, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_1004);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_209;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_210;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_211;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1004;

wire n_992;
wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_968;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_465;
wire n_367;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_933;
wire n_740;
wire n_578;
wire n_703;
wire n_1003;
wire n_365;
wire n_978;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_951;
wire n_783;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_994;
wire n_677;
wire n_969;
wire n_988;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_974;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_955;
wire n_865;
wire n_893;
wire n_214;
wire n_925;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_935;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_963;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_300;
wire n_222;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_996;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_923;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_948;
wire n_466;
wire n_704;
wire n_918;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_945;
wire n_977;
wire n_603;
wire n_991;
wire n_957;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_987;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_525;
wire n_842;
wire n_758;
wire n_611;
wire n_943;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_989;
wire n_797;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_795;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_953;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_930;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_947;
wire n_236;
wire n_653;
wire n_887;
wire n_908;
wire n_752;
wire n_944;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_976;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_926;
wire n_927;
wire n_839;
wire n_986;
wire n_734;
wire n_708;
wire n_919;
wire n_402;
wire n_352;
wire n_917;
wire n_668;
wire n_478;
wire n_626;
wire n_990;
wire n_574;
wire n_800;
wire n_779;
wire n_929;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_921;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_937;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_998;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_492;
wire n_972;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_962;
wire n_1000;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_936;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_984;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_916;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_934;
wire n_755;
wire n_931;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_958;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_942;
wire n_880;
wire n_792;
wire n_476;
wire n_981;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_985;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_939;
wire n_997;
wire n_821;
wire n_325;
wire n_938;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_964;
wire n_982;
wire n_561;
wire n_477;
wire n_549;
wire n_980;
wire n_533;
wire n_954;
wire n_408;
wire n_932;
wire n_806;
wire n_864;
wire n_879;
wire n_959;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_979;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_523;
wire n_322;
wire n_707;
wire n_993;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_966;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_941;
wire n_975;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_970;
wire n_560;
wire n_753;
wire n_642;
wire n_995;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_973;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_967;
wire n_775;
wire n_922;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_915;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_920;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_928;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_1002;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_965;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_983;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_688;
wire n_722;
wire n_961;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_295;
wire n_385;
wire n_701;
wire n_817;
wire n_950;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_960;
wire n_956;
wire n_531;
wire n_827;
wire n_1001;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_949;
wire n_678;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_37),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_203),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_165),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_84),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_127),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_102),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_105),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_110),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_6),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g222 ( 
.A(n_144),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_52),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_128),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_58),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_83),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_106),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_81),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_134),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_148),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_19),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_0),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_178),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_139),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_166),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_185),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_210),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_72),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_13),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_187),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_138),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_13),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_177),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_107),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g247 ( 
.A(n_183),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_184),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_55),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_172),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_77),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_111),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_173),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_20),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_193),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_6),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_3),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_201),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_133),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_153),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_195),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_51),
.Y(n_262)
);

INVx1_ASAP7_75t_SL g263 ( 
.A(n_1),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_117),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_3),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_176),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_5),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_46),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_180),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_98),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_169),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_130),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_108),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_190),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_206),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_186),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_11),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_156),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_189),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_119),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_49),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_33),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_32),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_171),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_9),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_71),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_89),
.Y(n_290)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_66),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_174),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_199),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_125),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_68),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_80),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_48),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_95),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_18),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_73),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_62),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_216),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_212),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_240),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_213),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_214),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_215),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_240),
.Y(n_308)
);

NAND2xp33_ASAP7_75t_R g309 ( 
.A(n_262),
.B(n_0),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_240),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_240),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_217),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_219),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g314 ( 
.A(n_293),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_218),
.Y(n_315)
);

HB1xp67_ASAP7_75t_L g316 ( 
.A(n_221),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_269),
.B(n_1),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_257),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_224),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_254),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_279),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_247),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g324 ( 
.A(n_216),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_220),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_225),
.Y(n_327)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_232),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_223),
.Y(n_329)
);

NOR2xp67_ASAP7_75t_L g330 ( 
.A(n_269),
.B(n_2),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_257),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_237),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_288),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_255),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_233),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_243),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_249),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_250),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_251),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_288),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_226),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_261),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_255),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_283),
.B(n_2),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_273),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_266),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_268),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_273),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_270),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g351 ( 
.A(n_242),
.Y(n_351)
);

INVxp67_ASAP7_75t_SL g352 ( 
.A(n_272),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_256),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_227),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_303),
.B(n_283),
.Y(n_355)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_304),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_342),
.Y(n_357)
);

INVx3_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

HB1xp67_ASAP7_75t_L g359 ( 
.A(n_316),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_310),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_311),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_326),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_329),
.Y(n_363)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_332),
.Y(n_364)
);

AND3x1_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_291),
.C(n_284),
.Y(n_365)
);

AND2x6_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_284),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_320),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_344),
.B(n_265),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_321),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_336),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_337),
.Y(n_371)
);

HB1xp67_ASAP7_75t_L g372 ( 
.A(n_328),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_322),
.Y(n_373)
);

AND2x4_ASAP7_75t_L g374 ( 
.A(n_352),
.B(n_291),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_305),
.B(n_285),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g376 ( 
.A(n_323),
.B(n_222),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_338),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_295),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_343),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_347),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g382 ( 
.A(n_302),
.B(n_222),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_348),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_350),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_325),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_335),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_330),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_307),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_314),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_312),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

BUFx2_ASAP7_75t_L g392 ( 
.A(n_351),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_319),
.B(n_297),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_327),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_341),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_351),
.B(n_298),
.Y(n_397)
);

BUFx6f_ASAP7_75t_L g398 ( 
.A(n_309),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_353),
.B(n_228),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_353),
.B(n_253),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_324),
.B(n_222),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_344),
.A2(n_267),
.B1(n_299),
.B2(n_274),
.Y(n_402)
);

INVx3_ASAP7_75t_L g403 ( 
.A(n_313),
.Y(n_403)
);

INVx3_ASAP7_75t_L g404 ( 
.A(n_334),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_346),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_346),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_349),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_349),
.B(n_4),
.Y(n_408)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_318),
.B(n_4),
.Y(n_409)
);

NAND2x1p5_ASAP7_75t_L g410 ( 
.A(n_318),
.B(n_229),
.Y(n_410)
);

INVx3_ASAP7_75t_L g411 ( 
.A(n_331),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_388),
.B(n_230),
.Y(n_412)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_357),
.B(n_231),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g414 ( 
.A1(n_366),
.A2(n_276),
.B1(n_235),
.B2(n_236),
.Y(n_414)
);

AND2x2_ASAP7_75t_SL g415 ( 
.A(n_365),
.B(n_7),
.Y(n_415)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_359),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_381),
.Y(n_417)
);

OAI22xp33_ASAP7_75t_L g418 ( 
.A1(n_382),
.A2(n_278),
.B1(n_238),
.B2(n_239),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_356),
.Y(n_419)
);

INVx8_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_381),
.Y(n_421)
);

INVx4_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

BUFx3_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_366),
.A2(n_280),
.B1(n_241),
.B2(n_245),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_234),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_367),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_356),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_367),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_388),
.B(n_246),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_398),
.B(n_7),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_390),
.B(n_394),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_369),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g433 ( 
.A(n_363),
.Y(n_433)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_398),
.Y(n_435)
);

NOR2xp67_ASAP7_75t_L g436 ( 
.A(n_400),
.B(n_248),
.Y(n_436)
);

INVx2_ASAP7_75t_SL g437 ( 
.A(n_372),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

BUFx3_ASAP7_75t_L g439 ( 
.A(n_363),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_373),
.Y(n_440)
);

NAND3x1_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_333),
.C(n_331),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_373),
.Y(n_442)
);

BUFx3_ASAP7_75t_L g443 ( 
.A(n_363),
.Y(n_443)
);

BUFx10_ASAP7_75t_L g444 ( 
.A(n_397),
.Y(n_444)
);

INVx5_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g446 ( 
.A(n_398),
.B(n_252),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_398),
.B(n_258),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_371),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_366),
.A2(n_374),
.B1(n_355),
.B2(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_371),
.Y(n_451)
);

INVx4_ASAP7_75t_L g452 ( 
.A(n_371),
.Y(n_452)
);

AND3x2_ASAP7_75t_L g453 ( 
.A(n_395),
.B(n_394),
.C(n_390),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_361),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_371),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_358),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_375),
.B(n_259),
.Y(n_457)
);

BUFx3_ASAP7_75t_L g458 ( 
.A(n_380),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_380),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_380),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_379),
.B(n_393),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_368),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_396),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_380),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_380),
.Y(n_465)
);

BUFx4f_ASAP7_75t_L g466 ( 
.A(n_395),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_386),
.B(n_260),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_358),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_383),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_358),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_392),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_383),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_383),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_376),
.B(n_264),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_396),
.B(n_376),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_374),
.B(n_271),
.Y(n_476)
);

INVxp67_ASAP7_75t_L g477 ( 
.A(n_387),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g478 ( 
.A(n_397),
.Y(n_478)
);

AND2x2_ASAP7_75t_SL g479 ( 
.A(n_374),
.B(n_8),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_383),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_383),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_366),
.B(n_275),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_391),
.B(n_277),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_366),
.B(n_281),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_384),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_362),
.B(n_282),
.Y(n_487)
);

HB1xp67_ASAP7_75t_L g488 ( 
.A(n_478),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_471),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_427),
.Y(n_490)
);

BUFx8_ASAP7_75t_L g491 ( 
.A(n_462),
.Y(n_491)
);

AND2x4_ASAP7_75t_L g492 ( 
.A(n_417),
.B(n_385),
.Y(n_492)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_471),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_427),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_419),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_434),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_421),
.B(n_385),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_L g498 ( 
.A1(n_461),
.A2(n_435),
.B1(n_475),
.B2(n_431),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_435),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_416),
.Y(n_500)
);

NAND2x1p5_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_403),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g502 ( 
.A(n_413),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_426),
.Y(n_503)
);

NAND2x1p5_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_403),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_461),
.B(n_384),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_454),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_428),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_432),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_438),
.Y(n_509)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_449),
.A2(n_362),
.B(n_364),
.C(n_397),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_449),
.B(n_384),
.Y(n_511)
);

AO22x2_ASAP7_75t_L g512 ( 
.A1(n_479),
.A2(n_409),
.B1(n_401),
.B2(n_402),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_457),
.B(n_384),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_440),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_468),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_468),
.Y(n_516)
);

AND2x4_ASAP7_75t_L g517 ( 
.A(n_442),
.B(n_370),
.Y(n_517)
);

AO22x2_ASAP7_75t_L g518 ( 
.A1(n_479),
.A2(n_409),
.B1(n_406),
.B2(n_407),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_470),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_457),
.B(n_362),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_425),
.B(n_387),
.Y(n_521)
);

OAI221xp5_ASAP7_75t_L g522 ( 
.A1(n_414),
.A2(n_370),
.B1(n_377),
.B2(n_378),
.C(n_364),
.Y(n_522)
);

NAND2x1p5_ASAP7_75t_L g523 ( 
.A(n_466),
.B(n_403),
.Y(n_523)
);

NOR2xp67_ASAP7_75t_L g524 ( 
.A(n_437),
.B(n_364),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_470),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_420),
.B(n_436),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_456),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_477),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_477),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_483),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_420),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_453),
.B(n_377),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_L g533 ( 
.A(n_420),
.B(n_286),
.Y(n_533)
);

NAND2x1p5_ASAP7_75t_L g534 ( 
.A(n_466),
.B(n_378),
.Y(n_534)
);

INVxp67_ASAP7_75t_L g535 ( 
.A(n_467),
.Y(n_535)
);

OAI221xp5_ASAP7_75t_L g536 ( 
.A1(n_414),
.A2(n_360),
.B1(n_287),
.B2(n_301),
.C(n_289),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g537 ( 
.A1(n_424),
.A2(n_360),
.B1(n_410),
.B2(n_292),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_L g538 ( 
.A(n_483),
.B(n_410),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_430),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_412),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_450),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_455),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_459),
.Y(n_543)
);

AO22x2_ASAP7_75t_L g544 ( 
.A1(n_430),
.A2(n_415),
.B1(n_406),
.B2(n_407),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_460),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_464),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVxp67_ASAP7_75t_L g548 ( 
.A(n_474),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_473),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g550 ( 
.A(n_444),
.Y(n_550)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_412),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_481),
.Y(n_552)
);

INVxp67_ASAP7_75t_L g553 ( 
.A(n_429),
.Y(n_553)
);

A2O1A1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_424),
.A2(n_290),
.B(n_294),
.C(n_296),
.Y(n_554)
);

BUFx8_ASAP7_75t_L g555 ( 
.A(n_429),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_423),
.Y(n_556)
);

BUFx8_ASAP7_75t_L g557 ( 
.A(n_441),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_485),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_486),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_476),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

NAND2x1p5_ASAP7_75t_L g562 ( 
.A(n_445),
.B(n_404),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_446),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_423),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_446),
.Y(n_565)
);

OAI22xp5_ASAP7_75t_L g566 ( 
.A1(n_447),
.A2(n_300),
.B1(n_410),
.B2(n_404),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

OAI221xp5_ASAP7_75t_L g568 ( 
.A1(n_447),
.A2(n_408),
.B1(n_368),
.B2(n_392),
.C(n_404),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_418),
.B(n_333),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_439),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_451),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_444),
.B(n_411),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_551),
.B(n_453),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_553),
.B(n_439),
.Y(n_574)
);

NAND2xp33_ASAP7_75t_SL g575 ( 
.A(n_540),
.B(n_408),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_498),
.B(n_530),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_538),
.B(n_415),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_521),
.B(n_411),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_539),
.B(n_411),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_535),
.B(n_418),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_560),
.B(n_405),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_443),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_548),
.B(n_445),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_505),
.B(n_487),
.Y(n_584)
);

AND2x4_ASAP7_75t_L g585 ( 
.A(n_503),
.B(n_443),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_561),
.B(n_445),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_563),
.B(n_445),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_482),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_528),
.B(n_529),
.Y(n_589)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_500),
.B(n_340),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_524),
.B(n_502),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_534),
.B(n_484),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_532),
.B(n_520),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_532),
.B(n_433),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_568),
.B(n_340),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_SL g596 ( 
.A(n_537),
.B(n_433),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_488),
.B(n_433),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_517),
.B(n_433),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_517),
.B(n_448),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_492),
.B(n_448),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_SL g601 ( 
.A(n_566),
.B(n_572),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g602 ( 
.A(n_492),
.B(n_448),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_507),
.B(n_458),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_508),
.B(n_458),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_497),
.B(n_448),
.Y(n_605)
);

NAND2xp33_ASAP7_75t_SL g606 ( 
.A(n_531),
.B(n_480),
.Y(n_606)
);

NAND2xp33_ASAP7_75t_SL g607 ( 
.A(n_526),
.B(n_480),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_497),
.B(n_523),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_509),
.B(n_472),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_514),
.B(n_472),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_SL g611 ( 
.A(n_501),
.B(n_480),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_504),
.B(n_513),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_SL g613 ( 
.A(n_550),
.B(n_480),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_SL g614 ( 
.A(n_511),
.B(n_489),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_SL g615 ( 
.A(n_569),
.B(n_422),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_510),
.B(n_422),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_SL g617 ( 
.A(n_555),
.B(n_452),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_555),
.B(n_452),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_554),
.B(n_469),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_SL g620 ( 
.A(n_495),
.B(n_469),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_496),
.B(n_30),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_494),
.B(n_8),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_SL g623 ( 
.A(n_506),
.B(n_31),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_562),
.B(n_34),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_527),
.B(n_36),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_556),
.B(n_39),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_564),
.B(n_40),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_570),
.B(n_41),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_494),
.B(n_42),
.Y(n_629)
);

NAND2xp33_ASAP7_75t_SL g630 ( 
.A(n_541),
.B(n_542),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_490),
.B(n_43),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_SL g632 ( 
.A(n_516),
.B(n_44),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_516),
.B(n_9),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_545),
.B(n_45),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_519),
.B(n_10),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_546),
.B(n_47),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_547),
.B(n_50),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_549),
.B(n_53),
.Y(n_638)
);

NAND2xp33_ASAP7_75t_SL g639 ( 
.A(n_541),
.B(n_10),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_576),
.B(n_544),
.Y(n_640)
);

O2A1O1Ixp5_ASAP7_75t_L g641 ( 
.A1(n_619),
.A2(n_542),
.B(n_543),
.C(n_559),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_584),
.B(n_544),
.Y(n_642)
);

AOI21xp5_ASAP7_75t_SL g643 ( 
.A1(n_616),
.A2(n_522),
.B(n_525),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_577),
.B(n_493),
.Y(n_644)
);

AO31x2_ASAP7_75t_L g645 ( 
.A1(n_633),
.A2(n_543),
.A3(n_552),
.B(n_558),
.Y(n_645)
);

OAI21x1_ASAP7_75t_L g646 ( 
.A1(n_588),
.A2(n_571),
.B(n_567),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_580),
.A2(n_536),
.B(n_515),
.C(n_567),
.Y(n_647)
);

AOI221x1_ASAP7_75t_L g648 ( 
.A1(n_601),
.A2(n_512),
.B1(n_518),
.B2(n_571),
.C(n_533),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_603),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_595),
.B(n_590),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_592),
.A2(n_512),
.B(n_518),
.Y(n_651)
);

OAI21x1_ASAP7_75t_L g652 ( 
.A1(n_604),
.A2(n_115),
.B(n_211),
.Y(n_652)
);

AOI21xp5_ASAP7_75t_L g653 ( 
.A1(n_612),
.A2(n_114),
.B(n_209),
.Y(n_653)
);

AOI21xp5_ASAP7_75t_L g654 ( 
.A1(n_596),
.A2(n_113),
.B(n_208),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_589),
.B(n_491),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_593),
.B(n_557),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_609),
.Y(n_657)
);

AOI221x1_ASAP7_75t_L g658 ( 
.A1(n_614),
.A2(n_557),
.B1(n_12),
.B2(n_14),
.C(n_15),
.Y(n_658)
);

BUFx6f_ASAP7_75t_L g659 ( 
.A(n_574),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_585),
.B(n_491),
.Y(n_660)
);

OAI21xp5_ASAP7_75t_L g661 ( 
.A1(n_587),
.A2(n_109),
.B(n_205),
.Y(n_661)
);

A2O1A1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_630),
.A2(n_11),
.B(n_12),
.C(n_14),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_573),
.B(n_54),
.Y(n_663)
);

AO22x2_ASAP7_75t_L g664 ( 
.A1(n_573),
.A2(n_615),
.B1(n_608),
.B2(n_617),
.Y(n_664)
);

A2O1A1Ixp33_ASAP7_75t_L g665 ( 
.A1(n_639),
.A2(n_15),
.B(n_16),
.C(n_17),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_607),
.A2(n_118),
.B(n_204),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_585),
.B(n_16),
.Y(n_667)
);

OAI21xp5_ASAP7_75t_L g668 ( 
.A1(n_586),
.A2(n_610),
.B(n_622),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_578),
.B(n_17),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_574),
.B(n_18),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_582),
.Y(n_671)
);

INVx2_ASAP7_75t_L g672 ( 
.A(n_582),
.Y(n_672)
);

NAND3xp33_ASAP7_75t_L g673 ( 
.A(n_579),
.B(n_19),
.C(n_20),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_591),
.B(n_21),
.Y(n_674)
);

OAI21xp5_ASAP7_75t_L g675 ( 
.A1(n_583),
.A2(n_121),
.B(n_202),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_594),
.B(n_21),
.Y(n_676)
);

O2A1O1Ixp5_ASAP7_75t_L g677 ( 
.A1(n_606),
.A2(n_122),
.B(n_200),
.C(n_198),
.Y(n_677)
);

AOI22xp5_ASAP7_75t_L g678 ( 
.A1(n_625),
.A2(n_116),
.B1(n_197),
.B2(n_194),
.Y(n_678)
);

AOI21xp5_ASAP7_75t_L g679 ( 
.A1(n_598),
.A2(n_112),
.B(n_191),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_635),
.Y(n_680)
);

BUFx6f_ASAP7_75t_L g681 ( 
.A(n_625),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_599),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_575),
.B(n_22),
.Y(n_683)
);

OAI21xp5_ASAP7_75t_L g684 ( 
.A1(n_632),
.A2(n_104),
.B(n_188),
.Y(n_684)
);

AOI21x1_ASAP7_75t_L g685 ( 
.A1(n_629),
.A2(n_103),
.B(n_182),
.Y(n_685)
);

NAND2x1p5_ASAP7_75t_L g686 ( 
.A(n_618),
.B(n_56),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_600),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_613),
.Y(n_688)
);

AO31x2_ASAP7_75t_L g689 ( 
.A1(n_620),
.A2(n_22),
.A3(n_23),
.B(n_24),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_602),
.B(n_23),
.Y(n_690)
);

OAI22xp5_ASAP7_75t_L g691 ( 
.A1(n_605),
.A2(n_120),
.B1(n_181),
.B2(n_175),
.Y(n_691)
);

AOI21xp5_ASAP7_75t_L g692 ( 
.A1(n_611),
.A2(n_101),
.B(n_170),
.Y(n_692)
);

INVx5_ASAP7_75t_L g693 ( 
.A(n_581),
.Y(n_693)
);

OAI21x1_ASAP7_75t_L g694 ( 
.A1(n_624),
.A2(n_597),
.B(n_631),
.Y(n_694)
);

AOI21xp5_ASAP7_75t_L g695 ( 
.A1(n_638),
.A2(n_100),
.B(n_168),
.Y(n_695)
);

BUFx3_ASAP7_75t_L g696 ( 
.A(n_626),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_646),
.Y(n_697)
);

AO21x2_ASAP7_75t_L g698 ( 
.A1(n_668),
.A2(n_637),
.B(n_636),
.Y(n_698)
);

OAI22xp5_ASAP7_75t_L g699 ( 
.A1(n_681),
.A2(n_634),
.B1(n_628),
.B2(n_627),
.Y(n_699)
);

AO21x2_ASAP7_75t_L g700 ( 
.A1(n_643),
.A2(n_623),
.B(n_621),
.Y(n_700)
);

NOR2xp67_ASAP7_75t_L g701 ( 
.A(n_693),
.B(n_57),
.Y(n_701)
);

OA21x2_ASAP7_75t_L g702 ( 
.A1(n_641),
.A2(n_99),
.B(n_167),
.Y(n_702)
);

OAI21x1_ASAP7_75t_L g703 ( 
.A1(n_694),
.A2(n_97),
.B(n_164),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_680),
.B(n_24),
.Y(n_704)
);

OAI222xp33_ASAP7_75t_L g705 ( 
.A1(n_678),
.A2(n_651),
.B1(n_640),
.B2(n_683),
.C1(n_642),
.C2(n_650),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_687),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_645),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_682),
.Y(n_708)
);

BUFx6f_ASAP7_75t_L g709 ( 
.A(n_659),
.Y(n_709)
);

NAND2x1p5_ASAP7_75t_L g710 ( 
.A(n_659),
.B(n_123),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_647),
.A2(n_96),
.B(n_163),
.Y(n_711)
);

OAI221xp5_ASAP7_75t_L g712 ( 
.A1(n_644),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.C(n_28),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_645),
.Y(n_713)
);

BUFx6f_ASAP7_75t_L g714 ( 
.A(n_659),
.Y(n_714)
);

BUFx6f_ASAP7_75t_L g715 ( 
.A(n_681),
.Y(n_715)
);

AND2x4_ASAP7_75t_L g716 ( 
.A(n_681),
.B(n_207),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_649),
.Y(n_717)
);

INVxp33_ASAP7_75t_L g718 ( 
.A(n_655),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_669),
.B(n_25),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_652),
.A2(n_94),
.B(n_161),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_657),
.B(n_671),
.Y(n_721)
);

AOI221xp5_ASAP7_75t_L g722 ( 
.A1(n_673),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.C(n_29),
.Y(n_722)
);

OR2x2_ASAP7_75t_L g723 ( 
.A(n_672),
.B(n_660),
.Y(n_723)
);

INVx1_ASAP7_75t_SL g724 ( 
.A(n_674),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_663),
.A2(n_29),
.B1(n_59),
.B2(n_60),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_648),
.B(n_61),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_685),
.Y(n_727)
);

OAI21x1_ASAP7_75t_L g728 ( 
.A1(n_654),
.A2(n_63),
.B(n_64),
.Y(n_728)
);

OAI21xp5_ASAP7_75t_L g729 ( 
.A1(n_690),
.A2(n_65),
.B(n_67),
.Y(n_729)
);

NAND3xp33_ASAP7_75t_L g730 ( 
.A(n_658),
.B(n_69),
.C(n_70),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_688),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_693),
.B(n_74),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_670),
.B(n_75),
.Y(n_733)
);

BUFx6f_ASAP7_75t_L g734 ( 
.A(n_693),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_656),
.B(n_76),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_667),
.Y(n_736)
);

AO31x2_ASAP7_75t_L g737 ( 
.A1(n_662),
.A2(n_665),
.A3(n_666),
.B(n_653),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_676),
.Y(n_738)
);

AND2x2_ASAP7_75t_L g739 ( 
.A(n_664),
.B(n_78),
.Y(n_739)
);

AOI21xp5_ASAP7_75t_L g740 ( 
.A1(n_684),
.A2(n_79),
.B(n_82),
.Y(n_740)
);

NAND2x1p5_ASAP7_75t_L g741 ( 
.A(n_696),
.B(n_85),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_673),
.Y(n_742)
);

AOI221xp5_ASAP7_75t_L g743 ( 
.A1(n_664),
.A2(n_86),
.B1(n_87),
.B2(n_88),
.C(n_90),
.Y(n_743)
);

AND2x4_ASAP7_75t_L g744 ( 
.A(n_678),
.B(n_162),
.Y(n_744)
);

BUFx3_ASAP7_75t_L g745 ( 
.A(n_686),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_675),
.A2(n_91),
.B1(n_92),
.B2(n_93),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_661),
.B(n_160),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_707),
.Y(n_748)
);

INVx3_ASAP7_75t_L g749 ( 
.A(n_728),
.Y(n_749)
);

NAND2x1_ASAP7_75t_L g750 ( 
.A(n_697),
.B(n_684),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_731),
.Y(n_751)
);

INVx3_ASAP7_75t_L g752 ( 
.A(n_703),
.Y(n_752)
);

OAI21x1_ASAP7_75t_L g753 ( 
.A1(n_720),
.A2(n_677),
.B(n_692),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_707),
.Y(n_754)
);

AND2x4_ASAP7_75t_L g755 ( 
.A(n_744),
.B(n_679),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_713),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_713),
.Y(n_757)
);

AOI211xp5_ASAP7_75t_L g758 ( 
.A1(n_712),
.A2(n_691),
.B(n_695),
.C(n_689),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_697),
.Y(n_759)
);

INVx4_ASAP7_75t_L g760 ( 
.A(n_744),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_742),
.B(n_689),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_706),
.Y(n_762)
);

OR2x2_ASAP7_75t_L g763 ( 
.A(n_724),
.B(n_689),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_717),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_708),
.Y(n_765)
);

INVx3_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

BUFx3_ASAP7_75t_L g767 ( 
.A(n_734),
.Y(n_767)
);

HB1xp67_ASAP7_75t_L g768 ( 
.A(n_723),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_727),
.Y(n_769)
);

BUFx3_ASAP7_75t_L g770 ( 
.A(n_734),
.Y(n_770)
);

OR2x2_ASAP7_75t_L g771 ( 
.A(n_738),
.B(n_124),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_737),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_721),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_734),
.Y(n_774)
);

AO31x2_ASAP7_75t_L g775 ( 
.A1(n_711),
.A2(n_126),
.A3(n_129),
.B(n_131),
.Y(n_775)
);

OAI21x1_ASAP7_75t_L g776 ( 
.A1(n_702),
.A2(n_132),
.B(n_135),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_739),
.B(n_136),
.Y(n_777)
);

BUFx2_ASAP7_75t_L g778 ( 
.A(n_737),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_726),
.Y(n_779)
);

OR2x2_ASAP7_75t_L g780 ( 
.A(n_736),
.B(n_704),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_737),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_716),
.Y(n_782)
);

OAI21x1_ASAP7_75t_L g783 ( 
.A1(n_740),
.A2(n_137),
.B(n_140),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_698),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_719),
.B(n_159),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_730),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_700),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_709),
.Y(n_788)
);

OR2x2_ASAP7_75t_L g789 ( 
.A(n_733),
.B(n_141),
.Y(n_789)
);

OA21x2_ASAP7_75t_L g790 ( 
.A1(n_705),
.A2(n_142),
.B(n_143),
.Y(n_790)
);

AND2x4_ASAP7_75t_L g791 ( 
.A(n_747),
.B(n_145),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_700),
.Y(n_792)
);

AOI21x1_ASAP7_75t_L g793 ( 
.A1(n_699),
.A2(n_146),
.B(n_147),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_747),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_709),
.Y(n_795)
);

BUFx12f_ASAP7_75t_L g796 ( 
.A(n_709),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_729),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_710),
.Y(n_798)
);

HB1xp67_ASAP7_75t_L g799 ( 
.A(n_714),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_732),
.Y(n_800)
);

OR2x2_ASAP7_75t_L g801 ( 
.A(n_718),
.B(n_149),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_732),
.Y(n_802)
);

INVx2_ASAP7_75t_L g803 ( 
.A(n_714),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_714),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_701),
.Y(n_805)
);

OR2x4_ASAP7_75t_L g806 ( 
.A(n_801),
.B(n_715),
.Y(n_806)
);

NAND2xp33_ASAP7_75t_R g807 ( 
.A(n_790),
.B(n_735),
.Y(n_807)
);

AND2x4_ASAP7_75t_L g808 ( 
.A(n_800),
.B(n_745),
.Y(n_808)
);

BUFx10_ASAP7_75t_L g809 ( 
.A(n_788),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_773),
.B(n_722),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_780),
.B(n_735),
.Y(n_811)
);

CKINVDCx11_ASAP7_75t_R g812 ( 
.A(n_751),
.Y(n_812)
);

AND2x4_ASAP7_75t_L g813 ( 
.A(n_800),
.B(n_715),
.Y(n_813)
);

INVxp67_ASAP7_75t_L g814 ( 
.A(n_768),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_R g815 ( 
.A(n_788),
.B(n_715),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_773),
.B(n_741),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_R g817 ( 
.A(n_790),
.B(n_150),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_780),
.B(n_764),
.Y(n_818)
);

AND2x4_ASAP7_75t_L g819 ( 
.A(n_802),
.B(n_725),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_R g820 ( 
.A(n_790),
.B(n_151),
.Y(n_820)
);

NAND2xp33_ASAP7_75t_R g821 ( 
.A(n_790),
.B(n_152),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_764),
.B(n_743),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_760),
.B(n_746),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_R g824 ( 
.A(n_791),
.B(n_154),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_777),
.B(n_155),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_771),
.B(n_157),
.Y(n_826)
);

AND2x4_ASAP7_75t_L g827 ( 
.A(n_802),
.B(n_760),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_777),
.B(n_158),
.Y(n_828)
);

BUFx3_ASAP7_75t_L g829 ( 
.A(n_751),
.Y(n_829)
);

NAND2xp33_ASAP7_75t_R g830 ( 
.A(n_791),
.B(n_766),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_760),
.B(n_782),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_760),
.B(n_782),
.Y(n_832)
);

CKINVDCx20_ASAP7_75t_R g833 ( 
.A(n_767),
.Y(n_833)
);

NOR2xp33_ASAP7_75t_R g834 ( 
.A(n_796),
.B(n_766),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_771),
.B(n_765),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_796),
.Y(n_836)
);

BUFx3_ASAP7_75t_L g837 ( 
.A(n_767),
.Y(n_837)
);

OR2x2_ASAP7_75t_L g838 ( 
.A(n_763),
.B(n_762),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_798),
.B(n_805),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_754),
.Y(n_840)
);

NAND2xp33_ASAP7_75t_R g841 ( 
.A(n_791),
.B(n_766),
.Y(n_841)
);

INVx2_ASAP7_75t_L g842 ( 
.A(n_762),
.Y(n_842)
);

NAND2xp33_ASAP7_75t_R g843 ( 
.A(n_791),
.B(n_782),
.Y(n_843)
);

OR2x2_ASAP7_75t_L g844 ( 
.A(n_763),
.B(n_779),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_779),
.B(n_794),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_765),
.Y(n_846)
);

INVxp67_ASAP7_75t_L g847 ( 
.A(n_799),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_798),
.B(n_794),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_805),
.B(n_755),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_755),
.B(n_801),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_769),
.Y(n_851)
);

AND2x2_ASAP7_75t_L g852 ( 
.A(n_840),
.B(n_778),
.Y(n_852)
);

OR2x2_ASAP7_75t_L g853 ( 
.A(n_844),
.B(n_772),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_818),
.B(n_761),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_842),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_816),
.B(n_755),
.Y(n_856)
);

INVx2_ASAP7_75t_L g857 ( 
.A(n_846),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_838),
.Y(n_858)
);

INVx2_ASAP7_75t_L g859 ( 
.A(n_851),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_814),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_845),
.B(n_778),
.Y(n_861)
);

OR2x2_ASAP7_75t_L g862 ( 
.A(n_850),
.B(n_772),
.Y(n_862)
);

INVx2_ASAP7_75t_L g863 ( 
.A(n_849),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_848),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_835),
.Y(n_865)
);

INVx1_ASAP7_75t_SL g866 ( 
.A(n_839),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_810),
.A2(n_797),
.B1(n_755),
.B2(n_758),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_848),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_827),
.B(n_761),
.Y(n_869)
);

AND2x2_ASAP7_75t_L g870 ( 
.A(n_827),
.B(n_781),
.Y(n_870)
);

INVx3_ASAP7_75t_L g871 ( 
.A(n_831),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_831),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_832),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_832),
.Y(n_874)
);

INVxp67_ASAP7_75t_SL g875 ( 
.A(n_830),
.Y(n_875)
);

NOR2x1_ASAP7_75t_L g876 ( 
.A(n_823),
.B(n_787),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_847),
.B(n_781),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_811),
.B(n_810),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_822),
.Y(n_879)
);

OR2x2_ASAP7_75t_L g880 ( 
.A(n_829),
.B(n_757),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_806),
.B(n_797),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_808),
.B(n_769),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_808),
.B(n_786),
.Y(n_883)
);

HB1xp67_ASAP7_75t_L g884 ( 
.A(n_877),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_857),
.Y(n_885)
);

INVx5_ASAP7_75t_L g886 ( 
.A(n_871),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_L g887 ( 
.A(n_865),
.B(n_786),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_857),
.Y(n_888)
);

OAI33xp33_ASAP7_75t_L g889 ( 
.A1(n_879),
.A2(n_878),
.A3(n_867),
.B1(n_865),
.B2(n_881),
.B3(n_880),
.Y(n_889)
);

OR2x2_ASAP7_75t_L g890 ( 
.A(n_858),
.B(n_757),
.Y(n_890)
);

INVx2_ASAP7_75t_SL g891 ( 
.A(n_880),
.Y(n_891)
);

HB1xp67_ASAP7_75t_L g892 ( 
.A(n_877),
.Y(n_892)
);

AOI22xp33_ASAP7_75t_L g893 ( 
.A1(n_867),
.A2(n_819),
.B1(n_812),
.B2(n_826),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_858),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_855),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_855),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_872),
.B(n_748),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_852),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_859),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_SL g900 ( 
.A(n_876),
.B(n_784),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_869),
.B(n_833),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_852),
.Y(n_902)
);

AND2x2_ASAP7_75t_L g903 ( 
.A(n_869),
.B(n_809),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_891),
.B(n_879),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_885),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_888),
.Y(n_906)
);

BUFx2_ASAP7_75t_L g907 ( 
.A(n_891),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_884),
.B(n_870),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_884),
.B(n_870),
.Y(n_909)
);

OR2x2_ASAP7_75t_L g910 ( 
.A(n_892),
.B(n_898),
.Y(n_910)
);

INVx6_ASAP7_75t_L g911 ( 
.A(n_886),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_903),
.B(n_871),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_899),
.Y(n_913)
);

AND2x2_ASAP7_75t_L g914 ( 
.A(n_892),
.B(n_861),
.Y(n_914)
);

AND2x4_ASAP7_75t_SL g915 ( 
.A(n_901),
.B(n_871),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_887),
.B(n_860),
.Y(n_916)
);

AOI22xp5_ASAP7_75t_L g917 ( 
.A1(n_916),
.A2(n_824),
.B1(n_889),
.B2(n_893),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_SL g918 ( 
.A(n_907),
.B(n_815),
.Y(n_918)
);

NOR2xp67_ASAP7_75t_L g919 ( 
.A(n_913),
.B(n_886),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_915),
.B(n_886),
.Y(n_920)
);

AOI22xp5_ASAP7_75t_L g921 ( 
.A1(n_915),
.A2(n_893),
.B1(n_843),
.B2(n_841),
.Y(n_921)
);

OAI221xp5_ASAP7_75t_L g922 ( 
.A1(n_904),
.A2(n_883),
.B1(n_875),
.B2(n_866),
.C(n_894),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_905),
.B(n_866),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_913),
.Y(n_924)
);

AND2x2_ASAP7_75t_L g925 ( 
.A(n_920),
.B(n_908),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_923),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_917),
.B(n_906),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_919),
.B(n_908),
.Y(n_928)
);

AOI21xp5_ASAP7_75t_L g929 ( 
.A1(n_918),
.A2(n_876),
.B(n_856),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_924),
.B(n_909),
.Y(n_930)
);

OAI22xp33_ASAP7_75t_L g931 ( 
.A1(n_927),
.A2(n_921),
.B1(n_922),
.B2(n_821),
.Y(n_931)
);

OAI22xp33_ASAP7_75t_L g932 ( 
.A1(n_927),
.A2(n_820),
.B1(n_817),
.B2(n_807),
.Y(n_932)
);

NAND3x2_ASAP7_75t_L g933 ( 
.A(n_925),
.B(n_890),
.C(n_910),
.Y(n_933)
);

OAI21xp33_ASAP7_75t_SL g934 ( 
.A1(n_928),
.A2(n_926),
.B(n_930),
.Y(n_934)
);

OAI221xp5_ASAP7_75t_L g935 ( 
.A1(n_934),
.A2(n_929),
.B1(n_931),
.B2(n_911),
.C(n_933),
.Y(n_935)
);

AOI22xp33_ASAP7_75t_L g936 ( 
.A1(n_932),
.A2(n_911),
.B1(n_863),
.B2(n_872),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_934),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_937),
.Y(n_938)
);

AND2x2_ASAP7_75t_L g939 ( 
.A(n_936),
.B(n_912),
.Y(n_939)
);

INVx1_ASAP7_75t_SL g940 ( 
.A(n_935),
.Y(n_940)
);

INVx2_ASAP7_75t_L g941 ( 
.A(n_937),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_938),
.A2(n_911),
.B1(n_836),
.B2(n_874),
.Y(n_942)
);

NAND4xp25_ASAP7_75t_L g943 ( 
.A(n_940),
.B(n_785),
.C(n_837),
.D(n_828),
.Y(n_943)
);

NOR4xp25_ASAP7_75t_L g944 ( 
.A(n_941),
.B(n_789),
.C(n_825),
.D(n_803),
.Y(n_944)
);

NOR2xp67_ASAP7_75t_SL g945 ( 
.A(n_939),
.B(n_770),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_938),
.B(n_886),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_941),
.Y(n_947)
);

AOI22xp5_ASAP7_75t_L g948 ( 
.A1(n_938),
.A2(n_874),
.B1(n_809),
.B2(n_863),
.Y(n_948)
);

OAI211xp5_ASAP7_75t_SL g949 ( 
.A1(n_947),
.A2(n_789),
.B(n_882),
.C(n_895),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_942),
.B(n_909),
.Y(n_950)
);

OAI311xp33_ASAP7_75t_L g951 ( 
.A1(n_943),
.A2(n_862),
.A3(n_914),
.B1(n_854),
.C1(n_896),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_944),
.B(n_914),
.Y(n_952)
);

NOR4xp25_ASAP7_75t_L g953 ( 
.A(n_946),
.B(n_945),
.C(n_948),
.D(n_795),
.Y(n_953)
);

NAND3xp33_ASAP7_75t_L g954 ( 
.A(n_947),
.B(n_774),
.C(n_770),
.Y(n_954)
);

OAI211xp5_ASAP7_75t_L g955 ( 
.A1(n_946),
.A2(n_834),
.B(n_793),
.C(n_774),
.Y(n_955)
);

INVxp33_ASAP7_75t_L g956 ( 
.A(n_950),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_954),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_953),
.B(n_902),
.Y(n_958)
);

NOR2x1_ASAP7_75t_L g959 ( 
.A(n_955),
.B(n_804),
.Y(n_959)
);

NOR2x1_ASAP7_75t_L g960 ( 
.A(n_952),
.B(n_804),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_949),
.Y(n_961)
);

NOR2xp33_ASAP7_75t_L g962 ( 
.A(n_951),
.B(n_899),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_957),
.B(n_774),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_960),
.B(n_774),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_961),
.B(n_774),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_L g966 ( 
.A(n_956),
.B(n_813),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_SL g967 ( 
.A(n_959),
.B(n_813),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_R g968 ( 
.A(n_958),
.B(n_793),
.Y(n_968)
);

XNOR2x1_ASAP7_75t_L g969 ( 
.A(n_962),
.B(n_783),
.Y(n_969)
);

NAND3xp33_ASAP7_75t_L g970 ( 
.A(n_957),
.B(n_803),
.C(n_795),
.Y(n_970)
);

XNOR2xp5_ASAP7_75t_L g971 ( 
.A(n_956),
.B(n_900),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_960),
.B(n_897),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_966),
.Y(n_973)
);

INVx1_ASAP7_75t_SL g974 ( 
.A(n_963),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_971),
.Y(n_975)
);

AOI221xp5_ASAP7_75t_L g976 ( 
.A1(n_965),
.A2(n_900),
.B1(n_897),
.B2(n_819),
.C(n_868),
.Y(n_976)
);

NAND4xp75_ASAP7_75t_L g977 ( 
.A(n_964),
.B(n_868),
.C(n_787),
.D(n_792),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_972),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_967),
.A2(n_783),
.B(n_776),
.Y(n_979)
);

NOR4xp25_ASAP7_75t_SL g980 ( 
.A(n_969),
.B(n_775),
.C(n_792),
.D(n_754),
.Y(n_980)
);

AOI222xp33_ASAP7_75t_L g981 ( 
.A1(n_970),
.A2(n_776),
.B1(n_897),
.B2(n_859),
.C1(n_753),
.C2(n_749),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_968),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_966),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_978),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_974),
.Y(n_985)
);

XNOR2xp5_ASAP7_75t_L g986 ( 
.A(n_973),
.B(n_873),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_983),
.Y(n_987)
);

NAND4xp25_ASAP7_75t_L g988 ( 
.A(n_975),
.B(n_873),
.C(n_862),
.D(n_864),
.Y(n_988)
);

AOI22xp5_ASAP7_75t_L g989 ( 
.A1(n_982),
.A2(n_864),
.B1(n_861),
.B2(n_749),
.Y(n_989)
);

XNOR2x1_ASAP7_75t_L g990 ( 
.A(n_977),
.B(n_753),
.Y(n_990)
);

INVx2_ASAP7_75t_L g991 ( 
.A(n_984),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_987),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_985),
.A2(n_976),
.B(n_980),
.Y(n_993)
);

AOI31xp33_ASAP7_75t_L g994 ( 
.A1(n_992),
.A2(n_986),
.A3(n_990),
.B(n_989),
.Y(n_994)
);

AOI31xp33_ASAP7_75t_L g995 ( 
.A1(n_991),
.A2(n_981),
.A3(n_988),
.B(n_979),
.Y(n_995)
);

XOR2xp5_ASAP7_75t_L g996 ( 
.A(n_994),
.B(n_991),
.Y(n_996)
);

INVxp67_ASAP7_75t_L g997 ( 
.A(n_995),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_R g998 ( 
.A1(n_997),
.A2(n_996),
.B1(n_993),
.B2(n_979),
.Y(n_998)
);

AOI22xp33_ASAP7_75t_SL g999 ( 
.A1(n_997),
.A2(n_749),
.B1(n_752),
.B2(n_756),
.Y(n_999)
);

INVx4_ASAP7_75t_L g1000 ( 
.A(n_998),
.Y(n_1000)
);

XOR2xp5_ASAP7_75t_L g1001 ( 
.A(n_999),
.B(n_853),
.Y(n_1001)
);

OAI221xp5_ASAP7_75t_R g1002 ( 
.A1(n_1001),
.A2(n_775),
.B1(n_750),
.B2(n_853),
.C(n_752),
.Y(n_1002)
);

OAI221xp5_ASAP7_75t_R g1003 ( 
.A1(n_1000),
.A2(n_775),
.B1(n_750),
.B2(n_752),
.C(n_756),
.Y(n_1003)
);

AOI211xp5_ASAP7_75t_L g1004 ( 
.A1(n_1002),
.A2(n_1003),
.B(n_759),
.C(n_784),
.Y(n_1004)
);


endmodule