module fake_jpeg_30722_n_520 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_520);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_520;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_SL g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx8_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_2),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_0),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx16f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx11_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_0),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_5),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_4),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_0),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_52),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g107 ( 
.A(n_54),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_55),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_56),
.Y(n_143)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_58),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx6_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx6_ASAP7_75t_L g148 ( 
.A(n_61),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g118 ( 
.A(n_62),
.Y(n_118)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_63),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

INVx8_ASAP7_75t_L g121 ( 
.A(n_65),
.Y(n_121)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_45),
.Y(n_66)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_66),
.Y(n_114)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_67),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_25),
.B(n_14),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_70),
.B(n_99),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_31),
.Y(n_71)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_71),
.Y(n_145)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_72),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_23),
.Y(n_74)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_75),
.Y(n_158)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_16),
.Y(n_76)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_76),
.Y(n_138)
);

BUFx4f_ASAP7_75t_L g77 ( 
.A(n_36),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_77),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g149 ( 
.A(n_78),
.Y(n_149)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_26),
.Y(n_79)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_79),
.Y(n_133)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_80),
.Y(n_135)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_36),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_97),
.Y(n_113)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx4_ASAP7_75t_SL g127 ( 
.A(n_83),
.Y(n_127)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_84),
.Y(n_141)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_36),
.Y(n_85)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_86),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_44),
.Y(n_87)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_87),
.Y(n_157)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_88),
.Y(n_159)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_21),
.Y(n_89)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_89),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_44),
.Y(n_90)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_90),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_91),
.Y(n_167)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_21),
.Y(n_92)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_92),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g147 ( 
.A(n_93),
.Y(n_147)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx4_ASAP7_75t_SL g156 ( 
.A(n_94),
.Y(n_156)
);

BUFx10_ASAP7_75t_L g95 ( 
.A(n_22),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_95),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g96 ( 
.A(n_22),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_96),
.Y(n_170)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_29),
.B(n_14),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_98),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_25),
.B(n_14),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_101),
.B(n_102),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g102 ( 
.A(n_24),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_33),
.B(n_14),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_27),
.Y(n_162)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_37),
.Y(n_104)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_104),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_105),
.Y(n_161)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_106),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_102),
.A2(n_18),
.B1(n_50),
.B2(n_47),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_110),
.A2(n_126),
.B1(n_131),
.B2(n_144),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_97),
.A2(n_33),
.B1(n_40),
.B2(n_35),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_70),
.B(n_51),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_130),
.B(n_136),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_102),
.A2(n_18),
.B1(n_50),
.B2(n_40),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_88),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_85),
.B(n_51),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_140),
.B(n_150),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_53),
.A2(n_40),
.B1(n_35),
.B2(n_39),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_55),
.A2(n_35),
.B1(n_50),
.B2(n_34),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_146),
.A2(n_62),
.B1(n_105),
.B2(n_91),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_77),
.B(n_34),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_67),
.B(n_27),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_154),
.B(n_37),
.Y(n_197)
);

OAI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_56),
.A2(n_18),
.B1(n_20),
.B2(n_32),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_155),
.A2(n_171),
.B1(n_19),
.B2(n_28),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_162),
.B(n_15),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_64),
.A2(n_20),
.B1(n_37),
.B2(n_39),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_169),
.B1(n_127),
.B2(n_24),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_59),
.A2(n_37),
.B1(n_29),
.B2(n_30),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_61),
.A2(n_15),
.B1(n_32),
.B2(n_30),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_173),
.A2(n_179),
.B1(n_180),
.B2(n_194),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_86),
.B1(n_65),
.B2(n_93),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_174),
.A2(n_128),
.B1(n_148),
.B2(n_120),
.Y(n_237)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_151),
.Y(n_176)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_176),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_112),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_177),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_113),
.B(n_69),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_178),
.B(n_194),
.C(n_170),
.Y(n_233)
);

OAI22xp33_ASAP7_75t_L g180 ( 
.A1(n_161),
.A2(n_75),
.B1(n_87),
.B2(n_71),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_132),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g251 ( 
.A(n_181),
.B(n_190),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_182),
.A2(n_207),
.B1(n_218),
.B2(n_219),
.Y(n_248)
);

INVx4_ASAP7_75t_L g183 ( 
.A(n_159),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g265 ( 
.A(n_183),
.Y(n_265)
);

BUFx2_ASAP7_75t_L g185 ( 
.A(n_132),
.Y(n_185)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_185),
.Y(n_232)
);

INVx11_ASAP7_75t_L g186 ( 
.A(n_116),
.Y(n_186)
);

INVx6_ASAP7_75t_L g226 ( 
.A(n_186),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_187),
.B(n_192),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_122),
.B(n_19),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_188),
.B(n_213),
.Y(n_230)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_189),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_155),
.A2(n_28),
.B1(n_72),
.B2(n_24),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_160),
.Y(n_191)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_191),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_149),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

INVx13_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_108),
.B(n_24),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_111),
.Y(n_195)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_195),
.Y(n_255)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_119),
.Y(n_196)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_196),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_197),
.B(n_199),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_37),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_119),
.Y(n_200)
);

CKINVDCx6p67_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

INVx4_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

INVx6_ASAP7_75t_L g254 ( 
.A(n_201),
.Y(n_254)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_138),
.Y(n_202)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_202),
.Y(n_258)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_135),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_203),
.B(n_205),
.Y(n_245)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_121),
.Y(n_204)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_204),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_117),
.B(n_101),
.Y(n_205)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_112),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g229 ( 
.A(n_206),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_118),
.A2(n_127),
.B1(n_156),
.B2(n_145),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_172),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_208),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_142),
.B(n_152),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_209),
.B(n_210),
.Y(n_247)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_147),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_114),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_211),
.Y(n_252)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_153),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_212),
.B(n_215),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_133),
.B(n_68),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_134),
.B(n_95),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_214),
.B(n_222),
.Y(n_264)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_225),
.Y(n_234)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_164),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_217),
.B(n_221),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_120),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_118),
.A2(n_90),
.B1(n_78),
.B2(n_96),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_156),
.A2(n_95),
.B1(n_13),
.B2(n_12),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_220),
.A2(n_224),
.B1(n_149),
.B2(n_107),
.Y(n_250)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_147),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_115),
.B(n_13),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_141),
.B(n_13),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_11),
.Y(n_257)
);

INVx4_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_167),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_233),
.B(n_240),
.Y(n_271)
);

O2A1O1Ixp33_ASAP7_75t_L g236 ( 
.A1(n_190),
.A2(n_170),
.B(n_169),
.C(n_165),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g266 ( 
.A(n_236),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_L g276 ( 
.A1(n_237),
.A2(n_218),
.B1(n_177),
.B2(n_206),
.Y(n_276)
);

O2A1O1Ixp33_ASAP7_75t_SL g239 ( 
.A1(n_184),
.A2(n_110),
.B(n_131),
.C(n_121),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_239),
.A2(n_243),
.B1(n_253),
.B2(n_262),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_188),
.A2(n_148),
.B1(n_143),
.B2(n_109),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_250),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_158),
.B1(n_145),
.B2(n_109),
.Y(n_253)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_198),
.B(n_168),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_256),
.B(n_175),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_263),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_223),
.A2(n_143),
.B1(n_158),
.B2(n_124),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_178),
.B(n_137),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_SL g323 ( 
.A(n_267),
.B(n_290),
.C(n_201),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_278),
.Y(n_298)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_238),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_238),
.Y(n_270)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_270),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_234),
.Y(n_273)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_273),
.Y(n_325)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_234),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_275),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_276),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_259),
.Y(n_278)
);

CKINVDCx16_ASAP7_75t_R g279 ( 
.A(n_228),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_279),
.B(n_280),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_247),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_251),
.A2(n_179),
.B1(n_180),
.B2(n_189),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_281),
.A2(n_296),
.B1(n_261),
.B2(n_249),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_239),
.A2(n_178),
.B1(n_194),
.B2(n_211),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g302 ( 
.A1(n_282),
.A2(n_246),
.B1(n_200),
.B2(n_181),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_283),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_230),
.B(n_216),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_284),
.B(n_292),
.C(n_227),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_230),
.B(n_208),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_285),
.B(n_288),
.Y(n_304)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_228),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_286),
.B(n_287),
.Y(n_316)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_228),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_257),
.B(n_191),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_264),
.B(n_224),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_289),
.B(n_291),
.Y(n_320)
);

OAI21xp33_ASAP7_75t_L g290 ( 
.A1(n_263),
.A2(n_176),
.B(n_183),
.Y(n_290)
);

INVx1_ASAP7_75t_SL g291 ( 
.A(n_251),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_233),
.B(n_225),
.C(n_196),
.Y(n_292)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_253),
.B(n_217),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_293),
.A2(n_261),
.B(n_202),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_244),
.B(n_215),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_297),
.Y(n_307)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_229),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_295),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_240),
.A2(n_204),
.B1(n_212),
.B2(n_200),
.Y(n_296)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_241),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_291),
.A2(n_251),
.B(n_236),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_299),
.A2(n_306),
.B(n_271),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_272),
.A2(n_239),
.B1(n_248),
.B2(n_262),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_300),
.Y(n_327)
);

OAI32xp33_ASAP7_75t_L g301 ( 
.A1(n_266),
.A2(n_243),
.A3(n_235),
.B1(n_264),
.B2(n_245),
.Y(n_301)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_301),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_302),
.A2(n_319),
.B1(n_324),
.B2(n_265),
.Y(n_346)
);

AOI22x1_ASAP7_75t_L g303 ( 
.A1(n_266),
.A2(n_246),
.B1(n_254),
.B2(n_258),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g332 ( 
.A(n_303),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_281),
.A2(n_256),
.B1(n_246),
.B2(n_255),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_255),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_314),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_273),
.B(n_252),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_284),
.B(n_260),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_315),
.B(n_326),
.C(n_232),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_SL g353 ( 
.A1(n_317),
.A2(n_323),
.B(n_232),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_318),
.A2(n_278),
.B1(n_296),
.B2(n_288),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_274),
.A2(n_252),
.B1(n_249),
.B2(n_241),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_322),
.B(n_231),
.C(n_139),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_274),
.A2(n_282),
.B1(n_271),
.B2(n_293),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_292),
.B(n_231),
.C(n_227),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_308),
.B(n_275),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_328),
.B(n_335),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_330),
.A2(n_334),
.B1(n_337),
.B2(n_345),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_331),
.A2(n_336),
.B(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_333),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_300),
.A2(n_271),
.B1(n_267),
.B2(n_277),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_316),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_299),
.A2(n_293),
.B(n_286),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_306),
.A2(n_277),
.B1(n_294),
.B2(n_269),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_307),
.Y(n_338)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_338),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_312),
.B(n_289),
.Y(n_339)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_339),
.Y(n_378)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_310),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_340),
.B(n_344),
.Y(n_356)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_310),
.Y(n_341)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_322),
.B(n_270),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_343),
.B(n_349),
.C(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_313),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_318),
.A2(n_287),
.B1(n_279),
.B2(n_268),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_346),
.A2(n_321),
.B1(n_325),
.B2(n_314),
.Y(n_357)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_313),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_352),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_312),
.B(n_265),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_348),
.Y(n_370)
);

CKINVDCx16_ASAP7_75t_R g350 ( 
.A(n_316),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_350),
.B(n_303),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_298),
.B(n_265),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_343),
.B(n_315),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_355),
.B(n_360),
.C(n_364),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_361),
.B1(n_363),
.B2(n_330),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_346),
.B1(n_327),
.B2(n_332),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_358),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g360 ( 
.A(n_343),
.B(n_326),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_329),
.A2(n_323),
.B1(n_324),
.B2(n_321),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_332),
.A2(n_321),
.B1(n_325),
.B2(n_304),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_351),
.B(n_320),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_320),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_372),
.Y(n_394)
);

INVx5_ASAP7_75t_L g369 ( 
.A(n_341),
.Y(n_369)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_369),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_331),
.B(n_304),
.Y(n_372)
);

OAI21xp33_ASAP7_75t_L g373 ( 
.A1(n_339),
.A2(n_298),
.B(n_301),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g408 ( 
.A(n_373),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_337),
.B(n_311),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_375),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_332),
.A2(n_319),
.B1(n_302),
.B2(n_303),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_376),
.A2(n_350),
.B1(n_335),
.B2(n_328),
.Y(n_390)
);

FAx1_ASAP7_75t_SL g377 ( 
.A(n_342),
.B(n_303),
.CI(n_317),
.CON(n_377),
.SN(n_377)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_338),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_342),
.B(n_311),
.Y(n_379)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_379),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g380 ( 
.A(n_334),
.B(n_349),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_380),
.B(n_381),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_374),
.A2(n_336),
.B(n_378),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_382),
.A2(n_383),
.B(n_392),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_374),
.A2(n_353),
.B(n_333),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_386),
.A2(n_395),
.B1(n_398),
.B2(n_404),
.Y(n_419)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_387),
.Y(n_410)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_356),
.Y(n_389)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_390),
.A2(n_397),
.B1(n_402),
.B2(n_369),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_367),
.B(n_352),
.Y(n_391)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_361),
.A2(n_345),
.B(n_348),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_356),
.Y(n_393)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_393),
.Y(n_432)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_357),
.A2(n_309),
.B1(n_344),
.B2(n_340),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_376),
.A2(n_347),
.B1(n_305),
.B2(n_297),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g398 ( 
.A1(n_363),
.A2(n_305),
.B1(n_297),
.B2(n_283),
.Y(n_398)
);

INVx1_ASAP7_75t_SL g399 ( 
.A(n_354),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_399),
.B(n_406),
.Y(n_430)
);

XOR2x1_ASAP7_75t_L g400 ( 
.A(n_380),
.B(n_258),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_400),
.B(n_242),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_371),
.A2(n_283),
.B1(n_295),
.B2(n_229),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_359),
.A2(n_362),
.B1(n_372),
.B2(n_370),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_379),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g423 ( 
.A(n_405),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_365),
.Y(n_406)
);

OR2x2_ASAP7_75t_L g407 ( 
.A(n_377),
.B(n_254),
.Y(n_407)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_407),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_365),
.B(n_10),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_409),
.A2(n_354),
.B(n_377),
.Y(n_416)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_360),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_411),
.B(n_414),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_368),
.C(n_366),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_412),
.B(n_413),
.C(n_421),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_368),
.C(n_364),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_403),
.B(n_355),
.Y(n_414)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_415),
.Y(n_437)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_416),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_401),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_420),
.Y(n_441)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_371),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_388),
.A2(n_226),
.B1(n_185),
.B2(n_210),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_424),
.B(n_402),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_425),
.B(n_426),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_408),
.A2(n_193),
.B(n_221),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_382),
.B(n_242),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_427),
.B(n_429),
.C(n_399),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_226),
.C(n_124),
.Y(n_429)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_401),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g436 ( 
.A(n_431),
.B(n_401),
.Y(n_436)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_433),
.Y(n_456)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_436),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_410),
.B(n_396),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_438),
.B(n_440),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g440 ( 
.A(n_428),
.B(n_396),
.Y(n_440)
);

FAx1_ASAP7_75t_SL g442 ( 
.A(n_421),
.B(n_386),
.CI(n_404),
.CON(n_442),
.SN(n_442)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_442),
.B(n_444),
.Y(n_459)
);

FAx1_ASAP7_75t_L g445 ( 
.A(n_422),
.B(n_407),
.CI(n_387),
.CON(n_445),
.SN(n_445)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_445),
.B(n_449),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_390),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_446),
.Y(n_462)
);

AOI21xp5_ASAP7_75t_L g447 ( 
.A1(n_418),
.A2(n_383),
.B(n_407),
.Y(n_447)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_447),
.A2(n_391),
.B(n_424),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_392),
.Y(n_448)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_448),
.A2(n_429),
.B(n_430),
.Y(n_458)
);

XOR2x1_ASAP7_75t_SL g449 ( 
.A(n_422),
.B(n_406),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_412),
.B(n_389),
.C(n_393),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_450),
.B(n_411),
.C(n_425),
.Y(n_454)
);

MAJx2_ASAP7_75t_L g451 ( 
.A(n_423),
.B(n_405),
.C(n_384),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_427),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_437),
.A2(n_415),
.B1(n_384),
.B2(n_432),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_452),
.A2(n_463),
.B1(n_447),
.B2(n_437),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g476 ( 
.A(n_453),
.B(n_457),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_464),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_435),
.B(n_450),
.C(n_434),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_455),
.B(n_460),
.C(n_461),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_434),
.B(n_414),
.Y(n_457)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_458),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_435),
.B(n_419),
.C(n_423),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_444),
.B(n_419),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_L g463 ( 
.A1(n_443),
.A2(n_417),
.B1(n_395),
.B2(n_398),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_442),
.B(n_397),
.C(n_420),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_442),
.C(n_433),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_462),
.B(n_441),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_469),
.B(n_473),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_467),
.B(n_441),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_465),
.B(n_409),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_474),
.B(n_466),
.Y(n_489)
);

OAI21xp33_ASAP7_75t_L g475 ( 
.A1(n_456),
.A2(n_449),
.B(n_439),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_475),
.B(n_242),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_477),
.B(n_483),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_454),
.Y(n_478)
);

OR2x2_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_479),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_439),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g492 ( 
.A(n_480),
.Y(n_492)
);

FAx1_ASAP7_75t_SL g481 ( 
.A(n_466),
.B(n_445),
.CI(n_451),
.CON(n_481),
.SN(n_481)
);

MAJIxp5_ASAP7_75t_L g484 ( 
.A(n_481),
.B(n_482),
.C(n_453),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_460),
.B(n_445),
.C(n_107),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_229),
.B1(n_186),
.B2(n_9),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_484),
.B(n_485),
.Y(n_504)
);

INVxp67_ASAP7_75t_L g485 ( 
.A(n_470),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_472),
.B(n_459),
.C(n_468),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_491),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_489),
.B(n_494),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_472),
.B(n_459),
.C(n_464),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_452),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g497 ( 
.A1(n_493),
.A2(n_495),
.B(n_490),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_471),
.B(n_229),
.C(n_12),
.Y(n_495)
);

NAND3xp33_ASAP7_75t_L g496 ( 
.A(n_481),
.B(n_11),
.C(n_9),
.Y(n_496)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_496),
.A2(n_475),
.B(n_123),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_497),
.B(n_0),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g498 ( 
.A1(n_488),
.A2(n_482),
.B(n_476),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g508 ( 
.A1(n_498),
.A2(n_503),
.B(n_7),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g499 ( 
.A(n_489),
.B(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_502),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_500),
.B(n_7),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_486),
.B(n_9),
.C(n_123),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_SL g503 ( 
.A1(n_493),
.A2(n_116),
.B(n_9),
.Y(n_503)
);

A2O1A1Ixp33_ASAP7_75t_L g506 ( 
.A1(n_505),
.A2(n_492),
.B(n_486),
.C(n_2),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_506),
.B(n_509),
.C(n_1),
.Y(n_511)
);

OAI21xp5_ASAP7_75t_L g512 ( 
.A1(n_508),
.A2(n_510),
.B(n_504),
.Y(n_512)
);

OR2x6_ASAP7_75t_L g514 ( 
.A(n_511),
.B(n_512),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_501),
.C(n_504),
.Y(n_513)
);

AOI21xp33_ASAP7_75t_L g515 ( 
.A1(n_513),
.A2(n_1),
.B(n_3),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_515),
.B(n_3),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_L g517 ( 
.A(n_516),
.B(n_514),
.Y(n_517)
);

AOI21xp5_ASAP7_75t_L g518 ( 
.A1(n_517),
.A2(n_4),
.B(n_5),
.Y(n_518)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_518),
.B(n_4),
.C(n_6),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_519),
.A2(n_4),
.B1(n_6),
.B2(n_485),
.Y(n_520)
);


endmodule