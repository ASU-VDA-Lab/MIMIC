module fake_jpeg_16143_n_360 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_360);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_360;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx4f_ASAP7_75t_SL g20 ( 
.A(n_7),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_37),
.Y(n_71)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_24),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_39),
.A2(n_26),
.B1(n_32),
.B2(n_27),
.Y(n_100)
);

BUFx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_45),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_15),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_44),
.B(n_26),
.Y(n_85)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_21),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_48),
.B(n_52),
.Y(n_86)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_51),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_21),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_14),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_53),
.B(n_62),
.Y(n_88)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_54),
.B(n_57),
.Y(n_96)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_58),
.Y(n_106)
);

INVx3_ASAP7_75t_SL g59 ( 
.A(n_22),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_20),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_16),
.Y(n_108)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_15),
.B(n_1),
.Y(n_61)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_36),
.B(n_26),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_14),
.B(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_66),
.B(n_82),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_15),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_76),
.B(n_113),
.C(n_114),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_34),
.B1(n_23),
.B2(n_19),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_80),
.A2(n_91),
.B1(n_95),
.B2(n_104),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_61),
.B(n_31),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_44),
.B(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_84),
.B(n_33),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_85),
.B(n_98),
.Y(n_133)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_37),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_59),
.A2(n_34),
.B1(n_23),
.B2(n_19),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_42),
.Y(n_92)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_46),
.Y(n_93)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_93),
.Y(n_148)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_94),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_43),
.A2(n_23),
.B1(n_19),
.B2(n_31),
.Y(n_95)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_97),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_50),
.B(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_41),
.Y(n_99)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_99),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_100),
.A2(n_33),
.B1(n_29),
.B2(n_65),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_45),
.B(n_35),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_101),
.B(n_109),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_54),
.A2(n_35),
.B1(n_30),
.B2(n_28),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_102),
.A2(n_112),
.B1(n_3),
.B2(n_4),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_36),
.B1(n_27),
.B2(n_32),
.Y(n_104)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_47),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_51),
.Y(n_107)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_107),
.Y(n_126)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_108),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_48),
.B(n_28),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_52),
.B(n_30),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_110),
.B(n_111),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_57),
.B(n_16),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_58),
.A2(n_36),
.B1(n_27),
.B2(n_29),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_60),
.B(n_56),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_49),
.B(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_115),
.B(n_88),
.Y(n_165)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_118),
.B(n_165),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_119),
.A2(n_144),
.B1(n_146),
.B2(n_154),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_76),
.B(n_64),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_120),
.B(n_124),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_103),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_121),
.A2(n_123),
.B1(n_138),
.B2(n_147),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_122),
.B(n_131),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_103),
.A2(n_33),
.B1(n_29),
.B2(n_25),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_76),
.B(n_25),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_68),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_125),
.Y(n_205)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_89),
.Y(n_128)
);

BUFx5_ASAP7_75t_L g194 ( 
.A(n_128),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_68),
.Y(n_131)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_134),
.Y(n_168)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_136),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_137),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_75),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g139 ( 
.A(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_139),
.B(n_74),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_140),
.B(n_72),
.Y(n_180)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_73),
.Y(n_141)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_114),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_94),
.A2(n_16),
.B1(n_4),
.B2(n_5),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_84),
.B(n_3),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_145),
.B(n_159),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_67),
.A2(n_16),
.B1(n_5),
.B2(n_6),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_3),
.B1(n_7),
.B2(n_8),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_81),
.Y(n_149)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_149),
.Y(n_203)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_96),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_114),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_154)
);

OAI22xp33_ASAP7_75t_L g156 ( 
.A1(n_67),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_156),
.A2(n_105),
.B1(n_106),
.B2(n_128),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_105),
.Y(n_157)
);

BUFx2_ASAP7_75t_SL g185 ( 
.A(n_157),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_97),
.B(n_8),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_158),
.B(n_83),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_100),
.B(n_10),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_113),
.B(n_10),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_162),
.B(n_163),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_70),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_83),
.A2(n_74),
.B1(n_77),
.B2(n_78),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_150),
.B(n_72),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_169),
.B(n_177),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_164),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_171),
.B(n_173),
.Y(n_215)
);

MAJx2_ASAP7_75t_L g211 ( 
.A(n_172),
.B(n_190),
.C(n_184),
.Y(n_211)
);

OAI32xp33_ASAP7_75t_L g174 ( 
.A1(n_120),
.A2(n_72),
.A3(n_92),
.B1(n_93),
.B2(n_90),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_174),
.A2(n_180),
.B1(n_204),
.B2(n_132),
.Y(n_226)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_157),
.Y(n_176)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_176),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_133),
.B(n_72),
.Y(n_177)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_127),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_179),
.B(n_197),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_118),
.B(n_145),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_183),
.B(n_187),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_SL g184 ( 
.A(n_160),
.B(n_124),
.C(n_162),
.Y(n_184)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_184),
.B(n_188),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_130),
.B(n_99),
.Y(n_187)
);

FAx1_ASAP7_75t_SL g188 ( 
.A(n_129),
.B(n_107),
.CI(n_78),
.CON(n_188),
.SN(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_153),
.B(n_77),
.Y(n_189)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_189),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_158),
.B(n_79),
.Y(n_190)
);

NOR3xp33_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_192),
.C(n_144),
.Y(n_241)
);

OAI21xp33_ASAP7_75t_L g192 ( 
.A1(n_143),
.A2(n_79),
.B(n_87),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_163),
.B(n_87),
.Y(n_193)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_193),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_196),
.A2(n_116),
.B1(n_126),
.B2(n_136),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_151),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_154),
.B(n_106),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_135),
.B(n_117),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_200),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_129),
.B(n_159),
.Y(n_204)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_134),
.Y(n_207)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_207),
.Y(n_220)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

BUFx2_ASAP7_75t_L g245 ( 
.A(n_208),
.Y(n_245)
);

OR2x2_ASAP7_75t_L g210 ( 
.A(n_171),
.B(n_202),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g250 ( 
.A1(n_210),
.A2(n_202),
.B(n_204),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_211),
.B(n_226),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_140),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_212),
.B(n_218),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_170),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_213),
.B(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_148),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_195),
.B(n_141),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_223),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_191),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_175),
.B(n_204),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_168),
.Y(n_225)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_225),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_168),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_227),
.B(n_232),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_156),
.Y(n_228)
);

NOR3xp33_ASAP7_75t_L g249 ( 
.A(n_228),
.B(n_178),
.C(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_186),
.Y(n_230)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_230),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_152),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_186),
.Y(n_233)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_233),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_234),
.A2(n_178),
.B1(n_189),
.B2(n_166),
.Y(n_261)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_206),
.Y(n_235)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_235),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_175),
.B(n_155),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_236),
.B(n_182),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_135),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_237),
.B(n_239),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_206),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_180),
.A2(n_161),
.B1(n_126),
.B2(n_146),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_205),
.B1(n_201),
.B2(n_203),
.Y(n_273)
);

NOR2xp67_ASAP7_75t_R g252 ( 
.A(n_241),
.B(n_174),
.Y(n_252)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_207),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g262 ( 
.A(n_242),
.Y(n_262)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_244),
.Y(n_269)
);

INVx2_ASAP7_75t_SL g246 ( 
.A(n_185),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_246),
.B(n_194),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_226),
.A2(n_198),
.B1(n_181),
.B2(n_180),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_247),
.A2(n_248),
.B1(n_261),
.B2(n_265),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_246),
.A2(n_243),
.B1(n_214),
.B2(n_209),
.Y(n_248)
);

AO21x1_ASAP7_75t_L g293 ( 
.A1(n_249),
.A2(n_250),
.B(n_252),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_172),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_253),
.B(n_231),
.C(n_211),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_257),
.B(n_218),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_216),
.A2(n_198),
.B(n_167),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g280 ( 
.A(n_258),
.B(n_266),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_212),
.A2(n_215),
.B1(n_217),
.B2(n_236),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_216),
.A2(n_167),
.B(n_188),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_217),
.A2(n_188),
.B1(n_177),
.B2(n_205),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_273),
.B1(n_214),
.B2(n_234),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_213),
.B(n_176),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_268),
.B(n_270),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_238),
.B(n_194),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g274 ( 
.A1(n_210),
.A2(n_201),
.B(n_203),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_258),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_246),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_277),
.B(n_245),
.Y(n_279)
);

NOR2x1_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_210),
.Y(n_278)
);

CKINVDCx14_ASAP7_75t_R g313 ( 
.A(n_278),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_284),
.B1(n_292),
.B2(n_294),
.Y(n_306)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_251),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_283),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_254),
.B(n_221),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_285),
.B(n_287),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_254),
.B(n_231),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_288),
.B(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_257),
.B(n_239),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_289),
.B(n_295),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_255),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_290),
.A2(n_262),
.B1(n_245),
.B2(n_149),
.Y(n_312)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_251),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_263),
.B(n_227),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_261),
.A2(n_240),
.B1(n_229),
.B2(n_222),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_297),
.A2(n_298),
.B1(n_302),
.B2(n_269),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_247),
.A2(n_244),
.B1(n_230),
.B2(n_242),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_219),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_300),
.Y(n_316)
);

A2O1A1Ixp33_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_225),
.B(n_235),
.C(n_233),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_266),
.C(n_250),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_263),
.A2(n_220),
.B1(n_243),
.B2(n_224),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_291),
.A2(n_273),
.B1(n_269),
.B2(n_275),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g326 ( 
.A1(n_303),
.A2(n_309),
.B1(n_310),
.B2(n_311),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_282),
.A2(n_267),
.B1(n_265),
.B2(n_274),
.Y(n_304)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g307 ( 
.A1(n_278),
.A2(n_270),
.A3(n_276),
.B1(n_275),
.B2(n_255),
.C1(n_260),
.C2(n_272),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_307),
.B(n_320),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_308),
.A2(n_287),
.B1(n_289),
.B2(n_285),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_297),
.A2(n_276),
.B1(n_259),
.B2(n_272),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_290),
.A2(n_256),
.B1(n_260),
.B2(n_259),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_298),
.A2(n_277),
.B1(n_262),
.B2(n_220),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_312),
.A2(n_302),
.B(n_280),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_295),
.A2(n_245),
.B1(n_125),
.B2(n_137),
.Y(n_319)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

AOI32xp33_ASAP7_75t_L g320 ( 
.A1(n_293),
.A2(n_300),
.A3(n_280),
.B1(n_286),
.B2(n_296),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_L g338 ( 
.A1(n_322),
.A2(n_327),
.B1(n_333),
.B2(n_303),
.Y(n_338)
);

NOR3xp33_ASAP7_75t_L g323 ( 
.A(n_306),
.B(n_293),
.C(n_284),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_323),
.B(n_328),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_305),
.B(n_281),
.Y(n_325)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_325),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_318),
.A2(n_292),
.B1(n_283),
.B2(n_294),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_321),
.B(n_281),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_329),
.A2(n_335),
.B(n_324),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_314),
.B(n_288),
.C(n_301),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_314),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_321),
.A2(n_317),
.B1(n_318),
.B2(n_313),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_332),
.A2(n_304),
.B1(n_319),
.B2(n_315),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_317),
.A2(n_299),
.B1(n_312),
.B2(n_311),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_315),
.B(n_310),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_SL g349 ( 
.A(n_336),
.B(n_330),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_316),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_337),
.B(n_339),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_338),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_316),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_340),
.B(n_342),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_324),
.A2(n_335),
.B(n_334),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_343),
.A2(n_322),
.B1(n_327),
.B2(n_344),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_334),
.B(n_326),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_344),
.B(n_340),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_348),
.A2(n_351),
.B1(n_342),
.B2(n_341),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_349),
.B(n_337),
.C(n_345),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_352),
.B(n_353),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_347),
.B(n_339),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_354),
.A2(n_347),
.B(n_348),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_356),
.A2(n_350),
.B1(n_346),
.B2(n_353),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_358),
.Y(n_359)
);

AO21x2_ASAP7_75t_L g360 ( 
.A1(n_359),
.A2(n_355),
.B(n_336),
.Y(n_360)
);


endmodule