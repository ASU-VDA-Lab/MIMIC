module fake_jpeg_15709_n_169 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_169);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_169;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

INVx2_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_21),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_22),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_26),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_4),
.Y(n_58)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_16),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_13),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_36),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx5_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_69),
.Y(n_81)
);

BUFx24_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_0),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_71),
.B(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_52),
.Y(n_72)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g74 ( 
.A(n_51),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_55),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_47),
.B(n_0),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_69),
.A2(n_46),
.B1(n_59),
.B2(n_57),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_77),
.A2(n_90),
.B(n_94),
.C(n_87),
.Y(n_110)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_68),
.B(n_67),
.Y(n_80)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_80),
.B(n_92),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_72),
.A2(n_46),
.B1(n_59),
.B2(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_83),
.A2(n_85),
.B1(n_90),
.B2(n_94),
.Y(n_106)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_84),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_70),
.A2(n_60),
.B1(n_65),
.B2(n_53),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_68),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_70),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_64),
.Y(n_95)
);

BUFx12f_ASAP7_75t_SL g92 ( 
.A(n_70),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_93),
.B(n_64),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_68),
.A2(n_49),
.B1(n_50),
.B2(n_53),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_95),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g96 ( 
.A(n_89),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_96),
.B(n_99),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_81),
.Y(n_99)
);

BUFx12_ASAP7_75t_L g101 ( 
.A(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_101),
.B(n_102),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_48),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_105),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_54),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_86),
.B(n_56),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_114),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_110),
.A2(n_113),
.B(n_115),
.Y(n_119)
);

BUFx8_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_92),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_1),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_78),
.B(n_1),
.Y(n_114)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_2),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_116),
.B(n_66),
.C(n_63),
.Y(n_127)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_79),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_117),
.A2(n_118),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_78),
.B(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_127),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_115),
.B(n_62),
.C(n_27),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_112),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_119),
.A2(n_106),
.B1(n_111),
.B2(n_100),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_132),
.B(n_135),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_133),
.B(n_136),
.Y(n_141)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_137),
.A2(n_97),
.B(n_104),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_121),
.C(n_134),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_138),
.B(n_140),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_137),
.A2(n_125),
.B(n_122),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_144),
.A2(n_145),
.B(n_124),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g145 ( 
.A1(n_142),
.A2(n_123),
.B(n_136),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_141),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_123),
.B(n_116),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_148),
.B(n_149),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_143),
.B(n_127),
.C(n_129),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_146),
.Y(n_150)
);

NOR2x1_ASAP7_75t_L g152 ( 
.A(n_150),
.B(n_151),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_113),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_154),
.A2(n_155),
.B1(n_152),
.B2(n_108),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_128),
.B(n_130),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_156),
.A2(n_3),
.B1(n_6),
.B2(n_7),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_7),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_158),
.B(n_8),
.Y(n_159)
);

AOI221xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_98),
.B1(n_31),
.B2(n_44),
.C(n_43),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_28),
.Y(n_161)
);

OAI21xp5_ASAP7_75t_SL g162 ( 
.A1(n_161),
.A2(n_29),
.B(n_35),
.Y(n_162)
);

AOI21x1_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_25),
.B(n_42),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_24),
.C(n_38),
.Y(n_164)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_164),
.Y(n_165)
);

AO22x1_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_23),
.B1(n_37),
.B2(n_34),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_95),
.B(n_12),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_167),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_10),
.C(n_33),
.Y(n_169)
);


endmodule