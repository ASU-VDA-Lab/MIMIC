module fake_jpeg_29371_n_438 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx16f_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_9),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_6),
.B(n_14),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_4),
.Y(n_42)
);

BUFx16f_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_45),
.B(n_58),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_46),
.B(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_0),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_48),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_51),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_26),
.Y(n_52)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_52),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_53),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_55),
.Y(n_111)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_16),
.B(n_0),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_57),
.B(n_59),
.Y(n_116)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_16),
.B(n_1),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_23),
.B(n_2),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_60),
.B(n_71),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g118 ( 
.A(n_61),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_62),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_63),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g65 ( 
.A(n_22),
.Y(n_65)
);

INVx6_ASAP7_75t_SL g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_69),
.Y(n_142)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_70),
.B(n_81),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_2),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_72),
.Y(n_100)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_73),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_80),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_75),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_35),
.B(n_2),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_76),
.B(n_79),
.Y(n_137)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_20),
.Y(n_77)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_21),
.Y(n_78)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_32),
.B(n_17),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_29),
.Y(n_80)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_83),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_29),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_32),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

BUFx16f_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_35),
.B(n_3),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_36),
.Y(n_107)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_41),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_89),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_44),
.B(n_3),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_91),
.Y(n_124)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

INVx11_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_92),
.B(n_28),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_48),
.A2(n_34),
.B1(n_18),
.B2(n_25),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_106),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_107),
.B(n_143),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_79),
.B(n_31),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_113),
.B(n_130),
.Y(n_163)
);

OAI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_67),
.A2(n_29),
.B1(n_17),
.B2(n_18),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_115),
.A2(n_132),
.B1(n_138),
.B2(n_72),
.Y(n_154)
);

AOI21xp33_ASAP7_75t_L g120 ( 
.A1(n_62),
.A2(n_17),
.B(n_44),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_68),
.C(n_82),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_49),
.A2(n_34),
.B1(n_18),
.B2(n_17),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_50),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g123 ( 
.A1(n_51),
.A2(n_40),
.B1(n_27),
.B2(n_37),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_126),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_58),
.B(n_37),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_128),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_58),
.B(n_36),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_62),
.B(n_33),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_129),
.B(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_52),
.B(n_31),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_92),
.A2(n_33),
.B1(n_30),
.B2(n_27),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_53),
.B(n_31),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_144),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_61),
.A2(n_30),
.B1(n_31),
.B2(n_6),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_134),
.A2(n_109),
.B1(n_93),
.B2(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_63),
.A2(n_31),
.B1(n_5),
.B2(n_7),
.Y(n_138)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g157 ( 
.A1(n_139),
.A2(n_75),
.B1(n_80),
.B2(n_83),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_86),
.B(n_73),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_64),
.B(n_4),
.Y(n_144)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_99),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_148),
.B(n_152),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_125),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_149),
.B(n_150),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_113),
.B(n_77),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_151),
.B(n_159),
.C(n_174),
.Y(n_201)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_98),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_153),
.B(n_156),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_154),
.A2(n_178),
.B1(n_103),
.B2(n_97),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_155),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_101),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_157),
.A2(n_188),
.B1(n_195),
.B2(n_147),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_138),
.A2(n_74),
.B1(n_69),
.B2(n_81),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_158),
.A2(n_176),
.B1(n_189),
.B2(n_93),
.Y(n_229)
);

AND2x2_ASAP7_75t_SL g159 ( 
.A(n_120),
.B(n_4),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_125),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g228 ( 
.A(n_160),
.B(n_175),
.Y(n_228)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_136),
.Y(n_161)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_161),
.Y(n_214)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_94),
.Y(n_162)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_162),
.Y(n_208)
);

INVxp33_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_164),
.B(n_168),
.Y(n_224)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_165),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_144),
.B(n_86),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_167),
.B(n_170),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_5),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_137),
.A2(n_114),
.A3(n_116),
.B1(n_117),
.B2(n_112),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_177),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_101),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_180),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_5),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_116),
.B(n_7),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_176)
);

OA22x2_ASAP7_75t_L g178 ( 
.A1(n_139),
.A2(n_11),
.B1(n_8),
.B2(n_10),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_133),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_179),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_117),
.B(n_8),
.Y(n_180)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_109),
.Y(n_181)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_181),
.Y(n_212)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_109),
.Y(n_182)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_96),
.Y(n_183)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_101),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_184),
.B(n_185),
.Y(n_230)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_186),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_112),
.B(n_8),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_187),
.Y(n_213)
);

OAI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_139),
.A2(n_11),
.B1(n_104),
.B2(n_136),
.Y(n_188)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_94),
.Y(n_191)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_191),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_142),
.B(n_145),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_192),
.B(n_197),
.Y(n_217)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_135),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_194),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_104),
.A2(n_140),
.B1(n_105),
.B2(n_96),
.Y(n_195)
);

INVx6_ASAP7_75t_L g196 ( 
.A(n_102),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_196),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_118),
.Y(n_197)
);

O2A1O1Ixp33_ASAP7_75t_L g198 ( 
.A1(n_130),
.A2(n_110),
.B(n_103),
.C(n_100),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_119),
.B(n_100),
.C(n_141),
.Y(n_218)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_198),
.B(n_110),
.Y(n_200)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_222),
.Y(n_247)
);

OAI22xp33_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_105),
.B1(n_147),
.B2(n_118),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_204),
.A2(n_216),
.B1(n_221),
.B2(n_229),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_156),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_206),
.B(n_215),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_163),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_227),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_181),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_218),
.A2(n_237),
.B(n_160),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_154),
.A2(n_119),
.B1(n_108),
.B2(n_145),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_166),
.B(n_103),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_179),
.B(n_142),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_232),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_179),
.B(n_108),
.Y(n_232)
);

AND2x2_ASAP7_75t_SL g235 ( 
.A(n_163),
.B(n_131),
.Y(n_235)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_235),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_159),
.A2(n_102),
.B1(n_141),
.B2(n_131),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_236),
.A2(n_158),
.B1(n_171),
.B2(n_157),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_151),
.A2(n_111),
.B(n_146),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_102),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_157),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_201),
.B(n_174),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_240),
.B(n_201),
.C(n_211),
.Y(n_276)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

INVx13_ASAP7_75t_L g286 ( 
.A(n_242),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_243),
.A2(n_267),
.B1(n_274),
.B2(n_210),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_220),
.B(n_159),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_248),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_202),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_246),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_169),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_220),
.B(n_170),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_249),
.B(n_252),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_210),
.B(n_150),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_250),
.B(n_268),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_175),
.Y(n_251)
);

NAND3xp33_ASAP7_75t_L g290 ( 
.A(n_251),
.B(n_233),
.C(n_213),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_209),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_224),
.B(n_190),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_253),
.B(n_271),
.Y(n_277)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_226),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

HB1xp67_ASAP7_75t_L g255 ( 
.A(n_212),
.Y(n_255)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_255),
.Y(n_289)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_226),
.Y(n_256)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_256),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_231),
.A2(n_150),
.B(n_193),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_257),
.A2(n_228),
.B(n_235),
.Y(n_300)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_214),
.Y(n_258)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_239),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

INVx8_ASAP7_75t_L g261 ( 
.A(n_202),
.Y(n_261)
);

INVx13_ASAP7_75t_L g291 ( 
.A(n_261),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_262),
.B(n_216),
.Y(n_280)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_239),
.Y(n_264)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_264),
.Y(n_307)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_265),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_209),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_266),
.B(n_269),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_199),
.A2(n_176),
.B1(n_178),
.B2(n_183),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_230),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_223),
.Y(n_270)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_270),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_225),
.B(n_149),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_225),
.B(n_193),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_272),
.B(n_273),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_224),
.B(n_161),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_222),
.A2(n_178),
.B1(n_109),
.B2(n_155),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_250),
.C(n_256),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_280),
.B(n_240),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_247),
.A2(n_229),
.B1(n_210),
.B2(n_221),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_282),
.A2(n_287),
.B(n_288),
.Y(n_308)
);

BUFx4f_ASAP7_75t_SL g284 ( 
.A(n_246),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_284),
.Y(n_311)
);

A2O1A1Ixp33_ASAP7_75t_SL g287 ( 
.A1(n_268),
.A2(n_237),
.B(n_200),
.C(n_218),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_247),
.A2(n_218),
.B(n_232),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_306),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_262),
.A2(n_235),
.B1(n_238),
.B2(n_227),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_292),
.A2(n_244),
.B1(n_249),
.B2(n_245),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_294),
.A2(n_296),
.B1(n_263),
.B2(n_275),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_274),
.A2(n_235),
.B1(n_236),
.B2(n_213),
.Y(n_296)
);

OAI21xp33_ASAP7_75t_SL g319 ( 
.A1(n_300),
.A2(n_305),
.B(n_259),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_247),
.A2(n_228),
.B(n_230),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_302),
.B(n_266),
.Y(n_315)
);

CKINVDCx12_ASAP7_75t_R g304 ( 
.A(n_241),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_304),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_257),
.A2(n_228),
.B(n_203),
.Y(n_305)
);

INVx13_ASAP7_75t_L g306 ( 
.A(n_261),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_277),
.B(n_252),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_310),
.Y(n_347)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_313),
.B(n_317),
.Y(n_357)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_314),
.B(n_315),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_320),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_244),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_283),
.A2(n_243),
.B1(n_269),
.B2(n_267),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_318),
.B(n_329),
.Y(n_341)
);

AOI21xp5_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_178),
.B(n_205),
.Y(n_354)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_298),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_278),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_321),
.B(n_325),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_283),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_322),
.B(n_331),
.C(n_332),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_297),
.B(n_259),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_324),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_279),
.B(n_253),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_303),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_326),
.B(n_327),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g327 ( 
.A(n_281),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_294),
.A2(n_263),
.B1(n_296),
.B2(n_282),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g355 ( 
.A(n_328),
.B(n_330),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_283),
.A2(n_250),
.B1(n_275),
.B2(n_254),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_278),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_300),
.B(n_264),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_303),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_335),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_280),
.B(n_260),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_334),
.B(n_302),
.Y(n_336)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_336),
.B(n_350),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_322),
.B(n_305),
.C(n_292),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_338),
.B(n_346),
.C(n_351),
.Y(n_363)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_309),
.B(n_287),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_SL g376 ( 
.A1(n_339),
.A2(n_354),
.B(n_356),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g342 ( 
.A1(n_318),
.A2(n_288),
.B1(n_287),
.B2(n_285),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_342),
.A2(n_343),
.B1(n_348),
.B2(n_332),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_329),
.A2(n_287),
.B1(n_295),
.B2(n_307),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_287),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_313),
.A2(n_307),
.B1(n_289),
.B2(n_277),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_334),
.B(n_279),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_289),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_325),
.B(n_207),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_323),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g356 ( 
.A1(n_308),
.A2(n_281),
.B(n_301),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_357),
.A2(n_317),
.B1(n_324),
.B2(n_308),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_360),
.A2(n_379),
.B1(n_344),
.B2(n_341),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_361),
.A2(n_370),
.B1(n_371),
.B2(n_374),
.Y(n_393)
);

AOI21xp33_ASAP7_75t_L g362 ( 
.A1(n_347),
.A2(n_323),
.B(n_312),
.Y(n_362)
);

AOI21xp5_ASAP7_75t_L g384 ( 
.A1(n_362),
.A2(n_369),
.B(n_354),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_364),
.B(n_365),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_207),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_349),
.B(n_320),
.Y(n_366)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_366),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_335),
.C(n_330),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_372),
.C(n_377),
.Y(n_381)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_359),
.Y(n_368)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_368),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_358),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_355),
.A2(n_311),
.B1(n_321),
.B2(n_326),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_348),
.A2(n_311),
.B1(n_333),
.B2(n_303),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_337),
.B(n_219),
.C(n_212),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_341),
.A2(n_356),
.B1(n_342),
.B2(n_343),
.Y(n_374)
);

INVx2_ASAP7_75t_L g375 ( 
.A(n_359),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_375),
.B(n_378),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_219),
.C(n_234),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_352),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_357),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_363),
.B(n_340),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_380),
.B(n_394),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_363),
.B(n_373),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g404 ( 
.A(n_382),
.B(n_383),
.Y(n_404)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_384),
.A2(n_299),
.B(n_284),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_360),
.A2(n_341),
.B1(n_339),
.B2(n_346),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_386),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_373),
.B(n_338),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_391),
.C(n_392),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g391 ( 
.A(n_361),
.B(n_340),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_367),
.B(n_350),
.C(n_336),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_SL g394 ( 
.A(n_366),
.B(n_301),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_234),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_395),
.B(n_370),
.C(n_371),
.Y(n_398)
);

A2O1A1O1Ixp25_ASAP7_75t_L g396 ( 
.A1(n_386),
.A2(n_376),
.B(n_374),
.C(n_369),
.D(n_372),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_396),
.B(n_398),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_382),
.B(n_376),
.C(n_375),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_399),
.B(n_400),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_387),
.A2(n_242),
.B1(n_299),
.B2(n_246),
.Y(n_400)
);

NOR3xp33_ASAP7_75t_L g402 ( 
.A(n_385),
.B(n_284),
.C(n_291),
.Y(n_402)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_402),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_388),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_403),
.B(n_406),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g411 ( 
.A1(n_405),
.A2(n_389),
.B(n_393),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_381),
.B(n_208),
.C(n_270),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_407),
.B(n_390),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_404),
.C(n_401),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g423 ( 
.A(n_411),
.B(n_417),
.Y(n_423)
);

AOI21x1_ASAP7_75t_L g412 ( 
.A1(n_396),
.A2(n_391),
.B(n_380),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_SL g420 ( 
.A1(n_412),
.A2(n_401),
.B(n_291),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_403),
.B(n_306),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_413),
.A2(n_414),
.B(n_404),
.Y(n_418)
);

AO21x1_ASAP7_75t_L g414 ( 
.A1(n_397),
.A2(n_395),
.B(n_392),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_407),
.B(n_381),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_418),
.B(n_425),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g430 ( 
.A(n_419),
.B(n_162),
.C(n_165),
.Y(n_430)
);

AOI21x1_ASAP7_75t_L g427 ( 
.A1(n_420),
.A2(n_414),
.B(n_146),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g421 ( 
.A1(n_417),
.A2(n_286),
.B(n_265),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_421),
.A2(n_413),
.B(n_415),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_208),
.C(n_223),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_422),
.B(n_424),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_416),
.B(n_286),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_410),
.B(n_258),
.Y(n_425)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_426),
.A2(n_430),
.B(n_423),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_427),
.Y(n_433)
);

BUFx24_ASAP7_75t_SL g431 ( 
.A(n_428),
.Y(n_431)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_432),
.A2(n_429),
.B(n_182),
.Y(n_434)
);

AOI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_434),
.A2(n_433),
.B(n_111),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_435),
.C(n_191),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g438 ( 
.A(n_437),
.B(n_196),
.Y(n_438)
);


endmodule