module fake_jpeg_333_n_396 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_11),
.B(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_3),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_47),
.Y(n_106)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_48),
.Y(n_113)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_49),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_29),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g129 ( 
.A1(n_50),
.A2(n_20),
.B1(n_39),
.B2(n_25),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_54),
.Y(n_95)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_55),
.Y(n_130)
);

AND2x2_ASAP7_75t_SL g56 ( 
.A(n_44),
.B(n_8),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_56),
.B(n_66),
.Y(n_122)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_57),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_58),
.Y(n_131)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_24),
.Y(n_60)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_61),
.Y(n_110)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_62),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_33),
.Y(n_63)
);

BUFx4f_ASAP7_75t_SL g97 ( 
.A(n_63),
.Y(n_97)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_64),
.Y(n_111)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_65),
.Y(n_133)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_67),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_33),
.Y(n_68)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_68),
.Y(n_136)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_70),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_42),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_71),
.Y(n_92)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_41),
.Y(n_72)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_72),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_45),
.Y(n_74)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_74),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_27),
.B(n_2),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_77),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

BUFx3_ASAP7_75t_L g77 ( 
.A(n_21),
.Y(n_77)
);

INVxp67_ASAP7_75t_SL g78 ( 
.A(n_30),
.Y(n_78)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_79),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_35),
.Y(n_80)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_82),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_35),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_83),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_84),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_86),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_18),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_87),
.B(n_88),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_18),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_45),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_89),
.B(n_19),
.C(n_20),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_21),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_90),
.A2(n_91),
.B1(n_45),
.B2(n_23),
.Y(n_94)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_32),
.C(n_43),
.Y(n_93)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_93),
.B(n_32),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_94),
.Y(n_152)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_90),
.A2(n_39),
.B1(n_25),
.B2(n_23),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_107),
.A2(n_127),
.B1(n_128),
.B2(n_66),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_27),
.B1(n_50),
.B2(n_53),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_78),
.A2(n_71),
.B1(n_28),
.B2(n_38),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_31),
.B1(n_26),
.B2(n_34),
.Y(n_147)
);

AND2x2_ASAP7_75t_SL g138 ( 
.A(n_135),
.B(n_19),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_137),
.A2(n_150),
.B1(n_158),
.B2(n_160),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_138),
.B(n_107),
.Y(n_182)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_95),
.Y(n_139)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_139),
.Y(n_184)
);

INVx13_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_140),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_141),
.B(n_145),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_142),
.Y(n_200)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

INVx3_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_144),
.B(n_157),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_36),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_132),
.A2(n_31),
.B1(n_40),
.B2(n_34),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_146),
.A2(n_147),
.B1(n_169),
.B2(n_128),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_122),
.B(n_43),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_148),
.B(n_156),
.Y(n_185)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_149),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_122),
.A2(n_28),
.B1(n_38),
.B2(n_36),
.Y(n_150)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_95),
.Y(n_151)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_151),
.Y(n_208)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_103),
.Y(n_153)
);

INVx3_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_102),
.Y(n_154)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_154),
.Y(n_202)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_108),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_22),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_99),
.A2(n_22),
.B1(n_40),
.B2(n_26),
.Y(n_158)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_105),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_161),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_113),
.A2(n_88),
.B1(n_87),
.B2(n_86),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_101),
.B(n_13),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_104),
.A2(n_85),
.B1(n_84),
.B2(n_80),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_162),
.A2(n_164),
.B1(n_173),
.B2(n_174),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_68),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_177),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_129),
.B(n_61),
.Y(n_164)
);

BUFx3_ASAP7_75t_L g165 ( 
.A(n_106),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_166),
.Y(n_201)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_109),
.B(n_10),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_167),
.B(n_168),
.Y(n_205)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_118),
.A2(n_51),
.B1(n_37),
.B2(n_4),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_123),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_110),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_126),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_172),
.Y(n_207)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_117),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_131),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_178),
.B2(n_120),
.Y(n_199)
);

INVx4_ASAP7_75t_L g176 ( 
.A(n_124),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_111),
.B(n_2),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_98),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_116),
.B(n_3),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_179),
.B(n_3),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_204),
.Y(n_216)
);

MAJx2_ASAP7_75t_L g209 ( 
.A(n_182),
.B(n_138),
.C(n_163),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_190),
.B(n_139),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_119),
.B1(n_129),
.B2(n_136),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_191),
.A2(n_206),
.B1(n_152),
.B2(n_97),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_156),
.B(n_134),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_195),
.B(n_179),
.Y(n_211)
);

CKINVDCx14_ASAP7_75t_R g227 ( 
.A(n_199),
.Y(n_227)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_152),
.A2(n_94),
.B1(n_136),
.B2(n_114),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_164),
.A2(n_125),
.B1(n_121),
.B2(n_97),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_185),
.C(n_195),
.Y(n_240)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_202),
.Y(n_210)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_210),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_211),
.B(n_221),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_196),
.B(n_177),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_214),
.Y(n_232)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_191),
.A2(n_164),
.B1(n_173),
.B2(n_168),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_217),
.A2(n_223),
.B1(n_197),
.B2(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_189),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_224),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_186),
.A2(n_148),
.B(n_138),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

AO22x1_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_151),
.B1(n_159),
.B2(n_143),
.Y(n_220)
);

NAND2x1_ASAP7_75t_L g237 ( 
.A(n_220),
.B(n_208),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_183),
.B(n_141),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_183),
.A2(n_125),
.B1(n_121),
.B2(n_133),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_229),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_182),
.A2(n_166),
.B1(n_155),
.B2(n_176),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_201),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_188),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_188),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_226),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_188),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_228),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_180),
.B(n_172),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_157),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_230),
.B(n_205),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_235),
.A2(n_241),
.B1(n_247),
.B2(n_216),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_229),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_237),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_221),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_204),
.B1(n_181),
.B2(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_243),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_185),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_223),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_245),
.B(n_215),
.Y(n_266)
);

OAI22xp33_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_204),
.B1(n_181),
.B2(n_194),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

CKINVDCx14_ASAP7_75t_R g257 ( 
.A(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_180),
.C(n_192),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_251),
.B(n_209),
.C(n_218),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_254),
.A2(n_231),
.B1(n_236),
.B2(n_246),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_255),
.B(n_258),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_256),
.B(n_271),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_261),
.B(n_265),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_217),
.B1(n_224),
.B2(n_216),
.Y(n_262)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_262),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_252),
.A2(n_216),
.B1(n_223),
.B2(n_212),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_267),
.B1(n_270),
.B2(n_241),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_237),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_264),
.B(n_269),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_243),
.B(n_219),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_266),
.B(n_235),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_252),
.A2(n_227),
.B1(n_214),
.B2(n_181),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_241),
.A2(n_227),
.B1(n_222),
.B2(n_204),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_268),
.A2(n_273),
.B(n_231),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_250),
.B(n_210),
.Y(n_269)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_269),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_245),
.A2(n_213),
.B1(n_226),
.B2(n_225),
.Y(n_270)
);

XNOR2x2_ASAP7_75t_L g271 ( 
.A(n_242),
.B(n_192),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_248),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g280 ( 
.A(n_272),
.B(n_248),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_234),
.A2(n_220),
.B(n_193),
.Y(n_273)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_273),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_275),
.B(n_277),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_232),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_279),
.A2(n_280),
.B1(n_268),
.B2(n_231),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_281),
.B(n_282),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_243),
.Y(n_282)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_284),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_242),
.Y(n_285)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_251),
.C(n_240),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_259),
.C(n_271),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_287),
.B(n_291),
.Y(n_316)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_288),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_289),
.A2(n_263),
.B1(n_253),
.B2(n_254),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_261),
.B(n_251),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_290),
.B(n_293),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_259),
.B(n_200),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_265),
.B(n_240),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_294),
.A2(n_237),
.B(n_239),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_296),
.B(n_311),
.C(n_307),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_298),
.A2(n_300),
.B1(n_303),
.B2(n_305),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_267),
.Y(n_299)
);

MAJx2_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_309),
.C(n_315),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_278),
.B(n_260),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_301),
.B(n_304),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g303 ( 
.A1(n_292),
.A2(n_249),
.B1(n_246),
.B2(n_238),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_278),
.B(n_260),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_289),
.A2(n_264),
.B1(n_249),
.B2(n_238),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_L g335 ( 
.A1(n_306),
.A2(n_193),
.B(n_207),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_244),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_307),
.B(n_311),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_293),
.B(n_244),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_287),
.A2(n_239),
.B1(n_220),
.B2(n_237),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_284),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_274),
.B(n_208),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_283),
.A2(n_228),
.B(n_207),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_312),
.B(n_288),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_274),
.B(n_220),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_309),
.B(n_283),
.Y(n_317)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_317),
.B(n_319),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_287),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_320),
.A2(n_298),
.B(n_310),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_294),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_321),
.B(n_329),
.Y(n_343)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_323),
.B(n_333),
.Y(n_347)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_308),
.Y(n_325)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_325),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_285),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_326),
.Y(n_337)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_314),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_327),
.B(n_328),
.Y(n_336)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_305),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_SL g329 ( 
.A(n_301),
.B(n_279),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_295),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_330),
.B(n_194),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_299),
.B(n_275),
.C(n_276),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_323),
.C(n_329),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_276),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_184),
.Y(n_349)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_335),
.A2(n_316),
.B(n_313),
.Y(n_339)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_339),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_331),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_340),
.B(n_341),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_317),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_344),
.B(n_324),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_345),
.B(n_318),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_SL g346 ( 
.A1(n_332),
.A2(n_315),
.B1(n_304),
.B2(n_198),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_346),
.A2(n_319),
.B1(n_321),
.B2(n_324),
.Y(n_350)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_348),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_175),
.Y(n_361)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_350),
.B(n_343),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_341),
.B(n_334),
.C(n_322),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_351),
.B(n_354),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_353),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_318),
.Y(n_355)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_355),
.A2(n_338),
.B(n_349),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_L g357 ( 
.A(n_343),
.B(n_165),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_357),
.B(n_361),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_347),
.B(n_198),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_358),
.B(n_200),
.Y(n_371)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_339),
.A2(n_187),
.B(n_184),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g370 ( 
.A1(n_360),
.A2(n_338),
.B1(n_187),
.B2(n_153),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_356),
.A2(n_342),
.B1(n_336),
.B2(n_347),
.Y(n_364)
);

OR2x2_ASAP7_75t_L g373 ( 
.A(n_364),
.B(n_366),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_370),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_359),
.B(n_352),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_368),
.B(n_369),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_355),
.B(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_371),
.B(n_360),
.Y(n_372)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_372),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_363),
.A2(n_351),
.B(n_354),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_SL g382 ( 
.A1(n_375),
.A2(n_379),
.B(n_14),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_365),
.B(n_361),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_378),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_371),
.B(n_357),
.Y(n_378)
);

A2O1A1O1Ixp25_ASAP7_75t_L g379 ( 
.A1(n_367),
.A2(n_140),
.B(n_12),
.C(n_13),
.D(n_15),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_9),
.Y(n_380)
);

OAI321xp33_ASAP7_75t_L g386 ( 
.A1(n_380),
.A2(n_14),
.A3(n_15),
.B1(n_6),
.B2(n_7),
.C(n_4),
.Y(n_386)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_382),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g383 ( 
.A(n_374),
.B(n_14),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_383),
.B(n_7),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_377),
.B(n_373),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g388 ( 
.A(n_385),
.B(n_5),
.Y(n_388)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_386),
.A2(n_372),
.B(n_15),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g391 ( 
.A1(n_387),
.A2(n_388),
.B(n_390),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_389),
.A2(n_381),
.B(n_384),
.Y(n_392)
);

AO21x1_ASAP7_75t_L g393 ( 
.A1(n_392),
.A2(n_5),
.B(n_6),
.Y(n_393)
);

AND2x2_ASAP7_75t_L g394 ( 
.A(n_393),
.B(n_6),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_391),
.C(n_6),
.Y(n_395)
);

BUFx24_ASAP7_75t_SL g396 ( 
.A(n_395),
.Y(n_396)
);


endmodule