module real_aes_2085_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_789, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_789;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g171 ( .A(n_0), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_1), .B(n_110), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_2), .B(n_177), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_3), .B(n_174), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_4), .A2(n_43), .B1(n_447), .B2(n_448), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g447 ( .A(n_4), .Y(n_447) );
INVx1_ASAP7_75t_L g137 ( .A(n_5), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_6), .B(n_177), .Y(n_199) );
NAND2xp33_ASAP7_75t_SL g157 ( .A(n_7), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g128 ( .A(n_8), .Y(n_128) );
CKINVDCx16_ASAP7_75t_R g110 ( .A(n_9), .Y(n_110) );
AND2x2_ASAP7_75t_L g197 ( .A(n_10), .B(n_180), .Y(n_197) );
AND2x2_ASAP7_75t_L g503 ( .A(n_11), .B(n_153), .Y(n_503) );
AND2x2_ASAP7_75t_L g554 ( .A(n_12), .B(n_208), .Y(n_554) );
INVx2_ASAP7_75t_L g131 ( .A(n_13), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_14), .B(n_174), .Y(n_527) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
AOI221x1_ASAP7_75t_L g149 ( .A1(n_16), .A2(n_150), .B1(n_152), .B2(n_153), .C(n_156), .Y(n_149) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_17), .B(n_177), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g559 ( .A(n_18), .B(n_177), .Y(n_559) );
INVx1_ASAP7_75t_L g114 ( .A(n_19), .Y(n_114) );
AOI22xp33_ASAP7_75t_L g507 ( .A1(n_20), .A2(n_92), .B1(n_132), .B2(n_177), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g200 ( .A1(n_21), .A2(n_152), .B(n_201), .Y(n_200) );
AOI221xp5_ASAP7_75t_SL g244 ( .A1(n_22), .A2(n_35), .B1(n_152), .B2(n_177), .C(n_245), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_23), .B(n_172), .Y(n_202) );
OR2x2_ASAP7_75t_L g130 ( .A(n_24), .B(n_91), .Y(n_130) );
OA21x2_ASAP7_75t_L g155 ( .A1(n_24), .A2(n_91), .B(n_131), .Y(n_155) );
INVxp67_ASAP7_75t_L g148 ( .A(n_25), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_26), .B(n_174), .Y(n_239) );
AND2x2_ASAP7_75t_L g191 ( .A(n_27), .B(n_179), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g169 ( .A1(n_28), .A2(n_152), .B(n_170), .Y(n_169) );
AO21x2_ASAP7_75t_L g522 ( .A1(n_29), .A2(n_153), .B(n_523), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_30), .B(n_174), .Y(n_246) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_31), .A2(n_152), .B(n_550), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_32), .B(n_174), .Y(n_535) );
AND2x2_ASAP7_75t_L g139 ( .A(n_33), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g143 ( .A(n_33), .Y(n_143) );
AND2x2_ASAP7_75t_L g158 ( .A(n_33), .B(n_137), .Y(n_158) );
NOR3xp33_ASAP7_75t_L g108 ( .A(n_34), .B(n_109), .C(n_111), .Y(n_108) );
OR2x6_ASAP7_75t_L g458 ( .A(n_34), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_36), .B(n_177), .Y(n_553) );
AOI22xp5_ASAP7_75t_L g211 ( .A1(n_37), .A2(n_84), .B1(n_141), .B2(n_152), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_38), .B(n_174), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_39), .A2(n_48), .B1(n_779), .B2(n_780), .Y(n_778) );
INVx1_ASAP7_75t_L g780 ( .A(n_39), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_40), .B(n_177), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_41), .B(n_172), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_42), .A2(n_152), .B(n_499), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_43), .Y(n_448) );
AND2x2_ASAP7_75t_L g178 ( .A(n_44), .B(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_45), .B(n_172), .Y(n_493) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_46), .B(n_179), .Y(n_248) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_47), .B(n_177), .Y(n_524) );
CKINVDCx20_ASAP7_75t_R g779 ( .A(n_48), .Y(n_779) );
INVx1_ASAP7_75t_L g135 ( .A(n_49), .Y(n_135) );
INVx1_ASAP7_75t_L g162 ( .A(n_49), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_50), .B(n_174), .Y(n_501) );
AND2x2_ASAP7_75t_L g513 ( .A(n_51), .B(n_179), .Y(n_513) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_52), .B(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_SL g189 ( .A(n_53), .B(n_177), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_54), .B(n_172), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_55), .B(n_172), .Y(n_534) );
AND2x2_ASAP7_75t_L g220 ( .A(n_56), .B(n_179), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_57), .B(n_177), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_58), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g515 ( .A(n_59), .B(n_177), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_60), .A2(n_152), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_61), .B(n_172), .Y(n_218) );
AND2x2_ASAP7_75t_SL g240 ( .A(n_62), .B(n_180), .Y(n_240) );
XNOR2xp5_ASAP7_75t_L g777 ( .A(n_63), .B(n_778), .Y(n_777) );
XNOR2x1_ASAP7_75t_SL g117 ( .A(n_64), .B(n_118), .Y(n_117) );
AND2x2_ASAP7_75t_L g565 ( .A(n_64), .B(n_180), .Y(n_565) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_65), .A2(n_152), .B(n_186), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_66), .B(n_174), .Y(n_203) );
AND2x2_ASAP7_75t_SL g212 ( .A(n_67), .B(n_208), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_68), .B(n_172), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_69), .B(n_172), .Y(n_528) );
AOI22xp5_ASAP7_75t_L g508 ( .A1(n_70), .A2(n_94), .B1(n_141), .B2(n_152), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_71), .B(n_466), .Y(n_465) );
XNOR2xp5_ASAP7_75t_L g776 ( .A(n_72), .B(n_777), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_73), .B(n_174), .Y(n_562) );
INVx1_ASAP7_75t_L g140 ( .A(n_74), .Y(n_140) );
INVx1_ASAP7_75t_L g164 ( .A(n_74), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_75), .B(n_172), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_76), .A2(n_152), .B(n_517), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_77), .A2(n_152), .B(n_491), .Y(n_490) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_78), .A2(n_152), .B(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g537 ( .A(n_79), .B(n_180), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g505 ( .A(n_80), .B(n_179), .Y(n_505) );
AOI22xp5_ASAP7_75t_L g210 ( .A1(n_81), .A2(n_86), .B1(n_132), .B2(n_177), .Y(n_210) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_82), .B(n_177), .Y(n_219) );
INVxp33_ASAP7_75t_L g785 ( .A(n_83), .Y(n_785) );
NOR2xp33_ASAP7_75t_L g113 ( .A(n_85), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g460 ( .A(n_85), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_87), .B(n_172), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_88), .B(n_172), .Y(n_247) );
AND2x2_ASAP7_75t_L g494 ( .A(n_89), .B(n_208), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_90), .A2(n_152), .B(n_216), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_93), .B(n_174), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_95), .A2(n_152), .B(n_561), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_96), .B(n_174), .Y(n_492) );
OAI22x1_ASAP7_75t_R g444 ( .A1(n_97), .A2(n_445), .B1(n_446), .B2(n_449), .Y(n_444) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_97), .Y(n_449) );
INVxp67_ASAP7_75t_L g151 ( .A(n_98), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_99), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_100), .B(n_174), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_101), .A2(n_152), .B(n_237), .Y(n_236) );
BUFx2_ASAP7_75t_L g564 ( .A(n_102), .Y(n_564) );
BUFx2_ASAP7_75t_L g451 ( .A(n_103), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_115), .B(n_784), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx20_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
BUFx4f_ASAP7_75t_SL g787 ( .A(n_107), .Y(n_787) );
NAND2xp5_ASAP7_75t_SL g107 ( .A(n_108), .B(n_113), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_112), .B(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g469 ( .A(n_112), .B(n_458), .Y(n_469) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_112), .B(n_458), .Y(n_477) );
OR2x6_ASAP7_75t_SL g481 ( .A(n_112), .B(n_457), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_114), .B(n_460), .Y(n_459) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_462), .Y(n_115) );
AOI22x1_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_450), .B1(n_453), .B2(n_461), .Y(n_116) );
OAI22x1_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_120), .B1(n_443), .B2(n_444), .Y(n_118) );
OAI22x1_ASAP7_75t_L g782 ( .A1(n_119), .A2(n_476), .B1(n_479), .B2(n_783), .Y(n_782) );
INVx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OA22x2_ASAP7_75t_L g475 ( .A1(n_120), .A2(n_476), .B1(n_478), .B2(n_482), .Y(n_475) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_320), .Y(n_120) );
NOR4xp25_ASAP7_75t_L g121 ( .A(n_122), .B(n_263), .C(n_302), .D(n_309), .Y(n_121) );
OAI221xp5_ASAP7_75t_L g122 ( .A1(n_123), .A2(n_181), .B1(n_221), .B2(n_230), .C(n_249), .Y(n_122) );
OR2x2_ASAP7_75t_L g393 ( .A(n_123), .B(n_255), .Y(n_393) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
AND2x2_ASAP7_75t_L g308 ( .A(n_124), .B(n_233), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_124), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_SL g373 ( .A(n_124), .B(n_374), .Y(n_373) );
AND2x4_ASAP7_75t_L g124 ( .A(n_125), .B(n_165), .Y(n_124) );
AND2x4_ASAP7_75t_SL g232 ( .A(n_125), .B(n_233), .Y(n_232) );
INVx3_ASAP7_75t_L g254 ( .A(n_125), .Y(n_254) );
AND2x2_ASAP7_75t_L g289 ( .A(n_125), .B(n_262), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_125), .B(n_166), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_125), .B(n_256), .Y(n_341) );
OR2x2_ASAP7_75t_L g419 ( .A(n_125), .B(n_233), .Y(n_419) );
AND2x4_ASAP7_75t_L g125 ( .A(n_126), .B(n_149), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_132), .B1(n_141), .B2(n_147), .Y(n_126) );
NOR2xp33_ASAP7_75t_L g127 ( .A(n_128), .B(n_129), .Y(n_127) );
NOR2xp33_ASAP7_75t_L g147 ( .A(n_129), .B(n_148), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g150 ( .A(n_129), .B(n_151), .Y(n_150) );
NOR3xp33_ASAP7_75t_L g156 ( .A(n_129), .B(n_157), .C(n_159), .Y(n_156) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_129), .A2(n_199), .B(n_200), .Y(n_198) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_129), .A2(n_515), .B(n_516), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_129), .A2(n_524), .B(n_525), .Y(n_523) );
AND2x4_ASAP7_75t_L g129 ( .A(n_130), .B(n_131), .Y(n_129) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_130), .B(n_131), .Y(n_180) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_138), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_136), .Y(n_133) );
INVx2_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
AND2x2_ASAP7_75t_L g146 ( .A(n_135), .B(n_137), .Y(n_146) );
AND2x4_ASAP7_75t_L g174 ( .A(n_135), .B(n_163), .Y(n_174) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g152 ( .A(n_139), .B(n_146), .Y(n_152) );
INVx2_ASAP7_75t_L g145 ( .A(n_140), .Y(n_145) );
AND2x6_ASAP7_75t_L g172 ( .A(n_140), .B(n_161), .Y(n_172) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NOR2x1p5_ASAP7_75t_L g142 ( .A(n_143), .B(n_144), .Y(n_142) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx3_ASAP7_75t_L g530 ( .A(n_153), .Y(n_530) );
INVx4_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AOI21x1_ASAP7_75t_L g167 ( .A1(n_154), .A2(n_168), .B(n_178), .Y(n_167) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_154), .A2(n_497), .B(n_503), .Y(n_496) );
INVx3_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
BUFx4f_ASAP7_75t_L g208 ( .A(n_155), .Y(n_208) );
INVx5_ASAP7_75t_L g175 ( .A(n_158), .Y(n_175) );
AND2x4_ASAP7_75t_L g177 ( .A(n_158), .B(n_160), .Y(n_177) );
INVx1_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g160 ( .A(n_161), .B(n_163), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx2_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
AND2x2_ASAP7_75t_L g241 ( .A(n_166), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_166), .B(n_262), .Y(n_261) );
INVx1_ASAP7_75t_L g267 ( .A(n_166), .Y(n_267) );
OR2x2_ASAP7_75t_L g272 ( .A(n_166), .B(n_256), .Y(n_272) );
AND2x2_ASAP7_75t_L g285 ( .A(n_166), .B(n_243), .Y(n_285) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_166), .Y(n_288) );
INVx1_ASAP7_75t_L g300 ( .A(n_166), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_166), .B(n_254), .Y(n_365) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_169), .B(n_176), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_173), .B(n_175), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_172), .B(n_564), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_175), .A2(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g201 ( .A1(n_175), .A2(n_202), .B(n_203), .Y(n_201) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_175), .A2(n_217), .B(n_218), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_175), .A2(n_238), .B(n_239), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_175), .A2(n_246), .B(n_247), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_175), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_175), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g517 ( .A1(n_175), .A2(n_518), .B(n_519), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_175), .A2(n_527), .B(n_528), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g533 ( .A1(n_175), .A2(n_534), .B(n_535), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_175), .A2(n_551), .B(n_552), .Y(n_550) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_175), .A2(n_562), .B(n_563), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g190 ( .A(n_179), .Y(n_190) );
OA21x2_ASAP7_75t_L g243 ( .A1(n_179), .A2(n_244), .B(n_248), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_179), .A2(n_489), .B(n_490), .Y(n_488) );
AO21x2_ASAP7_75t_L g506 ( .A1(n_179), .A2(n_507), .B(n_508), .Y(n_506) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_182), .B(n_192), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
OR2x2_ASAP7_75t_L g229 ( .A(n_183), .B(n_213), .Y(n_229) );
AND2x4_ASAP7_75t_L g259 ( .A(n_183), .B(n_196), .Y(n_259) );
INVx2_ASAP7_75t_L g293 ( .A(n_183), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g351 ( .A(n_183), .B(n_213), .Y(n_351) );
AND2x2_ASAP7_75t_L g398 ( .A(n_183), .B(n_227), .Y(n_398) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_184), .A2(n_190), .B(n_191), .Y(n_183) );
AO21x2_ASAP7_75t_L g251 ( .A1(n_184), .A2(n_190), .B(n_191), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_185), .B(n_189), .Y(n_184) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_190), .A2(n_214), .B(n_220), .Y(n_213) );
AOI21x1_ASAP7_75t_L g547 ( .A1(n_190), .A2(n_548), .B(n_554), .Y(n_547) );
AOI222xp33_ASAP7_75t_L g386 ( .A1(n_192), .A2(n_258), .B1(n_301), .B2(n_361), .C1(n_387), .C2(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_194), .B(n_204), .Y(n_193) );
AND2x2_ASAP7_75t_L g305 ( .A(n_194), .B(n_225), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g355 ( .A(n_194), .B(n_356), .Y(n_355) );
AND2x2_ASAP7_75t_L g434 ( .A(n_194), .B(n_274), .Y(n_434) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_195), .A2(n_265), .B(n_269), .Y(n_264) );
AND2x2_ASAP7_75t_L g345 ( .A(n_195), .B(n_228), .Y(n_345) );
OR2x2_ASAP7_75t_L g370 ( .A(n_195), .B(n_229), .Y(n_370) );
INVx2_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx5_ASAP7_75t_L g224 ( .A(n_196), .Y(n_224) );
AND2x2_ASAP7_75t_L g311 ( .A(n_196), .B(n_293), .Y(n_311) );
AND2x2_ASAP7_75t_L g337 ( .A(n_196), .B(n_213), .Y(n_337) );
OR2x2_ASAP7_75t_L g340 ( .A(n_196), .B(n_227), .Y(n_340) );
HB1xp67_ASAP7_75t_L g358 ( .A(n_196), .Y(n_358) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_196), .B(n_292), .Y(n_415) );
OR2x2_ASAP7_75t_L g424 ( .A(n_196), .B(n_251), .Y(n_424) );
OR2x6_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_L g257 ( .A(n_204), .Y(n_257) );
AOI221xp5_ASAP7_75t_SL g375 ( .A1(n_204), .A2(n_259), .B1(n_376), .B2(n_378), .C(n_379), .Y(n_375) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_213), .Y(n_204) );
OR2x2_ASAP7_75t_L g314 ( .A(n_205), .B(n_284), .Y(n_314) );
OR2x2_ASAP7_75t_L g324 ( .A(n_205), .B(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g350 ( .A(n_205), .B(n_351), .Y(n_350) );
AND2x4_ASAP7_75t_L g356 ( .A(n_205), .B(n_275), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g368 ( .A(n_205), .B(n_339), .Y(n_368) );
INVx2_ASAP7_75t_L g381 ( .A(n_205), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g402 ( .A(n_205), .B(n_259), .Y(n_402) );
AND2x2_ASAP7_75t_L g406 ( .A(n_205), .B(n_228), .Y(n_406) );
AND2x2_ASAP7_75t_L g414 ( .A(n_205), .B(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
INVx2_ASAP7_75t_L g227 ( .A(n_206), .Y(n_227) );
AOI21x1_ASAP7_75t_L g206 ( .A1(n_207), .A2(n_209), .B(n_212), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_208), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_208), .A2(n_235), .B(n_236), .Y(n_234) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_208), .A2(n_559), .B(n_560), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_210), .B(n_211), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_213), .B(n_224), .Y(n_223) );
AND2x2_ASAP7_75t_L g258 ( .A(n_213), .B(n_227), .Y(n_258) );
INVx2_ASAP7_75t_L g275 ( .A(n_213), .Y(n_275) );
AND2x4_ASAP7_75t_L g292 ( .A(n_213), .B(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g397 ( .A(n_213), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_219), .Y(n_214) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_222), .B(n_225), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g404 ( .A(n_223), .B(n_226), .Y(n_404) );
AND2x4_ASAP7_75t_L g250 ( .A(n_224), .B(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g291 ( .A(n_224), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g318 ( .A(n_224), .B(n_258), .Y(n_318) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_228), .Y(n_225) );
AND2x2_ASAP7_75t_L g422 ( .A(n_226), .B(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
AND2x2_ASAP7_75t_L g274 ( .A(n_227), .B(n_275), .Y(n_274) );
OAI21xp5_ASAP7_75t_SL g294 ( .A1(n_228), .A2(n_295), .B(n_301), .Y(n_294) );
INVx2_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
INVx1_ASAP7_75t_SL g230 ( .A(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_232), .B(n_241), .Y(n_231) );
INVx1_ASAP7_75t_SL g348 ( .A(n_232), .Y(n_348) );
AND2x2_ASAP7_75t_L g378 ( .A(n_232), .B(n_288), .Y(n_378) );
AND2x4_ASAP7_75t_L g389 ( .A(n_232), .B(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g255 ( .A(n_233), .B(n_256), .Y(n_255) );
INVx2_ASAP7_75t_L g262 ( .A(n_233), .Y(n_262) );
AND2x4_ASAP7_75t_L g268 ( .A(n_233), .B(n_254), .Y(n_268) );
INVx2_ASAP7_75t_L g279 ( .A(n_233), .Y(n_279) );
INVx1_ASAP7_75t_L g328 ( .A(n_233), .Y(n_328) );
OR2x2_ASAP7_75t_L g349 ( .A(n_233), .B(n_333), .Y(n_349) );
OR2x2_ASAP7_75t_L g363 ( .A(n_233), .B(n_243), .Y(n_363) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_233), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_233), .B(n_285), .Y(n_435) );
OR2x6_ASAP7_75t_L g233 ( .A(n_234), .B(n_240), .Y(n_233) );
INVx1_ASAP7_75t_L g280 ( .A(n_241), .Y(n_280) );
AND2x2_ASAP7_75t_L g413 ( .A(n_241), .B(n_279), .Y(n_413) );
AND2x2_ASAP7_75t_L g438 ( .A(n_241), .B(n_268), .Y(n_438) );
INVx2_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx2_ASAP7_75t_L g256 ( .A(n_243), .Y(n_256) );
BUFx3_ASAP7_75t_L g298 ( .A(n_243), .Y(n_298) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_243), .Y(n_325) );
INVx1_ASAP7_75t_L g334 ( .A(n_243), .Y(n_334) );
AOI33xp33_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_252), .A3(n_257), .B1(n_258), .B2(n_259), .B3(n_260), .Y(n_249) );
AOI21x1_ASAP7_75t_SL g352 ( .A1(n_250), .A2(n_274), .B(n_336), .Y(n_352) );
INVx2_ASAP7_75t_L g382 ( .A(n_250), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g388 ( .A(n_250), .B(n_381), .Y(n_388) );
AND2x2_ASAP7_75t_L g336 ( .A(n_251), .B(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g252 ( .A(n_253), .Y(n_252) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g299 ( .A(n_254), .B(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g400 ( .A(n_255), .Y(n_400) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_256), .Y(n_390) );
OAI32xp33_ASAP7_75t_L g439 ( .A1(n_257), .A2(n_259), .A3(n_435), .B1(n_440), .B2(n_442), .Y(n_439) );
AND2x2_ASAP7_75t_L g357 ( .A(n_258), .B(n_358), .Y(n_357) );
INVx2_ASAP7_75t_SL g347 ( .A(n_259), .Y(n_347) );
AND2x2_ASAP7_75t_L g412 ( .A(n_259), .B(n_356), .Y(n_412) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI221xp5_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_273), .B1(n_276), .B2(n_290), .C(n_294), .Y(n_263) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_268), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_267), .B(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_268), .B(n_271), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_268), .B(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_268), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR3xp33_ASAP7_75t_L g276 ( .A(n_277), .B(n_281), .C(n_286), .Y(n_276) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_278), .A2(n_340), .B1(n_380), .B2(n_383), .Y(n_379) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx1_ASAP7_75t_L g283 ( .A(n_279), .Y(n_283) );
NOR2x1p5_ASAP7_75t_L g297 ( .A(n_279), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g319 ( .A(n_279), .Y(n_319) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI322xp33_ASAP7_75t_L g346 ( .A1(n_282), .A2(n_324), .A3(n_347), .B1(n_348), .B2(n_349), .C1(n_350), .C2(n_352), .Y(n_346) );
OR2x2_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g302 ( .A1(n_284), .A2(n_303), .B(n_304), .C(n_306), .Y(n_302) );
OR2x2_ASAP7_75t_L g394 ( .A(n_284), .B(n_348), .Y(n_394) );
INVx2_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_L g301 ( .A(n_285), .B(n_289), .Y(n_301) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_288), .B(n_289), .Y(n_287) );
INVx2_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g307 ( .A(n_291), .B(n_308), .Y(n_307) );
INVx3_ASAP7_75t_SL g339 ( .A(n_292), .Y(n_339) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_296), .B(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_299), .Y(n_296) );
INVx1_ASAP7_75t_SL g343 ( .A(n_299), .Y(n_343) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_300), .Y(n_385) );
OR2x6_ASAP7_75t_SL g440 ( .A(n_303), .B(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVxp67_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
AOI211xp5_ASAP7_75t_L g430 ( .A1(n_308), .A2(n_431), .B(n_432), .C(n_439), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_312), .B(n_315), .C(n_319), .Y(n_309) );
OAI211xp5_ASAP7_75t_SL g321 ( .A1(n_310), .A2(n_322), .B(n_329), .C(n_353), .Y(n_321) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVxp67_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_318), .Y(n_316) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_321), .B(n_366), .C(n_410), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_323), .B(n_326), .Y(n_322) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g417 ( .A(n_325), .Y(n_417) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g372 ( .A(n_328), .Y(n_372) );
NOR3xp33_ASAP7_75t_SL g329 ( .A(n_330), .B(n_342), .C(n_346), .Y(n_329) );
OAI22xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_335), .B1(n_338), .B2(n_341), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
INVxp67_ASAP7_75t_SL g441 ( .A(n_334), .Y(n_441) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_340), .Y(n_338) );
INVx1_ASAP7_75t_SL g427 ( .A(n_340), .Y(n_427) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
OR2x2_ASAP7_75t_L g377 ( .A(n_343), .B(n_363), .Y(n_377) );
OR2x2_ASAP7_75t_L g428 ( .A(n_343), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g426 ( .A(n_351), .Y(n_426) );
OR2x2_ASAP7_75t_L g442 ( .A(n_351), .B(n_381), .Y(n_442) );
OAI21xp33_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_357), .B(n_359), .Y(n_353) );
OAI31xp33_ASAP7_75t_L g367 ( .A1(n_354), .A2(n_368), .A3(n_369), .B(n_371), .Y(n_367) );
INVx1_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
AND2x2_ASAP7_75t_L g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AND2x4_ASAP7_75t_L g399 ( .A(n_364), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
NAND4xp25_ASAP7_75t_SL g366 ( .A(n_367), .B(n_375), .C(n_386), .D(n_391), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_374), .Y(n_409) );
INVx1_ASAP7_75t_SL g376 ( .A(n_377), .Y(n_376) );
OR2x2_ASAP7_75t_L g380 ( .A(n_381), .B(n_382), .Y(n_380) );
INVxp67_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_395), .B1(n_399), .B2(n_401), .C(n_403), .Y(n_391) );
NAND2xp33_ASAP7_75t_SL g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g436 ( .A(n_395), .Y(n_436) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_396), .B(n_398), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
AOI21xp33_ASAP7_75t_L g403 ( .A1(n_404), .A2(n_405), .B(n_407), .Y(n_403) );
INVx1_ASAP7_75t_L g431 ( .A(n_405), .Y(n_431) );
INVx2_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_411), .B(n_430), .Y(n_410) );
AOI221xp5_ASAP7_75t_L g411 ( .A1(n_412), .A2(n_413), .B1(n_414), .B2(n_416), .C(n_420), .Y(n_411) );
AND2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx1_ASAP7_75t_SL g418 ( .A(n_419), .Y(n_418) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_425), .B(n_428), .Y(n_420) );
INVxp33_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_435), .B1(n_436), .B2(n_437), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVxp33_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NOR2x1_ASAP7_75t_R g461 ( .A(n_451), .B(n_456), .Y(n_461) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_451), .Y(n_473) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
NAND3xp33_ASAP7_75t_L g464 ( .A(n_453), .B(n_465), .C(n_470), .Y(n_464) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_458), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_463), .B(n_781), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx3_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
CKINVDCx5p33_ASAP7_75t_R g470 ( .A(n_471), .Y(n_470) );
BUFx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_473), .Y(n_472) );
NOR2xp33_ASAP7_75t_L g474 ( .A(n_475), .B(n_776), .Y(n_474) );
CKINVDCx11_ASAP7_75t_R g476 ( .A(n_477), .Y(n_476) );
BUFx4f_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
CKINVDCx20_ASAP7_75t_R g479 ( .A(n_480), .Y(n_479) );
CKINVDCx11_ASAP7_75t_R g480 ( .A(n_481), .Y(n_480) );
INVx3_ASAP7_75t_SL g783 ( .A(n_482), .Y(n_783) );
AND2x4_ASAP7_75t_SL g482 ( .A(n_483), .B(n_672), .Y(n_482) );
NOR3xp33_ASAP7_75t_SL g483 ( .A(n_484), .B(n_581), .C(n_613), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_509), .B1(n_538), .B2(n_555), .C(n_566), .Y(n_484) );
OR2x2_ASAP7_75t_L g485 ( .A(n_486), .B(n_495), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
AND2x2_ASAP7_75t_L g544 ( .A(n_487), .B(n_496), .Y(n_544) );
INVx4_ASAP7_75t_L g572 ( .A(n_487), .Y(n_572) );
AND2x4_ASAP7_75t_SL g612 ( .A(n_487), .B(n_546), .Y(n_612) );
BUFx2_ASAP7_75t_L g622 ( .A(n_487), .Y(n_622) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_487), .B(n_627), .Y(n_688) );
AND2x2_ASAP7_75t_L g697 ( .A(n_487), .B(n_625), .Y(n_697) );
OR2x2_ASAP7_75t_L g705 ( .A(n_487), .B(n_706), .Y(n_705) );
AND2x2_ASAP7_75t_L g731 ( .A(n_487), .B(n_570), .Y(n_731) );
AND2x4_ASAP7_75t_L g750 ( .A(n_487), .B(n_751), .Y(n_750) );
OR2x6_ASAP7_75t_L g487 ( .A(n_488), .B(n_494), .Y(n_487) );
INVx2_ASAP7_75t_SL g663 ( .A(n_495), .Y(n_663) );
OR2x2_ASAP7_75t_L g495 ( .A(n_496), .B(n_504), .Y(n_495) );
AND2x2_ASAP7_75t_L g570 ( .A(n_496), .B(n_547), .Y(n_570) );
INVx2_ASAP7_75t_L g597 ( .A(n_496), .Y(n_597) );
INVx2_ASAP7_75t_L g627 ( .A(n_496), .Y(n_627) );
AND2x2_ASAP7_75t_L g641 ( .A(n_496), .B(n_546), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_502), .Y(n_497) );
AND2x2_ASAP7_75t_L g571 ( .A(n_504), .B(n_572), .Y(n_571) );
INVx2_ASAP7_75t_L g594 ( .A(n_504), .Y(n_594) );
BUFx3_ASAP7_75t_L g608 ( .A(n_504), .Y(n_608) );
AND2x2_ASAP7_75t_L g637 ( .A(n_504), .B(n_638), .Y(n_637) );
AND2x4_ASAP7_75t_L g504 ( .A(n_505), .B(n_506), .Y(n_504) );
AND2x4_ASAP7_75t_L g542 ( .A(n_505), .B(n_506), .Y(n_542) );
INVx1_ASAP7_75t_L g643 ( .A(n_509), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_520), .Y(n_509) );
OR2x2_ASAP7_75t_L g754 ( .A(n_510), .B(n_555), .Y(n_754) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g610 ( .A(n_511), .B(n_611), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_511), .B(n_520), .Y(n_671) );
OR2x2_ASAP7_75t_L g769 ( .A(n_511), .B(n_691), .Y(n_769) );
INVx2_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
AND2x2_ASAP7_75t_L g580 ( .A(n_512), .B(n_556), .Y(n_580) );
OR2x2_ASAP7_75t_SL g590 ( .A(n_512), .B(n_591), .Y(n_590) );
INVx4_ASAP7_75t_L g601 ( .A(n_512), .Y(n_601) );
HB1xp67_ASAP7_75t_L g652 ( .A(n_512), .Y(n_652) );
NAND2x1_ASAP7_75t_L g658 ( .A(n_512), .B(n_557), .Y(n_658) );
AND2x2_ASAP7_75t_L g683 ( .A(n_512), .B(n_522), .Y(n_683) );
OR2x2_ASAP7_75t_L g704 ( .A(n_512), .B(n_587), .Y(n_704) );
OR2x6_ASAP7_75t_L g512 ( .A(n_513), .B(n_514), .Y(n_512) );
INVx1_ASAP7_75t_L g599 ( .A(n_520), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g692 ( .A1(n_520), .A2(n_693), .B(n_696), .C(n_698), .Y(n_692) );
AND2x2_ASAP7_75t_L g765 ( .A(n_520), .B(n_541), .Y(n_765) );
AND2x2_ASAP7_75t_L g520 ( .A(n_521), .B(n_529), .Y(n_520) );
INVx1_ASAP7_75t_L g632 ( .A(n_521), .Y(n_632) );
AND2x2_ASAP7_75t_L g702 ( .A(n_521), .B(n_557), .Y(n_702) );
INVx2_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g576 ( .A(n_522), .Y(n_576) );
OR2x2_ASAP7_75t_L g591 ( .A(n_522), .B(n_557), .Y(n_591) );
INVx1_ASAP7_75t_L g607 ( .A(n_522), .Y(n_607) );
AND2x2_ASAP7_75t_L g619 ( .A(n_522), .B(n_529), .Y(n_619) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_522), .Y(n_725) );
NOR2x1_ASAP7_75t_SL g556 ( .A(n_529), .B(n_557), .Y(n_556) );
AO21x1_ASAP7_75t_SL g529 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_529) );
AO21x2_ASAP7_75t_L g588 ( .A1(n_530), .A2(n_531), .B(n_537), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_536), .Y(n_531) );
INVxp67_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_543), .Y(n_539) );
OR2x2_ASAP7_75t_L g689 ( .A(n_540), .B(n_624), .Y(n_689) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_541), .B(n_707), .Y(n_706) );
OR2x2_ASAP7_75t_L g771 ( .A(n_541), .B(n_668), .Y(n_771) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g616 ( .A(n_542), .B(n_597), .Y(n_616) );
AND2x2_ASAP7_75t_L g712 ( .A(n_542), .B(n_625), .Y(n_712) );
INVx1_ASAP7_75t_L g629 ( .A(n_543), .Y(n_629) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
INVx1_ASAP7_75t_L g679 ( .A(n_544), .Y(n_679) );
INVx2_ASAP7_75t_L g646 ( .A(n_545), .Y(n_646) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g596 ( .A(n_546), .B(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g626 ( .A(n_546), .Y(n_626) );
INVx1_ASAP7_75t_L g751 ( .A(n_546), .Y(n_751) );
INVx3_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_547), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_549), .B(n_553), .Y(n_548) );
OR2x2_ASAP7_75t_L g722 ( .A(n_555), .B(n_723), .Y(n_722) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx2_ASAP7_75t_SL g577 ( .A(n_557), .Y(n_577) );
OR2x2_ASAP7_75t_L g600 ( .A(n_557), .B(n_601), .Y(n_600) );
AND2x2_ASAP7_75t_L g611 ( .A(n_557), .B(n_587), .Y(n_611) );
AND2x2_ASAP7_75t_L g685 ( .A(n_557), .B(n_601), .Y(n_685) );
BUFx2_ASAP7_75t_L g768 ( .A(n_557), .Y(n_768) );
OR2x6_ASAP7_75t_L g557 ( .A(n_558), .B(n_565), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_573), .B(n_578), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .Y(n_568) );
AND2x2_ASAP7_75t_L g720 ( .A(n_569), .B(n_642), .Y(n_720) );
BUFx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g579 ( .A(n_570), .B(n_572), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_571), .B(n_641), .Y(n_742) );
INVx1_ASAP7_75t_L g772 ( .A(n_571), .Y(n_772) );
NAND2x1p5_ASAP7_75t_L g668 ( .A(n_572), .B(n_669), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_572), .B(n_708), .Y(n_745) );
INVxp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_575), .B(n_577), .Y(n_574) );
AND2x4_ASAP7_75t_SL g609 ( .A(n_575), .B(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_575), .B(n_603), .Y(n_756) );
INVx3_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_576), .B(n_658), .Y(n_714) );
AND2x2_ASAP7_75t_L g732 ( .A(n_576), .B(n_685), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_577), .B(n_619), .Y(n_635) );
A2O1A1Ixp33_ASAP7_75t_L g664 ( .A1(n_577), .A2(n_623), .B(n_665), .C(n_670), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_577), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_580), .Y(n_578) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_579), .A2(n_652), .B1(n_760), .B2(n_766), .C(n_770), .Y(n_759) );
INVx1_ASAP7_75t_SL g747 ( .A(n_580), .Y(n_747) );
OAI221xp5_ASAP7_75t_L g581 ( .A1(n_582), .A2(n_592), .B1(n_598), .B2(n_602), .C(n_789), .Y(n_581) );
INVx2_ASAP7_75t_SL g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g657 ( .A(n_586), .Y(n_657) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
AND2x2_ASAP7_75t_L g631 ( .A(n_587), .B(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g662 ( .A(n_587), .B(n_607), .Y(n_662) );
INVx2_ASAP7_75t_L g695 ( .A(n_587), .Y(n_695) );
INVx3_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI32xp33_ASAP7_75t_L g746 ( .A1(n_590), .A2(n_637), .A3(n_668), .B1(n_747), .B2(n_748), .Y(n_746) );
OR2x2_ASAP7_75t_L g717 ( .A(n_591), .B(n_704), .Y(n_717) );
INVx1_ASAP7_75t_L g727 ( .A(n_592), .Y(n_727) );
OR2x2_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx2_ASAP7_75t_L g642 ( .A(n_593), .Y(n_642) );
AND2x2_ASAP7_75t_L g713 ( .A(n_593), .B(n_688), .Y(n_713) );
OR2x2_ASAP7_75t_L g744 ( .A(n_593), .B(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_594), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g638 ( .A(n_597), .Y(n_638) );
OR2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx2_ASAP7_75t_SL g603 ( .A(n_600), .Y(n_603) );
OR2x2_ASAP7_75t_L g690 ( .A(n_600), .B(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_601), .B(n_619), .Y(n_618) );
NOR2xp67_ASAP7_75t_L g724 ( .A(n_601), .B(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g737 ( .A(n_601), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_609), .C(n_612), .Y(n_602) );
AND2x2_ASAP7_75t_L g752 ( .A(n_604), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
BUFx2_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
OR2x2_ASAP7_75t_L g678 ( .A(n_608), .B(n_679), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_608), .B(n_612), .Y(n_699) );
AND2x2_ASAP7_75t_L g730 ( .A(n_608), .B(n_731), .Y(n_730) );
O2A1O1Ixp33_ASAP7_75t_L g740 ( .A1(n_610), .A2(n_741), .B(n_743), .C(n_746), .Y(n_740) );
AOI222xp33_ASAP7_75t_L g614 ( .A1(n_611), .A2(n_615), .B1(n_617), .B2(n_620), .C1(n_628), .C2(n_630), .Y(n_614) );
AND2x2_ASAP7_75t_L g682 ( .A(n_611), .B(n_683), .Y(n_682) );
AND2x2_ASAP7_75t_L g615 ( .A(n_612), .B(n_616), .Y(n_615) );
INVx2_ASAP7_75t_SL g636 ( .A(n_612), .Y(n_636) );
NAND4xp25_ASAP7_75t_L g613 ( .A(n_614), .B(n_633), .C(n_654), .D(n_664), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_616), .B(n_622), .Y(n_676) );
INVx1_ASAP7_75t_SL g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g684 ( .A(n_619), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g691 ( .A(n_619), .Y(n_691) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
A2O1A1Ixp33_ASAP7_75t_L g654 ( .A1(n_621), .A2(n_655), .B(n_659), .C(n_663), .Y(n_654) );
INVx2_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_622), .B(n_637), .Y(n_758) );
OR2x2_ASAP7_75t_L g762 ( .A(n_622), .B(n_648), .Y(n_762) );
INVx1_ASAP7_75t_L g735 ( .A(n_623), .Y(n_735) );
INVx2_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
INVx1_ASAP7_75t_SL g669 ( .A(n_626), .Y(n_669) );
INVx1_ASAP7_75t_L g649 ( .A(n_627), .Y(n_649) );
INVx2_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_629), .B(n_666), .Y(n_665) );
BUFx2_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g653 ( .A(n_631), .Y(n_653) );
AOI322xp5_ASAP7_75t_L g633 ( .A1(n_634), .A2(n_636), .A3(n_637), .B1(n_639), .B2(n_643), .C1(n_644), .C2(n_650), .Y(n_633) );
INVxp67_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
O2A1O1Ixp33_ASAP7_75t_SL g715 ( .A1(n_636), .A2(n_716), .B(n_717), .C(n_718), .Y(n_715) );
INVx1_ASAP7_75t_L g738 ( .A(n_637), .Y(n_738) );
NOR2xp67_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g696 ( .A(n_642), .B(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_647), .Y(n_644) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_648), .Y(n_718) );
INVx2_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
OR2x2_ASAP7_75t_L g651 ( .A(n_652), .B(n_653), .Y(n_651) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
OR2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
INVx3_ASAP7_75t_L g661 ( .A(n_658), .Y(n_661) );
OR2x2_ASAP7_75t_L g729 ( .A(n_658), .B(n_691), .Y(n_729) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_658), .B(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
INVx1_ASAP7_75t_SL g761 ( .A(n_662), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_663), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
NAND3xp33_ASAP7_75t_SL g766 ( .A(n_671), .B(n_767), .C(n_769), .Y(n_766) );
NOR3xp33_ASAP7_75t_SL g672 ( .A(n_673), .B(n_710), .C(n_739), .Y(n_672) );
NAND2xp5_ASAP7_75t_SL g673 ( .A(n_674), .B(n_692), .Y(n_673) );
O2A1O1Ixp33_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_677), .B(n_680), .C(n_686), .Y(n_674) );
OAI31xp33_ASAP7_75t_L g719 ( .A1(n_675), .A2(n_697), .A3(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_SL g675 ( .A(n_676), .Y(n_675) );
INVx1_ASAP7_75t_SL g677 ( .A(n_678), .Y(n_677) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g681 ( .A(n_682), .B(n_684), .Y(n_681) );
INVx2_ASAP7_75t_L g734 ( .A(n_682), .Y(n_734) );
INVx1_ASAP7_75t_L g709 ( .A(n_684), .Y(n_709) );
AOI21xp5_ASAP7_75t_L g686 ( .A1(n_687), .A2(n_689), .B(n_690), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
OR2x2_ASAP7_75t_L g736 ( .A(n_694), .B(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g775 ( .A(n_695), .Y(n_775) );
OAI22xp33_ASAP7_75t_SL g698 ( .A1(n_699), .A2(n_700), .B1(n_705), .B2(n_709), .Y(n_698) );
INVx3_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
AND2x4_ASAP7_75t_L g701 ( .A(n_702), .B(n_703), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g716 ( .A(n_704), .Y(n_716) );
OR2x2_ASAP7_75t_L g767 ( .A(n_704), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
NAND3xp33_ASAP7_75t_SL g710 ( .A(n_711), .B(n_719), .C(n_726), .Y(n_710) );
O2A1O1Ixp33_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B(n_714), .C(n_715), .Y(n_711) );
INVx2_ASAP7_75t_L g748 ( .A(n_712), .Y(n_748) );
INVx1_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_728), .B1(n_730), .B2(n_732), .C(n_733), .Y(n_726) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
OAI22xp33_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B1(n_736), .B2(n_738), .Y(n_733) );
NAND3xp33_ASAP7_75t_SL g739 ( .A(n_740), .B(n_749), .C(n_759), .Y(n_739) );
INVxp33_ASAP7_75t_SL g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_SL g743 ( .A(n_744), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_750), .A2(n_752), .B1(n_755), .B2(n_757), .Y(n_749) );
INVx2_ASAP7_75t_L g763 ( .A(n_750), .Y(n_763) );
INVx1_ASAP7_75t_L g753 ( .A(n_754), .Y(n_753) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
OAI22xp5_ASAP7_75t_L g760 ( .A1(n_761), .A2(n_762), .B1(n_763), .B2(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
OAI22xp33_ASAP7_75t_SL g770 ( .A1(n_769), .A2(n_771), .B1(n_772), .B2(n_773), .Y(n_770) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
NAND2xp33_ASAP7_75t_SL g781 ( .A(n_776), .B(n_782), .Y(n_781) );
NOR2xp33_ASAP7_75t_L g784 ( .A(n_785), .B(n_786), .Y(n_784) );
INVx1_ASAP7_75t_SL g786 ( .A(n_787), .Y(n_786) );
endmodule