module fake_netlist_6_4809_n_915 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_199, n_138, n_22, n_161, n_208, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_206, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_204, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_203, n_142, n_20, n_143, n_207, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_205, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_202, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_200, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_201, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_915);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_199;
input n_138;
input n_22;
input n_161;
input n_208;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_206;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_204;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_203;
input n_142;
input n_20;
input n_143;
input n_207;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_205;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_202;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_200;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_201;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_915;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_310;
wire n_509;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_400;
wire n_284;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_832;
wire n_280;
wire n_287;
wire n_685;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_447;
wire n_872;
wire n_222;
wire n_300;
wire n_248;
wire n_718;
wire n_517;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_901;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_343;
wire n_844;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_800;
wire n_779;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_859;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_286;
wire n_254;
wire n_834;
wire n_242;
wire n_835;
wire n_850;
wire n_690;
wire n_401;
wire n_324;
wire n_766;
wire n_743;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_862;
wire n_869;
wire n_351;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_858;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_900;
wire n_897;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_664;
wire n_678;
wire n_649;
wire n_283;

INVx1_ASAP7_75t_L g209 ( 
.A(n_171),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_14),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_198),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_202),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_69),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_131),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_184),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_154),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_78),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_23),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_201),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_122),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_16),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_13),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_12),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_14),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_41),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_178),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_87),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_185),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_17),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_40),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_128),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_68),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_16),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_117),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_90),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_164),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_199),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_134),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_104),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_193),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_13),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_123),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_186),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_196),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_45),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_65),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_82),
.Y(n_250)
);

BUFx3_ASAP7_75t_L g251 ( 
.A(n_190),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_52),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

BUFx3_ASAP7_75t_L g254 ( 
.A(n_34),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_187),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g256 ( 
.A(n_97),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_47),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_37),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_121),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_27),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_84),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_3),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_167),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_26),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_166),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_182),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_95),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_51),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_11),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_3),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_36),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_63),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_153),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_38),
.Y(n_277)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_62),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_130),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_168),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_139),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_32),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_64),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_175),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_93),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_30),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_49),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_6),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_33),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_200),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_151),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_120),
.Y(n_292)
);

INVx1_ASAP7_75t_SL g293 ( 
.A(n_25),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_102),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_188),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_125),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_21),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_212),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_243),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_275),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_228),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_231),
.Y(n_302)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_223),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_229),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_230),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_216),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_220),
.Y(n_307)
);

NOR2xp67_ASAP7_75t_L g308 ( 
.A(n_219),
.B(n_0),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_243),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_243),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_232),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_243),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_233),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_238),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_242),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_210),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

OR2x2_ASAP7_75t_L g318 ( 
.A(n_222),
.B(n_0),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_244),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g320 ( 
.A(n_225),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g323 ( 
.A(n_278),
.Y(n_323)
);

NOR2xp67_ASAP7_75t_L g324 ( 
.A(n_219),
.B(n_1),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_246),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_211),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_248),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_264),
.Y(n_328)
);

INVxp33_ASAP7_75t_SL g329 ( 
.A(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_272),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_288),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_251),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_250),
.Y(n_333)
);

INVxp33_ASAP7_75t_SL g334 ( 
.A(n_247),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_276),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_289),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_252),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_211),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_254),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_254),
.Y(n_340)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_239),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_209),
.Y(n_342)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_287),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g344 ( 
.A(n_273),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_214),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_215),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_257),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_218),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_217),
.B(n_1),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_256),
.Y(n_351)
);

BUFx2_ASAP7_75t_L g352 ( 
.A(n_239),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_240),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_259),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_262),
.Y(n_355)
);

INVxp67_ASAP7_75t_SL g356 ( 
.A(n_224),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_350),
.B(n_278),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_299),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_309),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_310),
.Y(n_361)
);

INVx3_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_298),
.B(n_287),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_318),
.B(n_240),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g365 ( 
.A(n_317),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_312),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_323),
.B(n_256),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_301),
.B(n_304),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_317),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_351),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_343),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_343),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_344),
.B(n_256),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_328),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_317),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_351),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_305),
.B(n_227),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_342),
.Y(n_378)
);

AND2x4_ASAP7_75t_L g379 ( 
.A(n_356),
.B(n_332),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_328),
.Y(n_380)
);

BUFx6f_ASAP7_75t_L g381 ( 
.A(n_316),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_311),
.B(n_234),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_345),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_348),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_338),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_322),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_300),
.B(n_245),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_349),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_330),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_339),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_340),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g393 ( 
.A(n_346),
.B(n_213),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_313),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_320),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_326),
.A2(n_245),
.B1(n_267),
.B2(n_293),
.Y(n_396)
);

OA21x2_ASAP7_75t_L g397 ( 
.A1(n_308),
.A2(n_237),
.B(n_236),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_314),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_324),
.B(n_263),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_315),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_319),
.Y(n_401)
);

BUFx6f_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g403 ( 
.A(n_352),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_327),
.Y(n_404)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_333),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_337),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_347),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_354),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_355),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_329),
.B(n_241),
.Y(n_410)
);

CKINVDCx8_ASAP7_75t_R g411 ( 
.A(n_306),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_334),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_307),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_335),
.Y(n_414)
);

INVx6_ASAP7_75t_L g415 ( 
.A(n_365),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_396),
.A2(n_353),
.B1(n_341),
.B2(n_326),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_265),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_362),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_390),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_362),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_249),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_378),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_365),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_365),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_365),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_371),
.B(n_253),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_372),
.B(n_255),
.Y(n_429)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_357),
.B(n_258),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_R g431 ( 
.A(n_398),
.B(n_336),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g432 ( 
.A(n_393),
.B(n_367),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_369),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_388),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_392),
.Y(n_435)
);

AND2x2_ASAP7_75t_L g436 ( 
.A(n_370),
.B(n_341),
.Y(n_436)
);

AOI22xp33_ASAP7_75t_L g437 ( 
.A1(n_397),
.A2(n_410),
.B1(n_357),
.B2(n_364),
.Y(n_437)
);

INVx4_ASAP7_75t_L g438 ( 
.A(n_369),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_R g439 ( 
.A(n_398),
.B(n_353),
.Y(n_439)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_394),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_381),
.Y(n_441)
);

INVx5_ASAP7_75t_L g442 ( 
.A(n_380),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g444 ( 
.A(n_376),
.B(n_268),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_381),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_397),
.A2(n_282),
.B1(n_261),
.B2(n_266),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_385),
.Y(n_447)
);

BUFx6f_ASAP7_75t_L g448 ( 
.A(n_369),
.Y(n_448)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_397),
.A2(n_260),
.B1(n_277),
.B2(n_285),
.Y(n_449)
);

OR2x2_ASAP7_75t_L g450 ( 
.A(n_364),
.B(n_286),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_358),
.B(n_269),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_411),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_381),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_410),
.A2(n_292),
.B1(n_294),
.B2(n_295),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_373),
.A2(n_283),
.B1(n_271),
.B2(n_296),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_394),
.B(n_270),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_381),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVx2_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_411),
.Y(n_460)
);

BUFx4f_ASAP7_75t_L g461 ( 
.A(n_394),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_384),
.Y(n_462)
);

INVx3_ASAP7_75t_L g463 ( 
.A(n_375),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_372),
.B(n_274),
.Y(n_464)
);

NAND2x1p5_ASAP7_75t_L g465 ( 
.A(n_394),
.B(n_279),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_379),
.B(n_280),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_384),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_375),
.Y(n_468)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_379),
.B(n_281),
.Y(n_469)
);

BUFx4f_ASAP7_75t_L g470 ( 
.A(n_400),
.Y(n_470)
);

AND2x6_ASAP7_75t_L g471 ( 
.A(n_401),
.B(n_28),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_359),
.Y(n_472)
);

CKINVDCx8_ASAP7_75t_R g473 ( 
.A(n_400),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_380),
.Y(n_474)
);

AND2x6_ASAP7_75t_L g475 ( 
.A(n_401),
.B(n_29),
.Y(n_475)
);

HB1xp67_ASAP7_75t_L g476 ( 
.A(n_395),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_406),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_360),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_361),
.Y(n_479)
);

BUFx6f_ASAP7_75t_L g480 ( 
.A(n_380),
.Y(n_480)
);

INVx2_ASAP7_75t_SL g481 ( 
.A(n_412),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx3_ASAP7_75t_L g483 ( 
.A(n_386),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_379),
.B(n_284),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_412),
.Y(n_485)
);

OR2x2_ASAP7_75t_L g486 ( 
.A(n_450),
.B(n_403),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_417),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_420),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g489 ( 
.A1(n_416),
.A2(n_387),
.B1(n_414),
.B2(n_413),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_423),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_426),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_434),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_432),
.B(n_400),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_461),
.B(n_400),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_435),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_437),
.A2(n_409),
.B1(n_405),
.B2(n_407),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_462),
.Y(n_498)
);

AND2x4_ASAP7_75t_L g499 ( 
.A(n_440),
.B(n_405),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_467),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_472),
.Y(n_501)
);

AO22x2_ASAP7_75t_L g502 ( 
.A1(n_454),
.A2(n_408),
.B1(n_409),
.B2(n_382),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_478),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_479),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_430),
.B(n_377),
.Y(n_505)
);

INVx2_ASAP7_75t_SL g506 ( 
.A(n_444),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_483),
.Y(n_507)
);

OAI221xp5_ASAP7_75t_L g508 ( 
.A1(n_454),
.A2(n_391),
.B1(n_386),
.B2(n_399),
.C(n_366),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_431),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_436),
.A2(n_399),
.B1(n_404),
.B2(n_368),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_430),
.B(n_402),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_483),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_476),
.B(n_402),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_437),
.A2(n_402),
.B1(n_291),
.B2(n_290),
.Y(n_514)
);

OR2x6_ASAP7_75t_L g515 ( 
.A(n_481),
.B(n_402),
.Y(n_515)
);

NAND2x1p5_ASAP7_75t_L g516 ( 
.A(n_461),
.B(n_391),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_466),
.A2(n_302),
.B1(n_321),
.B2(n_5),
.Y(n_517)
);

OR2x2_ASAP7_75t_SL g518 ( 
.A(n_447),
.B(n_476),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_469),
.A2(n_302),
.B1(n_321),
.B2(n_5),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

AO22x2_ASAP7_75t_L g521 ( 
.A1(n_484),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_521)
);

AO22x2_ASAP7_75t_L g522 ( 
.A1(n_456),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_421),
.Y(n_523)
);

AO22x2_ASAP7_75t_L g524 ( 
.A1(n_439),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_480),
.Y(n_525)
);

AND2x4_ASAP7_75t_L g526 ( 
.A(n_485),
.B(n_374),
.Y(n_526)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_473),
.Y(n_527)
);

AO22x2_ASAP7_75t_L g528 ( 
.A1(n_439),
.A2(n_464),
.B1(n_9),
.B2(n_10),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_422),
.Y(n_529)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_477),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_470),
.B(n_374),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_422),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_428),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_428),
.Y(n_534)
);

AO22x2_ASAP7_75t_L g535 ( 
.A1(n_464),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_429),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_429),
.Y(n_537)
);

NAND2x1p5_ASAP7_75t_L g538 ( 
.A(n_470),
.B(n_31),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_474),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_441),
.Y(n_540)
);

AND2x4_ASAP7_75t_L g541 ( 
.A(n_452),
.B(n_35),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_445),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_453),
.Y(n_543)
);

OR2x6_ASAP7_75t_L g544 ( 
.A(n_465),
.B(n_15),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_424),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_433),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_459),
.Y(n_548)
);

HB1xp67_ASAP7_75t_L g549 ( 
.A(n_460),
.Y(n_549)
);

AND2x4_ASAP7_75t_L g550 ( 
.A(n_468),
.B(n_482),
.Y(n_550)
);

BUFx3_ASAP7_75t_L g551 ( 
.A(n_465),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_418),
.B(n_15),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_482),
.Y(n_553)
);

AND2x4_ASAP7_75t_L g554 ( 
.A(n_455),
.B(n_39),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_513),
.B(n_418),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_511),
.B(n_431),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_529),
.B(n_446),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_505),
.B(n_446),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_493),
.B(n_480),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_554),
.B(n_506),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_554),
.B(n_480),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_499),
.B(n_449),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_497),
.B(n_449),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_486),
.B(n_427),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_532),
.B(n_463),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_533),
.B(n_534),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_551),
.B(n_427),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_536),
.B(n_427),
.Y(n_568)
);

AND2x4_ASAP7_75t_L g569 ( 
.A(n_503),
.B(n_471),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_537),
.B(n_443),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_514),
.B(n_443),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_518),
.B(n_463),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_494),
.B(n_443),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_495),
.B(n_448),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_487),
.B(n_448),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_488),
.B(n_448),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_490),
.B(n_458),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_491),
.B(n_458),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_509),
.B(n_458),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_492),
.B(n_442),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_496),
.B(n_442),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_501),
.B(n_442),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_504),
.B(n_541),
.Y(n_583)
);

NAND2xp33_ASAP7_75t_SL g584 ( 
.A(n_527),
.B(n_552),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_531),
.B(n_471),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_526),
.B(n_442),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_530),
.B(n_425),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_SL g588 ( 
.A(n_549),
.B(n_425),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_498),
.B(n_438),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_507),
.B(n_512),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_500),
.B(n_438),
.Y(n_591)
);

NAND2xp33_ASAP7_75t_SL g592 ( 
.A(n_540),
.B(n_471),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_SL g593 ( 
.A(n_542),
.B(n_543),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_516),
.B(n_471),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_SL g595 ( 
.A(n_520),
.B(n_471),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_502),
.B(n_475),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_502),
.B(n_475),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_523),
.B(n_475),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_545),
.B(n_550),
.Y(n_599)
);

NAND2xp33_ASAP7_75t_SL g600 ( 
.A(n_525),
.B(n_475),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_550),
.B(n_475),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_510),
.B(n_415),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_510),
.B(n_415),
.Y(n_603)
);

NAND2xp33_ASAP7_75t_SL g604 ( 
.A(n_553),
.B(n_546),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_SL g605 ( 
.A(n_538),
.B(n_415),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_539),
.B(n_42),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_547),
.B(n_43),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_548),
.B(n_44),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_515),
.B(n_46),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_SL g610 ( 
.A(n_515),
.B(n_48),
.Y(n_610)
);

OAI21x1_ASAP7_75t_L g611 ( 
.A1(n_601),
.A2(n_508),
.B(n_489),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_565),
.Y(n_612)
);

OAI21x1_ASAP7_75t_L g613 ( 
.A1(n_595),
.A2(n_598),
.B(n_594),
.Y(n_613)
);

INVxp67_ASAP7_75t_L g614 ( 
.A(n_572),
.Y(n_614)
);

NOR2xp67_ASAP7_75t_L g615 ( 
.A(n_556),
.B(n_53),
.Y(n_615)
);

OAI22xp5_ASAP7_75t_L g616 ( 
.A1(n_566),
.A2(n_521),
.B1(n_522),
.B2(n_524),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_585),
.A2(n_124),
.B(n_208),
.Y(n_617)
);

AOI221xp5_ASAP7_75t_L g618 ( 
.A1(n_560),
.A2(n_519),
.B1(n_517),
.B2(n_521),
.C(n_524),
.Y(n_618)
);

AOI21xp5_ASAP7_75t_L g619 ( 
.A1(n_563),
.A2(n_544),
.B(n_535),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_555),
.B(n_544),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_571),
.A2(n_116),
.B(n_207),
.Y(n_621)
);

OAI21x1_ASAP7_75t_L g622 ( 
.A1(n_568),
.A2(n_115),
.B(n_206),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_557),
.B(n_528),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_561),
.B(n_528),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_562),
.A2(n_535),
.B(n_519),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_569),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_599),
.Y(n_627)
);

OAI21xp5_ASAP7_75t_L g628 ( 
.A1(n_558),
.A2(n_517),
.B(n_113),
.Y(n_628)
);

AO31x2_ASAP7_75t_L g629 ( 
.A1(n_596),
.A2(n_17),
.A3(n_18),
.B(n_19),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g630 ( 
.A1(n_597),
.A2(n_205),
.B(n_112),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_564),
.B(n_559),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_570),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_573),
.A2(n_111),
.B(n_197),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_583),
.B(n_18),
.Y(n_634)
);

AND2x4_ASAP7_75t_L g635 ( 
.A(n_586),
.B(n_54),
.Y(n_635)
);

INVx1_ASAP7_75t_SL g636 ( 
.A(n_602),
.Y(n_636)
);

BUFx2_ASAP7_75t_L g637 ( 
.A(n_584),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_592),
.A2(n_114),
.B(n_195),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_569),
.B(n_55),
.Y(n_639)
);

INVxp67_ASAP7_75t_L g640 ( 
.A(n_603),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_574),
.B(n_19),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_589),
.A2(n_118),
.B(n_194),
.Y(n_642)
);

AND2x2_ASAP7_75t_L g643 ( 
.A(n_587),
.B(n_20),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_600),
.A2(n_110),
.B(n_192),
.Y(n_644)
);

A2O1A1Ixp33_ASAP7_75t_L g645 ( 
.A1(n_593),
.A2(n_590),
.B(n_569),
.C(n_588),
.Y(n_645)
);

CKINVDCx11_ASAP7_75t_R g646 ( 
.A(n_579),
.Y(n_646)
);

OAI21x1_ASAP7_75t_L g647 ( 
.A1(n_591),
.A2(n_109),
.B(n_191),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_609),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_605),
.A2(n_119),
.B(n_189),
.Y(n_649)
);

OAI21xp5_ASAP7_75t_L g650 ( 
.A1(n_606),
.A2(n_203),
.B(n_108),
.Y(n_650)
);

CKINVDCx5p33_ASAP7_75t_R g651 ( 
.A(n_610),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_567),
.B(n_22),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_SL g653 ( 
.A(n_604),
.B(n_56),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_575),
.B(n_23),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_576),
.B(n_24),
.Y(n_655)
);

AOI21xp5_ASAP7_75t_L g656 ( 
.A1(n_577),
.A2(n_127),
.B(n_57),
.Y(n_656)
);

AOI21xp5_ASAP7_75t_L g657 ( 
.A1(n_578),
.A2(n_129),
.B(n_58),
.Y(n_657)
);

OAI21xp5_ASAP7_75t_L g658 ( 
.A1(n_608),
.A2(n_132),
.B(n_59),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_612),
.B(n_580),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_627),
.Y(n_660)
);

O2A1O1Ixp33_ASAP7_75t_SL g661 ( 
.A1(n_645),
.A2(n_607),
.B(n_582),
.C(n_581),
.Y(n_661)
);

INVx3_ASAP7_75t_L g662 ( 
.A(n_626),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_628),
.A2(n_24),
.B1(n_60),
.B2(n_61),
.Y(n_663)
);

OAI22xp5_ASAP7_75t_SL g664 ( 
.A1(n_628),
.A2(n_66),
.B1(n_67),
.B2(n_70),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_626),
.Y(n_665)
);

OAI21x1_ASAP7_75t_L g666 ( 
.A1(n_613),
.A2(n_71),
.B(n_72),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_632),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_621),
.Y(n_669)
);

OAI21x1_ASAP7_75t_L g670 ( 
.A1(n_617),
.A2(n_647),
.B(n_642),
.Y(n_670)
);

OAI21x1_ASAP7_75t_L g671 ( 
.A1(n_622),
.A2(n_73),
.B(n_74),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_623),
.B(n_75),
.Y(n_672)
);

OAI21x1_ASAP7_75t_L g673 ( 
.A1(n_633),
.A2(n_76),
.B(n_77),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_646),
.Y(n_674)
);

AND2x4_ASAP7_75t_L g675 ( 
.A(n_635),
.B(n_79),
.Y(n_675)
);

OAI21x1_ASAP7_75t_L g676 ( 
.A1(n_649),
.A2(n_638),
.B(n_630),
.Y(n_676)
);

BUFx2_ASAP7_75t_L g677 ( 
.A(n_614),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_635),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_636),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_636),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_631),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_641),
.Y(n_682)
);

OAI21x1_ASAP7_75t_L g683 ( 
.A1(n_630),
.A2(n_80),
.B(n_81),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_640),
.Y(n_684)
);

OAI21x1_ASAP7_75t_L g685 ( 
.A1(n_644),
.A2(n_83),
.B(n_85),
.Y(n_685)
);

AND2x2_ASAP7_75t_SL g686 ( 
.A(n_618),
.B(n_86),
.Y(n_686)
);

OAI21x1_ASAP7_75t_L g687 ( 
.A1(n_619),
.A2(n_88),
.B(n_89),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_625),
.B(n_91),
.Y(n_688)
);

AOI21x1_ASAP7_75t_L g689 ( 
.A1(n_653),
.A2(n_92),
.B(n_94),
.Y(n_689)
);

OAI21x1_ASAP7_75t_L g690 ( 
.A1(n_656),
.A2(n_96),
.B(n_98),
.Y(n_690)
);

AO22x2_ASAP7_75t_L g691 ( 
.A1(n_616),
.A2(n_99),
.B1(n_100),
.B2(n_101),
.Y(n_691)
);

OAI21xp5_ASAP7_75t_L g692 ( 
.A1(n_615),
.A2(n_103),
.B(n_105),
.Y(n_692)
);

OAI21x1_ASAP7_75t_L g693 ( 
.A1(n_657),
.A2(n_106),
.B(n_107),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_629),
.Y(n_694)
);

NOR2xp67_ASAP7_75t_L g695 ( 
.A(n_651),
.B(n_183),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_655),
.Y(n_696)
);

OAI21x1_ASAP7_75t_L g697 ( 
.A1(n_650),
.A2(n_126),
.B(n_133),
.Y(n_697)
);

OA21x2_ASAP7_75t_L g698 ( 
.A1(n_658),
.A2(n_135),
.B(n_137),
.Y(n_698)
);

A2O1A1Ixp33_ASAP7_75t_L g699 ( 
.A1(n_620),
.A2(n_138),
.B(n_140),
.C(n_141),
.Y(n_699)
);

O2A1O1Ixp33_ASAP7_75t_L g700 ( 
.A1(n_648),
.A2(n_142),
.B(n_143),
.C(n_144),
.Y(n_700)
);

HB1xp67_ASAP7_75t_L g701 ( 
.A(n_677),
.Y(n_701)
);

OAI21x1_ASAP7_75t_L g702 ( 
.A1(n_670),
.A2(n_658),
.B(n_650),
.Y(n_702)
);

BUFx3_ASAP7_75t_L g703 ( 
.A(n_677),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_667),
.Y(n_704)
);

INVxp67_ASAP7_75t_L g705 ( 
.A(n_684),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_667),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_SL g707 ( 
.A1(n_686),
.A2(n_648),
.B1(n_616),
.B2(n_637),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_694),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_694),
.Y(n_709)
);

INVxp33_ASAP7_75t_L g710 ( 
.A(n_679),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_672),
.B(n_624),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_686),
.B(n_682),
.Y(n_712)
);

INVx2_ASAP7_75t_SL g713 ( 
.A(n_679),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_668),
.Y(n_714)
);

OAI21xp5_ASAP7_75t_L g715 ( 
.A1(n_683),
.A2(n_624),
.B(n_639),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_669),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_668),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_681),
.B(n_696),
.Y(n_718)
);

HB1xp67_ASAP7_75t_L g719 ( 
.A(n_680),
.Y(n_719)
);

OAI21x1_ASAP7_75t_L g720 ( 
.A1(n_670),
.A2(n_654),
.B(n_643),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_672),
.B(n_678),
.Y(n_721)
);

BUFx3_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

OAI21x1_ASAP7_75t_L g723 ( 
.A1(n_666),
.A2(n_652),
.B(n_634),
.Y(n_723)
);

AOI21x1_ASAP7_75t_L g724 ( 
.A1(n_676),
.A2(n_629),
.B(n_146),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_680),
.B(n_629),
.Y(n_725)
);

HB1xp67_ASAP7_75t_L g726 ( 
.A(n_660),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_687),
.Y(n_727)
);

AO21x2_ASAP7_75t_L g728 ( 
.A1(n_676),
.A2(n_145),
.B(n_147),
.Y(n_728)
);

BUFx2_ASAP7_75t_SL g729 ( 
.A(n_695),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_678),
.B(n_180),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_666),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_662),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_678),
.B(n_148),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_687),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_664),
.A2(n_149),
.B1(n_150),
.B2(n_152),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_691),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_691),
.Y(n_737)
);

HB1xp67_ASAP7_75t_L g738 ( 
.A(n_665),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_691),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_691),
.Y(n_740)
);

BUFx3_ASAP7_75t_L g741 ( 
.A(n_674),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_698),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_683),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_662),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_698),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_722),
.B(n_662),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_722),
.Y(n_747)
);

OR2x6_ASAP7_75t_L g748 ( 
.A(n_729),
.B(n_675),
.Y(n_748)
);

NAND2xp33_ASAP7_75t_R g749 ( 
.A(n_711),
.B(n_675),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_714),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_SL g751 ( 
.A(n_712),
.B(n_675),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_718),
.B(n_659),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_R g753 ( 
.A(n_722),
.B(n_741),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_714),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_R g755 ( 
.A(n_741),
.B(n_689),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_735),
.B(n_663),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_703),
.B(n_665),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_SL g758 ( 
.A(n_707),
.B(n_705),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_711),
.B(n_719),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_710),
.B(n_692),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_701),
.B(n_713),
.Y(n_761)
);

BUFx10_ASAP7_75t_L g762 ( 
.A(n_733),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_SL g763 ( 
.A(n_703),
.B(n_688),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_R g764 ( 
.A(n_741),
.B(n_689),
.Y(n_764)
);

OR2x6_ASAP7_75t_L g765 ( 
.A(n_729),
.B(n_700),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_713),
.B(n_659),
.Y(n_766)
);

NAND2xp33_ASAP7_75t_R g767 ( 
.A(n_721),
.B(n_698),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_717),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_703),
.B(n_697),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_717),
.Y(n_770)
);

BUFx3_ASAP7_75t_L g771 ( 
.A(n_744),
.Y(n_771)
);

CKINVDCx8_ASAP7_75t_R g772 ( 
.A(n_744),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_R g773 ( 
.A(n_732),
.B(n_155),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_R g774 ( 
.A(n_721),
.B(n_697),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_726),
.B(n_738),
.Y(n_775)
);

BUFx3_ASAP7_75t_L g776 ( 
.A(n_732),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_R g777 ( 
.A(n_724),
.B(n_156),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_R g778 ( 
.A(n_730),
.B(n_673),
.Y(n_778)
);

NAND2xp33_ASAP7_75t_R g779 ( 
.A(n_730),
.B(n_673),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_708),
.Y(n_780)
);

AND2x4_ASAP7_75t_L g781 ( 
.A(n_720),
.B(n_699),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_R g782 ( 
.A(n_725),
.B(n_671),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_715),
.B(n_661),
.Y(n_783)
);

NAND2xp5_ASAP7_75t_L g784 ( 
.A(n_715),
.B(n_693),
.Y(n_784)
);

HB1xp67_ASAP7_75t_L g785 ( 
.A(n_720),
.Y(n_785)
);

AND2x2_ASAP7_75t_L g786 ( 
.A(n_780),
.B(n_739),
.Y(n_786)
);

INVxp67_ASAP7_75t_L g787 ( 
.A(n_775),
.Y(n_787)
);

OR2x2_ASAP7_75t_L g788 ( 
.A(n_759),
.B(n_709),
.Y(n_788)
);

HB1xp67_ASAP7_75t_L g789 ( 
.A(n_761),
.Y(n_789)
);

AND2x2_ASAP7_75t_L g790 ( 
.A(n_750),
.B(n_739),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_754),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_768),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_770),
.Y(n_793)
);

OAI22xp5_ASAP7_75t_L g794 ( 
.A1(n_758),
.A2(n_737),
.B1(n_736),
.B2(n_740),
.Y(n_794)
);

AOI22xp33_ASAP7_75t_SL g795 ( 
.A1(n_773),
.A2(n_736),
.B1(n_740),
.B2(n_737),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_769),
.B(n_709),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_785),
.Y(n_797)
);

BUFx2_ASAP7_75t_L g798 ( 
.A(n_771),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_747),
.Y(n_799)
);

INVxp67_ASAP7_75t_L g800 ( 
.A(n_752),
.Y(n_800)
);

HB1xp67_ASAP7_75t_L g801 ( 
.A(n_772),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_766),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_783),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_776),
.Y(n_804)
);

NOR3xp33_ASAP7_75t_L g805 ( 
.A(n_756),
.B(n_723),
.C(n_743),
.Y(n_805)
);

HB1xp67_ASAP7_75t_L g806 ( 
.A(n_757),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_784),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_757),
.B(n_709),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_781),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_781),
.Y(n_810)
);

AND2x2_ASAP7_75t_L g811 ( 
.A(n_762),
.B(n_704),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_763),
.Y(n_812)
);

AOI22xp33_ASAP7_75t_SL g813 ( 
.A1(n_777),
.A2(n_762),
.B1(n_765),
.B2(n_753),
.Y(n_813)
);

HB1xp67_ASAP7_75t_L g814 ( 
.A(n_812),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_SL g815 ( 
.A1(n_805),
.A2(n_765),
.B1(n_748),
.B2(n_743),
.C(n_751),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_791),
.Y(n_816)
);

AOI22xp33_ASAP7_75t_L g817 ( 
.A1(n_813),
.A2(n_810),
.B1(n_809),
.B2(n_794),
.Y(n_817)
);

NAND2x1_ASAP7_75t_L g818 ( 
.A(n_797),
.B(n_708),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_799),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_796),
.B(n_706),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_791),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_792),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_792),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_796),
.B(n_706),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_793),
.Y(n_825)
);

NAND3xp33_ASAP7_75t_L g826 ( 
.A(n_803),
.B(n_760),
.C(n_782),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_786),
.B(n_704),
.Y(n_827)
);

INVx4_ASAP7_75t_L g828 ( 
.A(n_799),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_795),
.B(n_800),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_793),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_820),
.B(n_810),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_816),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_820),
.B(n_809),
.Y(n_833)
);

AND2x2_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_789),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_816),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_824),
.B(n_797),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_814),
.B(n_798),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_823),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_827),
.B(n_798),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_827),
.B(n_787),
.Y(n_840)
);

BUFx2_ASAP7_75t_L g841 ( 
.A(n_828),
.Y(n_841)
);

OAI22xp33_ASAP7_75t_L g842 ( 
.A1(n_841),
.A2(n_826),
.B1(n_749),
.B2(n_829),
.Y(n_842)
);

OAI221xp5_ASAP7_75t_L g843 ( 
.A1(n_837),
.A2(n_817),
.B1(n_815),
.B2(n_829),
.C(n_819),
.Y(n_843)
);

NOR4xp25_ASAP7_75t_SL g844 ( 
.A(n_832),
.B(n_767),
.C(n_779),
.D(n_778),
.Y(n_844)
);

CKINVDCx5p33_ASAP7_75t_R g845 ( 
.A(n_840),
.Y(n_845)
);

AOI22xp5_ASAP7_75t_L g846 ( 
.A1(n_840),
.A2(n_828),
.B1(n_748),
.B2(n_774),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_845),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_842),
.B(n_834),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_843),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_846),
.B(n_828),
.Y(n_850)
);

NOR2xp33_ASAP7_75t_L g851 ( 
.A(n_844),
.B(n_834),
.Y(n_851)
);

NAND2x1_ASAP7_75t_L g852 ( 
.A(n_846),
.B(n_839),
.Y(n_852)
);

INVx1_ASAP7_75t_SL g853 ( 
.A(n_847),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_850),
.B(n_849),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_848),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_851),
.A2(n_811),
.B1(n_801),
.B2(n_802),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_855),
.B(n_850),
.Y(n_857)
);

NOR2x1p5_ASAP7_75t_SL g858 ( 
.A(n_856),
.B(n_838),
.Y(n_858)
);

INVx1_ASAP7_75t_SL g859 ( 
.A(n_853),
.Y(n_859)
);

OAI21xp5_ASAP7_75t_L g860 ( 
.A1(n_854),
.A2(n_852),
.B(n_804),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_859),
.Y(n_861)
);

BUFx6f_ASAP7_75t_L g862 ( 
.A(n_857),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_860),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_858),
.Y(n_864)
);

AOI22xp5_ASAP7_75t_L g865 ( 
.A1(n_861),
.A2(n_864),
.B1(n_863),
.B2(n_862),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_862),
.B(n_831),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_861),
.B(n_839),
.Y(n_867)
);

OAI21xp5_ASAP7_75t_L g868 ( 
.A1(n_864),
.A2(n_811),
.B(n_802),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_861),
.B(n_831),
.Y(n_869)
);

NAND3xp33_ASAP7_75t_L g870 ( 
.A(n_861),
.B(n_806),
.C(n_807),
.Y(n_870)
);

NAND4xp25_ASAP7_75t_L g871 ( 
.A(n_861),
.B(n_807),
.C(n_788),
.D(n_822),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_867),
.A2(n_870),
.B1(n_865),
.B2(n_869),
.Y(n_872)
);

OAI211xp5_ASAP7_75t_SL g873 ( 
.A1(n_866),
.A2(n_835),
.B(n_821),
.C(n_830),
.Y(n_873)
);

HB1xp67_ASAP7_75t_L g874 ( 
.A(n_868),
.Y(n_874)
);

AOI221xp5_ASAP7_75t_L g875 ( 
.A1(n_871),
.A2(n_825),
.B1(n_764),
.B2(n_755),
.C(n_836),
.Y(n_875)
);

AOI211x1_ASAP7_75t_L g876 ( 
.A1(n_866),
.A2(n_836),
.B(n_833),
.C(n_786),
.Y(n_876)
);

NAND3xp33_ASAP7_75t_L g877 ( 
.A(n_865),
.B(n_818),
.C(n_823),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_867),
.A2(n_818),
.B1(n_833),
.B2(n_790),
.Y(n_878)
);

NAND2x1p5_ASAP7_75t_L g879 ( 
.A(n_865),
.B(n_746),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_879),
.B(n_808),
.Y(n_880)
);

INVxp67_ASAP7_75t_SL g881 ( 
.A(n_874),
.Y(n_881)
);

INVx2_ASAP7_75t_SL g882 ( 
.A(n_877),
.Y(n_882)
);

OAI22xp5_ASAP7_75t_L g883 ( 
.A1(n_872),
.A2(n_788),
.B1(n_790),
.B2(n_808),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_873),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_876),
.B(n_728),
.Y(n_885)
);

NOR2xp67_ASAP7_75t_L g886 ( 
.A(n_878),
.B(n_157),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_875),
.Y(n_887)
);

NOR4xp75_ASAP7_75t_L g888 ( 
.A(n_879),
.B(n_724),
.C(n_160),
.D(n_161),
.Y(n_888)
);

NAND2xp33_ASAP7_75t_SL g889 ( 
.A(n_882),
.B(n_884),
.Y(n_889)
);

NAND3xp33_ASAP7_75t_L g890 ( 
.A(n_881),
.B(n_727),
.C(n_734),
.Y(n_890)
);

NAND2xp33_ASAP7_75t_SL g891 ( 
.A(n_880),
.B(n_728),
.Y(n_891)
);

NAND2xp33_ASAP7_75t_SL g892 ( 
.A(n_887),
.B(n_883),
.Y(n_892)
);

NAND2xp33_ASAP7_75t_SL g893 ( 
.A(n_885),
.B(n_888),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_886),
.B(n_728),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_R g895 ( 
.A(n_887),
.B(n_158),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_SL g896 ( 
.A(n_882),
.B(n_728),
.Y(n_896)
);

OAI22xp5_ASAP7_75t_L g897 ( 
.A1(n_894),
.A2(n_727),
.B1(n_734),
.B2(n_731),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_889),
.Y(n_898)
);

AOI222xp33_ASAP7_75t_L g899 ( 
.A1(n_893),
.A2(n_723),
.B1(n_702),
.B2(n_685),
.C1(n_693),
.C2(n_690),
.Y(n_899)
);

NAND4xp25_ASAP7_75t_L g900 ( 
.A(n_892),
.B(n_734),
.C(n_731),
.D(n_745),
.Y(n_900)
);

HB1xp67_ASAP7_75t_L g901 ( 
.A(n_895),
.Y(n_901)
);

OAI221xp5_ASAP7_75t_L g902 ( 
.A1(n_896),
.A2(n_731),
.B1(n_745),
.B2(n_742),
.C(n_716),
.Y(n_902)
);

BUFx2_ASAP7_75t_L g903 ( 
.A(n_898),
.Y(n_903)
);

HB1xp67_ASAP7_75t_L g904 ( 
.A(n_901),
.Y(n_904)
);

AOI22xp5_ASAP7_75t_L g905 ( 
.A1(n_900),
.A2(n_891),
.B1(n_890),
.B2(n_897),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_902),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_903),
.B(n_904),
.Y(n_907)
);

XNOR2xp5_ASAP7_75t_L g908 ( 
.A(n_906),
.B(n_162),
.Y(n_908)
);

NOR2x1_ASAP7_75t_L g909 ( 
.A(n_905),
.B(n_163),
.Y(n_909)
);

AOI31xp33_ASAP7_75t_L g910 ( 
.A1(n_907),
.A2(n_899),
.A3(n_169),
.B(n_172),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_L g911 ( 
.A(n_910),
.B(n_909),
.C(n_908),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_L g912 ( 
.A1(n_911),
.A2(n_690),
.B(n_685),
.Y(n_912)
);

BUFx4_ASAP7_75t_R g913 ( 
.A(n_912),
.Y(n_913)
);

AOI221xp5_ASAP7_75t_L g914 ( 
.A1(n_913),
.A2(n_165),
.B1(n_173),
.B2(n_174),
.C(n_176),
.Y(n_914)
);

AOI211xp5_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_177),
.B(n_179),
.C(n_671),
.Y(n_915)
);


endmodule