module fake_aes_10190_n_17 (n_1, n_2, n_4, n_3, n_0, n_17);
input n_1;
input n_2;
input n_4;
input n_3;
input n_0;
output n_17;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
NOR2xp33_ASAP7_75t_L g5 ( .A(n_0), .B(n_2), .Y(n_5) );
INVx3_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
INVx2_ASAP7_75t_L g7 ( .A(n_1), .Y(n_7) );
NOR2xp33_ASAP7_75t_L g8 ( .A(n_4), .B(n_1), .Y(n_8) );
OAI21x1_ASAP7_75t_L g9 ( .A1(n_6), .A2(n_7), .B(n_5), .Y(n_9) );
OAI21x1_ASAP7_75t_SL g10 ( .A1(n_6), .A2(n_0), .B(n_1), .Y(n_10) );
AO31x2_ASAP7_75t_L g11 ( .A1(n_5), .A2(n_0), .A3(n_2), .B(n_3), .Y(n_11) );
OR2x2_ASAP7_75t_L g12 ( .A(n_9), .B(n_0), .Y(n_12) );
AOI211xp5_ASAP7_75t_L g13 ( .A1(n_9), .A2(n_8), .B(n_3), .C(n_4), .Y(n_13) );
OAI221xp5_ASAP7_75t_L g14 ( .A1(n_13), .A2(n_10), .B1(n_11), .B2(n_2), .C(n_4), .Y(n_14) );
AOI221xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_10), .B1(n_11), .B2(n_12), .C(n_13), .Y(n_15) );
HB1xp67_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
AOI21xp33_ASAP7_75t_L g17 ( .A1(n_16), .A2(n_11), .B(n_12), .Y(n_17) );
endmodule