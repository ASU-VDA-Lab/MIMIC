module real_jpeg_30346_n_19 (n_17, n_8, n_0, n_2, n_696, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_696;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_661;
wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_598;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_630;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_663;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_648;
wire n_541;
wire n_441;
wire n_657;
wire n_656;
wire n_643;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_669;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_679;
wire n_553;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_640;
wire n_666;
wire n_160;
wire n_211;
wire n_574;
wire n_627;
wire n_595;
wire n_490;
wire n_39;
wire n_685;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_680;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_678;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_578;
wire n_456;
wire n_620;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_623;
wire n_353;
wire n_668;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_605;
wire n_483;
wire n_367;
wire n_639;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_682;
wire n_317;
wire n_658;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_621;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_674;
wire n_252;
wire n_601;
wire n_655;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_611;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_634;
wire n_443;
wire n_599;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_607;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_684;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_646;
wire n_214;
wire n_671;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_673;
wire n_631;
wire n_175;
wire n_338;
wire n_653;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_650;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_652;
wire n_334;
wire n_647;
wire n_383;
wire n_593;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_612;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_614;
wire n_193;
wire n_651;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_689;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_615;
wire n_212;
wire n_284;
wire n_579;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_672;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_670;
wire n_524;
wire n_589;
wire n_25;
wire n_542;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_644;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_693;
wire n_419;
wire n_632;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_692;
wire n_49;
wire n_514;
wire n_68;
wire n_638;
wire n_497;
wire n_633;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_176;
wire n_166;
wire n_286;
wire n_596;
wire n_312;
wire n_617;
wire n_325;
wire n_316;
wire n_307;
wire n_594;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_604;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_688;
wire n_342;
wire n_120;
wire n_155;
wire n_572;
wire n_405;
wire n_412;
wire n_586;
wire n_548;
wire n_319;
wire n_664;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_637;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_613;
wire n_231;
wire n_44;
wire n_635;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_642;
wire n_106;
wire n_172;
wire n_546;
wire n_285;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_654;
wire n_377;
wire n_616;
wire n_109;
wire n_686;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_600;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_667;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_683;
wire n_159;
wire n_429;
wire n_347;
wire n_622;
wire n_183;
wire n_248;
wire n_192;
wire n_624;
wire n_537;
wire n_318;
wire n_603;
wire n_90;
wire n_336;
wire n_258;
wire n_691;
wire n_458;
wire n_677;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_628;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_675;
wire n_138;
wire n_662;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_649;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_545;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_608;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_681;
wire n_287;
wire n_400;
wire n_388;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_602;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_610;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_636;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_606;
wire n_245;
wire n_451;
wire n_626;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_597;
wire n_618;
wire n_609;
wire n_94;
wire n_645;
wire n_687;
wire n_547;
wire n_309;
wire n_294;
wire n_619;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_694;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_641;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_690;
wire n_63;
wire n_24;
wire n_92;
wire n_676;
wire n_187;
wire n_436;
wire n_629;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_659;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_660;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_625;
wire n_591;
wire n_96;
wire n_665;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_0),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_0),
.Y(n_285)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_0),
.Y(n_380)
);

BUFx12f_ASAP7_75t_L g523 ( 
.A(n_0),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_1),
.A2(n_122),
.B1(n_128),
.B2(n_129),
.Y(n_121)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g287 ( 
.A1(n_1),
.A2(n_128),
.B1(n_288),
.B2(n_292),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_1),
.A2(n_128),
.B1(n_312),
.B2(n_316),
.Y(n_311)
);

OAI22x1_ASAP7_75t_L g368 ( 
.A1(n_1),
.A2(n_128),
.B1(n_369),
.B2(n_374),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_2),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_3),
.A2(n_64),
.B1(n_65),
.B2(n_70),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_3),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_3),
.A2(n_64),
.B1(n_110),
.B2(n_114),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_3),
.A2(n_64),
.B1(n_172),
.B2(n_178),
.Y(n_171)
);

AO22x1_ASAP7_75t_SL g241 ( 
.A1(n_3),
.A2(n_64),
.B1(n_242),
.B2(n_244),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_L g297 ( 
.A1(n_4),
.A2(n_298),
.B1(n_299),
.B2(n_300),
.Y(n_297)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_4),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_4),
.A2(n_298),
.B1(n_398),
.B2(n_400),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_SL g552 ( 
.A1(n_4),
.A2(n_298),
.B1(n_553),
.B2(n_555),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_4),
.A2(n_298),
.B1(n_574),
.B2(n_577),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_5),
.B(n_131),
.Y(n_361)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_5),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g468 ( 
.A(n_5),
.B(n_74),
.Y(n_468)
);

OAI32xp33_ASAP7_75t_L g534 ( 
.A1(n_5),
.A2(n_535),
.A3(n_537),
.B1(n_542),
.B2(n_546),
.Y(n_534)
);

OAI21xp33_ASAP7_75t_L g610 ( 
.A1(n_5),
.A2(n_282),
.B(n_611),
.Y(n_610)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_5),
.A2(n_447),
.B1(n_661),
.B2(n_665),
.Y(n_660)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_201),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_6),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_6),
.A2(n_205),
.B1(n_306),
.B2(n_309),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_6),
.A2(n_205),
.B1(n_269),
.B2(n_418),
.Y(n_417)
);

AO22x1_ASAP7_75t_L g471 ( 
.A1(n_6),
.A2(n_205),
.B1(n_472),
.B2(n_475),
.Y(n_471)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_7),
.A2(n_389),
.B1(n_390),
.B2(n_392),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_7),
.A2(n_389),
.B1(n_451),
.B2(n_454),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_SL g566 ( 
.A1(n_7),
.A2(n_389),
.B1(n_567),
.B2(n_569),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_7),
.A2(n_389),
.B1(n_639),
.B2(n_642),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g689 ( 
.A(n_8),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_9),
.Y(n_62)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_10),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_10),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_11),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_11),
.Y(n_90)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_11),
.Y(n_240)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_11),
.Y(n_531)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_12),
.A2(n_53),
.B1(n_54),
.B2(n_59),
.Y(n_52)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_12),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_12),
.A2(n_53),
.B1(n_140),
.B2(n_145),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_12),
.A2(n_53),
.B1(n_260),
.B2(n_261),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g275 ( 
.A1(n_12),
.A2(n_53),
.B1(n_276),
.B2(n_279),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_13),
.A2(n_251),
.B1(n_254),
.B2(n_255),
.Y(n_250)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_13),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_13),
.A2(n_254),
.B1(n_407),
.B2(n_408),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_13),
.A2(n_254),
.B1(n_438),
.B2(n_440),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_L g526 ( 
.A1(n_13),
.A2(n_254),
.B1(n_527),
.B2(n_532),
.Y(n_526)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_14),
.Y(n_86)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_14),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_14),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_15),
.A2(n_59),
.B1(n_134),
.B2(n_135),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_15),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_15),
.A2(n_134),
.B1(n_216),
.B2(n_218),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_15),
.A2(n_134),
.B1(n_266),
.B2(n_269),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g381 ( 
.A1(n_15),
.A2(n_134),
.B1(n_382),
.B2(n_384),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_16),
.B(n_689),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_16),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g98 ( 
.A(n_17),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_17),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_17),
.Y(n_113)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_17),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_18),
.Y(n_144)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_18),
.Y(n_177)
);

OAI311xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_189),
.A3(n_688),
.B1(n_690),
.C1(n_693),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g694 ( 
.A(n_21),
.B(n_688),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_188),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_75),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_24),
.B(n_75),
.Y(n_188)
);

AOI22x1_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_52),
.B1(n_63),
.B2(n_73),
.Y(n_24)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_25),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_25),
.A2(n_52),
.B1(n_73),
.B2(n_186),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_25),
.A2(n_73),
.B1(n_121),
.B2(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2x1_ASAP7_75t_L g249 ( 
.A(n_26),
.B(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_26),
.B(n_297),
.Y(n_296)
);

AO22x1_ASAP7_75t_L g431 ( 
.A1(n_26),
.A2(n_74),
.B1(n_297),
.B2(n_388),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_26),
.B(n_445),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_42),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_34),
.B2(n_38),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_30),
.Y(n_127)
);

INVx3_ASAP7_75t_L g209 ( 
.A(n_30),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g256 ( 
.A(n_30),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_30),
.Y(n_360)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx2_ASAP7_75t_L g356 ( 
.A(n_32),
.Y(n_356)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_35),
.Y(n_299)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_37),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_SL g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_41),
.Y(n_366)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

AOI22x1_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_45),
.Y(n_217)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g363 ( 
.A(n_50),
.Y(n_363)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_51),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_51),
.Y(n_308)
);

INVx1_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_62),
.Y(n_253)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_62),
.Y(n_394)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_69),
.Y(n_131)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_71),
.Y(n_135)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_73),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_74),
.B(n_200),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_74),
.B(n_250),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_74),
.B(n_388),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_185),
.C(n_187),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_76),
.B(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_SL g76 ( 
.A(n_77),
.B(n_119),
.C(n_137),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_77),
.A2(n_78),
.B1(n_137),
.B2(n_138),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_77),
.A2(n_78),
.B1(n_213),
.B2(n_214),
.Y(n_331)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp33_ASAP7_75t_R g212 ( 
.A(n_78),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_78),
.B(n_213),
.Y(n_221)
);

OA21x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_93),
.B(n_109),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_79),
.A2(n_93),
.B1(n_109),
.B2(n_323),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g436 ( 
.A1(n_79),
.A2(n_93),
.B1(n_437),
.B2(n_442),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_79),
.B(n_437),
.Y(n_556)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_79),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g94 ( 
.A(n_80),
.B(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_80),
.Y(n_264)
);

OAI22x1_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_84),
.B1(n_87),
.B2(n_91),
.Y(n_80)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_81),
.Y(n_576)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_83),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_83),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g568 ( 
.A(n_83),
.Y(n_568)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_86),
.Y(n_92)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_89),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_89),
.Y(n_383)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_90),
.Y(n_598)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_93),
.B(n_603),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_93),
.B(n_437),
.Y(n_643)
);

AOI22xp5_ASAP7_75t_L g655 ( 
.A1(n_93),
.A2(n_656),
.B1(n_657),
.B2(n_658),
.Y(n_655)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_94),
.A2(n_259),
.B1(n_264),
.B2(n_265),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_94),
.A2(n_264),
.B1(n_265),
.B2(n_287),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_94),
.A2(n_264),
.B1(n_287),
.B2(n_417),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_94),
.A2(n_552),
.B(n_556),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_99),
.B1(n_103),
.B2(n_106),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_SL g97 ( 
.A(n_98),
.Y(n_97)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_98),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_98),
.Y(n_291)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_98),
.Y(n_421)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx6_ASAP7_75t_L g593 ( 
.A(n_101),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_108),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_108),
.Y(n_641)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g260 ( 
.A(n_112),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_112),
.Y(n_292)
);

INVx2_ASAP7_75t_SL g439 ( 
.A(n_112),
.Y(n_439)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_113),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_113),
.Y(n_270)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

HB1xp67_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_117),
.Y(n_554)
);

BUFx5_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_118),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_119),
.B(n_196),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_132),
.B1(n_133),
.B2(n_136),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

HB1xp67_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_127),
.Y(n_301)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_133),
.Y(n_186)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_148),
.B1(n_171),
.B2(n_182),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_139),
.A2(n_150),
.B1(n_182),
.B2(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_141),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_143),
.Y(n_147)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_143),
.Y(n_163)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_143),
.Y(n_410)
);

BUFx6f_ASAP7_75t_L g453 ( 
.A(n_143),
.Y(n_453)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_143),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g181 ( 
.A(n_144),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g354 ( 
.A(n_144),
.Y(n_354)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_144),
.Y(n_404)
);

BUFx6f_ASAP7_75t_L g664 ( 
.A(n_144),
.Y(n_664)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

OA21x2_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_171),
.B(n_182),
.Y(n_187)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_149),
.A2(n_397),
.B(n_405),
.Y(n_396)
);

OAI21x1_ASAP7_75t_L g426 ( 
.A1(n_149),
.A2(n_427),
.B(n_428),
.Y(n_426)
);

OA21x2_ASAP7_75t_L g659 ( 
.A1(n_149),
.A2(n_405),
.B(n_660),
.Y(n_659)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_150),
.A2(n_184),
.B1(n_305),
.B2(n_311),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_150),
.A2(n_182),
.B1(n_215),
.B2(n_311),
.Y(n_324)
);

AOI22x1_ASAP7_75t_L g449 ( 
.A1(n_150),
.A2(n_182),
.B1(n_450),
.B2(n_455),
.Y(n_449)
);

NAND2xp33_ASAP7_75t_SL g467 ( 
.A(n_150),
.B(n_406),
.Y(n_467)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_162),
.Y(n_150)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_151),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_153),
.Y(n_549)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_154),
.Y(n_607)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_157),
.Y(n_169)
);

INVx5_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_161),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_167),
.B2(n_170),
.Y(n_162)
);

INVx2_ASAP7_75t_SL g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g545 ( 
.A(n_166),
.Y(n_545)
);

INVx1_ASAP7_75t_SL g167 ( 
.A(n_168),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_174),
.B(n_543),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_176),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_177),
.Y(n_219)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_177),
.Y(n_315)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_180),
.Y(n_407)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g428 ( 
.A(n_183),
.B(n_429),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g465 ( 
.A1(n_183),
.A2(n_466),
.B(n_467),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_183),
.B(n_447),
.Y(n_636)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_184),
.B(n_406),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_185),
.B(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_189),
.B(n_694),
.Y(n_693)
);

OAI21x1_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_222),
.B(n_686),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g687 ( 
.A(n_192),
.B(n_194),
.Y(n_687)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.C(n_210),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_195),
.A2(n_335),
.B1(n_337),
.B2(n_338),
.Y(n_334)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_195),
.Y(n_337)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_197),
.A2(n_198),
.B1(n_211),
.B2(n_221),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

OA21x2_ASAP7_75t_SL g210 ( 
.A1(n_198),
.A2(n_211),
.B(n_220),
.Y(n_210)
);

OAI21xp33_ASAP7_75t_L g335 ( 
.A1(n_198),
.A2(n_212),
.B(n_336),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_198),
.B(n_221),
.Y(n_336)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_199),
.B(n_331),
.Y(n_330)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_219),
.Y(n_310)
);

INVx4_ASAP7_75t_L g319 ( 
.A(n_219),
.Y(n_319)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_219),
.Y(n_399)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21x1_ASAP7_75t_L g222 ( 
.A1(n_223),
.A2(n_342),
.B(n_680),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_333),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_326),
.Y(n_225)
);

NOR2xp67_ASAP7_75t_L g683 ( 
.A(n_226),
.B(n_326),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_271),
.C(n_320),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_227),
.B(n_320),
.Y(n_485)
);

XNOR2x1_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_257),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_247),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_229),
.A2(n_257),
.B1(n_328),
.B2(n_696),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_229),
.A2(n_230),
.B1(n_258),
.B2(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_230),
.B(n_258),
.Y(n_257)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B(n_241),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_234),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g616 ( 
.A(n_234),
.Y(n_616)
);

HB1xp67_ASAP7_75t_L g628 ( 
.A(n_234),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g653 ( 
.A(n_234),
.Y(n_653)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_235),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_235),
.A2(n_368),
.B1(n_377),
.B2(n_381),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_235),
.B(n_526),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g564 ( 
.A1(n_235),
.A2(n_477),
.B1(n_565),
.B2(n_572),
.Y(n_564)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_238),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g422 ( 
.A1(n_236),
.A2(n_275),
.B1(n_282),
.B2(n_423),
.Y(n_422)
);

INVx3_ASAP7_75t_SL g477 ( 
.A(n_236),
.Y(n_477)
);

INVx8_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_240),
.Y(n_246)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_240),
.Y(n_281)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_240),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g588 ( 
.A(n_240),
.Y(n_588)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_241),
.Y(n_283)
);

INVx4_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_244),
.Y(n_384)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx12f_ASAP7_75t_L g571 ( 
.A(n_246),
.Y(n_571)
);

HB1xp67_ASAP7_75t_L g328 ( 
.A(n_247),
.Y(n_328)
);

NAND2x1_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_249),
.B(n_387),
.Y(n_386)
);

INVx3_ASAP7_75t_SL g251 ( 
.A(n_252),
.Y(n_251)
);

INVx4_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx3_ASAP7_75t_L g446 ( 
.A(n_255),
.Y(n_446)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g491 ( 
.A(n_258),
.Y(n_491)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_259),
.Y(n_323)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g600 ( 
.A(n_262),
.Y(n_600)
);

INVx4_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_263),
.Y(n_441)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_264),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_266),
.Y(n_642)
);

INVx4_ASAP7_75t_SL g266 ( 
.A(n_267),
.Y(n_266)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_272),
.B(n_485),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_293),
.C(n_302),
.Y(n_272)
);

XNOR2x1_ASAP7_75t_L g494 ( 
.A(n_273),
.B(n_495),
.Y(n_494)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_286),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_274),
.B(n_286),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_275),
.A2(n_282),
.B1(n_283),
.B2(n_284),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g617 ( 
.A(n_276),
.B(n_618),
.Y(n_617)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g474 ( 
.A(n_281),
.Y(n_474)
);

OAI21xp5_ASAP7_75t_L g470 ( 
.A1(n_282),
.A2(n_471),
.B(n_476),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g634 ( 
.A1(n_282),
.A2(n_573),
.B(n_611),
.Y(n_634)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_291),
.Y(n_555)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g495 ( 
.A1(n_294),
.A2(n_303),
.B1(n_304),
.B2(n_496),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_294),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

AND2x2_ASAP7_75t_L g443 ( 
.A(n_295),
.B(n_444),
.Y(n_443)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

HB1xp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_305),
.Y(n_429)
);

INVx3_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

INVx8_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

NAND2x1_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_321),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g325 ( 
.A(n_322),
.B(n_324),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g326 ( 
.A(n_327),
.B(n_329),
.Y(n_326)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_327),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_330),
.B(n_332),
.Y(n_329)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_332),
.B(n_340),
.C(n_341),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_333),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_334),
.B(n_339),
.Y(n_685)
);

NAND2x1_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_507),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_344),
.A2(n_481),
.B(n_503),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_432),
.C(n_458),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_346),
.A2(n_510),
.B(n_511),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_411),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_348),
.B(n_413),
.C(n_502),
.Y(n_501)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_385),
.C(n_395),
.Y(n_348)
);

XNOR2x1_ASAP7_75t_L g433 ( 
.A(n_349),
.B(n_434),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_367),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_350),
.B(n_367),
.Y(n_462)
);

AOI32xp33_ASAP7_75t_L g350 ( 
.A1(n_351),
.A2(n_355),
.A3(n_357),
.B1(n_361),
.B2(n_362),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx4_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx11_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_SL g391 ( 
.A(n_360),
.Y(n_391)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_361),
.Y(n_448)
);

NAND2xp33_ASAP7_75t_R g362 ( 
.A(n_363),
.B(n_364),
.Y(n_362)
);

INVx3_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_368),
.B(n_477),
.Y(n_476)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx2_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

BUFx6f_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_379),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_380),
.Y(n_622)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_381),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g434 ( 
.A1(n_385),
.A2(n_386),
.B1(n_395),
.B2(n_396),
.Y(n_434)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_397),
.Y(n_455)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_399),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_406),
.Y(n_427)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_412),
.B(n_414),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_413),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g502 ( 
.A(n_414),
.Y(n_502)
);

XNOR2x1_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_424),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g488 ( 
.A(n_415),
.B(n_431),
.C(n_489),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_422),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_416),
.B(n_422),
.Y(n_457)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_417),
.Y(n_442)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

BUFx4f_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

AOI22x1_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_426),
.B1(n_430),
.B2(n_431),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_426),
.Y(n_489)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_432),
.Y(n_510)
);

MAJx2_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_456),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_433),
.B(n_479),
.Y(n_478)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_435),
.A2(n_456),
.B1(n_457),
.B2(n_480),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_435),
.Y(n_480)
);

MAJx2_ASAP7_75t_L g435 ( 
.A(n_436),
.B(n_443),
.C(n_449),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_436),
.B(n_449),
.Y(n_461)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_441),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_446),
.A2(n_447),
.B(n_448),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_447),
.B(n_547),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_447),
.B(n_540),
.Y(n_585)
);

OAI21xp33_ASAP7_75t_L g603 ( 
.A1(n_447),
.A2(n_585),
.B(n_604),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g618 ( 
.A(n_447),
.B(n_619),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_SL g624 ( 
.A(n_447),
.B(n_625),
.Y(n_624)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_450),
.Y(n_466)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx4_ASAP7_75t_L g454 ( 
.A(n_453),
.Y(n_454)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_457),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_478),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_459),
.B(n_478),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_462),
.C(n_463),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_460),
.B(n_515),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_462),
.A2(n_463),
.B1(n_464),
.B2(n_516),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_468),
.C(n_469),
.Y(n_464)
);

XOR2xp5_ASAP7_75t_L g558 ( 
.A(n_465),
.B(n_559),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_468),
.B(n_470),
.Y(n_559)
);

HB1xp67_ASAP7_75t_L g469 ( 
.A(n_470),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_R g520 ( 
.A(n_471),
.B(n_521),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g651 ( 
.A1(n_471),
.A2(n_525),
.B(n_652),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_474),
.Y(n_475)
);

INVxp67_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_509),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_L g482 ( 
.A1(n_483),
.A2(n_486),
.B(n_497),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_483),
.B(n_486),
.Y(n_506)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_484),
.B(n_487),
.Y(n_505)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_488),
.B(n_490),
.C(n_492),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_488),
.B(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_490),
.Y(n_500)
);

INVxp67_ASAP7_75t_SL g492 ( 
.A(n_493),
.Y(n_492)
);

INVxp67_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g499 ( 
.A(n_494),
.B(n_500),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_498),
.B(n_501),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_498),
.B(n_501),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_504),
.A2(n_505),
.B(n_506),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_508),
.B(n_512),
.Y(n_507)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_560),
.B(n_678),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_514),
.B(n_517),
.Y(n_513)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_514),
.Y(n_679)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_518),
.B(n_679),
.Y(n_678)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_550),
.C(n_557),
.Y(n_518)
);

OAI22xp5_ASAP7_75t_L g672 ( 
.A1(n_519),
.A2(n_550),
.B1(n_551),
.B2(n_673),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_519),
.Y(n_673)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_520),
.A2(n_524),
.B(n_534),
.Y(n_519)
);

BUFx3_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx8_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVxp67_ASAP7_75t_SL g524 ( 
.A(n_525),
.Y(n_524)
);

OAI21xp33_ASAP7_75t_SL g626 ( 
.A1(n_525),
.A2(n_566),
.B(n_627),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_526),
.B(n_612),
.Y(n_611)
);

INVx3_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

BUFx3_ASAP7_75t_L g528 ( 
.A(n_529),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_530),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);

INVx2_ASAP7_75t_L g581 ( 
.A(n_531),
.Y(n_581)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g650 ( 
.A(n_534),
.B(n_651),
.Y(n_650)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_536),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_539),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

INVx4_ASAP7_75t_L g540 ( 
.A(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_544),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_545),
.Y(n_544)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_548),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_551),
.Y(n_550)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_552),
.Y(n_658)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_556),
.B(n_602),
.Y(n_601)
);

HB1xp67_ASAP7_75t_L g557 ( 
.A(n_558),
.Y(n_557)
);

XNOR2xp5_ASAP7_75t_L g671 ( 
.A(n_558),
.B(n_672),
.Y(n_671)
);

OAI21xp5_ASAP7_75t_L g560 ( 
.A1(n_561),
.A2(n_669),
.B(n_677),
.Y(n_560)
);

O2A1O1Ixp5_ASAP7_75t_L g561 ( 
.A1(n_562),
.A2(n_631),
.B(n_644),
.C(n_645),
.Y(n_561)
);

AOI21x1_ASAP7_75t_L g562 ( 
.A1(n_563),
.A2(n_608),
.B(n_630),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_564),
.B(n_582),
.Y(n_563)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_564),
.B(n_582),
.Y(n_630)
);

INVxp67_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g567 ( 
.A(n_568),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g569 ( 
.A(n_570),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_571),
.Y(n_570)
);

INVxp33_ASAP7_75t_SL g572 ( 
.A(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_575),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_576),
.Y(n_575)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_578),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_579),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_580),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_581),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_601),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_583),
.B(n_601),
.Y(n_632)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_584),
.A2(n_586),
.B1(n_594),
.B2(n_599),
.Y(n_583)
);

INVxp67_ASAP7_75t_SL g584 ( 
.A(n_585),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_587),
.B(n_589),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_588),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g599 ( 
.A(n_589),
.B(n_600),
.Y(n_599)
);

BUFx2_ASAP7_75t_L g589 ( 
.A(n_590),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_591),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_592),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_593),
.Y(n_592)
);

INVx1_ASAP7_75t_SL g594 ( 
.A(n_595),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_596),
.Y(n_595)
);

HB1xp67_ASAP7_75t_L g596 ( 
.A(n_597),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_598),
.Y(n_597)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_605),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_606),
.Y(n_605)
);

INVx4_ASAP7_75t_L g606 ( 
.A(n_607),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_L g608 ( 
.A1(n_609),
.A2(n_623),
.B(n_629),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_610),
.B(n_617),
.Y(n_609)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_613),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_614),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_615),
.Y(n_614)
);

BUFx2_ASAP7_75t_L g615 ( 
.A(n_616),
.Y(n_615)
);

INVx4_ASAP7_75t_L g619 ( 
.A(n_620),
.Y(n_619)
);

INVx4_ASAP7_75t_L g620 ( 
.A(n_621),
.Y(n_620)
);

INVx2_ASAP7_75t_SL g621 ( 
.A(n_622),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g623 ( 
.A(n_624),
.B(n_626),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_624),
.B(n_626),
.Y(n_629)
);

OAI21xp5_ASAP7_75t_L g637 ( 
.A1(n_625),
.A2(n_638),
.B(n_643),
.Y(n_637)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_628),
.Y(n_627)
);

NOR2xp67_ASAP7_75t_L g631 ( 
.A(n_632),
.B(n_633),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_632),
.B(n_633),
.Y(n_644)
);

XNOR2xp5_ASAP7_75t_SL g633 ( 
.A(n_634),
.B(n_635),
.Y(n_633)
);

MAJIxp5_ASAP7_75t_L g646 ( 
.A(n_634),
.B(n_647),
.C(n_648),
.Y(n_646)
);

XNOR2xp5_ASAP7_75t_L g635 ( 
.A(n_636),
.B(n_637),
.Y(n_635)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_636),
.Y(n_648)
);

HB1xp67_ASAP7_75t_L g647 ( 
.A(n_637),
.Y(n_647)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_638),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g639 ( 
.A(n_640),
.Y(n_639)
);

BUFx6f_ASAP7_75t_L g640 ( 
.A(n_641),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g645 ( 
.A(n_646),
.B(n_649),
.Y(n_645)
);

OR2x2_ASAP7_75t_L g676 ( 
.A(n_646),
.B(n_649),
.Y(n_676)
);

XOR2xp5_ASAP7_75t_L g649 ( 
.A(n_650),
.B(n_654),
.Y(n_649)
);

INVxp67_ASAP7_75t_L g675 ( 
.A(n_650),
.Y(n_675)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_653),
.Y(n_652)
);

XNOR2xp5_ASAP7_75t_L g654 ( 
.A(n_655),
.B(n_659),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_655),
.B(n_659),
.C(n_675),
.Y(n_674)
);

INVx1_ASAP7_75t_L g661 ( 
.A(n_662),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_663),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_664),
.Y(n_663)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_666),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_667),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_668),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g669 ( 
.A(n_670),
.B(n_676),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_671),
.B(n_674),
.Y(n_670)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_671),
.B(n_674),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_L g680 ( 
.A1(n_681),
.A2(n_682),
.B(n_684),
.Y(n_680)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_683),
.Y(n_682)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_685),
.Y(n_684)
);

HB1xp67_ASAP7_75t_L g686 ( 
.A(n_687),
.Y(n_686)
);

INVxp33_ASAP7_75t_SL g692 ( 
.A(n_688),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_691),
.B(n_692),
.Y(n_690)
);


endmodule