module fake_jpeg_12256_n_66 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_66);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_66;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_15;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_7),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx5_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_19),
.B(n_23),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_16),
.A2(n_14),
.B1(n_15),
.B2(n_9),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g27 ( 
.A1(n_20),
.A2(n_21),
.B1(n_14),
.B2(n_15),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_16),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_17),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_22),
.B(n_9),
.Y(n_29)
);

INVx3_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_19),
.B(n_12),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_25),
.B(n_28),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_19),
.B(n_12),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_10),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_27),
.A2(n_18),
.B1(n_23),
.B2(n_10),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_30),
.A2(n_35),
.B(n_27),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_24),
.A2(n_20),
.B1(n_21),
.B2(n_18),
.Y(n_32)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_24),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_22),
.Y(n_37)
);

MAJx2_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_27),
.C(n_13),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_42),
.B(n_43),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_11),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_39),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_31),
.B(n_11),
.Y(n_40)
);

BUFx24_ASAP7_75t_SL g47 ( 
.A(n_40),
.Y(n_47)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g45 ( 
.A1(n_43),
.A2(n_33),
.B1(n_18),
.B2(n_26),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_45),
.A2(n_26),
.B1(n_17),
.B2(n_3),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_SL g46 ( 
.A(n_41),
.B(n_13),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_49),
.C(n_23),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_22),
.C(n_23),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_48),
.B(n_44),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_53),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_51),
.A2(n_17),
.B(n_1),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_47),
.A2(n_13),
.B(n_4),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_52),
.A2(n_50),
.B(n_6),
.Y(n_55)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

OA21x2_ASAP7_75t_L g57 ( 
.A1(n_54),
.A2(n_1),
.B(n_3),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_55),
.B(n_57),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_6),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_60),
.B(n_61),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_56),
.B(n_8),
.Y(n_61)
);

NAND2x1_ASAP7_75t_L g62 ( 
.A(n_59),
.B(n_60),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_62),
.A2(n_63),
.B(n_8),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_64),
.B(n_62),
.Y(n_65)
);

BUFx24_ASAP7_75t_SL g66 ( 
.A(n_65),
.Y(n_66)
);


endmodule