module real_jpeg_31085_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_288;
wire n_83;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_0),
.Y(n_210)
);

BUFx12f_ASAP7_75t_L g214 ( 
.A(n_0),
.Y(n_214)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_0),
.Y(n_254)
);

BUFx3_ASAP7_75t_L g327 ( 
.A(n_0),
.Y(n_327)
);

CKINVDCx11_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_1),
.B(n_20),
.Y(n_19)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_1),
.Y(n_529)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22x1_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_63),
.B1(n_107),
.B2(n_112),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_63),
.B1(n_135),
.B2(n_139),
.Y(n_134)
);

AO22x1_ASAP7_75t_SL g218 ( 
.A1(n_2),
.A2(n_63),
.B1(n_86),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_2),
.B(n_119),
.Y(n_436)
);

NAND2xp33_ASAP7_75t_SL g456 ( 
.A(n_2),
.B(n_451),
.Y(n_456)
);

OAI32xp33_ASAP7_75t_L g471 ( 
.A1(n_2),
.A2(n_472),
.A3(n_474),
.B1(n_477),
.B2(n_481),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_3),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_3),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_4),
.Y(n_126)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_4),
.Y(n_132)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_5),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_5),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_5),
.Y(n_219)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_6),
.A2(n_238),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_6),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_6),
.A2(n_240),
.B1(n_351),
.B2(n_353),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_6),
.A2(n_240),
.B1(n_429),
.B2(n_432),
.Y(n_428)
);

OAI22xp33_ASAP7_75t_SL g440 ( 
.A1(n_6),
.A2(n_240),
.B1(n_441),
.B2(n_443),
.Y(n_440)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_7),
.A2(n_15),
.B(n_18),
.Y(n_14)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_8),
.A2(n_73),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_8),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_8),
.A2(n_75),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_8),
.A2(n_75),
.B1(n_112),
.B2(n_226),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_8),
.A2(n_75),
.B1(n_308),
.B2(n_311),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_9),
.Y(n_115)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_9),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_11),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.Y(n_27)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

AO22x2_ASAP7_75t_SL g144 ( 
.A1(n_11),
.A2(n_31),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_11),
.A2(n_31),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_11),
.A2(n_31),
.B1(n_257),
.B2(n_260),
.Y(n_256)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_12),
.Y(n_85)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_12),
.Y(n_92)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_12),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_13),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_13),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_13),
.Y(n_160)
);

BUFx12f_ASAP7_75t_SL g15 ( 
.A(n_16),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22x1_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_288),
.B1(n_529),
.B2(n_530),
.Y(n_18)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_170),
.Y(n_20)
);

AOI21xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_67),
.B(n_68),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_22),
.B(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_23),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_23),
.B(n_231),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_55),
.Y(n_23)
);

INVxp33_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OA21x2_ASAP7_75t_SL g71 ( 
.A1(n_25),
.A2(n_58),
.B(n_72),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_26),
.B(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_37),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_27),
.B(n_57),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_37),
.A2(n_38),
.B(n_59),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_37),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_37),
.B(n_59),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_37),
.B(n_237),
.Y(n_236)
);

NOR2x1_ASAP7_75t_L g37 ( 
.A(n_38),
.B(n_47),
.Y(n_37)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

NAND2xp33_ASAP7_75t_L g304 ( 
.A(n_38),
.B(n_237),
.Y(n_304)
);

AO22x2_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_43),
.B2(n_44),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_40),
.Y(n_334)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_42),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g454 ( 
.A(n_42),
.Y(n_454)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_46),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_49),
.B1(n_51),
.B2(n_52),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_54),
.Y(n_343)
);

INVxp33_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_56),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp67_ASAP7_75t_SL g396 ( 
.A(n_58),
.B(n_63),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_63),
.B(n_64),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_62),
.Y(n_239)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_62),
.Y(n_243)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_62),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_63),
.B(n_65),
.Y(n_64)
);

AOI32xp33_ASAP7_75t_L g449 ( 
.A1(n_63),
.A2(n_450),
.A3(n_452),
.B1(n_455),
.B2(n_456),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_63),
.B(n_478),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_63),
.B(n_81),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g506 ( 
.A(n_63),
.B(n_206),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_64),
.Y(n_346)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_67),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_67),
.B(n_205),
.Y(n_265)
);

INVxp67_ASAP7_75t_SL g287 ( 
.A(n_69),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_162),
.C(n_166),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_70),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_78),
.C(n_116),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_71),
.B(n_271),
.Y(n_270)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_72),
.A2(n_163),
.B(n_165),
.Y(n_162)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

XNOR2x1_ASAP7_75t_L g177 ( 
.A(n_78),
.B(n_178),
.Y(n_177)
);

OAI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_78),
.A2(n_79),
.B1(n_116),
.B2(n_272),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_78),
.B(n_178),
.C(n_188),
.Y(n_275)
);

MAJx2_ASAP7_75t_L g379 ( 
.A(n_78),
.B(n_380),
.C(n_382),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_78),
.A2(n_79),
.B1(n_380),
.B2(n_392),
.Y(n_391)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21x1_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_96),
.B(n_106),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_80),
.B(n_106),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_80),
.B(n_225),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_80),
.B(n_428),
.Y(n_459)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_81),
.B(n_97),
.Y(n_96)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_82),
.B(n_197),
.Y(n_230)
);

OAI22x1_ASAP7_75t_L g82 ( 
.A1(n_83),
.A2(n_86),
.B1(n_89),
.B2(n_93),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_88),
.Y(n_216)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_95),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_95),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_96),
.B(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_96),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_96),
.B(n_106),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_96),
.B(n_428),
.Y(n_427)
);

OAI22xp33_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_101),
.B1(n_103),
.B2(n_104),
.Y(n_97)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_100),
.Y(n_105)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_111),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_113),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_115),
.Y(n_228)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_116),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_142),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_118),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_133),
.Y(n_118)
);

INVx1_ASAP7_75t_SL g169 ( 
.A(n_119),
.Y(n_169)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_119),
.B(n_144),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_119),
.A2(n_142),
.B(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_119),
.B(n_350),
.Y(n_381)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AO21x2_ASAP7_75t_L g150 ( 
.A1(n_120),
.A2(n_151),
.B(n_157),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_124),
.B1(n_127),
.B2(n_130),
.Y(n_120)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_121),
.Y(n_202)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_122),
.Y(n_483)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_123),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_123),
.Y(n_200)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_125),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_134),
.A2(n_150),
.B(n_169),
.Y(n_168)
);

NOR2x1_ASAP7_75t_L g246 ( 
.A(n_134),
.B(n_150),
.Y(n_246)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_138),
.Y(n_147)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx8_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_143),
.B(n_381),
.Y(n_380)
);

NAND2x1_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g345 ( 
.A(n_146),
.Y(n_345)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_147),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_149),
.B(n_350),
.Y(n_349)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g331 ( 
.A(n_153),
.Y(n_331)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp33_ASAP7_75t_L g455 ( 
.A(n_157),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_159),
.Y(n_352)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_162),
.A2(n_166),
.B1(n_167),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_162),
.Y(n_280)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

AND2x2_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_189),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_165),
.B(n_236),
.Y(n_356)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_167),
.B(n_366),
.C(n_367),
.Y(n_365)
);

HB1xp67_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2x2_ASAP7_75t_L g302 ( 
.A(n_168),
.B(n_303),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_171),
.A2(n_277),
.B(n_282),
.Y(n_170)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_267),
.B(n_276),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_232),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_173),
.B(n_232),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_204),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_176),
.B1(n_190),
.B2(n_203),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_176),
.B(n_190),
.C(n_204),
.Y(n_268)
);

XNOR2x1_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_187),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_184),
.B(n_185),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g395 ( 
.A(n_185),
.B(n_349),
.Y(n_395)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

NOR2x1_ASAP7_75t_L g245 ( 
.A(n_186),
.B(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_187),
.A2(n_188),
.B1(n_274),
.B2(n_275),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_187),
.B(n_270),
.C(n_274),
.Y(n_281)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_188),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_189),
.B(n_304),
.Y(n_382)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g203 ( 
.A(n_191),
.Y(n_203)
);

OA21x2_ASAP7_75t_L g262 ( 
.A1(n_191),
.A2(n_192),
.B(n_194),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_194),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_195),
.B(n_427),
.Y(n_519)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_196),
.A2(n_248),
.B(n_249),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_196),
.B(n_248),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_196),
.B(n_459),
.Y(n_458)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_200),
.Y(n_476)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_220),
.B(n_231),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_205),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_205),
.A2(n_222),
.B1(n_223),
.B2(n_363),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_SL g447 ( 
.A1(n_205),
.A2(n_222),
.B1(n_448),
.B2(n_449),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_205),
.B(n_449),
.Y(n_520)
);

AO21x1_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_217),
.Y(n_205)
);

INVx3_ASAP7_75t_SL g206 ( 
.A(n_207),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g306 ( 
.A1(n_211),
.A2(n_307),
.B(n_314),
.Y(n_306)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_212),
.B(n_256),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_212),
.B(n_218),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_212),
.B(n_440),
.Y(n_439)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_215),
.Y(n_212)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_213),
.Y(n_315)
);

INVx8_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

BUFx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_216),
.Y(n_310)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_218),
.B(n_251),
.Y(n_250)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_219),
.Y(n_313)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_219),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_219),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_220),
.A2(n_221),
.B1(n_265),
.B2(n_266),
.Y(n_264)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_223),
.Y(n_221)
);

INVxp33_ASAP7_75t_SL g363 ( 
.A(n_223),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_229),
.B(n_230),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx5_ASAP7_75t_L g434 ( 
.A(n_228),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g451 ( 
.A(n_228),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_230),
.B(n_317),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_230),
.B(n_427),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_262),
.C(n_263),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_233),
.B(n_415),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_244),
.C(n_247),
.Y(n_233)
);

HB1xp67_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_235),
.B(n_245),
.Y(n_361)
);

BUFx12f_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx3_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g462 ( 
.A(n_246),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_247),
.B(n_361),
.Y(n_360)
);

XNOR2x2_ASAP7_75t_SL g320 ( 
.A(n_249),
.B(n_321),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_255),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_250),
.B(n_439),
.Y(n_438)
);

INVx4_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_253),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_255),
.A2(n_307),
.B(n_326),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g493 ( 
.A(n_255),
.B(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_256),
.B(n_315),
.Y(n_314)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g445 ( 
.A(n_259),
.Y(n_445)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g415 ( 
.A1(n_262),
.A2(n_263),
.B1(n_264),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_262),
.Y(n_416)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_265),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_292),
.Y(n_291)
);

NOR2xp67_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_268),
.B(n_269),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_277),
.Y(n_283)
);

NOR2x1_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_281),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_281),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B(n_286),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_286),
.C(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_293),
.Y(n_288)
);

INVxp67_ASAP7_75t_SL g290 ( 
.A(n_291),
.Y(n_290)
);

NAND2x1p5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_417),
.Y(n_293)
);

OAI21x1_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_370),
.B(n_407),
.Y(n_294)
);

NOR2x1_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_357),
.Y(n_295)
);

INVxp33_ASAP7_75t_SL g296 ( 
.A(n_297),
.Y(n_296)
);

AOI21x1_ASAP7_75t_L g405 ( 
.A1(n_297),
.A2(n_369),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_319),
.C(n_322),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_300),
.B(n_320),
.Y(n_387)
);

OAI22x1_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_302),
.B1(n_305),
.B2(n_318),
.Y(n_300)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_303),
.Y(n_368)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_305),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g366 ( 
.A(n_305),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_316),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_316),
.Y(n_384)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

BUFx3_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

INVx4_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

AND2x2_ASAP7_75t_SL g398 ( 
.A(n_314),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_314),
.B(n_439),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_317),
.B(n_459),
.Y(n_490)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVxp33_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_323),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_347),
.C(n_355),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_324),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g393 ( 
.A(n_325),
.B(n_328),
.Y(n_393)
);

INVx5_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_327),
.Y(n_495)
);

OAI31xp33_ASAP7_75t_L g328 ( 
.A1(n_329),
.A2(n_332),
.A3(n_335),
.B(n_339),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

BUFx4f_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

BUFx2_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_336),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_340),
.A2(n_344),
.B(n_346),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_341),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_345),
.Y(n_344)
);

INVxp67_ASAP7_75t_SL g347 ( 
.A(n_348),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_348),
.A2(n_355),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_377),
.Y(n_376)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_356),
.Y(n_377)
);

OAI21xp33_ASAP7_75t_SL g357 ( 
.A1(n_358),
.A2(n_364),
.B(n_369),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g369 ( 
.A(n_359),
.B(n_364),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_364),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_362),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_360),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_362),
.Y(n_412)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_365),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_365),
.B(n_410),
.C(n_412),
.Y(n_409)
);

INVxp33_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g370 ( 
.A1(n_371),
.A2(n_402),
.B(n_405),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_372),
.B(n_388),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g418 ( 
.A(n_372),
.B(n_419),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_385),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_373),
.Y(n_404)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_378),
.C(n_383),
.Y(n_373)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_374),
.B(n_401),
.Y(n_400)
);

HB1xp67_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_379),
.B(n_384),
.Y(n_401)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_380),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_381),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_391),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g403 ( 
.A(n_385),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_400),
.Y(n_388)
);

OR2x2_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_400),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_393),
.C(n_394),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_390),
.B(n_524),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_393),
.B(n_394),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g515 ( 
.A(n_395),
.B(n_516),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_396),
.A2(n_397),
.B1(n_398),
.B2(n_517),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_396),
.Y(n_517)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_399),
.B(n_494),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g527 ( 
.A1(n_405),
.A2(n_408),
.B(n_413),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_408),
.B(n_413),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g528 ( 
.A(n_409),
.B(n_414),
.Y(n_528)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

AOI31xp67_ASAP7_75t_L g417 ( 
.A1(n_418),
.A2(n_420),
.A3(n_527),
.B(n_528),
.Y(n_417)
);

OAI21x1_ASAP7_75t_L g420 ( 
.A1(n_421),
.A2(n_522),
.B(n_526),
.Y(n_420)
);

AOI21x1_ASAP7_75t_L g421 ( 
.A1(n_422),
.A2(n_511),
.B(n_521),
.Y(n_421)
);

AO21x1_ASAP7_75t_L g422 ( 
.A1(n_423),
.A2(n_464),
.B(n_510),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_424),
.B(n_446),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_424),
.B(n_446),
.Y(n_510)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_425),
.B(n_435),
.C(n_437),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g467 ( 
.A1(n_426),
.A2(n_435),
.B1(n_436),
.B2(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_426),
.Y(n_468)
);

INVx2_ASAP7_75t_SL g429 ( 
.A(n_430),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_433),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_438),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g466 ( 
.A(n_438),
.B(n_467),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_440),
.B(n_495),
.Y(n_494)
);

INVx4_ASAP7_75t_L g441 ( 
.A(n_442),
.Y(n_441)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_457),
.Y(n_446)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_447),
.Y(n_513)
);

INVxp67_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx3_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_454),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_458),
.A2(n_460),
.B1(n_461),
.B2(n_463),
.Y(n_457)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_458),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_460),
.B(n_463),
.C(n_513),
.Y(n_512)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_465),
.A2(n_491),
.B(n_509),
.Y(n_464)
);

NOR2x1_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_469),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_466),
.B(n_469),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_470),
.B(n_489),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_470),
.A2(n_471),
.B1(n_489),
.B2(n_490),
.Y(n_496)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_471),
.Y(n_470)
);

BUFx2_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx3_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

INVx4_ASAP7_75t_L g475 ( 
.A(n_476),
.Y(n_475)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_480),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_482),
.B(n_484),
.Y(n_481)
);

HB1xp67_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx2_ASAP7_75t_SL g485 ( 
.A(n_486),
.Y(n_485)
);

INVx3_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

AOI21xp5_ASAP7_75t_SL g491 ( 
.A1(n_492),
.A2(n_497),
.B(n_508),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_496),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g497 ( 
.A1(n_498),
.A2(n_501),
.B(n_507),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_499),
.B(n_500),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_499),
.B(n_500),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_504),
.B(n_506),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_505),
.Y(n_504)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_514),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_512),
.B(n_514),
.Y(n_521)
);

XOR2xp5_ASAP7_75t_L g514 ( 
.A(n_515),
.B(n_518),
.Y(n_514)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_515),
.B(n_519),
.C(n_520),
.Y(n_525)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_519),
.B(n_520),
.Y(n_518)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_523),
.B(n_525),
.Y(n_522)
);

OR2x2_ASAP7_75t_L g526 ( 
.A(n_523),
.B(n_525),
.Y(n_526)
);


endmodule