module real_jpeg_15277_n_4 (n_3, n_1, n_0, n_2, n_4);

input n_3;
input n_1;
input n_0;
input n_2;

output n_4;

wire n_5;
wire n_12;
wire n_8;
wire n_11;
wire n_6;
wire n_7;
wire n_10;
wire n_9;

AOI21xp5_ASAP7_75t_SL g5 ( 
.A1(n_0),
.A2(n_6),
.B(n_10),
.Y(n_5)
);

INVx2_ASAP7_75t_R g9 ( 
.A(n_1),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_L g4 ( 
.A1(n_2),
.A2(n_5),
.B1(n_11),
.B2(n_12),
.Y(n_4)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_2),
.Y(n_11)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_7),
.B(n_9),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_SL g10 ( 
.A(n_7),
.B(n_9),
.Y(n_10)
);

INVx2_ASAP7_75t_R g7 ( 
.A(n_8),
.Y(n_7)
);


endmodule