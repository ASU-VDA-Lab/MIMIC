module fake_netlist_1_3367_n_674 (n_44, n_81, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_87, n_74, n_7, n_29, n_45, n_85, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_82, n_15, n_61, n_21, n_51, n_39, n_674);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_87;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_82;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_674;
wire n_117;
wire n_663;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_476;
wire n_384;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_482;
wire n_394;
wire n_415;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_428;
wire n_364;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_570;
wire n_508;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g88 ( .A(n_46), .Y(n_88) );
CKINVDCx20_ASAP7_75t_R g89 ( .A(n_48), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_28), .Y(n_90) );
CKINVDCx20_ASAP7_75t_R g91 ( .A(n_22), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_53), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_66), .Y(n_93) );
BUFx2_ASAP7_75t_L g94 ( .A(n_80), .Y(n_94) );
CKINVDCx16_ASAP7_75t_R g95 ( .A(n_31), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_59), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_82), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_54), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_38), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_24), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_49), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_73), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_45), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_50), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_7), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_36), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_52), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_43), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
CKINVDCx16_ASAP7_75t_R g111 ( .A(n_44), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_69), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_81), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_67), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_47), .Y(n_116) );
NOR2xp67_ASAP7_75t_L g117 ( .A(n_40), .B(n_14), .Y(n_117) );
BUFx2_ASAP7_75t_L g118 ( .A(n_55), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_14), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_41), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_75), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_3), .Y(n_122) );
INVx2_ASAP7_75t_L g123 ( .A(n_35), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_110), .Y(n_124) );
INVx3_ASAP7_75t_L g125 ( .A(n_110), .Y(n_125) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_108), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_98), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_98), .Y(n_128) );
INVx4_ASAP7_75t_L g129 ( .A(n_94), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_89), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_90), .Y(n_132) );
OAI21x1_ASAP7_75t_L g133 ( .A1(n_102), .A2(n_42), .B(n_86), .Y(n_133) );
NAND2xp33_ASAP7_75t_R g134 ( .A(n_94), .B(n_0), .Y(n_134) );
AND2x4_ASAP7_75t_L g135 ( .A(n_118), .B(n_1), .Y(n_135) );
XNOR2x2_ASAP7_75t_L g136 ( .A(n_105), .B(n_3), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_118), .B(n_4), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_102), .Y(n_138) );
AND2x4_ASAP7_75t_L g139 ( .A(n_113), .B(n_4), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_96), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_113), .Y(n_141) );
OA21x2_ASAP7_75t_L g142 ( .A1(n_96), .A2(n_56), .B(n_85), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_108), .B(n_5), .Y(n_143) );
INVx1_ASAP7_75t_L g144 ( .A(n_97), .Y(n_144) );
INVx4_ASAP7_75t_L g145 ( .A(n_99), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_127), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_129), .B(n_95), .Y(n_147) );
BUFx10_ASAP7_75t_L g148 ( .A(n_135), .Y(n_148) );
INVx3_ASAP7_75t_L g149 ( .A(n_139), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_139), .Y(n_150) );
AND2x4_ASAP7_75t_L g151 ( .A(n_129), .B(n_119), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_127), .Y(n_152) );
INVx3_ASAP7_75t_L g153 ( .A(n_139), .Y(n_153) );
AOI22xp33_ASAP7_75t_L g154 ( .A1(n_135), .A2(n_122), .B1(n_112), .B2(n_97), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_127), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_139), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_133), .Y(n_157) );
NAND2xp33_ASAP7_75t_R g158 ( .A(n_131), .B(n_112), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_133), .Y(n_159) );
CKINVDCx11_ASAP7_75t_R g160 ( .A(n_129), .Y(n_160) );
AOI22xp5_ASAP7_75t_L g161 ( .A1(n_134), .A2(n_122), .B1(n_91), .B2(n_111), .Y(n_161) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_129), .B(n_88), .Y(n_162) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_129), .B(n_99), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_145), .B(n_100), .Y(n_164) );
BUFx10_ASAP7_75t_L g165 ( .A(n_135), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_145), .B(n_100), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
AOI22xp33_ASAP7_75t_L g168 ( .A1(n_135), .A2(n_107), .B1(n_121), .B2(n_109), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_128), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_145), .B(n_130), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_137), .Y(n_171) );
INVx2_ASAP7_75t_SL g172 ( .A(n_145), .Y(n_172) );
NOR2x1p5_ASAP7_75t_L g173 ( .A(n_143), .B(n_103), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_135), .A2(n_107), .B1(n_92), .B2(n_106), .Y(n_174) );
INVx4_ASAP7_75t_L g175 ( .A(n_139), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_145), .B(n_130), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_128), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_133), .Y(n_178) );
BUFx2_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_132), .B(n_103), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_138), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_165), .B(n_132), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_179), .B(n_140), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_179), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_146), .Y(n_185) );
OR2x6_ASAP7_75t_L g186 ( .A(n_175), .B(n_143), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_151), .B(n_173), .Y(n_187) );
CKINVDCx5p33_ASAP7_75t_R g188 ( .A(n_160), .Y(n_188) );
AOI22xp33_ASAP7_75t_L g189 ( .A1(n_151), .A2(n_136), .B1(n_144), .B2(n_140), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_146), .Y(n_190) );
NOR2x1p5_ASAP7_75t_L g191 ( .A(n_147), .B(n_134), .Y(n_191) );
O2A1O1Ixp33_ASAP7_75t_L g192 ( .A1(n_171), .A2(n_144), .B(n_141), .C(n_138), .Y(n_192) );
NAND2x1p5_ASAP7_75t_L g193 ( .A(n_175), .B(n_126), .Y(n_193) );
INVx2_ASAP7_75t_SL g194 ( .A(n_165), .Y(n_194) );
INVx2_ASAP7_75t_SL g195 ( .A(n_165), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_161), .B(n_126), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_155), .Y(n_197) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_151), .A2(n_136), .B1(n_141), .B2(n_138), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_163), .B(n_114), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_165), .B(n_93), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_155), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_151), .B(n_124), .Y(n_203) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_175), .B(n_124), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_162), .B(n_114), .Y(n_205) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_148), .B(n_101), .Y(n_206) );
INVx3_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
NAND2xp5_ASAP7_75t_SL g208 ( .A(n_148), .B(n_104), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_173), .Y(n_209) );
AOI22xp33_ASAP7_75t_L g210 ( .A1(n_149), .A2(n_136), .B1(n_141), .B2(n_125), .Y(n_210) );
INVx3_ASAP7_75t_L g211 ( .A(n_149), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_167), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_170), .B(n_124), .Y(n_213) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_157), .B(n_115), .Y(n_214) );
AOI22xp5_ASAP7_75t_SL g215 ( .A1(n_161), .A2(n_158), .B1(n_149), .B2(n_153), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_166), .B(n_168), .Y(n_216) );
OAI22xp5_ASAP7_75t_SL g217 ( .A1(n_154), .A2(n_142), .B1(n_116), .B2(n_124), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_167), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_174), .B(n_125), .Y(n_219) );
OAI221xp5_ASAP7_75t_L g220 ( .A1(n_180), .A2(n_125), .B1(n_117), .B2(n_123), .C(n_120), .Y(n_220) );
NOR2xp33_ASAP7_75t_L g221 ( .A(n_164), .B(n_125), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_150), .B(n_123), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_200), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_194), .Y(n_224) );
O2A1O1Ixp33_ASAP7_75t_L g225 ( .A1(n_216), .A2(n_156), .B(n_150), .C(n_153), .Y(n_225) );
O2A1O1Ixp33_ASAP7_75t_L g226 ( .A1(n_183), .A2(n_156), .B(n_150), .C(n_153), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g227 ( .A(n_184), .B(n_209), .Y(n_227) );
O2A1O1Ixp33_ASAP7_75t_L g228 ( .A1(n_219), .A2(n_156), .B(n_176), .C(n_177), .Y(n_228) );
OAI21xp5_ASAP7_75t_L g229 ( .A1(n_214), .A2(n_172), .B(n_142), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_187), .B(n_177), .Y(n_230) );
NOR2xp33_ASAP7_75t_L g231 ( .A(n_209), .B(n_172), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_194), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_195), .B(n_157), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_196), .B(n_181), .Y(n_234) );
INVx2_ASAP7_75t_L g235 ( .A(n_200), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_182), .A2(n_157), .B(n_178), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_193), .B(n_181), .Y(n_237) );
AOI22xp33_ASAP7_75t_L g238 ( .A1(n_193), .A2(n_191), .B1(n_187), .B2(n_189), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_182), .A2(n_178), .B(n_159), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_203), .Y(n_240) );
NOR2xp33_ASAP7_75t_SL g241 ( .A(n_188), .B(n_178), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g242 ( .A1(n_192), .A2(n_169), .B(n_152), .C(n_159), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_195), .B(n_178), .Y(n_243) );
O2A1O1Ixp33_ASAP7_75t_L g244 ( .A1(n_210), .A2(n_169), .B(n_120), .C(n_142), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_187), .B(n_178), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_186), .B(n_159), .Y(n_246) );
CKINVDCx5p33_ASAP7_75t_R g247 ( .A(n_188), .Y(n_247) );
A2O1A1Ixp33_ASAP7_75t_SL g248 ( .A1(n_221), .A2(n_198), .B(n_220), .C(n_199), .Y(n_248) );
OAI22xp5_ASAP7_75t_L g249 ( .A1(n_186), .A2(n_159), .B1(n_157), .B2(n_142), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_186), .B(n_159), .Y(n_250) );
CKINVDCx16_ASAP7_75t_R g251 ( .A(n_215), .Y(n_251) );
BUFx2_ASAP7_75t_L g252 ( .A(n_186), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g253 ( .A(n_205), .B(n_157), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_203), .B(n_142), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g255 ( .A(n_204), .B(n_5), .Y(n_255) );
OAI21x1_ASAP7_75t_L g256 ( .A1(n_249), .A2(n_214), .B(n_222), .Y(n_256) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_236), .A2(n_201), .B(n_206), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_234), .B(n_211), .Y(n_258) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_239), .A2(n_201), .B(n_206), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g260 ( .A1(n_238), .A2(n_208), .B1(n_207), .B2(n_217), .Y(n_260) );
OA21x2_ASAP7_75t_L g261 ( .A1(n_229), .A2(n_242), .B(n_254), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_223), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_233), .A2(n_208), .B(n_213), .Y(n_263) );
AND2x2_ASAP7_75t_L g264 ( .A(n_237), .B(n_185), .Y(n_264) );
AOI21xp5_ASAP7_75t_L g265 ( .A1(n_233), .A2(n_218), .B(n_212), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_223), .Y(n_266) );
OAI21xp5_ASAP7_75t_L g267 ( .A1(n_242), .A2(n_202), .B(n_197), .Y(n_267) );
OAI21x1_ASAP7_75t_L g268 ( .A1(n_244), .A2(n_204), .B(n_190), .Y(n_268) );
INVx3_ASAP7_75t_L g269 ( .A(n_224), .Y(n_269) );
AOI21xp5_ASAP7_75t_SL g270 ( .A1(n_246), .A2(n_207), .B(n_57), .Y(n_270) );
BUFx3_ASAP7_75t_L g271 ( .A(n_224), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_235), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_235), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_251), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g275 ( .A1(n_243), .A2(n_211), .B(n_207), .Y(n_275) );
AO31x2_ASAP7_75t_L g276 ( .A1(n_253), .A2(n_211), .A3(n_7), .B(n_8), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_243), .A2(n_51), .B(n_84), .Y(n_277) );
OAI21x1_ASAP7_75t_L g278 ( .A1(n_268), .A2(n_250), .B(n_225), .Y(n_278) );
AND2x4_ASAP7_75t_L g279 ( .A(n_264), .B(n_252), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_264), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_266), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_262), .Y(n_282) );
AOI222xp33_ASAP7_75t_L g283 ( .A1(n_258), .A2(n_240), .B1(n_227), .B2(n_247), .C1(n_230), .C2(n_255), .Y(n_283) );
AOI21xp33_ASAP7_75t_SL g284 ( .A1(n_274), .A2(n_247), .B(n_8), .Y(n_284) );
OAI21x1_ASAP7_75t_L g285 ( .A1(n_268), .A2(n_245), .B(n_226), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_262), .Y(n_286) );
AND2x4_ASAP7_75t_L g287 ( .A(n_266), .B(n_224), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g288 ( .A1(n_257), .A2(n_248), .B(n_228), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_272), .Y(n_289) );
AO31x2_ASAP7_75t_L g290 ( .A1(n_265), .A2(n_231), .A3(n_248), .B(n_241), .Y(n_290) );
OAI21x1_ASAP7_75t_L g291 ( .A1(n_256), .A2(n_232), .B(n_224), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_272), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_260), .B(n_232), .C(n_9), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_273), .Y(n_294) );
OAI21x1_ASAP7_75t_L g295 ( .A1(n_256), .A2(n_232), .B(n_58), .Y(n_295) );
OA21x2_ASAP7_75t_L g296 ( .A1(n_267), .A2(n_232), .B(n_60), .Y(n_296) );
BUFx10_ASAP7_75t_L g297 ( .A(n_274), .Y(n_297) );
AO21x2_ASAP7_75t_L g298 ( .A1(n_270), .A2(n_6), .B(n_9), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_273), .B(n_6), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_271), .B(n_10), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_276), .Y(n_301) );
OA21x2_ASAP7_75t_L g302 ( .A1(n_291), .A2(n_259), .B(n_263), .Y(n_302) );
OA21x2_ASAP7_75t_L g303 ( .A1(n_291), .A2(n_301), .B(n_295), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_282), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_286), .Y(n_305) );
AO21x2_ASAP7_75t_L g306 ( .A1(n_301), .A2(n_270), .B(n_277), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_286), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_287), .Y(n_308) );
INVx2_ASAP7_75t_SL g309 ( .A(n_287), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_281), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_287), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_289), .Y(n_312) );
AOI21xp5_ASAP7_75t_L g313 ( .A1(n_288), .A2(n_261), .B(n_275), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_280), .B(n_289), .Y(n_314) );
INVx2_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
INVx2_ASAP7_75t_SL g316 ( .A(n_287), .Y(n_316) );
OA21x2_ASAP7_75t_L g317 ( .A1(n_295), .A2(n_261), .B(n_276), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_280), .B(n_269), .Y(n_318) );
AO21x2_ASAP7_75t_L g319 ( .A1(n_293), .A2(n_261), .B(n_276), .Y(n_319) );
OA21x2_ASAP7_75t_L g320 ( .A1(n_278), .A2(n_261), .B(n_276), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_294), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_281), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_292), .Y(n_323) );
OR2x6_ASAP7_75t_L g324 ( .A(n_293), .B(n_271), .Y(n_324) );
AO21x2_ASAP7_75t_L g325 ( .A1(n_278), .A2(n_276), .B(n_269), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_292), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_279), .B(n_269), .Y(n_327) );
AO21x2_ASAP7_75t_L g328 ( .A1(n_285), .A2(n_10), .B(n_11), .Y(n_328) );
INVx2_ASAP7_75t_SL g329 ( .A(n_279), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
OR2x2_ASAP7_75t_L g331 ( .A(n_279), .B(n_11), .Y(n_331) );
INVxp67_ASAP7_75t_L g332 ( .A(n_279), .Y(n_332) );
INVx3_ASAP7_75t_L g333 ( .A(n_285), .Y(n_333) );
INVxp67_ASAP7_75t_SL g334 ( .A(n_283), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_296), .Y(n_335) );
AO21x2_ASAP7_75t_L g336 ( .A1(n_298), .A2(n_12), .B(n_13), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_298), .Y(n_337) );
INVx6_ASAP7_75t_L g338 ( .A(n_297), .Y(n_338) );
BUFx3_ASAP7_75t_L g339 ( .A(n_338), .Y(n_339) );
INVx5_ASAP7_75t_L g340 ( .A(n_338), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_331), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_310), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_310), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_310), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_334), .B(n_284), .Y(n_345) );
BUFx2_ASAP7_75t_L g346 ( .A(n_315), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_315), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_322), .B(n_298), .Y(n_348) );
AND2x2_ASAP7_75t_L g349 ( .A(n_322), .B(n_315), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_323), .B(n_296), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND2x4_ASAP7_75t_L g352 ( .A(n_308), .B(n_290), .Y(n_352) );
OR2x2_ASAP7_75t_L g353 ( .A(n_312), .B(n_300), .Y(n_353) );
AND2x4_ASAP7_75t_SL g354 ( .A(n_314), .B(n_297), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_331), .Y(n_355) );
HB1xp67_ASAP7_75t_L g356 ( .A(n_314), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_323), .Y(n_357) );
AND2x2_ASAP7_75t_L g358 ( .A(n_326), .B(n_296), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_304), .B(n_284), .Y(n_359) );
AND2x2_ASAP7_75t_L g360 ( .A(n_326), .B(n_296), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_304), .B(n_297), .Y(n_361) );
AND2x2_ASAP7_75t_L g362 ( .A(n_305), .B(n_290), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_312), .Y(n_363) );
AND2x4_ASAP7_75t_SL g364 ( .A(n_327), .B(n_297), .Y(n_364) );
INVx1_ASAP7_75t_SL g365 ( .A(n_338), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_305), .B(n_290), .Y(n_366) );
AND2x4_ASAP7_75t_L g367 ( .A(n_308), .B(n_290), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_307), .B(n_290), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_338), .Y(n_369) );
AND2x2_ASAP7_75t_L g370 ( .A(n_307), .B(n_290), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_321), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_321), .B(n_308), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g373 ( .A1(n_330), .A2(n_13), .B1(n_15), .B2(n_16), .Y(n_373) );
HB1xp67_ASAP7_75t_L g374 ( .A(n_311), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_337), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_303), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_303), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_325), .Y(n_378) );
BUFx3_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_330), .B(n_16), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_332), .B(n_17), .Y(n_381) );
INVx5_ASAP7_75t_L g382 ( .A(n_324), .Y(n_382) );
BUFx2_ASAP7_75t_L g383 ( .A(n_308), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_303), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_329), .B(n_18), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_319), .B(n_19), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_303), .Y(n_387) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_329), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_325), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_329), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_332), .B(n_87), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_320), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_319), .B(n_20), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_318), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_309), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_309), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_319), .B(n_21), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_309), .Y(n_398) );
OR2x6_ASAP7_75t_L g399 ( .A(n_324), .B(n_23), .Y(n_399) );
BUFx3_ASAP7_75t_L g400 ( .A(n_316), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_362), .B(n_320), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_362), .B(n_320), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_366), .B(n_320), .Y(n_403) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_345), .B(n_336), .Y(n_404) );
INVx2_ASAP7_75t_L g405 ( .A(n_346), .Y(n_405) );
OR2x2_ASAP7_75t_L g406 ( .A(n_356), .B(n_316), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_341), .B(n_327), .Y(n_407) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_346), .Y(n_408) );
INVxp33_ASAP7_75t_L g409 ( .A(n_349), .Y(n_409) );
AND2x2_ASAP7_75t_L g410 ( .A(n_366), .B(n_325), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g411 ( .A(n_359), .B(n_336), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_370), .B(n_325), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_370), .B(n_319), .Y(n_413) );
OR2x2_ASAP7_75t_L g414 ( .A(n_357), .B(n_316), .Y(n_414) );
OR2x2_ASAP7_75t_L g415 ( .A(n_357), .B(n_336), .Y(n_415) );
AND2x2_ASAP7_75t_L g416 ( .A(n_348), .B(n_317), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_348), .B(n_317), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_372), .B(n_317), .Y(n_418) );
NOR2x1_ASAP7_75t_SL g419 ( .A(n_399), .B(n_336), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_355), .B(n_328), .Y(n_420) );
AND2x4_ASAP7_75t_SL g421 ( .A(n_399), .B(n_324), .Y(n_421) );
AND2x2_ASAP7_75t_L g422 ( .A(n_372), .B(n_317), .Y(n_422) );
AND2x2_ASAP7_75t_L g423 ( .A(n_352), .B(n_328), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_352), .B(n_328), .Y(n_424) );
INVx3_ASAP7_75t_SL g425 ( .A(n_340), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_363), .B(n_328), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_352), .B(n_333), .Y(n_427) );
INVxp67_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
OR2x2_ASAP7_75t_L g429 ( .A(n_371), .B(n_313), .Y(n_429) );
INVxp67_ASAP7_75t_SL g430 ( .A(n_342), .Y(n_430) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_349), .B(n_313), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_352), .B(n_333), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_342), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_361), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_353), .Y(n_435) );
INVx3_ASAP7_75t_L g436 ( .A(n_382), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_353), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_367), .B(n_333), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_343), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_343), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_367), .B(n_333), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_367), .B(n_302), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_367), .B(n_302), .Y(n_443) );
HB1xp67_ASAP7_75t_L g444 ( .A(n_374), .Y(n_444) );
INVx1_ASAP7_75t_SL g445 ( .A(n_354), .Y(n_445) );
INVxp67_ASAP7_75t_L g446 ( .A(n_380), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_351), .B(n_324), .Y(n_447) );
INVxp67_ASAP7_75t_SL g448 ( .A(n_344), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_368), .B(n_302), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_354), .B(n_324), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_375), .B(n_302), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_375), .B(n_302), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_378), .B(n_335), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_354), .B(n_306), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_351), .B(n_306), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_344), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_347), .Y(n_457) );
OR2x2_ASAP7_75t_L g458 ( .A(n_347), .B(n_335), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_392), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_398), .B(n_306), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_378), .B(n_306), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_388), .B(n_25), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_390), .B(n_26), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_389), .B(n_27), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_392), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_383), .Y(n_466) );
NOR2xp67_ASAP7_75t_L g467 ( .A(n_382), .B(n_29), .Y(n_467) );
INVx1_ASAP7_75t_SL g468 ( .A(n_365), .Y(n_468) );
BUFx3_ASAP7_75t_L g469 ( .A(n_340), .Y(n_469) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_373), .B(n_30), .Y(n_470) );
INVx1_ASAP7_75t_SL g471 ( .A(n_369), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_389), .B(n_32), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_350), .B(n_360), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_395), .B(n_33), .Y(n_474) );
NOR2x1_ASAP7_75t_SL g475 ( .A(n_399), .B(n_34), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_340), .Y(n_476) );
BUFx2_ASAP7_75t_SL g477 ( .A(n_340), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_350), .B(n_37), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_395), .Y(n_479) );
INVx2_ASAP7_75t_L g480 ( .A(n_376), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g481 ( .A(n_340), .B(n_39), .Y(n_481) );
NAND2x1_ASAP7_75t_L g482 ( .A(n_436), .B(n_399), .Y(n_482) );
INVxp67_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_409), .B(n_400), .Y(n_484) );
NAND2xp67_ASAP7_75t_SL g485 ( .A(n_478), .B(n_393), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_409), .B(n_400), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_473), .B(n_400), .Y(n_487) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_436), .B(n_399), .Y(n_488) );
INVx2_ASAP7_75t_SL g489 ( .A(n_425), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_473), .B(n_396), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_428), .B(n_396), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_468), .B(n_396), .Y(n_492) );
INVx1_ASAP7_75t_SL g493 ( .A(n_425), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_471), .B(n_395), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_404), .B(n_393), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_435), .B(n_382), .Y(n_496) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_404), .B(n_386), .Y(n_497) );
AND2x2_ASAP7_75t_L g498 ( .A(n_437), .B(n_382), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_406), .B(n_379), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_434), .B(n_382), .Y(n_500) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_446), .B(n_339), .Y(n_501) );
NOR2xp33_ASAP7_75t_L g502 ( .A(n_407), .B(n_339), .Y(n_502) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_411), .B(n_373), .C(n_386), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_408), .B(n_414), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_405), .Y(n_505) );
INVxp67_ASAP7_75t_SL g506 ( .A(n_430), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_469), .Y(n_507) );
INVx2_ASAP7_75t_L g508 ( .A(n_405), .Y(n_508) );
INVx2_ASAP7_75t_L g509 ( .A(n_459), .Y(n_509) );
AND2x4_ASAP7_75t_L g510 ( .A(n_421), .B(n_379), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_401), .B(n_402), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_402), .B(n_379), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_411), .B(n_358), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
INVx1_ASAP7_75t_SL g515 ( .A(n_476), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_466), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_410), .B(n_358), .Y(n_517) );
INVx1_ASAP7_75t_SL g518 ( .A(n_477), .Y(n_518) );
BUFx2_ASAP7_75t_L g519 ( .A(n_469), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_448), .Y(n_520) );
INVx3_ASAP7_75t_SL g521 ( .A(n_445), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_403), .B(n_339), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_465), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_451), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_410), .B(n_360), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_427), .B(n_384), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_412), .B(n_384), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_403), .B(n_364), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_413), .B(n_387), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_413), .B(n_387), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_433), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_451), .B(n_377), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_452), .B(n_377), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_449), .B(n_397), .Y(n_534) );
OR2x2_ASAP7_75t_L g535 ( .A(n_431), .B(n_397), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_452), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_427), .B(n_376), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_449), .B(n_385), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_433), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_432), .B(n_385), .Y(n_540) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_416), .B(n_391), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_416), .B(n_381), .Y(n_542) );
OAI21xp33_ASAP7_75t_L g543 ( .A1(n_420), .A2(n_61), .B(n_62), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_438), .B(n_63), .Y(n_544) );
OAI211xp5_ASAP7_75t_L g545 ( .A1(n_454), .A2(n_64), .B(n_65), .C(n_68), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_439), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_439), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_440), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_441), .B(n_70), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_440), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_417), .B(n_418), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_417), .B(n_71), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_479), .B(n_72), .Y(n_553) );
NAND2x1_ASAP7_75t_L g554 ( .A(n_467), .B(n_74), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_418), .B(n_76), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_456), .Y(n_556) );
INVx1_ASAP7_75t_L g557 ( .A(n_456), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_513), .B(n_461), .Y(n_558) );
HB1xp67_ASAP7_75t_L g559 ( .A(n_506), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_513), .B(n_461), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_551), .B(n_422), .Y(n_561) );
BUFx2_ASAP7_75t_L g562 ( .A(n_521), .Y(n_562) );
INVx2_ASAP7_75t_L g563 ( .A(n_520), .Y(n_563) );
INVx1_ASAP7_75t_SL g564 ( .A(n_493), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_551), .B(n_422), .Y(n_565) );
INVxp67_ASAP7_75t_SL g566 ( .A(n_482), .Y(n_566) );
INVxp67_ASAP7_75t_L g567 ( .A(n_501), .Y(n_567) );
INVxp67_ASAP7_75t_L g568 ( .A(n_519), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_524), .B(n_426), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g570 ( .A(n_483), .B(n_470), .Y(n_570) );
INVx2_ASAP7_75t_L g571 ( .A(n_522), .Y(n_571) );
AND2x4_ASAP7_75t_L g572 ( .A(n_528), .B(n_443), .Y(n_572) );
INVx1_ASAP7_75t_SL g573 ( .A(n_493), .Y(n_573) );
NOR2xp33_ASAP7_75t_L g574 ( .A(n_491), .B(n_470), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_511), .B(n_441), .Y(n_575) );
AND2x2_ASAP7_75t_SL g576 ( .A(n_510), .B(n_450), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_492), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_536), .B(n_429), .Y(n_578) );
INVx2_ASAP7_75t_L g579 ( .A(n_509), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_517), .B(n_423), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_517), .B(n_415), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_525), .B(n_423), .Y(n_582) );
INVx3_ASAP7_75t_L g583 ( .A(n_488), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_512), .B(n_443), .Y(n_584) );
INVxp67_ASAP7_75t_SL g585 ( .A(n_532), .Y(n_585) );
OAI22xp5_ASAP7_75t_L g586 ( .A1(n_503), .A2(n_447), .B1(n_462), .B2(n_474), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_516), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_527), .B(n_457), .Y(n_588) );
OAI21xp33_ASAP7_75t_L g589 ( .A1(n_495), .A2(n_424), .B(n_455), .Y(n_589) );
AND2x4_ASAP7_75t_L g590 ( .A(n_510), .B(n_442), .Y(n_590) );
AND2x2_ASAP7_75t_L g591 ( .A(n_487), .B(n_442), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_490), .B(n_419), .Y(n_592) );
OR2x2_ASAP7_75t_L g593 ( .A(n_529), .B(n_457), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_529), .B(n_453), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_514), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_484), .B(n_460), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_530), .B(n_480), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_530), .B(n_480), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_504), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_532), .B(n_458), .Y(n_600) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_503), .A2(n_472), .B1(n_464), .B2(n_481), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_533), .B(n_472), .Y(n_602) );
INVx1_ASAP7_75t_SL g603 ( .A(n_518), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_523), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_533), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_531), .Y(n_606) );
OA22x2_ASAP7_75t_L g607 ( .A1(n_562), .A2(n_489), .B1(n_507), .B2(n_515), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_570), .A2(n_502), .B1(n_497), .B2(n_495), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_559), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_585), .B(n_497), .Y(n_610) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_574), .A2(n_500), .B1(n_542), .B2(n_541), .Y(n_611) );
INVx1_ASAP7_75t_SL g612 ( .A(n_603), .Y(n_612) );
AOI322xp5_ASAP7_75t_L g613 ( .A1(n_566), .A2(n_534), .A3(n_538), .B1(n_486), .B2(n_540), .C1(n_542), .C2(n_541), .Y(n_613) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_552), .B(n_555), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_605), .B(n_537), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_584), .B(n_494), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_591), .B(n_526), .Y(n_617) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_576), .A2(n_499), .B1(n_515), .B2(n_538), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_558), .B(n_505), .Y(n_619) );
OAI31xp33_ASAP7_75t_L g620 ( .A1(n_583), .A2(n_545), .A3(n_549), .B(n_544), .Y(n_620) );
OAI33xp33_ASAP7_75t_L g621 ( .A1(n_567), .A2(n_485), .A3(n_552), .B1(n_535), .B2(n_556), .B3(n_548), .Y(n_621) );
OR2x2_ASAP7_75t_L g622 ( .A(n_561), .B(n_508), .Y(n_622) );
AOI222xp33_ASAP7_75t_L g623 ( .A1(n_589), .A2(n_526), .B1(n_496), .B2(n_498), .C1(n_475), .C2(n_549), .Y(n_623) );
O2A1O1Ixp33_ASAP7_75t_L g624 ( .A1(n_586), .A2(n_481), .B(n_554), .C(n_543), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_588), .Y(n_625) );
AOI21xp33_ASAP7_75t_SL g626 ( .A1(n_583), .A2(n_553), .B(n_463), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_575), .B(n_557), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_558), .B(n_547), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_601), .A2(n_546), .B1(n_550), .B2(n_539), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_560), .B(n_464), .Y(n_630) );
INVx1_ASAP7_75t_SL g631 ( .A(n_564), .Y(n_631) );
OR2x2_ASAP7_75t_L g632 ( .A(n_565), .B(n_77), .Y(n_632) );
INVx1_ASAP7_75t_SL g633 ( .A(n_564), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g634 ( .A(n_573), .B(n_78), .Y(n_634) );
HB1xp67_ASAP7_75t_L g635 ( .A(n_573), .Y(n_635) );
NOR2xp33_ASAP7_75t_R g636 ( .A(n_568), .B(n_79), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_609), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g638 ( .A1(n_607), .A2(n_596), .B1(n_599), .B2(n_592), .Y(n_638) );
AOI21xp33_ASAP7_75t_L g639 ( .A1(n_620), .A2(n_586), .B(n_587), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_613), .B(n_560), .Y(n_640) );
AOI22xp5_ASAP7_75t_L g641 ( .A1(n_607), .A2(n_577), .B1(n_590), .B2(n_578), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_623), .A2(n_590), .B1(n_602), .B2(n_571), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g643 ( .A1(n_618), .A2(n_629), .B1(n_608), .B2(n_611), .Y(n_643) );
OAI221xp5_ASAP7_75t_L g644 ( .A1(n_624), .A2(n_578), .B1(n_569), .B2(n_563), .C(n_580), .Y(n_644) );
AOI21xp33_ASAP7_75t_L g645 ( .A1(n_624), .A2(n_602), .B(n_581), .Y(n_645) );
OAI311xp33_ASAP7_75t_L g646 ( .A1(n_611), .A2(n_582), .A3(n_597), .B1(n_598), .C1(n_593), .Y(n_646) );
OAI322xp33_ASAP7_75t_SL g647 ( .A1(n_615), .A2(n_594), .A3(n_600), .B1(n_606), .B2(n_604), .C1(n_579), .C2(n_595), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_635), .B(n_572), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_635), .B(n_83), .Y(n_649) );
AOI211xp5_ASAP7_75t_SL g650 ( .A1(n_614), .A2(n_632), .B(n_636), .C(n_630), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g651 ( .A1(n_631), .A2(n_633), .B1(n_628), .B2(n_619), .C(n_625), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_626), .A2(n_627), .B1(n_636), .B2(n_616), .C(n_622), .Y(n_652) );
NOR3xp33_ASAP7_75t_L g653 ( .A(n_634), .B(n_621), .C(n_624), .Y(n_653) );
NOR3x1_ASAP7_75t_L g654 ( .A(n_617), .B(n_562), .C(n_566), .Y(n_654) );
OAI322xp33_ASAP7_75t_L g655 ( .A1(n_607), .A2(n_608), .A3(n_610), .B1(n_609), .B2(n_483), .C1(n_612), .C2(n_618), .Y(n_655) );
NOR2x1_ASAP7_75t_L g656 ( .A(n_655), .B(n_644), .Y(n_656) );
AOI21xp5_ASAP7_75t_L g657 ( .A1(n_647), .A2(n_644), .B(n_653), .Y(n_657) );
NOR2xp33_ASAP7_75t_SL g658 ( .A(n_639), .B(n_645), .Y(n_658) );
HB1xp67_ASAP7_75t_L g659 ( .A(n_637), .Y(n_659) );
NOR4xp25_ASAP7_75t_L g660 ( .A(n_646), .B(n_640), .C(n_651), .D(n_642), .Y(n_660) );
NAND2x1p5_ASAP7_75t_L g661 ( .A(n_656), .B(n_654), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_659), .Y(n_662) );
NAND3xp33_ASAP7_75t_L g663 ( .A(n_657), .B(n_650), .C(n_652), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_662), .Y(n_664) );
NOR2x1_ASAP7_75t_L g665 ( .A(n_663), .B(n_649), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_664), .Y(n_666) );
BUFx2_ASAP7_75t_L g667 ( .A(n_665), .Y(n_667) );
AND2x4_ASAP7_75t_L g668 ( .A(n_666), .B(n_643), .Y(n_668) );
AND2x4_ASAP7_75t_L g669 ( .A(n_667), .B(n_648), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_668), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_670), .B(n_669), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_671), .B(n_660), .Y(n_672) );
OR2x6_ASAP7_75t_L g673 ( .A(n_672), .B(n_661), .Y(n_673) );
AOI22xp5_ASAP7_75t_L g674 ( .A1(n_673), .A2(n_658), .B1(n_638), .B2(n_641), .Y(n_674) );
endmodule