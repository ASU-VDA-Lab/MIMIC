module fake_jpeg_8491_n_42 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_42);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_42;

wire n_21;
wire n_33;
wire n_23;
wire n_27;
wire n_22;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_36;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_32;
wire n_15;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_19),
.A2(n_20),
.B1(n_16),
.B2(n_17),
.Y(n_21)
);

AOI21xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_24),
.B(n_8),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_0),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_13),
.B1(n_5),
.B2(n_6),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

INVxp67_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_26),
.B(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

AND2x6_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_21),
.Y(n_30)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_21),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_31),
.B(n_33),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_39),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_SL g39 ( 
.A(n_35),
.B(n_34),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g41 ( 
.A1(n_40),
.A2(n_36),
.B(n_32),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g42 ( 
.A1(n_41),
.A2(n_27),
.B(n_12),
.Y(n_42)
);


endmodule