module real_jpeg_20996_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_288;
wire n_166;
wire n_176;
wire n_249;
wire n_215;
wire n_221;
wire n_292;
wire n_286;
wire n_194;
wire n_153;
wire n_104;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_40;
wire n_105;
wire n_299;
wire n_173;
wire n_243;
wire n_115;
wire n_197;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_178;
wire n_79;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_258;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_297;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_240;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

INVx13_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_1),
.A2(n_42),
.B1(n_43),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_2),
.A2(n_29),
.B1(n_30),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_2),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_2),
.A2(n_25),
.B1(n_27),
.B2(n_149),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_2),
.A2(n_42),
.B1(n_43),
.B2(n_149),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_149),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g142 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_3),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_143),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_143),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_3),
.A2(n_42),
.B1(n_43),
.B2(n_143),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_4),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_24),
.Y(n_176)
);

AOI21xp33_ASAP7_75t_L g198 ( 
.A1(n_4),
.A2(n_14),
.B(n_49),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_4),
.A2(n_42),
.B1(n_43),
.B2(n_147),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_4),
.A2(n_80),
.B1(n_134),
.B2(n_207),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_180),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_4),
.B(n_27),
.Y(n_231)
);

AOI21xp33_ASAP7_75t_L g235 ( 
.A1(n_4),
.A2(n_27),
.B(n_231),
.Y(n_235)
);

BUFx16f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_6),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_42),
.B1(n_43),
.B2(n_64),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_64),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_31),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_7),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_7),
.A2(n_25),
.B1(n_27),
.B2(n_31),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_7),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_7),
.A2(n_31),
.B1(n_48),
.B2(n_49),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_8),
.B(n_48),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_8),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_8),
.B(n_84),
.Y(n_107)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_8),
.Y(n_134)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_10),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_10),
.A2(n_25),
.B1(n_27),
.B2(n_113),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_10),
.A2(n_48),
.B1(n_49),
.B2(n_113),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_10),
.A2(n_42),
.B1(n_43),
.B2(n_113),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_34),
.Y(n_33)
);

CKINVDCx14_ASAP7_75t_R g34 ( 
.A(n_13),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_13),
.A2(n_25),
.B1(n_27),
.B2(n_34),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_13),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_13),
.A2(n_34),
.B1(n_48),
.B2(n_49),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g41 ( 
.A1(n_14),
.A2(n_42),
.B(n_46),
.C(n_47),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_14),
.B(n_42),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_14),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_14),
.Y(n_50)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_121),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_119),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_94),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_19),
.B(n_94),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g300 ( 
.A(n_19),
.Y(n_300)
);

FAx1_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_67),
.CI(n_76),
.CON(n_19),
.SN(n_19)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_37),
.B2(n_38),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_32),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_23),
.A2(n_90),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_23),
.A2(n_90),
.B1(n_112),
.B2(n_160),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g35 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_24),
.B(n_33),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_24),
.B(n_92),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_24),
.A2(n_35),
.B1(n_146),
.B2(n_148),
.Y(n_145)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_25),
.A2(n_36),
.B1(n_146),
.B2(n_153),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g230 ( 
.A1(n_25),
.A2(n_42),
.A3(n_59),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_26),
.B(n_27),
.Y(n_153)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_58),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g146 ( 
.A(n_30),
.B(n_147),
.CON(n_146),
.SN(n_146)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_35),
.Y(n_32)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_54),
.B2(n_55),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_47),
.B(n_51),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_41),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g85 ( 
.A1(n_41),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_41),
.A2(n_47),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_41),
.A2(n_51),
.B(n_87),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_41),
.A2(n_47),
.B1(n_201),
.B2(n_202),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_41),
.A2(n_47),
.B1(n_202),
.B2(n_222),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_41),
.A2(n_47),
.B1(n_222),
.B2(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_41),
.A2(n_71),
.B(n_238),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_43),
.B1(n_58),
.B2(n_59),
.Y(n_61)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

A2O1A1Ixp33_ASAP7_75t_L g197 ( 
.A1(n_43),
.A2(n_50),
.B(n_147),
.C(n_198),
.Y(n_197)
);

NAND2xp33_ASAP7_75t_SL g232 ( 
.A(n_43),
.B(n_58),
.Y(n_232)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_47),
.A2(n_73),
.B(n_109),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_47),
.B(n_147),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_48),
.B(n_211),
.Y(n_210)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_52),
.B(n_72),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_65),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_56),
.B(n_118),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_56),
.A2(n_163),
.B(n_164),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_56),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_56),
.A2(n_65),
.B(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_57),
.A2(n_61),
.B1(n_63),
.B2(n_69),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_57),
.A2(n_61),
.B1(n_142),
.B2(n_144),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_57),
.A2(n_61),
.B1(n_179),
.B2(n_235),
.Y(n_234)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_61),
.B(n_66),
.Y(n_65)
);

OAI21xp5_ASAP7_75t_L g116 ( 
.A1(n_61),
.A2(n_69),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_61),
.B(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_61),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_66),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_67),
.A2(n_68),
.B(n_70),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_70),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_73),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_72),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_75),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_89),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_77),
.A2(n_78),
.B1(n_96),
.B2(n_97),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_85),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_79),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_79),
.A2(n_88),
.B1(n_89),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_79),
.A2(n_85),
.B1(n_88),
.B2(n_291),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_82),
.B(n_83),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_80),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_80),
.A2(n_131),
.B1(n_134),
.B2(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_80),
.A2(n_82),
.B1(n_191),
.B2(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_80),
.A2(n_107),
.B(n_194),
.Y(n_223)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_81),
.A2(n_190),
.B1(n_192),
.B2(n_193),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_81),
.A2(n_84),
.B(n_133),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_85),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_89),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_112),
.B(n_114),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_99),
.C(n_100),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_95),
.B(n_99),
.Y(n_298)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_100),
.A2(n_101),
.B1(n_297),
.B2(n_298),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_101),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_110),
.C(n_115),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_102),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_108),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_103),
.B(n_108),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_107),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_104),
.A2(n_134),
.B(n_155),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_110),
.A2(n_111),
.B1(n_115),
.B2(n_116),
.Y(n_288)
);

CKINVDCx14_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_116),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_294),
.B(n_299),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_123),
.A2(n_282),
.B(n_293),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_SL g123 ( 
.A1(n_124),
.A2(n_182),
.B(n_261),
.C(n_281),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_167),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_125),
.B(n_167),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_150),
.B2(n_166),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_137),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_128),
.B(n_137),
.C(n_166),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_130),
.B1(n_135),
.B2(n_136),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_129),
.B(n_136),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_134),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_134),
.B(n_147),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_145),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_142),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_144),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_145),
.B(n_169),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_148),
.Y(n_159)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_150),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_156),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_151),
.B(n_157),
.C(n_162),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_152),
.B(n_154),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_156)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_165),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_168),
.B(n_258),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_170),
.A2(n_171),
.B1(n_172),
.B2(n_173),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_173),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_176),
.C(n_177),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_174),
.A2(n_175),
.B1(n_176),
.B2(n_249),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_177),
.B(n_248),
.Y(n_247)
);

CKINVDCx16_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_260),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_255),
.B(n_259),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_185),
.A2(n_243),
.B(n_254),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_225),
.B(n_242),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_214),
.B(n_224),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g187 ( 
.A1(n_188),
.A2(n_203),
.B(n_213),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_195),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_195),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g215 ( 
.A(n_197),
.B(n_199),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_208),
.B(n_212),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_206),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_210),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_216),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_216),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_218),
.B(n_221),
.C(n_223),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_227),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_233),
.B1(n_240),
.B2(n_241),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_228),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_230),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_229),
.B(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_233),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_236),
.B1(n_237),
.B2(n_239),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_234),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_236),
.B(n_239),
.C(n_240),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_237),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_245),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_244),
.B(n_245),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_246),
.A2(n_247),
.B1(n_250),
.B2(n_251),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_252),
.C(n_253),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g246 ( 
.A(n_247),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_253),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_256),
.B(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_262),
.B(n_263),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_279),
.B2(n_280),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_266),
.B(n_269),
.C(n_280),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_272),
.B2(n_278),
.Y(n_269)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_270),
.Y(n_278)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_276),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_273),
.B(n_276),
.C(n_278),
.Y(n_292)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_279),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_290),
.C(n_292),
.Y(n_295)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx14_ASAP7_75t_R g289 ( 
.A(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);


endmodule