module fake_jpeg_9832_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_37),
.Y(n_52)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_40),
.Y(n_53)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_17),
.Y(n_59)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_41),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_43),
.B(n_45),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_42),
.A2(n_16),
.B1(n_24),
.B2(n_21),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_49),
.B1(n_54),
.B2(n_55),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_36),
.B(n_31),
.C(n_29),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_47),
.B(n_18),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_16),
.B1(n_24),
.B2(n_21),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_42),
.A2(n_16),
.B1(n_24),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_63),
.B1(n_34),
.B2(n_40),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_24),
.B1(n_33),
.B2(n_21),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_33),
.B1(n_31),
.B2(n_17),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx11_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_59),
.Y(n_67)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_60),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_17),
.B1(n_25),
.B2(n_32),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_61),
.A2(n_26),
.B1(n_19),
.B2(n_27),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_30),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_26),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_30),
.B1(n_25),
.B2(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_25),
.Y(n_64)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_65),
.B(n_76),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_0),
.Y(n_66)
);

XNOR2xp5_ASAP7_75t_SL g102 ( 
.A(n_66),
.B(n_69),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_82),
.B1(n_87),
.B2(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_62),
.B(n_43),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_72),
.B(n_77),
.Y(n_107)
);

BUFx4f_ASAP7_75t_SL g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_75),
.B(n_36),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_56),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_28),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_45),
.A2(n_27),
.B1(n_19),
.B2(n_28),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_79),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_0),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_80),
.A2(n_18),
.B(n_22),
.Y(n_108)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_44),
.Y(n_81)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_81),
.Y(n_92)
);

INVx1_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g104 ( 
.A1(n_83),
.A2(n_86),
.B1(n_35),
.B2(n_48),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_64),
.B(n_36),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_58),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_56),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_39),
.B1(n_35),
.B2(n_23),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_67),
.B(n_63),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_89),
.B(n_91),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_52),
.Y(n_91)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_93),
.B(n_94),
.Y(n_129)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_72),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g95 ( 
.A(n_73),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_103),
.Y(n_123)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_69),
.A2(n_55),
.B(n_52),
.C(n_53),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_SL g124 ( 
.A(n_96),
.B(n_108),
.C(n_77),
.Y(n_124)
);

OA22x2_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_60),
.B1(n_51),
.B2(n_49),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_98),
.A2(n_111),
.B1(n_65),
.B2(n_81),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_100),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_101),
.A2(n_74),
.B1(n_70),
.B2(n_67),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_84),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_104),
.A2(n_73),
.B(n_58),
.Y(n_127)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_78),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_110),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_29),
.B(n_53),
.C(n_56),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_106),
.A2(n_71),
.B(n_66),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_109),
.B(n_71),
.C(n_83),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_85),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_70),
.A2(n_48),
.B1(n_51),
.B2(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_112),
.B(n_22),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_113),
.B(n_66),
.Y(n_119)
);

AO21x2_ASAP7_75t_L g114 ( 
.A1(n_111),
.A2(n_87),
.B(n_57),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_114),
.A2(n_96),
.B1(n_105),
.B2(n_92),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_115),
.A2(n_118),
.B1(n_131),
.B2(n_136),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_75),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_116),
.B(n_125),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_99),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_117),
.B(n_121),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_79),
.B1(n_68),
.B2(n_48),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_130),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_120),
.A2(n_122),
.B(n_92),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_113),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_94),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_124),
.A2(n_127),
.B(n_134),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_128),
.B(n_138),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_77),
.Y(n_130)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_106),
.B(n_18),
.CON(n_133),
.SN(n_133)
);

AO32x1_ASAP7_75t_L g153 ( 
.A1(n_133),
.A2(n_98),
.A3(n_108),
.B1(n_22),
.B2(n_29),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_107),
.B(n_57),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_139),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_90),
.A2(n_78),
.B1(n_58),
.B2(n_57),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_98),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_103),
.B(n_73),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_132),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_141),
.B(n_145),
.Y(n_169)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_91),
.Y(n_146)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_93),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_147),
.B(n_156),
.Y(n_172)
);

AND2x6_ASAP7_75t_L g148 ( 
.A(n_124),
.B(n_102),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_117),
.B(n_97),
.Y(n_151)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_151),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_152),
.A2(n_153),
.B(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_139),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_158),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_138),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_155),
.A2(n_126),
.B(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_123),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_137),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_157),
.Y(n_179)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_129),
.Y(n_158)
);

AND2x6_ASAP7_75t_L g159 ( 
.A(n_116),
.B(n_102),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_159),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_129),
.B(n_97),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_161),
.Y(n_174)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_136),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_127),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_100),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_134),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_165),
.A2(n_114),
.B1(n_22),
.B2(n_76),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_166),
.A2(n_114),
.B(n_22),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_125),
.C(n_119),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_171),
.C(n_180),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_142),
.B(n_120),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_176),
.A2(n_143),
.B(n_140),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_166),
.B(n_126),
.Y(n_180)
);

A2O1A1O1Ixp25_ASAP7_75t_L g181 ( 
.A1(n_150),
.A2(n_122),
.B(n_114),
.C(n_118),
.D(n_131),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_181),
.B(n_160),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_144),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_182),
.B(n_164),
.Y(n_200)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_183),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_149),
.B(n_114),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_190),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_186),
.A2(n_153),
.B(n_155),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_159),
.B(n_114),
.C(n_86),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_187),
.B(n_9),
.Y(n_211)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_157),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_188),
.B(n_156),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_163),
.A2(n_23),
.B1(n_20),
.B2(n_22),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g207 ( 
.A1(n_189),
.A2(n_23),
.B1(n_147),
.B2(n_146),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_23),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_188),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_191),
.B(n_194),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_175),
.Y(n_192)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g194 ( 
.A(n_179),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_195),
.B(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_186),
.A2(n_162),
.B1(n_141),
.B2(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_197),
.Y(n_225)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_200),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_180),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_201),
.A2(n_206),
.B1(n_208),
.B2(n_177),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_174),
.A2(n_165),
.B1(n_155),
.B2(n_152),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_202),
.A2(n_207),
.B1(n_209),
.B2(n_210),
.Y(n_224)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_169),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_203),
.B(n_172),
.Y(n_226)
);

OA21x2_ASAP7_75t_SL g204 ( 
.A1(n_171),
.A2(n_148),
.B(n_140),
.Y(n_204)
);

OAI21x1_ASAP7_75t_L g214 ( 
.A1(n_204),
.A2(n_168),
.B(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_185),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_181),
.A2(n_143),
.B1(n_2),
.B2(n_1),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_211),
.B(n_187),
.C(n_178),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_209),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_212),
.B(n_2),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_218),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_191),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_219),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_206),
.B1(n_205),
.B2(n_170),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_222),
.B1(n_199),
.B2(n_3),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_190),
.C(n_172),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_228),
.C(n_10),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_189),
.B1(n_177),
.B2(n_170),
.Y(n_222)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_226),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_193),
.B(n_185),
.C(n_173),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_225),
.B(n_210),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_229),
.B(n_239),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_224),
.A2(n_201),
.B1(n_211),
.B2(n_173),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_231),
.A2(n_232),
.B1(n_238),
.B2(n_223),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_212),
.A2(n_199),
.B1(n_195),
.B2(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_233),
.Y(n_246)
);

O2A1O1Ixp33_ASAP7_75t_L g245 ( 
.A1(n_234),
.A2(n_238),
.B(n_216),
.C(n_6),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_237),
.B(n_241),
.C(n_228),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_213),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_10),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_240),
.B(n_5),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_2),
.C(n_4),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_220),
.B(n_219),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_242),
.A2(n_231),
.B(n_230),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_236),
.B(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_243),
.B(n_247),
.Y(n_261)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_245),
.Y(n_253)
);

HB1xp67_ASAP7_75t_L g248 ( 
.A(n_241),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_248),
.B(n_5),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_249),
.B(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_237),
.B(n_218),
.C(n_223),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_9),
.C(n_10),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_251),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_5),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_254),
.A2(n_244),
.B(n_246),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_242),
.A2(n_230),
.B1(n_6),
.B2(n_8),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_255),
.B(n_259),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_256),
.A2(n_260),
.B(n_261),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_13),
.C(n_14),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_12),
.B(n_13),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_250),
.C(n_249),
.Y(n_262)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_262),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_263),
.A2(n_257),
.B1(n_258),
.B2(n_255),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_265),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_253),
.B(n_245),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_266),
.B(n_259),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_268),
.B(n_267),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_270),
.B(n_13),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_273),
.B(n_271),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_274),
.A2(n_269),
.B(n_270),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_14),
.B(n_15),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_15),
.Y(n_277)
);


endmodule