module fake_jpeg_12749_n_202 (n_13, n_21, n_53, n_33, n_54, n_1, n_45, n_10, n_23, n_27, n_55, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_56, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_202);

input n_13;
input n_21;
input n_53;
input n_33;
input n_54;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_55;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_56;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_202;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_182;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_51),
.Y(n_57)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_29),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_43),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_45),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_18),
.Y(n_62)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_37),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_49),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_50),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_36),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_33),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_32),
.Y(n_73)
);

BUFx12_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

BUFx5_ASAP7_75t_L g75 ( 
.A(n_9),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_14),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_0),
.Y(n_78)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_25),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_0),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_14),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_2),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_78),
.B(n_1),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_87),
.B(n_88),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_19),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_SL g90 ( 
.A(n_61),
.Y(n_90)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_84),
.B(n_1),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_92),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_93),
.Y(n_102)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_79),
.Y(n_95)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_95),
.Y(n_101)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_92),
.Y(n_97)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_97),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_88),
.A2(n_58),
.B(n_66),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_100),
.A2(n_75),
.B(n_74),
.C(n_4),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_96),
.A2(n_77),
.B1(n_73),
.B2(n_66),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_63),
.B1(n_76),
.B2(n_72),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_95),
.A2(n_79),
.B1(n_58),
.B2(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_105),
.A2(n_110),
.B1(n_75),
.B2(n_74),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_70),
.Y(n_107)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_94),
.Y(n_109)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_90),
.A2(n_85),
.B1(n_73),
.B2(n_77),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_110),
.A2(n_90),
.B1(n_93),
.B2(n_65),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_113),
.A2(n_134),
.B1(n_120),
.B2(n_133),
.Y(n_156)
);

BUFx8_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_114),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_98),
.B(n_68),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_115),
.B(n_118),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_116),
.A2(n_129),
.B1(n_133),
.B2(n_6),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_82),
.B1(n_57),
.B2(n_80),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_119),
.B1(n_3),
.B2(n_5),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_108),
.B(n_81),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_120),
.B(n_3),
.Y(n_136)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_103),
.B(n_26),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g135 ( 
.A(n_121),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_101),
.B(n_59),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_126),
.Y(n_155)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_112),
.Y(n_125)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_60),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_112),
.Y(n_127)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_127),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_97),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_128),
.B(n_131),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_99),
.A2(n_71),
.B1(n_69),
.B2(n_67),
.Y(n_129)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_99),
.Y(n_130)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_130),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_64),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_102),
.B(n_2),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_132),
.B(n_23),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_105),
.A2(n_74),
.B1(n_4),
.B2(n_5),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_136),
.A2(n_145),
.B(n_11),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g137 ( 
.A(n_121),
.B(n_22),
.C(n_53),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_114),
.C(n_10),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_140),
.A2(n_156),
.B1(n_9),
.B2(n_10),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_142),
.B(n_146),
.Y(n_163)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_56),
.Y(n_144)
);

A2O1A1O1Ixp25_ASAP7_75t_L g167 ( 
.A1(n_144),
.A2(n_15),
.B(n_52),
.C(n_21),
.D(n_24),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_116),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_7),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_148),
.B(n_154),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_119),
.B(n_8),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_149),
.B(n_17),
.Y(n_169)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_129),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_157),
.B(n_167),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_168),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_160)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_165),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_145),
.B(n_147),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_135),
.B(n_12),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_170),
.C(n_163),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_156),
.A2(n_13),
.B1(n_15),
.B2(n_16),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_139),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g178 ( 
.A1(n_169),
.A2(n_170),
.B(n_137),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_31),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_172),
.Y(n_175)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_136),
.B(n_141),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_178),
.B(n_182),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_158),
.Y(n_180)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_180),
.Y(n_189)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_181),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_183),
.A2(n_171),
.B1(n_164),
.B2(n_151),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_171),
.C(n_151),
.Y(n_188)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_176),
.A2(n_167),
.A3(n_152),
.B1(n_143),
.B2(n_44),
.C1(n_46),
.C2(n_35),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_190),
.A2(n_184),
.B1(n_179),
.B2(n_182),
.Y(n_193)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_186),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_194),
.A2(n_192),
.B(n_189),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_188),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_196),
.A2(n_174),
.B(n_191),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_197),
.B(n_191),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_187),
.B1(n_177),
.B2(n_152),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_199),
.A2(n_187),
.B1(n_184),
.B2(n_48),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_38),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_40),
.Y(n_202)
);


endmodule