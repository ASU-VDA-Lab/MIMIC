module fake_netlist_5_968_n_1810 (n_137, n_210, n_168, n_260, n_164, n_191, n_286, n_91, n_208, n_82, n_122, n_194, n_282, n_142, n_176, n_10, n_214, n_140, n_24, n_248, n_124, n_86, n_136, n_146, n_268, n_182, n_143, n_83, n_132, n_61, n_237, n_90, n_241, n_127, n_75, n_101, n_180, n_184, n_226, n_235, n_65, n_78, n_74, n_144, n_281, n_207, n_240, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_229, n_108, n_231, n_257, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_236, n_18, n_116, n_195, n_42, n_22, n_227, n_1, n_45, n_117, n_249, n_271, n_284, n_46, n_233, n_21, n_94, n_203, n_245, n_274, n_205, n_113, n_38, n_123, n_139, n_105, n_280, n_246, n_80, n_4, n_179, n_125, n_35, n_269, n_167, n_128, n_73, n_234, n_277, n_17, n_92, n_19, n_267, n_149, n_120, n_285, n_232, n_135, n_30, n_156, n_5, n_33, n_126, n_254, n_14, n_225, n_84, n_23, n_202, n_130, n_266, n_272, n_219, n_157, n_258, n_265, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_244, n_251, n_25, n_53, n_160, n_198, n_223, n_288, n_247, n_188, n_190, n_8, n_201, n_158, n_263, n_44, n_224, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_228, n_264, n_283, n_109, n_112, n_212, n_85, n_159, n_163, n_276, n_95, n_119, n_183, n_185, n_243, n_239, n_275, n_175, n_252, n_169, n_59, n_262, n_26, n_255, n_133, n_238, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_242, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_259, n_273, n_287, n_270, n_222, n_230, n_81, n_118, n_28, n_89, n_279, n_70, n_115, n_68, n_93, n_253, n_261, n_72, n_174, n_186, n_199, n_289, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_256, n_48, n_204, n_50, n_250, n_52, n_278, n_88, n_110, n_216, n_1810);

input n_137;
input n_210;
input n_168;
input n_260;
input n_164;
input n_191;
input n_286;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_282;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_268;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_237;
input n_90;
input n_241;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_226;
input n_235;
input n_65;
input n_78;
input n_74;
input n_144;
input n_281;
input n_207;
input n_240;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_229;
input n_108;
input n_231;
input n_257;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_236;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_227;
input n_1;
input n_45;
input n_117;
input n_249;
input n_271;
input n_284;
input n_46;
input n_233;
input n_21;
input n_94;
input n_203;
input n_245;
input n_274;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_280;
input n_246;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_269;
input n_167;
input n_128;
input n_73;
input n_234;
input n_277;
input n_17;
input n_92;
input n_19;
input n_267;
input n_149;
input n_120;
input n_285;
input n_232;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_254;
input n_14;
input n_225;
input n_84;
input n_23;
input n_202;
input n_130;
input n_266;
input n_272;
input n_219;
input n_157;
input n_258;
input n_265;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_244;
input n_251;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_288;
input n_247;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_228;
input n_264;
input n_283;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_276;
input n_95;
input n_119;
input n_183;
input n_185;
input n_243;
input n_239;
input n_275;
input n_175;
input n_252;
input n_169;
input n_59;
input n_262;
input n_26;
input n_255;
input n_133;
input n_238;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_242;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_259;
input n_273;
input n_287;
input n_270;
input n_222;
input n_230;
input n_81;
input n_118;
input n_28;
input n_89;
input n_279;
input n_70;
input n_115;
input n_68;
input n_93;
input n_253;
input n_261;
input n_72;
input n_174;
input n_186;
input n_199;
input n_289;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_256;
input n_48;
input n_204;
input n_50;
input n_250;
input n_52;
input n_278;
input n_88;
input n_110;
input n_216;

output n_1810;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1677;
wire n_1150;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1607;
wire n_1563;
wire n_606;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_929;
wire n_1124;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_291;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_1598;
wire n_1723;
wire n_955;
wire n_339;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1565;
wire n_1809;
wire n_647;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_1538;
wire n_1162;
wire n_1199;
wire n_1779;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1660;
wire n_887;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1710;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1614;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_1551;
wire n_545;
wire n_860;
wire n_441;
wire n_450;
wire n_1805;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1205;
wire n_1044;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_1553;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_1307;
wire n_988;
wire n_814;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_770;
wire n_458;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_707;
wire n_1168;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1440;
wire n_421;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1313;
wire n_1136;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1747;
wire n_714;
wire n_1683;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1792;
wire n_1564;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_934;
wire n_1618;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1619;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_1739;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_187),
.Y(n_290)
);

BUFx2_ASAP7_75t_SL g291 ( 
.A(n_136),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_253),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_90),
.Y(n_293)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_107),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_62),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_155),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_252),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_204),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_192),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_41),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_173),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_287),
.Y(n_302)
);

BUFx3_ASAP7_75t_L g303 ( 
.A(n_249),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_72),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_67),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_273),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_5),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_146),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_271),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_14),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_169),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_123),
.Y(n_313)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_103),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_89),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_158),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_183),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_130),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_23),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_17),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_120),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_266),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_34),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_214),
.Y(n_325)
);

BUFx2_ASAP7_75t_L g326 ( 
.A(n_244),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_91),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_64),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_129),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_106),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_228),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_145),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_94),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_113),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_65),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_156),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_213),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_236),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_161),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_251),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_256),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g342 ( 
.A(n_53),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_93),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_229),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_261),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_223),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_152),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_190),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_198),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_85),
.Y(n_350)
);

BUFx2_ASAP7_75t_SL g351 ( 
.A(n_61),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_235),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_246),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_80),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g355 ( 
.A(n_112),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_245),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_2),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_33),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_224),
.Y(n_360)
);

BUFx2_ASAP7_75t_SL g361 ( 
.A(n_79),
.Y(n_361)
);

BUFx5_ASAP7_75t_L g362 ( 
.A(n_92),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_50),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_47),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_176),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_149),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_134),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_260),
.Y(n_368)
);

BUFx5_ASAP7_75t_L g369 ( 
.A(n_191),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_241),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_128),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_248),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_95),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_65),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_185),
.Y(n_375)
);

BUFx3_ASAP7_75t_L g376 ( 
.A(n_8),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_186),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_232),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_280),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_62),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g381 ( 
.A(n_227),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_53),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_0),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_68),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_147),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_121),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_270),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_288),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_284),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_70),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_164),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_219),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_3),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_60),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_76),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_1),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_200),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_255),
.Y(n_398)
);

CKINVDCx5p33_ASAP7_75t_R g399 ( 
.A(n_19),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_80),
.Y(n_400)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_184),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_172),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_182),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_265),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_197),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_166),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_49),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_85),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_139),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_0),
.Y(n_410)
);

BUFx8_ASAP7_75t_SL g411 ( 
.A(n_58),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_37),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_268),
.Y(n_413)
);

CKINVDCx16_ASAP7_75t_R g414 ( 
.A(n_199),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_48),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_272),
.Y(n_416)
);

INVxp67_ASAP7_75t_SL g417 ( 
.A(n_151),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_82),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_10),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_3),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_215),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_88),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_56),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_100),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_119),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_148),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_159),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_278),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_234),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_276),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g431 ( 
.A(n_140),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_76),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_133),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_17),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_231),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_63),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_1),
.Y(n_437)
);

BUFx2_ASAP7_75t_L g438 ( 
.A(n_179),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_99),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_194),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_240),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_180),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_54),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_258),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_201),
.Y(n_445)
);

HB1xp67_ASAP7_75t_L g446 ( 
.A(n_289),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_207),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_78),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_142),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_8),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_7),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_32),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_277),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_243),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_208),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_114),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_44),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_49),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_195),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_73),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_45),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_41),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_97),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_218),
.Y(n_464)
);

INVx1_ASAP7_75t_SL g465 ( 
.A(n_36),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_22),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_13),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_286),
.Y(n_468)
);

CKINVDCx5p33_ASAP7_75t_R g469 ( 
.A(n_174),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_89),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_144),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_154),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_84),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_32),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_84),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_6),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g477 ( 
.A(n_329),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_411),
.Y(n_478)
);

CKINVDCx16_ASAP7_75t_R g479 ( 
.A(n_314),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_411),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_326),
.B(n_2),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_295),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_329),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_308),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_376),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_376),
.Y(n_486)
);

INVxp67_ASAP7_75t_SL g487 ( 
.A(n_446),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_467),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_381),
.B(n_4),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_438),
.B(n_4),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_304),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_333),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_304),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_319),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_321),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_304),
.Y(n_497)
);

INVxp67_ASAP7_75t_SL g498 ( 
.A(n_303),
.Y(n_498)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_333),
.Y(n_499)
);

BUFx2_ASAP7_75t_L g500 ( 
.A(n_305),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_304),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_R g502 ( 
.A(n_302),
.B(n_5),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_328),
.Y(n_503)
);

BUFx3_ASAP7_75t_L g504 ( 
.A(n_303),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_371),
.Y(n_505)
);

HB1xp67_ASAP7_75t_L g506 ( 
.A(n_305),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_371),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_294),
.B(n_6),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_290),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_372),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_350),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_372),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_405),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_342),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_342),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_354),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_342),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g518 ( 
.A(n_467),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_357),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_342),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_405),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_380),
.Y(n_522)
);

CKINVDCx5p33_ASAP7_75t_R g523 ( 
.A(n_358),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_363),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_380),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_309),
.B(n_7),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_364),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g528 ( 
.A(n_467),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_380),
.Y(n_529)
);

INVxp33_ASAP7_75t_SL g530 ( 
.A(n_390),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_380),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_410),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g533 ( 
.A(n_300),
.B(n_9),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_410),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_410),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_410),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_432),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_435),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_432),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_432),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_374),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_394),
.Y(n_542)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_432),
.Y(n_543)
);

CKINVDCx16_ASAP7_75t_R g544 ( 
.A(n_414),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_395),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_435),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_396),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_306),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_355),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_320),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_399),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_390),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_324),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_407),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_355),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_335),
.Y(n_556)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_292),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_408),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_382),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_453),
.B(n_9),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_383),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_431),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_418),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_294),
.B(n_10),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_498),
.B(n_302),
.Y(n_565)
);

INVxp67_ASAP7_75t_L g566 ( 
.A(n_506),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_492),
.B(n_336),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_494),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_SL g569 ( 
.A(n_478),
.B(n_11),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_497),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_501),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_504),
.B(n_336),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_562),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_488),
.A2(n_311),
.B1(n_436),
.B2(n_315),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_562),
.Y(n_575)
);

OA21x2_ASAP7_75t_L g576 ( 
.A1(n_549),
.A2(n_450),
.B(n_359),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_562),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_562),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_514),
.Y(n_579)
);

OAI22xp5_ASAP7_75t_L g580 ( 
.A1(n_481),
.A2(n_311),
.B1(n_436),
.B2(n_315),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_515),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_517),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_520),
.B(n_307),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_522),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_529),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_562),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_531),
.Y(n_588)
);

INVx3_ASAP7_75t_L g589 ( 
.A(n_549),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_534),
.Y(n_591)
);

XNOR2xp5_ASAP7_75t_L g592 ( 
.A(n_477),
.B(n_461),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_535),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_555),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_555),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_482),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_536),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_537),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_539),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_540),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_543),
.B(n_307),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_548),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_550),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_553),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_564),
.B(n_403),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_556),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_508),
.Y(n_607)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_559),
.Y(n_608)
);

INVx3_ASAP7_75t_L g609 ( 
.A(n_561),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_563),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_504),
.B(n_403),
.Y(n_611)
);

INVx3_ASAP7_75t_L g612 ( 
.A(n_533),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_485),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_486),
.B(n_293),
.Y(n_614)
);

AND2x2_ASAP7_75t_L g615 ( 
.A(n_487),
.B(n_332),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_490),
.B(n_296),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_560),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_526),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_491),
.Y(n_619)
);

AND2x6_ASAP7_75t_L g620 ( 
.A(n_489),
.B(n_332),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_509),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_552),
.B(n_334),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_500),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_518),
.B(n_334),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_482),
.Y(n_625)
);

INVx3_ASAP7_75t_L g626 ( 
.A(n_484),
.Y(n_626)
);

NAND2xp5_ASAP7_75t_L g627 ( 
.A(n_484),
.B(n_297),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_495),
.Y(n_628)
);

INVx3_ASAP7_75t_L g629 ( 
.A(n_495),
.Y(n_629)
);

BUFx6f_ASAP7_75t_L g630 ( 
.A(n_496),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_496),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g632 ( 
.A(n_530),
.B(n_310),
.Y(n_632)
);

BUFx8_ASAP7_75t_L g633 ( 
.A(n_479),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_503),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_528),
.B(n_401),
.Y(n_635)
);

BUFx3_ASAP7_75t_L g636 ( 
.A(n_576),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_576),
.Y(n_637)
);

INVx4_ASAP7_75t_L g638 ( 
.A(n_576),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_576),
.Y(n_639)
);

BUFx3_ASAP7_75t_L g640 ( 
.A(n_576),
.Y(n_640)
);

INVx3_ASAP7_75t_L g641 ( 
.A(n_576),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_609),
.Y(n_642)
);

NOR2x1p5_ASAP7_75t_L g643 ( 
.A(n_621),
.B(n_478),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_619),
.B(n_503),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_567),
.B(n_619),
.Y(n_645)
);

INVx3_ASAP7_75t_L g646 ( 
.A(n_589),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_567),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_589),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_SL g649 ( 
.A(n_632),
.B(n_544),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_598),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_567),
.B(n_417),
.Y(n_651)
);

INVx1_ASAP7_75t_SL g652 ( 
.A(n_592),
.Y(n_652)
);

INVx4_ASAP7_75t_L g653 ( 
.A(n_598),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_609),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_616),
.B(n_530),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_609),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_598),
.Y(n_657)
);

NAND2xp33_ASAP7_75t_L g658 ( 
.A(n_630),
.B(n_511),
.Y(n_658)
);

INVx4_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

AND2x6_ASAP7_75t_L g660 ( 
.A(n_607),
.B(n_401),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_594),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_598),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_619),
.B(n_511),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_609),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_619),
.B(n_516),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_567),
.Y(n_666)
);

INVxp33_ASAP7_75t_L g667 ( 
.A(n_592),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_594),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_616),
.B(n_557),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_609),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_594),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_618),
.B(n_516),
.Y(n_672)
);

INVx5_ASAP7_75t_L g673 ( 
.A(n_589),
.Y(n_673)
);

INVxp67_ASAP7_75t_L g674 ( 
.A(n_632),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_594),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_595),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_567),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_618),
.B(n_519),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_572),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_595),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_595),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_595),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_618),
.B(n_519),
.Y(n_683)
);

AND2x6_ASAP7_75t_L g684 ( 
.A(n_607),
.B(n_431),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_627),
.B(n_523),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_589),
.Y(n_686)
);

BUFx3_ASAP7_75t_L g687 ( 
.A(n_607),
.Y(n_687)
);

INVx4_ASAP7_75t_L g688 ( 
.A(n_598),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_627),
.B(n_523),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_589),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_568),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_618),
.B(n_524),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_568),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_573),
.Y(n_694)
);

AND2x4_ASAP7_75t_L g695 ( 
.A(n_572),
.B(n_298),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_572),
.B(n_316),
.Y(n_696)
);

OR2x2_ASAP7_75t_L g697 ( 
.A(n_623),
.B(n_524),
.Y(n_697)
);

AND2x4_ASAP7_75t_L g698 ( 
.A(n_612),
.B(n_317),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_630),
.B(n_527),
.Y(n_699)
);

NOR2x1p5_ASAP7_75t_L g700 ( 
.A(n_621),
.B(n_480),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_645),
.Y(n_701)
);

AO22x2_ASAP7_75t_L g702 ( 
.A1(n_674),
.A2(n_580),
.B1(n_574),
.B2(n_617),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_645),
.B(n_607),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_645),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_645),
.Y(n_705)
);

AO22x2_ASAP7_75t_L g706 ( 
.A1(n_649),
.A2(n_580),
.B1(n_574),
.B2(n_617),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_666),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_691),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_691),
.Y(n_709)
);

AO22x2_ASAP7_75t_L g710 ( 
.A1(n_652),
.A2(n_623),
.B1(n_634),
.B2(n_631),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_655),
.Y(n_711)
);

AO22x2_ASAP7_75t_L g712 ( 
.A1(n_697),
.A2(n_623),
.B1(n_634),
.B2(n_631),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_693),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_679),
.B(n_612),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_679),
.B(n_612),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_693),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_697),
.B(n_623),
.Y(n_717)
);

OAI22xp5_ASAP7_75t_L g718 ( 
.A1(n_672),
.A2(n_612),
.B1(n_625),
.B2(n_628),
.Y(n_718)
);

INVxp67_ASAP7_75t_L g719 ( 
.A(n_669),
.Y(n_719)
);

AO22x2_ASAP7_75t_L g720 ( 
.A1(n_678),
.A2(n_566),
.B1(n_569),
.B2(n_361),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_644),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_647),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_647),
.B(n_612),
.Y(n_723)
);

BUFx2_ASAP7_75t_L g724 ( 
.A(n_663),
.Y(n_724)
);

AO22x2_ASAP7_75t_L g725 ( 
.A1(n_683),
.A2(n_566),
.B1(n_569),
.B2(n_351),
.Y(n_725)
);

AND2x4_ASAP7_75t_L g726 ( 
.A(n_666),
.B(n_621),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_666),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_677),
.Y(n_728)
);

AND2x4_ASAP7_75t_L g729 ( 
.A(n_677),
.B(n_621),
.Y(n_729)
);

NAND2x1p5_ASAP7_75t_L g730 ( 
.A(n_677),
.B(n_621),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_685),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_689),
.B(n_630),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_692),
.B(n_625),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_642),
.Y(n_734)
);

AND2x4_ASAP7_75t_L g735 ( 
.A(n_695),
.B(n_625),
.Y(n_735)
);

NAND2x1p5_ASAP7_75t_L g736 ( 
.A(n_687),
.B(n_626),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_642),
.Y(n_737)
);

OAI221xp5_ASAP7_75t_L g738 ( 
.A1(n_665),
.A2(n_605),
.B1(n_393),
.B2(n_615),
.C(n_466),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_654),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_654),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_656),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_656),
.Y(n_742)
);

AND2x4_ASAP7_75t_L g743 ( 
.A(n_695),
.B(n_625),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_664),
.Y(n_744)
);

AO22x2_ASAP7_75t_L g745 ( 
.A1(n_698),
.A2(n_569),
.B1(n_400),
.B2(n_465),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_661),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_664),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_643),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_670),
.Y(n_749)
);

AO22x2_ASAP7_75t_L g750 ( 
.A1(n_698),
.A2(n_628),
.B1(n_622),
.B2(n_450),
.Y(n_750)
);

INVxp67_ASAP7_75t_L g751 ( 
.A(n_695),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_687),
.B(n_607),
.Y(n_752)
);

NOR2xp33_ASAP7_75t_L g753 ( 
.A(n_699),
.B(n_628),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_687),
.B(n_607),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_661),
.Y(n_755)
);

OR2x2_ASAP7_75t_SL g756 ( 
.A(n_667),
.B(n_630),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_698),
.B(n_607),
.Y(n_757)
);

BUFx8_ASAP7_75t_L g758 ( 
.A(n_695),
.Y(n_758)
);

BUFx8_ASAP7_75t_L g759 ( 
.A(n_696),
.Y(n_759)
);

AO22x2_ASAP7_75t_L g760 ( 
.A1(n_698),
.A2(n_622),
.B1(n_359),
.B2(n_626),
.Y(n_760)
);

AO22x2_ASAP7_75t_L g761 ( 
.A1(n_696),
.A2(n_622),
.B1(n_629),
.B2(n_626),
.Y(n_761)
);

AOI22xp33_ASAP7_75t_L g762 ( 
.A1(n_638),
.A2(n_607),
.B1(n_620),
.B2(n_605),
.Y(n_762)
);

CKINVDCx14_ASAP7_75t_R g763 ( 
.A(n_696),
.Y(n_763)
);

AND2x4_ASAP7_75t_L g764 ( 
.A(n_696),
.B(n_643),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_670),
.Y(n_765)
);

AO22x2_ASAP7_75t_L g766 ( 
.A1(n_639),
.A2(n_629),
.B1(n_626),
.B2(n_624),
.Y(n_766)
);

HB1xp67_ASAP7_75t_L g767 ( 
.A(n_700),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_700),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_646),
.Y(n_769)
);

AO22x2_ASAP7_75t_L g770 ( 
.A1(n_639),
.A2(n_629),
.B1(n_626),
.B2(n_624),
.Y(n_770)
);

OAI221xp5_ASAP7_75t_L g771 ( 
.A1(n_658),
.A2(n_615),
.B1(n_565),
.B2(n_614),
.C(n_601),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_646),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_651),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_646),
.Y(n_774)
);

CKINVDCx20_ASAP7_75t_R g775 ( 
.A(n_636),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_646),
.Y(n_776)
);

NAND3xp33_ASAP7_75t_L g777 ( 
.A(n_651),
.B(n_565),
.C(n_611),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_668),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_686),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_636),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_SL g781 ( 
.A(n_651),
.B(n_630),
.Y(n_781)
);

AO22x2_ASAP7_75t_L g782 ( 
.A1(n_638),
.A2(n_629),
.B1(n_635),
.B2(n_624),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_636),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_640),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_651),
.Y(n_785)
);

HB1xp67_ASAP7_75t_L g786 ( 
.A(n_640),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_640),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_731),
.B(n_630),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_711),
.B(n_630),
.Y(n_789)
);

NAND2xp5_ASAP7_75t_SL g790 ( 
.A(n_735),
.B(n_743),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_785),
.B(n_630),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_733),
.B(n_629),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_SL g793 ( 
.A(n_735),
.B(n_638),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_714),
.B(n_638),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_719),
.B(n_483),
.Y(n_795)
);

AND2x2_ASAP7_75t_SL g796 ( 
.A(n_753),
.B(n_431),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_SL g797 ( 
.A(n_724),
.B(n_596),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_SL g798 ( 
.A(n_743),
.B(n_596),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_721),
.B(n_596),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_726),
.B(n_633),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_726),
.B(n_633),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_729),
.B(n_633),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_729),
.B(n_633),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_714),
.B(n_633),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_717),
.B(n_635),
.Y(n_805)
);

AND2x4_ASAP7_75t_L g806 ( 
.A(n_764),
.B(n_613),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_715),
.B(n_611),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_715),
.B(n_723),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_723),
.B(n_614),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_718),
.B(n_637),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_764),
.B(n_615),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_707),
.B(n_493),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_707),
.B(n_499),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_701),
.B(n_505),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_701),
.B(n_507),
.Y(n_815)
);

NAND2xp5_ASAP7_75t_L g816 ( 
.A(n_708),
.B(n_637),
.Y(n_816)
);

NAND2xp33_ASAP7_75t_SL g817 ( 
.A(n_768),
.B(n_510),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_704),
.B(n_512),
.Y(n_818)
);

NAND2xp33_ASAP7_75t_R g819 ( 
.A(n_748),
.B(n_480),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_712),
.B(n_635),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_704),
.B(n_513),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_705),
.B(n_521),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_705),
.B(n_538),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_SL g824 ( 
.A(n_777),
.B(n_546),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_773),
.B(n_583),
.Y(n_825)
);

NAND2xp33_ASAP7_75t_SL g826 ( 
.A(n_775),
.B(n_767),
.Y(n_826)
);

NAND2xp33_ASAP7_75t_SL g827 ( 
.A(n_732),
.B(n_709),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_SL g828 ( 
.A(n_751),
.B(n_583),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_713),
.B(n_637),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_716),
.B(n_722),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_727),
.B(n_613),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_SL g832 ( 
.A(n_728),
.B(n_601),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_781),
.B(n_527),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_SL g834 ( 
.A(n_780),
.B(n_541),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_786),
.B(n_637),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_780),
.B(n_641),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_783),
.B(n_784),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_783),
.B(n_641),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_784),
.B(n_541),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_787),
.B(n_542),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_712),
.B(n_542),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_787),
.B(n_545),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_SL g843 ( 
.A(n_730),
.B(n_545),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_703),
.B(n_547),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_762),
.B(n_641),
.Y(n_845)
);

AND2x4_ASAP7_75t_L g846 ( 
.A(n_769),
.B(n_641),
.Y(n_846)
);

NAND2xp33_ASAP7_75t_SL g847 ( 
.A(n_757),
.B(n_461),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_750),
.B(n_620),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_758),
.B(n_547),
.Y(n_849)
);

NOR2xp33_ASAP7_75t_L g850 ( 
.A(n_738),
.B(n_592),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_SL g851 ( 
.A(n_758),
.B(n_551),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_SL g852 ( 
.A(n_734),
.B(n_473),
.Y(n_852)
);

NAND2xp33_ASAP7_75t_SL g853 ( 
.A(n_737),
.B(n_473),
.Y(n_853)
);

NAND2xp33_ASAP7_75t_SL g854 ( 
.A(n_739),
.B(n_502),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_759),
.B(n_551),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_710),
.B(n_554),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_710),
.B(n_554),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_759),
.B(n_558),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_736),
.B(n_558),
.Y(n_859)
);

AND2x2_ASAP7_75t_L g860 ( 
.A(n_706),
.B(n_602),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_SL g861 ( 
.A(n_772),
.B(n_312),
.Y(n_861)
);

NAND2xp33_ASAP7_75t_SL g862 ( 
.A(n_740),
.B(n_299),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_706),
.B(n_602),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_774),
.B(n_330),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_776),
.B(n_301),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_741),
.B(n_603),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_752),
.B(n_686),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_754),
.B(n_313),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_SL g869 ( 
.A(n_742),
.B(n_744),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_750),
.B(n_620),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_SL g871 ( 
.A(n_747),
.B(n_318),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_SL g872 ( 
.A(n_749),
.B(n_322),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_765),
.B(n_620),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_779),
.B(n_327),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_SL g875 ( 
.A(n_746),
.B(n_331),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_760),
.B(n_620),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_SL g877 ( 
.A(n_756),
.B(n_337),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_763),
.B(n_412),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_755),
.B(n_339),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_782),
.B(n_620),
.Y(n_880)
);

NAND2xp33_ASAP7_75t_SL g881 ( 
.A(n_745),
.B(n_343),
.Y(n_881)
);

NAND2xp33_ASAP7_75t_SL g882 ( 
.A(n_745),
.B(n_344),
.Y(n_882)
);

NAND2xp33_ASAP7_75t_SL g883 ( 
.A(n_778),
.B(n_346),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_761),
.B(n_347),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_761),
.B(n_348),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_782),
.B(n_620),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_850),
.A2(n_771),
.B(n_323),
.C(n_338),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_866),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_795),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_SL g890 ( 
.A(n_796),
.B(n_620),
.Y(n_890)
);

OAI21x1_ASAP7_75t_L g891 ( 
.A1(n_867),
.A2(n_694),
.B(n_690),
.Y(n_891)
);

INVxp67_ASAP7_75t_L g892 ( 
.A(n_799),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_810),
.A2(n_845),
.B(n_880),
.Y(n_893)
);

OA21x2_ASAP7_75t_L g894 ( 
.A1(n_886),
.A2(n_690),
.B(n_694),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_816),
.A2(n_675),
.B(n_671),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_846),
.Y(n_896)
);

INVx2_ASAP7_75t_L g897 ( 
.A(n_846),
.Y(n_897)
);

OAI21xp5_ASAP7_75t_L g898 ( 
.A1(n_829),
.A2(n_675),
.B(n_671),
.Y(n_898)
);

OA22x2_ASAP7_75t_L g899 ( 
.A1(n_856),
.A2(n_702),
.B1(n_725),
.B2(n_720),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_866),
.Y(n_900)
);

AND2x2_ASAP7_75t_L g901 ( 
.A(n_805),
.B(n_857),
.Y(n_901)
);

OAI21x1_ASAP7_75t_L g902 ( 
.A1(n_867),
.A2(n_680),
.B(n_676),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_796),
.A2(n_702),
.B1(n_770),
.B2(n_766),
.Y(n_903)
);

AOI21xp5_ASAP7_75t_L g904 ( 
.A1(n_794),
.A2(n_657),
.B(n_653),
.Y(n_904)
);

OAI21x1_ASAP7_75t_L g905 ( 
.A1(n_873),
.A2(n_838),
.B(n_836),
.Y(n_905)
);

OAI21x1_ASAP7_75t_L g906 ( 
.A1(n_837),
.A2(n_680),
.B(n_676),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_792),
.B(n_766),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_866),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_860),
.B(n_770),
.Y(n_909)
);

O2A1O1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_824),
.A2(n_340),
.B(n_341),
.C(n_325),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_863),
.B(n_620),
.Y(n_911)
);

BUFx10_ASAP7_75t_L g912 ( 
.A(n_878),
.Y(n_912)
);

AND2x4_ASAP7_75t_L g913 ( 
.A(n_806),
.B(n_603),
.Y(n_913)
);

A2O1A1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_847),
.A2(n_345),
.B(n_356),
.C(n_353),
.Y(n_914)
);

AOI211x1_ASAP7_75t_L g915 ( 
.A1(n_820),
.A2(n_443),
.B(n_448),
.C(n_419),
.Y(n_915)
);

NOR2xp67_ASAP7_75t_L g916 ( 
.A(n_797),
.B(n_606),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_854),
.A2(n_360),
.B(n_366),
.C(n_365),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_831),
.Y(n_918)
);

NAND3xp33_ASAP7_75t_SL g919 ( 
.A(n_852),
.B(n_475),
.C(n_420),
.Y(n_919)
);

AND2x4_ASAP7_75t_L g920 ( 
.A(n_806),
.B(n_606),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_819),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_806),
.Y(n_922)
);

OA21x2_ASAP7_75t_L g923 ( 
.A1(n_848),
.A2(n_870),
.B(n_876),
.Y(n_923)
);

OAI21xp5_ASAP7_75t_L g924 ( 
.A1(n_793),
.A2(n_660),
.B(n_668),
.Y(n_924)
);

OAI21x1_ASAP7_75t_L g925 ( 
.A1(n_869),
.A2(n_682),
.B(n_681),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_831),
.Y(n_926)
);

HB1xp67_ASAP7_75t_L g927 ( 
.A(n_812),
.Y(n_927)
);

OAI22xp5_ASAP7_75t_L g928 ( 
.A1(n_790),
.A2(n_725),
.B1(n_720),
.B2(n_452),
.Y(n_928)
);

AO21x1_ASAP7_75t_L g929 ( 
.A1(n_827),
.A2(n_387),
.B(n_373),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_846),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_793),
.A2(n_657),
.B(n_653),
.Y(n_931)
);

OR2x2_ASAP7_75t_SL g932 ( 
.A(n_817),
.B(n_451),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_835),
.A2(n_657),
.B(n_653),
.Y(n_933)
);

O2A1O1Ixp5_ASAP7_75t_L g934 ( 
.A1(n_788),
.A2(n_389),
.B(n_421),
.C(n_409),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_807),
.B(n_684),
.Y(n_935)
);

OAI21x1_ASAP7_75t_L g936 ( 
.A1(n_830),
.A2(n_575),
.B(n_573),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_831),
.Y(n_937)
);

AOI211x1_ASAP7_75t_L g938 ( 
.A1(n_811),
.A2(n_462),
.B(n_460),
.C(n_427),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_SL g939 ( 
.A1(n_790),
.A2(n_657),
.B(n_653),
.Y(n_939)
);

AOI31xp33_ASAP7_75t_L g940 ( 
.A1(n_804),
.A2(n_475),
.A3(n_422),
.B(n_423),
.Y(n_940)
);

AO31x2_ASAP7_75t_L g941 ( 
.A1(n_884),
.A2(n_430),
.A3(n_433),
.B(n_424),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_813),
.B(n_608),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_808),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_809),
.A2(n_662),
.B(n_659),
.Y(n_944)
);

AO32x2_ASAP7_75t_L g945 ( 
.A1(n_885),
.A2(n_688),
.A3(n_662),
.B1(n_659),
.B2(n_660),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_832),
.Y(n_946)
);

OAI21x1_ASAP7_75t_L g947 ( 
.A1(n_868),
.A2(n_575),
.B(n_573),
.Y(n_947)
);

INVx5_ASAP7_75t_L g948 ( 
.A(n_841),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_789),
.B(n_684),
.Y(n_949)
);

OAI21x1_ASAP7_75t_L g950 ( 
.A1(n_825),
.A2(n_575),
.B(n_573),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_828),
.B(n_684),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_844),
.B(n_660),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_798),
.Y(n_953)
);

OAI22xp5_ASAP7_75t_L g954 ( 
.A1(n_814),
.A2(n_415),
.B1(n_437),
.B2(n_434),
.Y(n_954)
);

AOI21x1_ASAP7_75t_SL g955 ( 
.A1(n_881),
.A2(n_882),
.B(n_877),
.Y(n_955)
);

OA22x2_ASAP7_75t_L g956 ( 
.A1(n_815),
.A2(n_458),
.B1(n_470),
.B2(n_457),
.Y(n_956)
);

AO31x2_ASAP7_75t_L g957 ( 
.A1(n_791),
.A2(n_442),
.A3(n_445),
.B(n_440),
.Y(n_957)
);

OA21x2_ASAP7_75t_L g958 ( 
.A1(n_865),
.A2(n_455),
.B(n_454),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_834),
.B(n_660),
.Y(n_959)
);

INVx4_ASAP7_75t_L g960 ( 
.A(n_826),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_818),
.A2(n_660),
.B1(n_349),
.B2(n_367),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_853),
.B(n_608),
.Y(n_962)
);

A2O1A1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_833),
.A2(n_463),
.B(n_472),
.C(n_468),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_839),
.B(n_840),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_871),
.A2(n_577),
.B(n_575),
.Y(n_965)
);

OAI21x1_ASAP7_75t_L g966 ( 
.A1(n_875),
.A2(n_578),
.B(n_577),
.Y(n_966)
);

AOI21x1_ASAP7_75t_L g967 ( 
.A1(n_872),
.A2(n_578),
.B(n_577),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_842),
.B(n_684),
.Y(n_968)
);

A2O1A1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_862),
.A2(n_610),
.B(n_604),
.C(n_291),
.Y(n_969)
);

AND2x4_ASAP7_75t_L g970 ( 
.A(n_800),
.B(n_604),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_859),
.B(n_352),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_874),
.A2(n_662),
.B(n_659),
.Y(n_972)
);

OAI21x1_ASAP7_75t_L g973 ( 
.A1(n_879),
.A2(n_578),
.B(n_577),
.Y(n_973)
);

OAI21xp5_ASAP7_75t_L g974 ( 
.A1(n_821),
.A2(n_660),
.B(n_684),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_822),
.A2(n_660),
.B(n_684),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_861),
.B(n_684),
.Y(n_976)
);

AO31x2_ASAP7_75t_L g977 ( 
.A1(n_883),
.A2(n_662),
.A3(n_688),
.B(n_659),
.Y(n_977)
);

OAI21x1_ASAP7_75t_L g978 ( 
.A1(n_864),
.A2(n_587),
.B(n_578),
.Y(n_978)
);

OA21x2_ASAP7_75t_L g979 ( 
.A1(n_843),
.A2(n_587),
.B(n_571),
.Y(n_979)
);

AND2x2_ASAP7_75t_L g980 ( 
.A(n_823),
.B(n_604),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_801),
.Y(n_981)
);

OAI21x1_ASAP7_75t_L g982 ( 
.A1(n_802),
.A2(n_803),
.B(n_587),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_849),
.A2(n_688),
.B(n_650),
.Y(n_983)
);

OA21x2_ASAP7_75t_L g984 ( 
.A1(n_893),
.A2(n_571),
.B(n_570),
.Y(n_984)
);

BUFx12f_ASAP7_75t_L g985 ( 
.A(n_912),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_939),
.A2(n_688),
.B(n_650),
.Y(n_986)
);

AND2x4_ASAP7_75t_L g987 ( 
.A(n_888),
.B(n_851),
.Y(n_987)
);

INVx2_ASAP7_75t_L g988 ( 
.A(n_930),
.Y(n_988)
);

AOI22xp33_ASAP7_75t_SL g989 ( 
.A1(n_956),
.A2(n_397),
.B1(n_296),
.B2(n_474),
.Y(n_989)
);

NOR2xp33_ASAP7_75t_L g990 ( 
.A(n_889),
.B(n_855),
.Y(n_990)
);

OAI21x1_ASAP7_75t_L g991 ( 
.A1(n_905),
.A2(n_579),
.B(n_570),
.Y(n_991)
);

INVx1_ASAP7_75t_SL g992 ( 
.A(n_927),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_891),
.A2(n_582),
.B(n_581),
.Y(n_993)
);

AOI21x1_ASAP7_75t_L g994 ( 
.A1(n_907),
.A2(n_582),
.B(n_581),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_901),
.B(n_858),
.Y(n_995)
);

BUFx2_ASAP7_75t_L g996 ( 
.A(n_913),
.Y(n_996)
);

CKINVDCx20_ASAP7_75t_R g997 ( 
.A(n_921),
.Y(n_997)
);

NOR2xp33_ASAP7_75t_L g998 ( 
.A(n_892),
.B(n_476),
.Y(n_998)
);

OAI21x1_ASAP7_75t_L g999 ( 
.A1(n_902),
.A2(n_585),
.B(n_584),
.Y(n_999)
);

AOI22xp33_ASAP7_75t_L g1000 ( 
.A1(n_899),
.A2(n_397),
.B1(n_296),
.B2(n_362),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_943),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_930),
.Y(n_1002)
);

OAI21x1_ASAP7_75t_L g1003 ( 
.A1(n_965),
.A2(n_967),
.B(n_947),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_913),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_887),
.A2(n_610),
.B(n_584),
.C(n_586),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_L g1006 ( 
.A(n_953),
.B(n_610),
.Y(n_1006)
);

OAI21x1_ASAP7_75t_L g1007 ( 
.A1(n_966),
.A2(n_586),
.B(n_585),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_946),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_894),
.Y(n_1009)
);

AND2x2_ASAP7_75t_L g1010 ( 
.A(n_980),
.B(n_397),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_893),
.A2(n_951),
.B(n_911),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_900),
.Y(n_1012)
);

OAI21x1_ASAP7_75t_L g1013 ( 
.A1(n_973),
.A2(n_590),
.B(n_588),
.Y(n_1013)
);

AOI22xp33_ASAP7_75t_L g1014 ( 
.A1(n_899),
.A2(n_928),
.B1(n_956),
.B2(n_919),
.Y(n_1014)
);

AOI32xp33_ASAP7_75t_L g1015 ( 
.A1(n_928),
.A2(n_954),
.A3(n_890),
.B1(n_981),
.B2(n_964),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_908),
.Y(n_1016)
);

INVx3_ASAP7_75t_L g1017 ( 
.A(n_896),
.Y(n_1017)
);

NOR3xp33_ASAP7_75t_L g1018 ( 
.A(n_940),
.B(n_610),
.C(n_819),
.Y(n_1018)
);

OAI21x1_ASAP7_75t_L g1019 ( 
.A1(n_950),
.A2(n_590),
.B(n_588),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_982),
.A2(n_593),
.B(n_591),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_918),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_926),
.B(n_591),
.Y(n_1022)
);

AOI22xp33_ASAP7_75t_L g1023 ( 
.A1(n_909),
.A2(n_362),
.B1(n_369),
.B2(n_355),
.Y(n_1023)
);

OAI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_935),
.A2(n_597),
.B(n_593),
.Y(n_1024)
);

OAI21x1_ASAP7_75t_L g1025 ( 
.A1(n_906),
.A2(n_599),
.B(n_597),
.Y(n_1025)
);

OAI22xp33_ASAP7_75t_L g1026 ( 
.A1(n_890),
.A2(n_940),
.B1(n_948),
.B2(n_942),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_937),
.B(n_948),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_922),
.Y(n_1028)
);

OAI21x1_ASAP7_75t_L g1029 ( 
.A1(n_925),
.A2(n_600),
.B(n_599),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_897),
.B(n_600),
.Y(n_1030)
);

OAI22xp5_ASAP7_75t_L g1031 ( 
.A1(n_981),
.A2(n_425),
.B1(n_370),
.B2(n_375),
.Y(n_1031)
);

AOI222xp33_ASAP7_75t_L g1032 ( 
.A1(n_954),
.A2(n_368),
.B1(n_377),
.B2(n_378),
.C1(n_379),
.C2(n_385),
.Y(n_1032)
);

OR2x2_ASAP7_75t_L g1033 ( 
.A(n_920),
.B(n_386),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_960),
.B(n_388),
.Y(n_1034)
);

OAI222xp33_ASAP7_75t_L g1035 ( 
.A1(n_960),
.A2(n_391),
.B1(n_392),
.B2(n_398),
.C1(n_402),
.C2(n_404),
.Y(n_1035)
);

OAI21x1_ASAP7_75t_L g1036 ( 
.A1(n_936),
.A2(n_650),
.B(n_362),
.Y(n_1036)
);

OA21x2_ASAP7_75t_L g1037 ( 
.A1(n_895),
.A2(n_413),
.B(n_406),
.Y(n_1037)
);

OAI21x1_ASAP7_75t_L g1038 ( 
.A1(n_904),
.A2(n_933),
.B(n_978),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_895),
.A2(n_650),
.B(n_648),
.Y(n_1039)
);

OAI21x1_ASAP7_75t_L g1040 ( 
.A1(n_931),
.A2(n_944),
.B(n_924),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_894),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_920),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_912),
.Y(n_1043)
);

OAI21x1_ASAP7_75t_SL g1044 ( 
.A1(n_929),
.A2(n_362),
.B(n_355),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_SL g1045 ( 
.A1(n_903),
.A2(n_362),
.B(n_355),
.Y(n_1045)
);

AOI21x1_ASAP7_75t_L g1046 ( 
.A1(n_898),
.A2(n_650),
.B(n_598),
.Y(n_1046)
);

INVxp67_ASAP7_75t_SL g1047 ( 
.A(n_923),
.Y(n_1047)
);

NOR2xp33_ASAP7_75t_L g1048 ( 
.A(n_948),
.B(n_416),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_898),
.A2(n_650),
.B(n_648),
.Y(n_1049)
);

AO31x2_ASAP7_75t_L g1050 ( 
.A1(n_903),
.A2(n_355),
.A3(n_362),
.B(n_369),
.Y(n_1050)
);

AND2x2_ASAP7_75t_L g1051 ( 
.A(n_948),
.B(n_426),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_916),
.B(n_428),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_971),
.Y(n_1053)
);

AOI21x1_ASAP7_75t_L g1054 ( 
.A1(n_972),
.A2(n_598),
.B(n_362),
.Y(n_1054)
);

OAI222xp33_ASAP7_75t_L g1055 ( 
.A1(n_962),
.A2(n_429),
.B1(n_439),
.B2(n_444),
.C1(n_447),
.C2(n_449),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_923),
.Y(n_1056)
);

AOI22xp33_ASAP7_75t_L g1057 ( 
.A1(n_970),
.A2(n_355),
.B1(n_369),
.B2(n_431),
.Y(n_1057)
);

INVx2_ASAP7_75t_SL g1058 ( 
.A(n_970),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_924),
.A2(n_369),
.B(n_441),
.Y(n_1059)
);

AND2x4_ASAP7_75t_L g1060 ( 
.A(n_983),
.B(n_96),
.Y(n_1060)
);

INVx6_ASAP7_75t_L g1061 ( 
.A(n_955),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_917),
.B(n_914),
.Y(n_1062)
);

INVxp67_ASAP7_75t_L g1063 ( 
.A(n_959),
.Y(n_1063)
);

OAI21x1_ASAP7_75t_L g1064 ( 
.A1(n_979),
.A2(n_369),
.B(n_441),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_941),
.Y(n_1065)
);

INVx4_ASAP7_75t_L g1066 ( 
.A(n_958),
.Y(n_1066)
);

BUFx2_ASAP7_75t_L g1067 ( 
.A(n_932),
.Y(n_1067)
);

OAI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_952),
.A2(n_459),
.B(n_456),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_958),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_938),
.B(n_464),
.Y(n_1070)
);

OAI21x1_ASAP7_75t_L g1071 ( 
.A1(n_952),
.A2(n_369),
.B(n_441),
.Y(n_1071)
);

A2O1A1Ixp33_ASAP7_75t_L g1072 ( 
.A1(n_910),
.A2(n_469),
.B(n_471),
.C(n_13),
.Y(n_1072)
);

OAI21x1_ASAP7_75t_SL g1073 ( 
.A1(n_974),
.A2(n_101),
.B(n_98),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_977),
.Y(n_1074)
);

OAI21x1_ASAP7_75t_L g1075 ( 
.A1(n_975),
.A2(n_673),
.B(n_648),
.Y(n_1075)
);

INVx5_ASAP7_75t_SL g1076 ( 
.A(n_915),
.Y(n_1076)
);

INVxp67_ASAP7_75t_SL g1077 ( 
.A(n_959),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_975),
.A2(n_11),
.B1(n_12),
.B2(n_14),
.Y(n_1078)
);

BUFx8_ASAP7_75t_L g1079 ( 
.A(n_945),
.Y(n_1079)
);

AND2x2_ASAP7_75t_L g1080 ( 
.A(n_941),
.B(n_12),
.Y(n_1080)
);

INVx3_ASAP7_75t_L g1081 ( 
.A(n_941),
.Y(n_1081)
);

OAI21x1_ASAP7_75t_L g1082 ( 
.A1(n_934),
.A2(n_104),
.B(n_102),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_968),
.B(n_15),
.Y(n_1083)
);

OA21x2_ASAP7_75t_L g1084 ( 
.A1(n_969),
.A2(n_673),
.B(n_648),
.Y(n_1084)
);

INVxp67_ASAP7_75t_L g1085 ( 
.A(n_963),
.Y(n_1085)
);

OAI221xp5_ASAP7_75t_L g1086 ( 
.A1(n_961),
.A2(n_673),
.B1(n_648),
.B2(n_18),
.C(n_19),
.Y(n_1086)
);

O2A1O1Ixp33_ASAP7_75t_SL g1087 ( 
.A1(n_976),
.A2(n_15),
.B(n_16),
.C(n_18),
.Y(n_1087)
);

OAI21x1_ASAP7_75t_L g1088 ( 
.A1(n_949),
.A2(n_108),
.B(n_105),
.Y(n_1088)
);

OAI21x1_ASAP7_75t_L g1089 ( 
.A1(n_945),
.A2(n_110),
.B(n_109),
.Y(n_1089)
);

INVx2_ASAP7_75t_L g1090 ( 
.A(n_977),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_957),
.Y(n_1091)
);

OR2x2_ASAP7_75t_L g1092 ( 
.A(n_1056),
.B(n_957),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_1009),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_1009),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_1041),
.Y(n_1095)
);

INVx1_ASAP7_75t_L g1096 ( 
.A(n_1041),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_1050),
.Y(n_1097)
);

BUFx2_ASAP7_75t_L g1098 ( 
.A(n_1077),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_1050),
.Y(n_1099)
);

AOI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_1018),
.A2(n_945),
.B1(n_673),
.B2(n_957),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_1000),
.A2(n_1026),
.B1(n_1078),
.B2(n_1014),
.Y(n_1101)
);

BUFx6f_ASAP7_75t_L g1102 ( 
.A(n_1060),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_1050),
.Y(n_1103)
);

AOI21x1_ASAP7_75t_L g1104 ( 
.A1(n_1054),
.A2(n_977),
.B(n_673),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1015),
.B(n_16),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_1061),
.Y(n_1106)
);

AOI22xp33_ASAP7_75t_L g1107 ( 
.A1(n_1026),
.A2(n_20),
.B1(n_21),
.B2(n_22),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_1050),
.Y(n_1108)
);

INVx1_ASAP7_75t_L g1109 ( 
.A(n_1047),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1091),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_992),
.Y(n_1111)
);

AND2x2_ASAP7_75t_L g1112 ( 
.A(n_1083),
.B(n_1063),
.Y(n_1112)
);

INVx2_ASAP7_75t_L g1113 ( 
.A(n_1074),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1074),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_L g1115 ( 
.A(n_1008),
.B(n_20),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_1081),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1090),
.Y(n_1117)
);

AO21x2_ASAP7_75t_L g1118 ( 
.A1(n_1046),
.A2(n_115),
.B(n_111),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1081),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_1090),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_984),
.Y(n_1121)
);

OAI22xp5_ASAP7_75t_L g1122 ( 
.A1(n_1000),
.A2(n_21),
.B1(n_23),
.B2(n_24),
.Y(n_1122)
);

OR2x2_ASAP7_75t_L g1123 ( 
.A(n_1011),
.B(n_24),
.Y(n_1123)
);

INVx2_ASAP7_75t_L g1124 ( 
.A(n_984),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_996),
.Y(n_1125)
);

INVx2_ASAP7_75t_L g1126 ( 
.A(n_984),
.Y(n_1126)
);

CKINVDCx6p67_ASAP7_75t_R g1127 ( 
.A(n_985),
.Y(n_1127)
);

BUFx3_ASAP7_75t_L g1128 ( 
.A(n_985),
.Y(n_1128)
);

OA21x2_ASAP7_75t_L g1129 ( 
.A1(n_1089),
.A2(n_25),
.B(n_26),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_1065),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_991),
.Y(n_1131)
);

AO21x2_ASAP7_75t_L g1132 ( 
.A1(n_1089),
.A2(n_135),
.B(n_283),
.Y(n_1132)
);

BUFx2_ASAP7_75t_L g1133 ( 
.A(n_1004),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_1014),
.B(n_26),
.Y(n_1134)
);

HB1xp67_ASAP7_75t_L g1135 ( 
.A(n_1001),
.Y(n_1135)
);

AOI22xp33_ASAP7_75t_L g1136 ( 
.A1(n_1067),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1136)
);

INVx2_ASAP7_75t_SL g1137 ( 
.A(n_1061),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_991),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_1083),
.B(n_116),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1020),
.Y(n_1140)
);

INVx2_ASAP7_75t_L g1141 ( 
.A(n_1064),
.Y(n_1141)
);

INVx2_ASAP7_75t_L g1142 ( 
.A(n_1059),
.Y(n_1142)
);

BUFx3_ASAP7_75t_L g1143 ( 
.A(n_1028),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1020),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_993),
.Y(n_1145)
);

INVx2_ASAP7_75t_L g1146 ( 
.A(n_1069),
.Y(n_1146)
);

AND2x2_ASAP7_75t_L g1147 ( 
.A(n_1080),
.B(n_285),
.Y(n_1147)
);

OAI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_989),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_999),
.Y(n_1149)
);

INVx3_ASAP7_75t_L g1150 ( 
.A(n_1060),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1019),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_1069),
.Y(n_1152)
);

BUFx3_ASAP7_75t_L g1153 ( 
.A(n_1028),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_1019),
.Y(n_1154)
);

HB1xp67_ASAP7_75t_L g1155 ( 
.A(n_1012),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1025),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_1038),
.A2(n_138),
.B(n_281),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1071),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1061),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_1076),
.B(n_30),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1029),
.Y(n_1161)
);

INVx2_ASAP7_75t_L g1162 ( 
.A(n_1036),
.Y(n_1162)
);

BUFx3_ASAP7_75t_L g1163 ( 
.A(n_1028),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1016),
.Y(n_1164)
);

AND2x6_ASAP7_75t_L g1165 ( 
.A(n_1076),
.B(n_117),
.Y(n_1165)
);

OR2x6_ASAP7_75t_L g1166 ( 
.A(n_1040),
.B(n_118),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_1021),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1042),
.Y(n_1168)
);

OA21x2_ASAP7_75t_L g1169 ( 
.A1(n_1003),
.A2(n_30),
.B(n_31),
.Y(n_1169)
);

BUFx2_ASAP7_75t_L g1170 ( 
.A(n_1027),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1036),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_986),
.A2(n_143),
.B(n_279),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1076),
.B(n_1062),
.Y(n_1173)
);

OAI21x1_ASAP7_75t_L g1174 ( 
.A1(n_1003),
.A2(n_141),
.B(n_275),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_1032),
.A2(n_33),
.B1(n_34),
.B2(n_35),
.Y(n_1175)
);

INVx2_ASAP7_75t_L g1176 ( 
.A(n_1084),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1084),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_1013),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_1013),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_1127),
.Y(n_1180)
);

NAND2xp33_ASAP7_75t_R g1181 ( 
.A(n_1133),
.B(n_1043),
.Y(n_1181)
);

OR2x6_ASAP7_75t_L g1182 ( 
.A(n_1128),
.B(n_987),
.Y(n_1182)
);

INVxp67_ASAP7_75t_L g1183 ( 
.A(n_1111),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_R g1184 ( 
.A(n_1127),
.B(n_997),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_1143),
.B(n_1028),
.Y(n_1185)
);

OR2x6_ASAP7_75t_L g1186 ( 
.A(n_1128),
.B(n_987),
.Y(n_1186)
);

AND2x4_ASAP7_75t_L g1187 ( 
.A(n_1143),
.B(n_987),
.Y(n_1187)
);

BUFx10_ASAP7_75t_L g1188 ( 
.A(n_1125),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_1112),
.B(n_1010),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_R g1190 ( 
.A(n_1127),
.B(n_997),
.Y(n_1190)
);

INVxp67_ASAP7_75t_L g1191 ( 
.A(n_1133),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1112),
.B(n_1105),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1105),
.B(n_1053),
.Y(n_1193)
);

NOR2xp33_ASAP7_75t_R g1194 ( 
.A(n_1128),
.B(n_1043),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1170),
.B(n_995),
.Y(n_1195)
);

AND2x4_ASAP7_75t_L g1196 ( 
.A(n_1143),
.B(n_988),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1135),
.Y(n_1197)
);

AND2x4_ASAP7_75t_L g1198 ( 
.A(n_1153),
.B(n_988),
.Y(n_1198)
);

NOR2xp33_ASAP7_75t_L g1199 ( 
.A(n_1173),
.B(n_1034),
.Y(n_1199)
);

AND2x4_ASAP7_75t_L g1200 ( 
.A(n_1153),
.B(n_1163),
.Y(n_1200)
);

OR2x6_ASAP7_75t_L g1201 ( 
.A(n_1102),
.B(n_1058),
.Y(n_1201)
);

OR2x6_ASAP7_75t_L g1202 ( 
.A(n_1102),
.B(n_1045),
.Y(n_1202)
);

XOR2xp5_ASAP7_75t_L g1203 ( 
.A(n_1173),
.B(n_1053),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1160),
.B(n_1034),
.Y(n_1204)
);

AND2x2_ASAP7_75t_L g1205 ( 
.A(n_1170),
.B(n_1051),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_R g1206 ( 
.A(n_1153),
.B(n_990),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1135),
.Y(n_1207)
);

NAND2xp33_ASAP7_75t_R g1208 ( 
.A(n_1139),
.B(n_990),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_R g1209 ( 
.A(n_1139),
.B(n_1048),
.Y(n_1209)
);

NAND2xp5_ASAP7_75t_L g1210 ( 
.A(n_1134),
.B(n_1048),
.Y(n_1210)
);

NAND2xp33_ASAP7_75t_R g1211 ( 
.A(n_1160),
.B(n_1147),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_R g1212 ( 
.A(n_1163),
.B(n_1033),
.Y(n_1212)
);

AND2x4_ASAP7_75t_L g1213 ( 
.A(n_1163),
.B(n_1002),
.Y(n_1213)
);

NAND2xp33_ASAP7_75t_R g1214 ( 
.A(n_1147),
.B(n_1037),
.Y(n_1214)
);

NAND2xp33_ASAP7_75t_R g1215 ( 
.A(n_1123),
.B(n_1037),
.Y(n_1215)
);

NOR2xp33_ASAP7_75t_R g1216 ( 
.A(n_1106),
.B(n_1017),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_SL g1217 ( 
.A(n_1102),
.B(n_1060),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1106),
.Y(n_1218)
);

AND2x2_ASAP7_75t_L g1219 ( 
.A(n_1168),
.B(n_1002),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1106),
.Y(n_1220)
);

CKINVDCx5p33_ASAP7_75t_R g1221 ( 
.A(n_1137),
.Y(n_1221)
);

INVxp67_ASAP7_75t_L g1222 ( 
.A(n_1155),
.Y(n_1222)
);

XOR2xp5_ASAP7_75t_L g1223 ( 
.A(n_1102),
.B(n_1031),
.Y(n_1223)
);

NOR2xp33_ASAP7_75t_R g1224 ( 
.A(n_1137),
.B(n_1017),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1102),
.B(n_1072),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_1137),
.Y(n_1226)
);

CKINVDCx12_ASAP7_75t_R g1227 ( 
.A(n_1123),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_SL g1228 ( 
.A(n_1102),
.B(n_1072),
.Y(n_1228)
);

BUFx3_ASAP7_75t_L g1229 ( 
.A(n_1159),
.Y(n_1229)
);

NAND2xp33_ASAP7_75t_SL g1230 ( 
.A(n_1101),
.B(n_1052),
.Y(n_1230)
);

NOR2x1_ASAP7_75t_L g1231 ( 
.A(n_1115),
.B(n_1134),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1155),
.B(n_1030),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1164),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1164),
.Y(n_1234)
);

NAND2xp33_ASAP7_75t_R g1235 ( 
.A(n_1098),
.B(n_1037),
.Y(n_1235)
);

XNOR2xp5_ASAP7_75t_L g1236 ( 
.A(n_1148),
.B(n_1030),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1110),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_R g1238 ( 
.A(n_1159),
.B(n_998),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1115),
.B(n_1030),
.Y(n_1239)
);

AND2x4_ASAP7_75t_L g1240 ( 
.A(n_1159),
.B(n_1150),
.Y(n_1240)
);

INVxp67_ASAP7_75t_L g1241 ( 
.A(n_1167),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1167),
.Y(n_1242)
);

NAND2xp33_ASAP7_75t_R g1243 ( 
.A(n_1098),
.B(n_998),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1166),
.B(n_1073),
.Y(n_1244)
);

NAND2xp5_ASAP7_75t_L g1245 ( 
.A(n_1107),
.B(n_1006),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1233),
.B(n_1097),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1197),
.Y(n_1247)
);

INVxp67_ASAP7_75t_SL g1248 ( 
.A(n_1222),
.Y(n_1248)
);

AOI22xp33_ASAP7_75t_L g1249 ( 
.A1(n_1230),
.A2(n_1101),
.B1(n_1175),
.B2(n_1148),
.Y(n_1249)
);

AND2x2_ASAP7_75t_L g1250 ( 
.A(n_1234),
.B(n_1097),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1243),
.Y(n_1251)
);

INVx3_ASAP7_75t_SL g1252 ( 
.A(n_1221),
.Y(n_1252)
);

AND2x4_ASAP7_75t_L g1253 ( 
.A(n_1240),
.B(n_1166),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1237),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1207),
.B(n_1241),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1237),
.Y(n_1256)
);

AND2x2_ASAP7_75t_SL g1257 ( 
.A(n_1211),
.B(n_1129),
.Y(n_1257)
);

BUFx3_ASAP7_75t_L g1258 ( 
.A(n_1218),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1242),
.B(n_1109),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1199),
.B(n_1035),
.Y(n_1260)
);

OR2x2_ASAP7_75t_L g1261 ( 
.A(n_1195),
.B(n_1099),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1189),
.B(n_1099),
.Y(n_1262)
);

AND2x2_ASAP7_75t_L g1263 ( 
.A(n_1240),
.B(n_1103),
.Y(n_1263)
);

OR2x2_ASAP7_75t_L g1264 ( 
.A(n_1192),
.B(n_1103),
.Y(n_1264)
);

INVxp67_ASAP7_75t_L g1265 ( 
.A(n_1235),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1232),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1204),
.A2(n_1165),
.B1(n_1231),
.B2(n_1210),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1205),
.B(n_1109),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1239),
.B(n_1093),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1219),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1187),
.B(n_1108),
.Y(n_1271)
);

AND2x2_ASAP7_75t_L g1272 ( 
.A(n_1187),
.B(n_1108),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1220),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1191),
.B(n_1110),
.Y(n_1274)
);

AND2x4_ASAP7_75t_L g1275 ( 
.A(n_1244),
.B(n_1166),
.Y(n_1275)
);

NOR2x1_ASAP7_75t_L g1276 ( 
.A(n_1229),
.B(n_1169),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1225),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1228),
.Y(n_1278)
);

AND2x2_ASAP7_75t_L g1279 ( 
.A(n_1244),
.B(n_1116),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_1200),
.B(n_1116),
.Y(n_1280)
);

AND2x2_ASAP7_75t_L g1281 ( 
.A(n_1200),
.B(n_1119),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1196),
.B(n_1119),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1202),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1227),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1202),
.B(n_1166),
.Y(n_1285)
);

HB1xp67_ASAP7_75t_L g1286 ( 
.A(n_1183),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_1196),
.Y(n_1287)
);

OR2x2_ASAP7_75t_L g1288 ( 
.A(n_1193),
.B(n_1121),
.Y(n_1288)
);

AND2x2_ASAP7_75t_L g1289 ( 
.A(n_1198),
.B(n_1113),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1198),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1213),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1213),
.Y(n_1292)
);

AND2x2_ASAP7_75t_L g1293 ( 
.A(n_1182),
.B(n_1113),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1182),
.Y(n_1294)
);

OR2x2_ASAP7_75t_L g1295 ( 
.A(n_1186),
.B(n_1121),
.Y(n_1295)
);

AOI22xp33_ASAP7_75t_SL g1296 ( 
.A1(n_1245),
.A2(n_1122),
.B1(n_1165),
.B2(n_1079),
.Y(n_1296)
);

OR2x2_ASAP7_75t_L g1297 ( 
.A(n_1186),
.B(n_1124),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1247),
.Y(n_1298)
);

INVx3_ASAP7_75t_L g1299 ( 
.A(n_1253),
.Y(n_1299)
);

NAND2xp5_ASAP7_75t_L g1300 ( 
.A(n_1288),
.B(n_1124),
.Y(n_1300)
);

XNOR2x2_ASAP7_75t_L g1301 ( 
.A(n_1260),
.B(n_1122),
.Y(n_1301)
);

INVx2_ASAP7_75t_L g1302 ( 
.A(n_1254),
.Y(n_1302)
);

AND2x2_ASAP7_75t_SL g1303 ( 
.A(n_1257),
.B(n_1129),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1254),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_1256),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1263),
.B(n_1176),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1263),
.B(n_1176),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_L g1308 ( 
.A(n_1288),
.B(n_1124),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1257),
.B(n_1176),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1256),
.Y(n_1310)
);

HB1xp67_ASAP7_75t_L g1311 ( 
.A(n_1247),
.Y(n_1311)
);

AOI31xp33_ASAP7_75t_SL g1312 ( 
.A1(n_1251),
.A2(n_1236),
.A3(n_1209),
.B(n_1208),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1255),
.Y(n_1313)
);

INVx2_ASAP7_75t_L g1314 ( 
.A(n_1246),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1255),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1246),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1250),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1264),
.B(n_1126),
.Y(n_1318)
);

OAI33xp33_ASAP7_75t_L g1319 ( 
.A1(n_1277),
.A2(n_1226),
.A3(n_1180),
.B1(n_37),
.B2(n_38),
.B3(n_39),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_1250),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1259),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1252),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1257),
.B(n_1177),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1264),
.B(n_1126),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1259),
.Y(n_1325)
);

NAND3xp33_ASAP7_75t_L g1326 ( 
.A(n_1249),
.B(n_1215),
.C(n_1136),
.Y(n_1326)
);

AND2x4_ASAP7_75t_L g1327 ( 
.A(n_1253),
.B(n_1177),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1276),
.B(n_1262),
.Y(n_1328)
);

NAND2xp5_ASAP7_75t_SL g1329 ( 
.A(n_1251),
.B(n_1212),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1253),
.B(n_1177),
.Y(n_1330)
);

HB1xp67_ASAP7_75t_L g1331 ( 
.A(n_1277),
.Y(n_1331)
);

INVx1_ASAP7_75t_SL g1332 ( 
.A(n_1295),
.Y(n_1332)
);

INVx3_ASAP7_75t_L g1333 ( 
.A(n_1253),
.Y(n_1333)
);

OAI33xp33_ASAP7_75t_L g1334 ( 
.A1(n_1278),
.A2(n_35),
.A3(n_36),
.B1(n_38),
.B2(n_39),
.B3(n_40),
.Y(n_1334)
);

NOR2xp33_ASAP7_75t_L g1335 ( 
.A(n_1284),
.B(n_1203),
.Y(n_1335)
);

OR2x2_ASAP7_75t_L g1336 ( 
.A(n_1261),
.B(n_1126),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1276),
.B(n_1169),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1262),
.B(n_1169),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1274),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1283),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1271),
.B(n_1169),
.Y(n_1341)
);

NOR2x1_ASAP7_75t_L g1342 ( 
.A(n_1258),
.B(n_1169),
.Y(n_1342)
);

OR2x2_ASAP7_75t_L g1343 ( 
.A(n_1261),
.B(n_1113),
.Y(n_1343)
);

AND2x2_ASAP7_75t_L g1344 ( 
.A(n_1271),
.B(n_1131),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1272),
.B(n_1131),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1275),
.B(n_1166),
.Y(n_1346)
);

AND2x2_ASAP7_75t_L g1347 ( 
.A(n_1272),
.B(n_1138),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1275),
.B(n_1265),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1275),
.B(n_1138),
.Y(n_1349)
);

AND2x2_ASAP7_75t_L g1350 ( 
.A(n_1275),
.B(n_1130),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1265),
.B(n_1130),
.Y(n_1351)
);

INVx2_ASAP7_75t_L g1352 ( 
.A(n_1289),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1279),
.B(n_1114),
.Y(n_1353)
);

AND2x2_ASAP7_75t_L g1354 ( 
.A(n_1348),
.B(n_1279),
.Y(n_1354)
);

AND2x4_ASAP7_75t_L g1355 ( 
.A(n_1299),
.B(n_1285),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1348),
.B(n_1283),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1302),
.Y(n_1357)
);

AND2x2_ASAP7_75t_L g1358 ( 
.A(n_1348),
.B(n_1283),
.Y(n_1358)
);

AND2x2_ASAP7_75t_L g1359 ( 
.A(n_1328),
.B(n_1299),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1328),
.B(n_1285),
.Y(n_1360)
);

AND2x2_ASAP7_75t_L g1361 ( 
.A(n_1328),
.B(n_1285),
.Y(n_1361)
);

OR2x2_ASAP7_75t_L g1362 ( 
.A(n_1332),
.B(n_1295),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1302),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1332),
.B(n_1297),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1302),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1310),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1310),
.Y(n_1367)
);

OR2x2_ASAP7_75t_L g1368 ( 
.A(n_1352),
.B(n_1297),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1299),
.B(n_1285),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1310),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1304),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1313),
.B(n_1286),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1304),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1301),
.A2(n_1296),
.B1(n_1165),
.B2(n_1284),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1305),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1322),
.B(n_1252),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1305),
.Y(n_1377)
);

NAND2xp5_ASAP7_75t_L g1378 ( 
.A(n_1313),
.B(n_1268),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1315),
.B(n_1268),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1299),
.B(n_1266),
.Y(n_1380)
);

NOR2xp33_ASAP7_75t_SL g1381 ( 
.A(n_1319),
.B(n_1252),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1315),
.B(n_1270),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1333),
.B(n_1266),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1298),
.Y(n_1384)
);

INVxp67_ASAP7_75t_L g1385 ( 
.A(n_1331),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1321),
.B(n_1248),
.Y(n_1386)
);

OR2x2_ASAP7_75t_L g1387 ( 
.A(n_1364),
.B(n_1352),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1372),
.B(n_1321),
.Y(n_1388)
);

INVxp67_ASAP7_75t_L g1389 ( 
.A(n_1381),
.Y(n_1389)
);

OAI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1381),
.A2(n_1326),
.B1(n_1346),
.B2(n_1214),
.Y(n_1390)
);

NAND2xp5_ASAP7_75t_L g1391 ( 
.A(n_1378),
.B(n_1325),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1379),
.B(n_1325),
.Y(n_1392)
);

NOR2xp33_ASAP7_75t_R g1393 ( 
.A(n_1376),
.B(n_1181),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1362),
.A2(n_1326),
.B1(n_1346),
.B2(n_1301),
.Y(n_1394)
);

INVx3_ASAP7_75t_L g1395 ( 
.A(n_1355),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1385),
.B(n_1309),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1386),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1362),
.A2(n_1346),
.B1(n_1301),
.B2(n_1278),
.Y(n_1398)
);

NAND2xp33_ASAP7_75t_SL g1399 ( 
.A(n_1374),
.B(n_1184),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_SL g1400 ( 
.A(n_1386),
.B(n_1329),
.Y(n_1400)
);

OAI22xp33_ASAP7_75t_L g1401 ( 
.A1(n_1364),
.A2(n_1346),
.B1(n_1333),
.B2(n_1294),
.Y(n_1401)
);

NAND2xp5_ASAP7_75t_L g1402 ( 
.A(n_1354),
.B(n_1309),
.Y(n_1402)
);

CKINVDCx5p33_ASAP7_75t_R g1403 ( 
.A(n_1382),
.Y(n_1403)
);

AOI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1355),
.A2(n_1319),
.B1(n_1334),
.B2(n_1296),
.Y(n_1404)
);

OR2x6_ASAP7_75t_L g1405 ( 
.A(n_1355),
.B(n_1346),
.Y(n_1405)
);

AO221x2_ASAP7_75t_L g1406 ( 
.A1(n_1384),
.A2(n_1312),
.B1(n_1339),
.B2(n_1334),
.C(n_1223),
.Y(n_1406)
);

INVx3_ASAP7_75t_L g1407 ( 
.A(n_1355),
.Y(n_1407)
);

OAI221xp5_ASAP7_75t_L g1408 ( 
.A1(n_1384),
.A2(n_1312),
.B1(n_1267),
.B2(n_1335),
.C(n_1346),
.Y(n_1408)
);

BUFx3_ASAP7_75t_L g1409 ( 
.A(n_1354),
.Y(n_1409)
);

AOI22xp5_ASAP7_75t_L g1410 ( 
.A1(n_1369),
.A2(n_1303),
.B1(n_1349),
.B2(n_1333),
.Y(n_1410)
);

OAI22xp5_ASAP7_75t_L g1411 ( 
.A1(n_1360),
.A2(n_1303),
.B1(n_1294),
.B2(n_1333),
.Y(n_1411)
);

AO221x2_ASAP7_75t_L g1412 ( 
.A1(n_1373),
.A2(n_1339),
.B1(n_1303),
.B2(n_1317),
.C(n_1316),
.Y(n_1412)
);

AO221x2_ASAP7_75t_L g1413 ( 
.A1(n_1373),
.A2(n_1317),
.B1(n_1316),
.B2(n_1273),
.C(n_1314),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1360),
.B(n_1352),
.Y(n_1414)
);

AO221x2_ASAP7_75t_L g1415 ( 
.A1(n_1375),
.A2(n_1273),
.B1(n_1314),
.B2(n_1320),
.C(n_1270),
.Y(n_1415)
);

AO221x2_ASAP7_75t_L g1416 ( 
.A1(n_1375),
.A2(n_1314),
.B1(n_1320),
.B2(n_1318),
.C(n_1324),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1356),
.B(n_1309),
.Y(n_1417)
);

OAI221xp5_ASAP7_75t_L g1418 ( 
.A1(n_1368),
.A2(n_1248),
.B1(n_1340),
.B2(n_1300),
.C(n_1308),
.Y(n_1418)
);

NAND2x1_ASAP7_75t_L g1419 ( 
.A(n_1405),
.B(n_1359),
.Y(n_1419)
);

INVx1_ASAP7_75t_SL g1420 ( 
.A(n_1393),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1406),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1413),
.Y(n_1422)
);

NAND2xp5_ASAP7_75t_L g1423 ( 
.A(n_1389),
.B(n_1356),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1405),
.B(n_1361),
.Y(n_1424)
);

BUFx3_ASAP7_75t_L g1425 ( 
.A(n_1406),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1403),
.B(n_1397),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1395),
.B(n_1361),
.Y(n_1427)
);

NOR2xp33_ASAP7_75t_L g1428 ( 
.A(n_1400),
.B(n_1358),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1416),
.B(n_1368),
.Y(n_1429)
);

INVx3_ASAP7_75t_L g1430 ( 
.A(n_1413),
.Y(n_1430)
);

INVx1_ASAP7_75t_SL g1431 ( 
.A(n_1388),
.Y(n_1431)
);

NOR2xp33_ASAP7_75t_L g1432 ( 
.A(n_1408),
.B(n_1358),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1415),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1396),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1416),
.B(n_1371),
.Y(n_1435)
);

NAND3xp33_ASAP7_75t_L g1436 ( 
.A(n_1394),
.B(n_1337),
.C(n_1342),
.Y(n_1436)
);

INVx2_ASAP7_75t_SL g1437 ( 
.A(n_1415),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1391),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1392),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1387),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1412),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1407),
.B(n_1369),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_L g1443 ( 
.A(n_1412),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1414),
.Y(n_1444)
);

BUFx6f_ASAP7_75t_L g1445 ( 
.A(n_1409),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1410),
.B(n_1359),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1402),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1411),
.B(n_1380),
.Y(n_1448)
);

OR2x2_ASAP7_75t_L g1449 ( 
.A(n_1417),
.B(n_1371),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_L g1450 ( 
.A1(n_1390),
.A2(n_1165),
.B1(n_1350),
.B2(n_1349),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1418),
.Y(n_1451)
);

INVx2_ASAP7_75t_L g1452 ( 
.A(n_1404),
.Y(n_1452)
);

NOR2xp33_ASAP7_75t_L g1453 ( 
.A(n_1420),
.B(n_1398),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1421),
.A2(n_1399),
.B1(n_1401),
.B2(n_1350),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1421),
.A2(n_1342),
.B1(n_1337),
.B2(n_1323),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1452),
.B(n_1380),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1421),
.A2(n_1350),
.B1(n_1349),
.B2(n_1323),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1440),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1452),
.B(n_1383),
.Y(n_1459)
);

OR2x2_ASAP7_75t_L g1460 ( 
.A(n_1431),
.B(n_1311),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1440),
.Y(n_1461)
);

NAND2xp33_ASAP7_75t_L g1462 ( 
.A(n_1436),
.B(n_1190),
.Y(n_1462)
);

INVx1_ASAP7_75t_SL g1463 ( 
.A(n_1445),
.Y(n_1463)
);

NAND2x1_ASAP7_75t_L g1464 ( 
.A(n_1430),
.B(n_1383),
.Y(n_1464)
);

INVx2_ASAP7_75t_L g1465 ( 
.A(n_1445),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1436),
.A2(n_1337),
.B(n_1351),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1424),
.B(n_1445),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_SL g1468 ( 
.A1(n_1425),
.A2(n_1238),
.B1(n_1165),
.B2(n_1323),
.Y(n_1468)
);

OAI322xp33_ASAP7_75t_L g1469 ( 
.A1(n_1452),
.A2(n_1377),
.A3(n_1371),
.B1(n_1370),
.B2(n_1367),
.C1(n_1366),
.C2(n_1365),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1419),
.Y(n_1470)
);

INVx1_ASAP7_75t_SL g1471 ( 
.A(n_1445),
.Y(n_1471)
);

INVx2_ASAP7_75t_SL g1472 ( 
.A(n_1445),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1424),
.B(n_1340),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_L g1474 ( 
.A1(n_1425),
.A2(n_1055),
.B(n_1087),
.C(n_1086),
.Y(n_1474)
);

AOI31xp33_ASAP7_75t_L g1475 ( 
.A1(n_1443),
.A2(n_1194),
.A3(n_1217),
.B(n_1351),
.Y(n_1475)
);

AOI31xp33_ASAP7_75t_SL g1476 ( 
.A1(n_1432),
.A2(n_1308),
.A3(n_1300),
.B(n_1318),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1438),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1438),
.Y(n_1478)
);

OAI22xp33_ASAP7_75t_L g1479 ( 
.A1(n_1425),
.A2(n_1294),
.B1(n_1258),
.B2(n_1166),
.Y(n_1479)
);

HB1xp67_ASAP7_75t_L g1480 ( 
.A(n_1430),
.Y(n_1480)
);

OAI22xp33_ASAP7_75t_SL g1481 ( 
.A1(n_1430),
.A2(n_1377),
.B1(n_1357),
.B2(n_1365),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1439),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1445),
.Y(n_1483)
);

OAI322xp33_ASAP7_75t_L g1484 ( 
.A1(n_1441),
.A2(n_1370),
.A3(n_1367),
.B1(n_1366),
.B2(n_1363),
.C1(n_1357),
.C2(n_1324),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1467),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1480),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1453),
.B(n_1441),
.Y(n_1487)
);

AND2x2_ASAP7_75t_L g1488 ( 
.A(n_1470),
.B(n_1430),
.Y(n_1488)
);

AND2x4_ASAP7_75t_L g1489 ( 
.A(n_1472),
.B(n_1437),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1480),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1470),
.B(n_1433),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1458),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1463),
.B(n_1451),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1461),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1471),
.B(n_1465),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_L g1496 ( 
.A1(n_1454),
.A2(n_1450),
.B1(n_1451),
.B2(n_1433),
.Y(n_1496)
);

NAND2xp5_ASAP7_75t_L g1497 ( 
.A(n_1483),
.B(n_1439),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1462),
.B(n_1426),
.Y(n_1498)
);

INVx3_ASAP7_75t_L g1499 ( 
.A(n_1464),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1483),
.B(n_1422),
.Y(n_1500)
);

NOR2x1_ASAP7_75t_L g1501 ( 
.A(n_1475),
.B(n_1422),
.Y(n_1501)
);

INVx2_ASAP7_75t_SL g1502 ( 
.A(n_1460),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1477),
.B(n_1419),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1478),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_1456),
.Y(n_1505)
);

OR2x2_ASAP7_75t_L g1506 ( 
.A(n_1459),
.B(n_1429),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1473),
.B(n_1437),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1482),
.B(n_1428),
.Y(n_1508)
);

INVxp67_ASAP7_75t_L g1509 ( 
.A(n_1466),
.Y(n_1509)
);

INVx2_ASAP7_75t_L g1510 ( 
.A(n_1457),
.Y(n_1510)
);

INVxp67_ASAP7_75t_SL g1511 ( 
.A(n_1481),
.Y(n_1511)
);

NAND2x1_ASAP7_75t_L g1512 ( 
.A(n_1455),
.B(n_1435),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1479),
.B(n_1429),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1468),
.B(n_1434),
.Y(n_1514)
);

INVxp67_ASAP7_75t_L g1515 ( 
.A(n_1468),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1469),
.B(n_1423),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1476),
.Y(n_1517)
);

NOR2xp67_ASAP7_75t_SL g1518 ( 
.A(n_1474),
.B(n_1435),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1484),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1474),
.B(n_1446),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1486),
.Y(n_1521)
);

NAND2xp5_ASAP7_75t_L g1522 ( 
.A(n_1485),
.B(n_1444),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1490),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1499),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1490),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1499),
.Y(n_1526)
);

INVxp67_ASAP7_75t_SL g1527 ( 
.A(n_1499),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1492),
.Y(n_1528)
);

BUFx2_ASAP7_75t_L g1529 ( 
.A(n_1488),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1488),
.Y(n_1530)
);

INVxp67_ASAP7_75t_SL g1531 ( 
.A(n_1512),
.Y(n_1531)
);

INVx1_ASAP7_75t_SL g1532 ( 
.A(n_1495),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1492),
.Y(n_1533)
);

BUFx4f_ASAP7_75t_SL g1534 ( 
.A(n_1495),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1500),
.Y(n_1535)
);

INVx1_ASAP7_75t_SL g1536 ( 
.A(n_1491),
.Y(n_1536)
);

HB1xp67_ASAP7_75t_L g1537 ( 
.A(n_1502),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1500),
.Y(n_1538)
);

INVx2_ASAP7_75t_SL g1539 ( 
.A(n_1503),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1497),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1494),
.Y(n_1541)
);

BUFx2_ASAP7_75t_L g1542 ( 
.A(n_1511),
.Y(n_1542)
);

INVxp33_ASAP7_75t_SL g1543 ( 
.A(n_1498),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_1512),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

NOR2x1_ASAP7_75t_L g1546 ( 
.A(n_1501),
.B(n_1446),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1502),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1491),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1505),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1489),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1489),
.Y(n_1551)
);

INVxp33_ASAP7_75t_SL g1552 ( 
.A(n_1518),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1507),
.B(n_1442),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1518),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1489),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_L g1556 ( 
.A(n_1487),
.B(n_1447),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1517),
.Y(n_1557)
);

HB1xp67_ASAP7_75t_L g1558 ( 
.A(n_1507),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1520),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1517),
.B(n_1444),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1513),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_1493),
.Y(n_1562)
);

INVx1_ASAP7_75t_L g1563 ( 
.A(n_1506),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1506),
.Y(n_1564)
);

INVx2_ASAP7_75t_SL g1565 ( 
.A(n_1513),
.Y(n_1565)
);

NAND4xp25_ASAP7_75t_SL g1566 ( 
.A(n_1546),
.B(n_1519),
.C(n_1514),
.D(n_1510),
.Y(n_1566)
);

NOR3xp33_ASAP7_75t_L g1567 ( 
.A(n_1542),
.B(n_1515),
.C(n_1509),
.Y(n_1567)
);

AOI322xp5_ASAP7_75t_L g1568 ( 
.A1(n_1542),
.A2(n_1516),
.A3(n_1510),
.B1(n_1508),
.B2(n_1447),
.C1(n_1496),
.C2(n_1448),
.Y(n_1568)
);

OAI32xp33_ASAP7_75t_L g1569 ( 
.A1(n_1544),
.A2(n_1448),
.A3(n_1449),
.B1(n_1427),
.B2(n_1298),
.Y(n_1569)
);

NOR3x1_ASAP7_75t_L g1570 ( 
.A(n_1565),
.B(n_1449),
.C(n_1363),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_SL g1571 ( 
.A1(n_1531),
.A2(n_1427),
.B(n_1442),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1572)
);

O2A1O1Ixp33_ASAP7_75t_L g1573 ( 
.A1(n_1552),
.A2(n_1087),
.B(n_1172),
.C(n_1442),
.Y(n_1573)
);

NOR3xp33_ASAP7_75t_L g1574 ( 
.A(n_1557),
.B(n_1070),
.C(n_1006),
.Y(n_1574)
);

AND3x1_ASAP7_75t_L g1575 ( 
.A(n_1544),
.B(n_1351),
.C(n_1294),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_L g1576 ( 
.A(n_1554),
.B(n_1172),
.C(n_1057),
.Y(n_1576)
);

NAND4xp75_ASAP7_75t_L g1577 ( 
.A(n_1554),
.B(n_1129),
.C(n_1274),
.D(n_1341),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1552),
.A2(n_1085),
.B(n_1068),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1536),
.B(n_1188),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1537),
.Y(n_1580)
);

NOR3xp33_ASAP7_75t_L g1581 ( 
.A(n_1559),
.B(n_1022),
.C(n_1185),
.Y(n_1581)
);

AOI221xp5_ASAP7_75t_L g1582 ( 
.A1(n_1565),
.A2(n_1206),
.B1(n_1338),
.B2(n_1341),
.C(n_1057),
.Y(n_1582)
);

OAI21xp33_ASAP7_75t_L g1583 ( 
.A1(n_1543),
.A2(n_1258),
.B(n_1280),
.Y(n_1583)
);

NAND2xp33_ASAP7_75t_L g1584 ( 
.A(n_1558),
.B(n_1216),
.Y(n_1584)
);

NOR3xp33_ASAP7_75t_L g1585 ( 
.A(n_1562),
.B(n_1185),
.C(n_1005),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1530),
.B(n_1188),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1543),
.A2(n_1165),
.B1(n_1330),
.B2(n_1327),
.Y(n_1587)
);

O2A1O1Ixp5_ASAP7_75t_L g1588 ( 
.A1(n_1544),
.A2(n_1327),
.B(n_1330),
.C(n_1341),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1529),
.B(n_1344),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1529),
.B(n_1344),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1344),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1539),
.A2(n_1023),
.B(n_1044),
.Y(n_1592)
);

NOR2xp33_ASAP7_75t_L g1593 ( 
.A(n_1534),
.B(n_42),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1535),
.B(n_1345),
.Y(n_1594)
);

NAND3xp33_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1023),
.C(n_1129),
.Y(n_1595)
);

NAND4xp25_ASAP7_75t_L g1596 ( 
.A(n_1556),
.B(n_1269),
.C(n_1280),
.D(n_1281),
.Y(n_1596)
);

NAND4xp25_ASAP7_75t_L g1597 ( 
.A(n_1561),
.B(n_1269),
.C(n_1281),
.D(n_1100),
.Y(n_1597)
);

OAI211xp5_ASAP7_75t_L g1598 ( 
.A1(n_1561),
.A2(n_1224),
.B(n_1129),
.C(n_1338),
.Y(n_1598)
);

NOR4xp25_ASAP7_75t_L g1599 ( 
.A(n_1555),
.B(n_42),
.C(n_43),
.D(n_44),
.Y(n_1599)
);

NAND4xp25_ASAP7_75t_L g1600 ( 
.A(n_1549),
.B(n_43),
.C(n_45),
.D(n_46),
.Y(n_1600)
);

AND2x4_ASAP7_75t_L g1601 ( 
.A(n_1550),
.B(n_1320),
.Y(n_1601)
);

AOI211xp5_ASAP7_75t_L g1602 ( 
.A1(n_1539),
.A2(n_1338),
.B(n_47),
.C(n_48),
.Y(n_1602)
);

OAI21xp33_ASAP7_75t_L g1603 ( 
.A1(n_1560),
.A2(n_1522),
.B(n_1553),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_SL g1604 ( 
.A(n_1548),
.B(n_1165),
.Y(n_1604)
);

NAND4xp75_ASAP7_75t_L g1605 ( 
.A(n_1555),
.B(n_1524),
.C(n_1535),
.D(n_1564),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1524),
.Y(n_1606)
);

AO21x1_ASAP7_75t_L g1607 ( 
.A1(n_1527),
.A2(n_1525),
.B(n_1528),
.Y(n_1607)
);

NAND4xp25_ASAP7_75t_L g1608 ( 
.A(n_1563),
.B(n_1330),
.C(n_1327),
.D(n_1292),
.Y(n_1608)
);

NAND3xp33_ASAP7_75t_L g1609 ( 
.A(n_1563),
.B(n_1291),
.C(n_1290),
.Y(n_1609)
);

AOI221xp5_ASAP7_75t_L g1610 ( 
.A1(n_1564),
.A2(n_1290),
.B1(n_1291),
.B2(n_1292),
.C(n_1347),
.Y(n_1610)
);

NAND5xp2_ASAP7_75t_L g1611 ( 
.A(n_1538),
.B(n_1540),
.C(n_1553),
.D(n_1523),
.E(n_1525),
.Y(n_1611)
);

NAND2x1_ASAP7_75t_SL g1612 ( 
.A(n_1521),
.B(n_1345),
.Y(n_1612)
);

NAND5xp2_ASAP7_75t_L g1613 ( 
.A(n_1541),
.B(n_994),
.C(n_1293),
.D(n_1282),
.E(n_1353),
.Y(n_1613)
);

AOI221x1_ASAP7_75t_L g1614 ( 
.A1(n_1567),
.A2(n_1526),
.B1(n_1550),
.B2(n_1533),
.C(n_1528),
.Y(n_1614)
);

OAI22xp33_ASAP7_75t_SL g1615 ( 
.A1(n_1580),
.A2(n_1533),
.B1(n_1526),
.B2(n_1545),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1605),
.A2(n_1330),
.B1(n_1327),
.B2(n_1336),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1611),
.B(n_46),
.Y(n_1617)
);

AO22x2_ASAP7_75t_L g1618 ( 
.A1(n_1606),
.A2(n_1165),
.B1(n_51),
.B2(n_52),
.Y(n_1618)
);

AOI322xp5_ASAP7_75t_L g1619 ( 
.A1(n_1603),
.A2(n_1593),
.A3(n_1566),
.B1(n_1568),
.B2(n_1571),
.C1(n_1572),
.C2(n_1584),
.Y(n_1619)
);

AOI21xp33_ASAP7_75t_L g1620 ( 
.A1(n_1586),
.A2(n_50),
.B(n_51),
.Y(n_1620)
);

NOR3xp33_ASAP7_75t_L g1621 ( 
.A(n_1579),
.B(n_1088),
.C(n_1157),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1607),
.A2(n_1613),
.B1(n_1583),
.B2(n_1581),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1599),
.A2(n_1201),
.B(n_1132),
.Y(n_1623)
);

INVx2_ASAP7_75t_SL g1624 ( 
.A(n_1612),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1570),
.Y(n_1625)
);

OAI211xp5_ASAP7_75t_L g1626 ( 
.A1(n_1602),
.A2(n_52),
.B(n_54),
.C(n_55),
.Y(n_1626)
);

XNOR2x1_ASAP7_75t_L g1627 ( 
.A(n_1576),
.B(n_55),
.Y(n_1627)
);

OA211x2_ASAP7_75t_L g1628 ( 
.A1(n_1604),
.A2(n_56),
.B(n_57),
.C(n_58),
.Y(n_1628)
);

O2A1O1Ixp33_ASAP7_75t_L g1629 ( 
.A1(n_1600),
.A2(n_1132),
.B(n_59),
.C(n_60),
.Y(n_1629)
);

OAI21xp33_ASAP7_75t_L g1630 ( 
.A1(n_1591),
.A2(n_1347),
.B(n_1345),
.Y(n_1630)
);

OAI22xp5_ASAP7_75t_L g1631 ( 
.A1(n_1575),
.A2(n_1330),
.B1(n_1327),
.B2(n_1336),
.Y(n_1631)
);

INVxp33_ASAP7_75t_L g1632 ( 
.A(n_1600),
.Y(n_1632)
);

NAND3xp33_ASAP7_75t_SL g1633 ( 
.A(n_1578),
.B(n_1165),
.C(n_57),
.Y(n_1633)
);

NAND3xp33_ASAP7_75t_SL g1634 ( 
.A(n_1573),
.B(n_1574),
.C(n_1585),
.Y(n_1634)
);

NOR2xp67_ASAP7_75t_L g1635 ( 
.A(n_1609),
.B(n_59),
.Y(n_1635)
);

NOR4xp25_ASAP7_75t_L g1636 ( 
.A(n_1598),
.B(n_61),
.C(n_63),
.D(n_64),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1569),
.A2(n_1347),
.B1(n_1353),
.B2(n_1287),
.C(n_1282),
.Y(n_1637)
);

AOI22xp5_ASAP7_75t_L g1638 ( 
.A1(n_1589),
.A2(n_1353),
.B1(n_1287),
.B2(n_1293),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1590),
.B(n_1306),
.Y(n_1639)
);

AOI21x1_ASAP7_75t_L g1640 ( 
.A1(n_1601),
.A2(n_1174),
.B(n_1157),
.Y(n_1640)
);

OAI211xp5_ASAP7_75t_L g1641 ( 
.A1(n_1594),
.A2(n_1582),
.B(n_1592),
.C(n_1608),
.Y(n_1641)
);

NAND3xp33_ASAP7_75t_SL g1642 ( 
.A(n_1587),
.B(n_1588),
.C(n_1610),
.Y(n_1642)
);

OAI21xp33_ASAP7_75t_L g1643 ( 
.A1(n_1596),
.A2(n_1287),
.B(n_1306),
.Y(n_1643)
);

OAI211xp5_ASAP7_75t_L g1644 ( 
.A1(n_1595),
.A2(n_66),
.B(n_67),
.C(n_68),
.Y(n_1644)
);

AOI222xp33_ASAP7_75t_L g1645 ( 
.A1(n_1601),
.A2(n_1079),
.B1(n_69),
.B2(n_70),
.C1(n_71),
.C2(n_72),
.Y(n_1645)
);

AOI21xp33_ASAP7_75t_L g1646 ( 
.A1(n_1577),
.A2(n_66),
.B(n_69),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1597),
.Y(n_1647)
);

NAND3xp33_ASAP7_75t_L g1648 ( 
.A(n_1567),
.B(n_1201),
.C(n_73),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1607),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1605),
.A2(n_1343),
.B1(n_1307),
.B2(n_1306),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1605),
.Y(n_1651)
);

AOI21xp5_ASAP7_75t_L g1652 ( 
.A1(n_1566),
.A2(n_1132),
.B(n_1174),
.Y(n_1652)
);

AOI222xp33_ASAP7_75t_L g1653 ( 
.A1(n_1580),
.A2(n_1079),
.B1(n_74),
.B2(n_75),
.C1(n_77),
.C2(n_78),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1566),
.A2(n_1307),
.B1(n_1150),
.B2(n_1289),
.Y(n_1654)
);

OAI211xp5_ASAP7_75t_SL g1655 ( 
.A1(n_1568),
.A2(n_71),
.B(n_74),
.C(n_75),
.Y(n_1655)
);

OAI22xp33_ASAP7_75t_L g1656 ( 
.A1(n_1604),
.A2(n_1343),
.B1(n_1150),
.B2(n_1307),
.Y(n_1656)
);

OAI211xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1568),
.A2(n_77),
.B(n_79),
.C(n_81),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_SL g1658 ( 
.A1(n_1567),
.A2(n_1150),
.B(n_82),
.Y(n_1658)
);

BUFx2_ASAP7_75t_L g1659 ( 
.A(n_1571),
.Y(n_1659)
);

AOI221xp5_ASAP7_75t_L g1660 ( 
.A1(n_1566),
.A2(n_81),
.B1(n_83),
.B2(n_86),
.C(n_87),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1568),
.A2(n_1174),
.B(n_1157),
.Y(n_1661)
);

AOI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1566),
.A2(n_83),
.B1(n_86),
.B2(n_87),
.C(n_88),
.Y(n_1662)
);

OAI211xp5_ASAP7_75t_L g1663 ( 
.A1(n_1568),
.A2(n_1088),
.B(n_1066),
.C(n_1092),
.Y(n_1663)
);

AOI221x1_ASAP7_75t_SL g1664 ( 
.A1(n_1603),
.A2(n_1093),
.B1(n_1094),
.B2(n_1096),
.C(n_1145),
.Y(n_1664)
);

AOI321xp33_ASAP7_75t_L g1665 ( 
.A1(n_1567),
.A2(n_1158),
.A3(n_1156),
.B1(n_1142),
.B2(n_1149),
.C(n_1145),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1607),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1566),
.A2(n_1132),
.B1(n_1118),
.B2(n_1094),
.C(n_1096),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1605),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1649),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_SL g1670 ( 
.A(n_1666),
.B(n_1066),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1624),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1617),
.B(n_1118),
.Y(n_1672)
);

INVx2_ASAP7_75t_L g1673 ( 
.A(n_1659),
.Y(n_1673)
);

NOR2x1_ASAP7_75t_L g1674 ( 
.A(n_1651),
.B(n_1118),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1615),
.Y(n_1675)
);

NAND4xp75_ASAP7_75t_L g1676 ( 
.A(n_1614),
.B(n_1024),
.C(n_1084),
.D(n_1049),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1618),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1615),
.Y(n_1678)
);

NOR2x1_ASAP7_75t_L g1679 ( 
.A(n_1668),
.B(n_1118),
.Y(n_1679)
);

NAND4xp75_ASAP7_75t_L g1680 ( 
.A(n_1660),
.B(n_1039),
.C(n_1156),
.D(n_1149),
.Y(n_1680)
);

NAND4xp75_ASAP7_75t_L g1681 ( 
.A(n_1662),
.B(n_1161),
.C(n_124),
.D(n_125),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1625),
.Y(n_1682)
);

NAND4xp75_ASAP7_75t_L g1683 ( 
.A(n_1646),
.B(n_1628),
.C(n_1667),
.D(n_1635),
.Y(n_1683)
);

AOI211xp5_ASAP7_75t_SL g1684 ( 
.A1(n_1655),
.A2(n_122),
.B(n_126),
.C(n_127),
.Y(n_1684)
);

INVx2_ASAP7_75t_L g1685 ( 
.A(n_1618),
.Y(n_1685)
);

NAND2x1p5_ASAP7_75t_L g1686 ( 
.A(n_1627),
.B(n_1082),
.Y(n_1686)
);

AOI221xp5_ASAP7_75t_L g1687 ( 
.A1(n_1657),
.A2(n_1142),
.B1(n_1158),
.B2(n_1092),
.C(n_1161),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1626),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1636),
.B(n_131),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1639),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1647),
.Y(n_1691)
);

INVx1_ASAP7_75t_L g1692 ( 
.A(n_1632),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1648),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1629),
.Y(n_1694)
);

NAND4xp75_ASAP7_75t_L g1695 ( 
.A(n_1620),
.B(n_132),
.C(n_137),
.D(n_150),
.Y(n_1695)
);

NAND4xp75_ASAP7_75t_L g1696 ( 
.A(n_1652),
.B(n_153),
.C(n_157),
.D(n_160),
.Y(n_1696)
);

NOR2x1_ASAP7_75t_L g1697 ( 
.A(n_1644),
.B(n_162),
.Y(n_1697)
);

NAND2xp33_ASAP7_75t_L g1698 ( 
.A(n_1622),
.B(n_1158),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1634),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1641),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1664),
.Y(n_1701)
);

NOR2xp33_ASAP7_75t_L g1702 ( 
.A(n_1658),
.B(n_163),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1673),
.B(n_1619),
.Y(n_1703)
);

NOR3xp33_ASAP7_75t_SL g1704 ( 
.A(n_1682),
.B(n_1663),
.C(n_1642),
.Y(n_1704)
);

NAND2xp33_ASAP7_75t_SL g1705 ( 
.A(n_1675),
.B(n_1616),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_R g1706 ( 
.A(n_1689),
.B(n_1633),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_R g1707 ( 
.A(n_1692),
.B(n_1653),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1671),
.B(n_1645),
.Y(n_1708)
);

NAND2xp33_ASAP7_75t_SL g1709 ( 
.A(n_1678),
.B(n_1650),
.Y(n_1709)
);

NAND2xp33_ASAP7_75t_SL g1710 ( 
.A(n_1677),
.B(n_1661),
.Y(n_1710)
);

NOR2xp33_ASAP7_75t_R g1711 ( 
.A(n_1699),
.B(n_165),
.Y(n_1711)
);

NAND3xp33_ASAP7_75t_L g1712 ( 
.A(n_1669),
.B(n_1665),
.C(n_1637),
.Y(n_1712)
);

NAND2x1_ASAP7_75t_SL g1713 ( 
.A(n_1697),
.B(n_1654),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_SL g1714 ( 
.A(n_1685),
.B(n_1631),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_SL g1715 ( 
.A(n_1687),
.B(n_1623),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_SL g1716 ( 
.A(n_1684),
.B(n_1638),
.C(n_1630),
.Y(n_1716)
);

NAND3xp33_ASAP7_75t_L g1717 ( 
.A(n_1700),
.B(n_1621),
.C(n_1656),
.Y(n_1717)
);

NOR3xp33_ASAP7_75t_SL g1718 ( 
.A(n_1693),
.B(n_1643),
.C(n_168),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1688),
.B(n_1640),
.C(n_1142),
.Y(n_1719)
);

NAND2xp33_ASAP7_75t_SL g1720 ( 
.A(n_1694),
.B(n_1140),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1688),
.B(n_167),
.Y(n_1721)
);

NAND2xp33_ASAP7_75t_SL g1722 ( 
.A(n_1691),
.B(n_1140),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_R g1723 ( 
.A(n_1702),
.B(n_170),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1684),
.B(n_171),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_R g1725 ( 
.A(n_1702),
.B(n_175),
.Y(n_1725)
);

NOR2xp33_ASAP7_75t_R g1726 ( 
.A(n_1691),
.B(n_177),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_SL g1727 ( 
.A(n_1687),
.B(n_1146),
.Y(n_1727)
);

NOR2xp33_ASAP7_75t_R g1728 ( 
.A(n_1698),
.B(n_178),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_R g1729 ( 
.A(n_1698),
.B(n_181),
.Y(n_1729)
);

NOR2xp33_ASAP7_75t_R g1730 ( 
.A(n_1701),
.B(n_188),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_SL g1731 ( 
.A(n_1690),
.B(n_1146),
.Y(n_1731)
);

NAND3xp33_ASAP7_75t_L g1732 ( 
.A(n_1672),
.B(n_1144),
.C(n_1178),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_SL g1733 ( 
.A(n_1674),
.B(n_1679),
.Y(n_1733)
);

NOR3xp33_ASAP7_75t_SL g1734 ( 
.A(n_1683),
.B(n_189),
.C(n_193),
.Y(n_1734)
);

XNOR2xp5_ASAP7_75t_L g1735 ( 
.A(n_1681),
.B(n_1695),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1670),
.B(n_1696),
.C(n_1676),
.Y(n_1736)
);

NOR2xp33_ASAP7_75t_R g1737 ( 
.A(n_1680),
.B(n_196),
.Y(n_1737)
);

NAND2xp33_ASAP7_75t_SL g1738 ( 
.A(n_1670),
.B(n_1686),
.Y(n_1738)
);

NAND2xp33_ASAP7_75t_SL g1739 ( 
.A(n_1686),
.B(n_1144),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_R g1740 ( 
.A(n_1673),
.B(n_202),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1673),
.B(n_203),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1687),
.B(n_1146),
.Y(n_1742)
);

OAI22x1_ASAP7_75t_L g1743 ( 
.A1(n_1735),
.A2(n_1104),
.B1(n_1152),
.B2(n_1120),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1703),
.A2(n_1114),
.B1(n_1117),
.B2(n_1120),
.Y(n_1744)
);

OAI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1712),
.A2(n_1082),
.B(n_1007),
.Y(n_1745)
);

NAND3xp33_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1179),
.C(n_1178),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1708),
.B(n_205),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1734),
.B(n_206),
.Y(n_1748)
);

AOI211xp5_ASAP7_75t_L g1749 ( 
.A1(n_1709),
.A2(n_209),
.B(n_210),
.C(n_211),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1713),
.B(n_212),
.Y(n_1750)
);

NAND4xp25_ASAP7_75t_SL g1751 ( 
.A(n_1717),
.B(n_1179),
.C(n_1151),
.D(n_1154),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1728),
.B(n_1152),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1721),
.Y(n_1753)
);

INVx2_ASAP7_75t_L g1754 ( 
.A(n_1741),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1704),
.B(n_216),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1724),
.B(n_217),
.Y(n_1756)
);

XNOR2x1_ASAP7_75t_L g1757 ( 
.A(n_1736),
.B(n_220),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1733),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1706),
.Y(n_1759)
);

NOR3xp33_ASAP7_75t_L g1760 ( 
.A(n_1710),
.B(n_1104),
.C(n_1075),
.Y(n_1760)
);

AO22x2_ASAP7_75t_L g1761 ( 
.A1(n_1715),
.A2(n_1154),
.B1(n_1151),
.B2(n_1152),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1707),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1719),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1723),
.B(n_1725),
.Y(n_1764)
);

OAI22xp5_ASAP7_75t_SL g1765 ( 
.A1(n_1740),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_L g1766 ( 
.A(n_1726),
.B(n_226),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1762),
.Y(n_1767)
);

CKINVDCx20_ASAP7_75t_R g1768 ( 
.A(n_1759),
.Y(n_1768)
);

AOI22xp33_ASAP7_75t_SL g1769 ( 
.A1(n_1758),
.A2(n_1730),
.B1(n_1729),
.B2(n_1737),
.Y(n_1769)
);

INVx2_ASAP7_75t_SL g1770 ( 
.A(n_1750),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1748),
.B(n_1718),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1747),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1756),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1766),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1757),
.Y(n_1775)
);

AOI21xp33_ASAP7_75t_L g1776 ( 
.A1(n_1764),
.A2(n_1731),
.B(n_1732),
.Y(n_1776)
);

AND2x2_ASAP7_75t_SL g1777 ( 
.A(n_1755),
.B(n_1711),
.Y(n_1777)
);

HB1xp67_ASAP7_75t_L g1778 ( 
.A(n_1765),
.Y(n_1778)
);

AND2x4_ASAP7_75t_L g1779 ( 
.A(n_1754),
.B(n_1742),
.Y(n_1779)
);

OAI21xp5_ASAP7_75t_L g1780 ( 
.A1(n_1746),
.A2(n_1714),
.B(n_1716),
.Y(n_1780)
);

NAND4xp25_ASAP7_75t_L g1781 ( 
.A(n_1749),
.B(n_1763),
.C(n_1753),
.D(n_1745),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1744),
.A2(n_1752),
.B1(n_1761),
.B2(n_1727),
.Y(n_1782)
);

AOI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1751),
.A2(n_1738),
.B1(n_1720),
.B2(n_1739),
.Y(n_1783)
);

INVx1_ASAP7_75t_L g1784 ( 
.A(n_1761),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1769),
.B(n_1760),
.C(n_1722),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1768),
.Y(n_1786)
);

OAI22xp5_ASAP7_75t_L g1787 ( 
.A1(n_1767),
.A2(n_1737),
.B1(n_1743),
.B2(n_1114),
.Y(n_1787)
);

OR2x2_ASAP7_75t_L g1788 ( 
.A(n_1771),
.B(n_230),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1778),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1770),
.A2(n_1117),
.B1(n_1120),
.B2(n_1162),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1780),
.Y(n_1791)
);

AO22x2_ASAP7_75t_L g1792 ( 
.A1(n_1775),
.A2(n_1772),
.B1(n_1774),
.B2(n_1773),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1777),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_SL g1794 ( 
.A1(n_1786),
.A2(n_1789),
.B1(n_1791),
.B2(n_1793),
.Y(n_1794)
);

AOI31xp33_ASAP7_75t_L g1795 ( 
.A1(n_1788),
.A2(n_1776),
.A3(n_1779),
.B(n_1784),
.Y(n_1795)
);

AOI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1792),
.A2(n_1779),
.B1(n_1781),
.B2(n_1782),
.Y(n_1796)
);

AOI31xp33_ASAP7_75t_L g1797 ( 
.A1(n_1785),
.A2(n_1783),
.A3(n_237),
.B(n_238),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_SL g1798 ( 
.A1(n_1795),
.A2(n_1787),
.B1(n_1792),
.B2(n_1790),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1794),
.B(n_233),
.Y(n_1799)
);

XOR2xp5_ASAP7_75t_L g1800 ( 
.A(n_1796),
.B(n_239),
.Y(n_1800)
);

AO22x2_ASAP7_75t_L g1801 ( 
.A1(n_1797),
.A2(n_242),
.B1(n_247),
.B2(n_250),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1799),
.A2(n_254),
.B(n_257),
.Y(n_1802)
);

OAI31xp33_ASAP7_75t_SL g1803 ( 
.A1(n_1800),
.A2(n_259),
.A3(n_262),
.B(n_263),
.Y(n_1803)
);

OR2x2_ASAP7_75t_L g1804 ( 
.A(n_1798),
.B(n_264),
.Y(n_1804)
);

OAI222xp33_ASAP7_75t_L g1805 ( 
.A1(n_1801),
.A2(n_1117),
.B1(n_1171),
.B2(n_1162),
.C1(n_1095),
.C2(n_1141),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1804),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1802),
.Y(n_1807)
);

HB1xp67_ASAP7_75t_L g1808 ( 
.A(n_1803),
.Y(n_1808)
);

OAI221xp5_ASAP7_75t_R g1809 ( 
.A1(n_1808),
.A2(n_1805),
.B1(n_267),
.B2(n_269),
.C(n_274),
.Y(n_1809)
);

AOI211xp5_ASAP7_75t_L g1810 ( 
.A1(n_1809),
.A2(n_1806),
.B(n_1807),
.C(n_282),
.Y(n_1810)
);


endmodule