module fake_jpeg_11888_n_172 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_172);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_172;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g49 ( 
.A(n_16),
.Y(n_49)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_1),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_26),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_0),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_31),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_19),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_32),
.B(n_43),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_27),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_6),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_14),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_17),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_11),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_48),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_67),
.B(n_0),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_76),
.B(n_80),
.Y(n_90)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_78),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_79),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_56),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g81 ( 
.A(n_70),
.B(n_1),
.CON(n_81),
.SN(n_81)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_81),
.B(n_82),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_2),
.Y(n_82)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_50),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_84),
.Y(n_88)
);

OA22x2_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_73),
.B1(n_52),
.B2(n_62),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_54),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_73),
.B1(n_50),
.B2(n_51),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_92),
.A2(n_99),
.B1(n_63),
.B2(n_54),
.Y(n_107)
);

CKINVDCx12_ASAP7_75t_R g93 ( 
.A(n_80),
.Y(n_93)
);

INVx4_ASAP7_75t_SL g102 ( 
.A(n_93),
.Y(n_102)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_81),
.Y(n_94)
);

OR2x2_ASAP7_75t_L g105 ( 
.A(n_94),
.B(n_61),
.Y(n_105)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_77),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_96),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_84),
.A2(n_63),
.B1(n_51),
.B2(n_70),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_100),
.A2(n_59),
.B1(n_113),
.B2(n_109),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_90),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_106),
.Y(n_120)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_103),
.Y(n_126)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_95),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_104),
.B(n_108),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_72),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_107),
.A2(n_116),
.B1(n_4),
.B2(n_5),
.Y(n_131)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_111),
.B(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_86),
.A2(n_88),
.B1(n_89),
.B2(n_99),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_113),
.A2(n_59),
.B1(n_68),
.B2(n_66),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_74),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_114),
.B(n_117),
.Y(n_123)
);

OAI22x1_ASAP7_75t_SL g116 ( 
.A1(n_86),
.A2(n_49),
.B1(n_71),
.B2(n_69),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_60),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_119),
.Y(n_130)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_122),
.A2(n_133),
.B1(n_8),
.B2(n_9),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_105),
.B(n_65),
.C(n_64),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_129),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g125 ( 
.A1(n_109),
.A2(n_21),
.B(n_46),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_115),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_128),
.A2(n_131),
.B1(n_10),
.B2(n_11),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_102),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_113),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_10),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_130),
.A2(n_126),
.B1(n_121),
.B2(n_127),
.Y(n_137)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_127),
.Y(n_138)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_132),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_140),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_135),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_143),
.A2(n_124),
.B1(n_13),
.B2(n_30),
.Y(n_148)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_144),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_120),
.B(n_12),
.Y(n_145)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_145),
.Y(n_156)
);

INVx13_ASAP7_75t_L g146 ( 
.A(n_125),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_146),
.A2(n_147),
.B1(n_29),
.B2(n_33),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_13),
.B(n_22),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_149),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_137),
.A2(n_45),
.B1(n_37),
.B2(n_39),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

OA22x2_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_34),
.B1(n_41),
.B2(n_42),
.Y(n_153)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_153),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_160),
.B(n_161),
.Y(n_162)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_154),
.Y(n_161)
);

INVx13_ASAP7_75t_L g163 ( 
.A(n_159),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_163),
.B(n_164),
.C(n_142),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_142),
.Y(n_164)
);

O2A1O1Ixp33_ASAP7_75t_L g166 ( 
.A1(n_165),
.A2(n_155),
.B(n_157),
.C(n_158),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_166),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_167),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_168),
.B(n_162),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_169),
.A2(n_152),
.B1(n_156),
.B2(n_149),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_153),
.C(n_148),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_150),
.Y(n_172)
);


endmodule