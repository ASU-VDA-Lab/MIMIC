module real_aes_109_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_503;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_753;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_0), .B(n_140), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_1), .A2(n_148), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g772 ( .A(n_2), .B(n_773), .Y(n_772) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_3), .B(n_140), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_4), .B(n_167), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g493 ( .A(n_5), .B(n_167), .Y(n_493) );
INVx1_ASAP7_75t_L g136 ( .A(n_6), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_7), .B(n_167), .Y(n_542) );
CKINVDCx16_ASAP7_75t_R g773 ( .A(n_8), .Y(n_773) );
OAI22xp33_ASAP7_75t_SL g761 ( .A1(n_9), .A2(n_115), .B1(n_745), .B2(n_762), .Y(n_761) );
CKINVDCx20_ASAP7_75t_R g762 ( .A(n_9), .Y(n_762) );
NAND2xp33_ASAP7_75t_L g534 ( .A(n_10), .B(n_165), .Y(n_534) );
AND2x2_ASAP7_75t_L g170 ( .A(n_11), .B(n_171), .Y(n_170) );
AND2x2_ASAP7_75t_L g181 ( .A(n_12), .B(n_182), .Y(n_181) );
INVx2_ASAP7_75t_L g127 ( .A(n_13), .Y(n_127) );
AOI221x1_ASAP7_75t_L g478 ( .A1(n_14), .A2(n_25), .B1(n_140), .B2(n_148), .C(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_15), .B(n_167), .Y(n_207) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_16), .Y(n_107) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_17), .B(n_140), .Y(n_530) );
AO21x2_ASAP7_75t_L g528 ( .A1(n_18), .A2(n_182), .B(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_19), .B(n_125), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_20), .B(n_167), .Y(n_467) );
AO21x1_ASAP7_75t_L g488 ( .A1(n_21), .A2(n_140), .B(n_489), .Y(n_488) );
NAND2xp5_ASAP7_75t_SL g223 ( .A(n_22), .B(n_140), .Y(n_223) );
INVx1_ASAP7_75t_L g111 ( .A(n_23), .Y(n_111) );
AOI22xp33_ASAP7_75t_L g130 ( .A1(n_24), .A2(n_88), .B1(n_131), .B2(n_140), .Y(n_130) );
NAND2x1_ASAP7_75t_L g509 ( .A(n_26), .B(n_167), .Y(n_509) );
NAND2x1_ASAP7_75t_L g541 ( .A(n_27), .B(n_165), .Y(n_541) );
OR2x2_ASAP7_75t_L g128 ( .A(n_28), .B(n_85), .Y(n_128) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_28), .A2(n_85), .B(n_127), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_29), .B(n_165), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_30), .B(n_167), .Y(n_533) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_31), .A2(n_171), .B(n_203), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_32), .B(n_165), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_33), .A2(n_148), .B(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_34), .B(n_167), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_35), .A2(n_148), .B(n_499), .Y(n_498) );
AND2x2_ASAP7_75t_L g138 ( .A(n_36), .B(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g146 ( .A(n_36), .B(n_136), .Y(n_146) );
INVx1_ASAP7_75t_L g152 ( .A(n_36), .Y(n_152) );
OR2x6_ASAP7_75t_L g109 ( .A(n_37), .B(n_110), .Y(n_109) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_37), .B(n_772), .C(n_774), .Y(n_771) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_38), .B(n_140), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_39), .B(n_140), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_40), .B(n_167), .Y(n_218) );
CKINVDCx20_ASAP7_75t_R g471 ( .A(n_41), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_42), .B(n_165), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_43), .B(n_140), .Y(n_189) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_44), .Y(n_104) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_45), .A2(n_148), .B(n_163), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_46), .A2(n_148), .B(n_540), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_47), .B(n_165), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_48), .B(n_165), .Y(n_510) );
NAND2xp5_ASAP7_75t_SL g204 ( .A(n_49), .B(n_140), .Y(n_204) );
INVx1_ASAP7_75t_L g134 ( .A(n_50), .Y(n_134) );
INVx1_ASAP7_75t_L g143 ( .A(n_50), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_51), .B(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g213 ( .A(n_52), .B(n_125), .Y(n_213) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_53), .B(n_165), .Y(n_164) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_54), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_55), .B(n_167), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_56), .B(n_165), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g507 ( .A1(n_57), .A2(n_148), .B(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_58), .B(n_140), .Y(n_169) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_59), .B(n_140), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g234 ( .A1(n_60), .A2(n_148), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g229 ( .A(n_61), .B(n_126), .Y(n_229) );
AO21x1_ASAP7_75t_L g490 ( .A1(n_62), .A2(n_148), .B(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_63), .B(n_140), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_64), .B(n_165), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g543 ( .A(n_65), .B(n_140), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_66), .B(n_165), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g147 ( .A1(n_67), .A2(n_92), .B1(n_148), .B2(n_150), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g777 ( .A(n_68), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_69), .B(n_167), .Y(n_226) );
AND2x2_ASAP7_75t_L g503 ( .A(n_70), .B(n_126), .Y(n_503) );
INVx1_ASAP7_75t_L g139 ( .A(n_71), .Y(n_139) );
INVx1_ASAP7_75t_L g145 ( .A(n_71), .Y(n_145) );
AND2x2_ASAP7_75t_L g544 ( .A(n_72), .B(n_171), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_73), .B(n_165), .Y(n_178) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_74), .A2(n_148), .B(n_217), .Y(n_216) );
AOI221xp5_ASAP7_75t_L g113 ( .A1(n_75), .A2(n_114), .B1(n_743), .B2(n_744), .C(n_748), .Y(n_113) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_75), .Y(n_743) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_76), .A2(n_148), .B(n_191), .Y(n_190) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_77), .A2(n_148), .B(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_L g239 ( .A(n_78), .B(n_126), .Y(n_239) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_79), .B(n_125), .Y(n_124) );
INVx1_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
NOR2xp33_ASAP7_75t_L g775 ( .A(n_80), .B(n_111), .Y(n_775) );
AND2x2_ASAP7_75t_L g455 ( .A(n_81), .B(n_171), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g469 ( .A(n_82), .B(n_140), .Y(n_469) );
AND2x2_ASAP7_75t_L g194 ( .A(n_83), .B(n_182), .Y(n_194) );
AND2x2_ASAP7_75t_L g489 ( .A(n_84), .B(n_209), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_86), .B(n_165), .Y(n_468) );
AND2x2_ASAP7_75t_L g512 ( .A(n_87), .B(n_171), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_89), .B(n_167), .Y(n_501) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_90), .A2(n_148), .B(n_466), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_91), .B(n_165), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_93), .A2(n_148), .B(n_225), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_94), .B(n_167), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_95), .B(n_167), .Y(n_460) );
BUFx2_ASAP7_75t_L g228 ( .A(n_96), .Y(n_228) );
BUFx2_ASAP7_75t_L g757 ( .A(n_97), .Y(n_757) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_98), .A2(n_148), .B(n_532), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g99 ( .A1(n_100), .A2(n_766), .B(n_776), .Y(n_99) );
AO21x2_ASAP7_75t_L g100 ( .A1(n_101), .A2(n_753), .B(n_758), .Y(n_100) );
NAND2xp5_ASAP7_75t_L g101 ( .A(n_102), .B(n_113), .Y(n_101) );
CKINVDCx16_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
AOI21xp5_ASAP7_75t_L g760 ( .A1(n_103), .A2(n_761), .B(n_763), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
BUFx3_ASAP7_75t_L g765 ( .A(n_106), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_108), .Y(n_106) );
AND2x6_ASAP7_75t_SL g447 ( .A(n_107), .B(n_109), .Y(n_447) );
OR2x6_ASAP7_75t_SL g742 ( .A(n_107), .B(n_108), .Y(n_742) );
OR2x2_ASAP7_75t_L g752 ( .A(n_107), .B(n_109), .Y(n_752) );
CKINVDCx16_ASAP7_75t_R g774 ( .A(n_107), .Y(n_774) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_112), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_444), .B1(n_448), .B2(n_740), .Y(n_114) );
INVx3_ASAP7_75t_L g745 ( .A(n_115), .Y(n_745) );
AND2x4_ASAP7_75t_L g115 ( .A(n_116), .B(n_369), .Y(n_115) );
NOR3xp33_ASAP7_75t_L g116 ( .A(n_117), .B(n_305), .C(n_352), .Y(n_116) );
NAND4xp25_ASAP7_75t_SL g117 ( .A(n_118), .B(n_240), .C(n_258), .D(n_284), .Y(n_117) );
OAI21xp33_ASAP7_75t_SL g118 ( .A1(n_119), .A2(n_198), .B(n_199), .Y(n_118) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_120), .B(n_183), .Y(n_119) );
INVx1_ASAP7_75t_L g420 ( .A(n_120), .Y(n_420) );
OR2x2_ASAP7_75t_L g120 ( .A(n_121), .B(n_155), .Y(n_120) );
INVx2_ASAP7_75t_L g244 ( .A(n_121), .Y(n_244) );
AND2x2_ASAP7_75t_L g264 ( .A(n_121), .B(n_265), .Y(n_264) );
OR2x2_ASAP7_75t_L g366 ( .A(n_121), .B(n_185), .Y(n_366) );
AND2x2_ASAP7_75t_L g426 ( .A(n_121), .B(n_245), .Y(n_426) );
INVx2_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_122), .B(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
OR2x2_ASAP7_75t_L g310 ( .A(n_123), .B(n_158), .Y(n_310) );
BUFx3_ASAP7_75t_L g320 ( .A(n_123), .Y(n_320) );
AND2x2_ASAP7_75t_L g383 ( .A(n_123), .B(n_384), .Y(n_383) );
AND2x4_ASAP7_75t_L g123 ( .A(n_124), .B(n_129), .Y(n_123) );
AND2x4_ASAP7_75t_L g197 ( .A(n_124), .B(n_129), .Y(n_197) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_125), .A2(n_130), .B(n_147), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_125), .Y(n_174) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_125), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g456 ( .A1(n_125), .A2(n_457), .B(n_458), .Y(n_456) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_125), .A2(n_478), .B(n_482), .Y(n_477) );
OA21x2_ASAP7_75t_L g548 ( .A1(n_125), .A2(n_478), .B(n_482), .Y(n_548) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
AND2x2_ASAP7_75t_SL g126 ( .A(n_127), .B(n_128), .Y(n_126) );
AND2x4_ASAP7_75t_L g209 ( .A(n_127), .B(n_128), .Y(n_209) );
AND2x4_ASAP7_75t_L g131 ( .A(n_132), .B(n_137), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g149 ( .A(n_134), .B(n_136), .Y(n_149) );
AND2x4_ASAP7_75t_L g167 ( .A(n_134), .B(n_144), .Y(n_167) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
BUFx3_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x6_ASAP7_75t_L g148 ( .A(n_138), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g154 ( .A(n_139), .Y(n_154) );
AND2x6_ASAP7_75t_L g165 ( .A(n_139), .B(n_142), .Y(n_165) );
AND2x4_ASAP7_75t_L g140 ( .A(n_141), .B(n_146), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx5_ASAP7_75t_L g168 ( .A(n_146), .Y(n_168) );
AND2x4_ASAP7_75t_L g150 ( .A(n_149), .B(n_151), .Y(n_150) );
NOR2x1p5_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
INVx3_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_SL g155 ( .A(n_156), .Y(n_155) );
INVx1_ASAP7_75t_L g429 ( .A(n_156), .Y(n_429) );
AND2x2_ASAP7_75t_L g156 ( .A(n_157), .B(n_172), .Y(n_156) );
AND2x2_ASAP7_75t_L g196 ( .A(n_157), .B(n_197), .Y(n_196) );
INVx1_ASAP7_75t_L g384 ( .A(n_157), .Y(n_384) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g198 ( .A(n_158), .B(n_187), .Y(n_198) );
AND2x2_ASAP7_75t_L g261 ( .A(n_158), .B(n_172), .Y(n_261) );
INVx2_ASAP7_75t_L g266 ( .A(n_158), .Y(n_266) );
AND2x2_ASAP7_75t_L g268 ( .A(n_158), .B(n_173), .Y(n_268) );
AO21x2_ASAP7_75t_L g158 ( .A1(n_159), .A2(n_161), .B(n_170), .Y(n_158) );
INVx4_ASAP7_75t_L g171 ( .A(n_159), .Y(n_171) );
INVx3_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
BUFx4f_ASAP7_75t_L g182 ( .A(n_160), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_162), .B(n_169), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_168), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_165), .B(n_228), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g177 ( .A1(n_168), .A2(n_178), .B(n_179), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_168), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_168), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_168), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g225 ( .A1(n_168), .A2(n_226), .B(n_227), .Y(n_225) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_168), .A2(n_236), .B(n_237), .Y(n_235) );
AOI21xp5_ASAP7_75t_L g459 ( .A1(n_168), .A2(n_460), .B(n_461), .Y(n_459) );
AOI21xp5_ASAP7_75t_L g466 ( .A1(n_168), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_168), .A2(n_480), .B(n_481), .Y(n_479) );
AOI21xp5_ASAP7_75t_L g491 ( .A1(n_168), .A2(n_492), .B(n_493), .Y(n_491) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_168), .A2(n_500), .B(n_501), .Y(n_499) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_168), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_168), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_168), .A2(n_541), .B(n_542), .Y(n_540) );
INVx3_ASAP7_75t_L g232 ( .A(n_171), .Y(n_232) );
INVx1_ASAP7_75t_L g246 ( .A(n_172), .Y(n_246) );
INVx2_ASAP7_75t_L g250 ( .A(n_172), .Y(n_250) );
AND2x4_ASAP7_75t_SL g281 ( .A(n_172), .B(n_187), .Y(n_281) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_172), .Y(n_313) );
INVx3_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
HB1xp67_ASAP7_75t_L g195 ( .A(n_173), .Y(n_195) );
AOI21x1_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_181), .Y(n_173) );
AO21x2_ASAP7_75t_L g537 ( .A1(n_174), .A2(n_538), .B(n_544), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_176), .B(n_180), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g222 ( .A1(n_182), .A2(n_223), .B(n_224), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_184), .B(n_196), .Y(n_183) );
AND2x2_ASAP7_75t_L g347 ( .A(n_184), .B(n_292), .Y(n_347) );
INVx2_ASAP7_75t_SL g435 ( .A(n_184), .Y(n_435) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_186), .B(n_195), .Y(n_185) );
NAND2x1p5_ASAP7_75t_L g248 ( .A(n_186), .B(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g355 ( .A(n_186), .B(n_268), .Y(n_355) );
INVx4_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx2_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
AND2x4_ASAP7_75t_L g245 ( .A(n_187), .B(n_246), .Y(n_245) );
NOR2x1_ASAP7_75t_L g265 ( .A(n_187), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_L g338 ( .A(n_187), .Y(n_338) );
AND2x2_ASAP7_75t_L g357 ( .A(n_187), .B(n_296), .Y(n_357) );
AND2x2_ASAP7_75t_L g388 ( .A(n_187), .B(n_297), .Y(n_388) );
OR2x6_ASAP7_75t_L g187 ( .A(n_188), .B(n_194), .Y(n_187) );
AND2x2_ASAP7_75t_L g327 ( .A(n_196), .B(n_281), .Y(n_327) );
NAND2xp5_ASAP7_75t_SL g363 ( .A(n_196), .B(n_338), .Y(n_363) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_196), .A2(n_438), .B1(n_440), .B2(n_441), .Y(n_437) );
AND2x2_ASAP7_75t_L g440 ( .A(n_196), .B(n_247), .Y(n_440) );
INVx3_ASAP7_75t_L g293 ( .A(n_197), .Y(n_293) );
AND2x2_ASAP7_75t_L g296 ( .A(n_197), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g312 ( .A(n_198), .B(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g321 ( .A(n_198), .Y(n_321) );
AND2x4_ASAP7_75t_SL g199 ( .A(n_200), .B(n_210), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_200), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g372 ( .A(n_200), .B(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_200), .B(n_334), .C(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g442 ( .A(n_200), .B(n_336), .Y(n_442) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g257 ( .A(n_202), .B(n_221), .Y(n_257) );
INVx1_ASAP7_75t_L g274 ( .A(n_202), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_202), .Y(n_287) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_202), .Y(n_302) );
AND2x2_ASAP7_75t_L g316 ( .A(n_202), .B(n_289), .Y(n_316) );
AND2x2_ASAP7_75t_L g395 ( .A(n_202), .B(n_212), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_204), .A2(n_205), .B(n_209), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_209), .A2(n_215), .B(n_216), .Y(n_214) );
INVx1_ASAP7_75t_SL g463 ( .A(n_209), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g494 ( .A(n_209), .B(n_495), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_209), .A2(n_530), .B(n_531), .Y(n_529) );
AOI221xp5_ASAP7_75t_L g258 ( .A1(n_210), .A2(n_259), .B1(n_262), .B2(n_269), .C(n_275), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g387 ( .A1(n_210), .A2(n_388), .B1(n_389), .B2(n_390), .C(n_391), .Y(n_387) );
AND2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_220), .Y(n_210) );
INVx2_ASAP7_75t_L g329 ( .A(n_211), .Y(n_329) );
AND2x2_ASAP7_75t_L g389 ( .A(n_211), .B(n_273), .Y(n_389) );
AND2x2_ASAP7_75t_L g399 ( .A(n_211), .B(n_285), .Y(n_399) );
OR2x2_ASAP7_75t_L g439 ( .A(n_211), .B(n_323), .Y(n_439) );
INVx2_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
OR2x2_ASAP7_75t_SL g256 ( .A(n_212), .B(n_257), .Y(n_256) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_212), .B(n_221), .Y(n_272) );
INVx4_ASAP7_75t_L g301 ( .A(n_212), .Y(n_301) );
OR2x2_ASAP7_75t_L g343 ( .A(n_212), .B(n_230), .Y(n_343) );
OR2x6_ASAP7_75t_L g212 ( .A(n_213), .B(n_214), .Y(n_212) );
AND2x2_ASAP7_75t_L g394 ( .A(n_220), .B(n_395), .Y(n_394) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_230), .Y(n_220) );
INVx2_ASAP7_75t_SL g282 ( .A(n_221), .Y(n_282) );
NOR2x1_ASAP7_75t_SL g288 ( .A(n_221), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g303 ( .A(n_221), .B(n_304), .Y(n_303) );
OR2x2_ASAP7_75t_L g334 ( .A(n_221), .B(n_301), .Y(n_334) );
AND2x2_ASAP7_75t_L g341 ( .A(n_221), .B(n_287), .Y(n_341) );
BUFx2_ASAP7_75t_L g375 ( .A(n_221), .Y(n_375) );
AND2x2_ASAP7_75t_L g386 ( .A(n_221), .B(n_301), .Y(n_386) );
OR2x6_ASAP7_75t_L g221 ( .A(n_222), .B(n_229), .Y(n_221) );
HB1xp67_ASAP7_75t_L g254 ( .A(n_230), .Y(n_254) );
AND2x2_ASAP7_75t_L g273 ( .A(n_230), .B(n_274), .Y(n_273) );
INVx2_ASAP7_75t_L g304 ( .A(n_230), .Y(n_304) );
AND2x2_ASAP7_75t_L g330 ( .A(n_230), .B(n_286), .Y(n_330) );
INVx3_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
AO21x2_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_231) );
AO21x1_ASAP7_75t_SL g289 ( .A1(n_232), .A2(n_233), .B(n_239), .Y(n_289) );
AO21x2_ASAP7_75t_L g496 ( .A1(n_232), .A2(n_497), .B(n_503), .Y(n_496) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_232), .A2(n_506), .B(n_512), .Y(n_505) );
AO21x2_ASAP7_75t_L g518 ( .A1(n_232), .A2(n_506), .B(n_512), .Y(n_518) );
AO21x2_ASAP7_75t_L g521 ( .A1(n_232), .A2(n_497), .B(n_503), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_234), .B(n_238), .Y(n_233) );
OAI31xp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_245), .A3(n_247), .B(n_251), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
INVx2_ASAP7_75t_L g349 ( .A(n_243), .Y(n_349) );
NOR2xp67_ASAP7_75t_L g259 ( .A(n_244), .B(n_260), .Y(n_259) );
AOI322xp5_ASAP7_75t_L g339 ( .A1(n_244), .A2(n_333), .A3(n_340), .B1(n_344), .B2(n_345), .C1(n_347), .C2(n_348), .Y(n_339) );
AND2x2_ASAP7_75t_L g411 ( .A(n_244), .B(n_388), .Y(n_411) );
AOI221xp5_ASAP7_75t_SL g324 ( .A1(n_245), .A2(n_325), .B1(n_327), .B2(n_328), .C(n_331), .Y(n_324) );
INVx2_ASAP7_75t_L g344 ( .A(n_245), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_247), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_247), .B(n_340), .Y(n_443) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
OR2x2_ASAP7_75t_L g318 ( .A(n_248), .B(n_293), .Y(n_318) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
AND2x2_ASAP7_75t_L g297 ( .A(n_250), .B(n_266), .Y(n_297) );
AND2x4_ASAP7_75t_L g251 ( .A(n_252), .B(n_255), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
INVx1_ASAP7_75t_L g368 ( .A(n_254), .Y(n_368) );
O2A1O1Ixp5_ASAP7_75t_L g359 ( .A1(n_255), .A2(n_360), .B(n_362), .C(n_364), .Y(n_359) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_256), .A2(n_392), .B1(n_393), .B2(n_396), .Y(n_391) );
OR2x2_ASAP7_75t_L g346 ( .A(n_257), .B(n_343), .Y(n_346) );
INVx1_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g262 ( .A(n_263), .B(n_267), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g279 ( .A(n_266), .Y(n_279) );
INVx1_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_268), .B(n_292), .Y(n_291) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx3_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g322 ( .A(n_272), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_272), .B(n_273), .Y(n_365) );
OR2x2_ASAP7_75t_L g367 ( .A(n_272), .B(n_368), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g415 ( .A(n_272), .B(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g283 ( .A(n_274), .Y(n_283) );
NOR4xp25_ASAP7_75t_L g275 ( .A(n_276), .B(n_280), .C(n_282), .D(n_283), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g403 ( .A(n_277), .B(n_404), .Y(n_403) );
AND2x2_ASAP7_75t_L g431 ( .A(n_277), .B(n_280), .Y(n_431) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g361 ( .A(n_279), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_280), .B(n_309), .Y(n_396) );
AOI321xp33_ASAP7_75t_L g398 ( .A1(n_280), .A2(n_399), .A3(n_400), .B1(n_401), .B2(n_403), .C(n_406), .Y(n_398) );
INVx2_ASAP7_75t_SL g280 ( .A(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_SL g360 ( .A(n_281), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_281), .B(n_320), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_282), .B(n_304), .Y(n_409) );
OR2x2_ASAP7_75t_L g436 ( .A(n_283), .B(n_320), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_285), .A2(n_290), .B(n_294), .Y(n_284) );
AND2x2_ASAP7_75t_L g325 ( .A(n_285), .B(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g351 ( .A(n_287), .B(n_289), .Y(n_351) );
INVx2_ASAP7_75t_L g336 ( .A(n_288), .Y(n_336) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_291), .B(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g392 ( .A(n_292), .B(n_344), .Y(n_392) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
AND2x2_ASAP7_75t_L g350 ( .A(n_293), .B(n_351), .Y(n_350) );
NOR2x1_ASAP7_75t_L g428 ( .A(n_293), .B(n_429), .Y(n_428) );
NOR2xp67_ASAP7_75t_L g294 ( .A(n_295), .B(n_298), .Y(n_294) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g379 ( .A(n_297), .Y(n_379) );
INVx2_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .Y(n_299) );
NOR2xp67_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_301), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g326 ( .A(n_301), .Y(n_326) );
BUFx2_ASAP7_75t_L g408 ( .A(n_301), .Y(n_408) );
INVxp67_ASAP7_75t_L g416 ( .A(n_304), .Y(n_416) );
NAND3xp33_ASAP7_75t_L g305 ( .A(n_306), .B(n_324), .C(n_339), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_307), .A2(n_314), .B(n_317), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_308), .B(n_311), .Y(n_307) );
INVx2_ASAP7_75t_SL g309 ( .A(n_310), .Y(n_309) );
OR2x2_ASAP7_75t_L g337 ( .A(n_310), .B(n_338), .Y(n_337) );
INVx2_ASAP7_75t_L g390 ( .A(n_311), .Y(n_390) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx2_ASAP7_75t_L g405 ( .A(n_313), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_314), .A2(n_411), .B(n_412), .Y(n_410) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
INVx2_ASAP7_75t_SL g323 ( .A(n_316), .Y(n_323) );
AND2x2_ASAP7_75t_L g385 ( .A(n_316), .B(n_386), .Y(n_385) );
AOI21xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B(n_322), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_318), .A2(n_365), .B1(n_366), .B2(n_367), .Y(n_364) );
OR2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_321), .Y(n_319) );
INVx1_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
OR2x2_ASAP7_75t_L g402 ( .A(n_323), .B(n_334), .Y(n_402) );
NOR4xp25_ASAP7_75t_L g434 ( .A(n_326), .B(n_375), .C(n_435), .D(n_436), .Y(n_434) );
AND2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
OR2x2_ASAP7_75t_L g335 ( .A(n_329), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_329), .B(n_351), .Y(n_433) );
AOI21xp33_ASAP7_75t_SL g331 ( .A1(n_332), .A2(n_335), .B(n_337), .Y(n_331) );
INVx2_ASAP7_75t_SL g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g422 ( .A(n_334), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g430 ( .A(n_336), .Y(n_430) );
AND2x4_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
INVxp67_ASAP7_75t_L g358 ( .A(n_341), .Y(n_358) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g374 ( .A(n_343), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AND2x2_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
AND2x2_ASAP7_75t_L g377 ( .A(n_349), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g423 ( .A(n_351), .Y(n_423) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_356), .B(n_358), .C(n_359), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g413 ( .A(n_355), .Y(n_413) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVxp67_ASAP7_75t_L g417 ( .A(n_360), .Y(n_417) );
INVx1_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
NOR3xp33_ASAP7_75t_L g369 ( .A(n_370), .B(n_397), .C(n_418), .Y(n_369) );
OAI211xp5_ASAP7_75t_SL g370 ( .A1(n_371), .A2(n_376), .B(n_380), .C(n_387), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
INVxp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g380 ( .A1(n_381), .A2(n_383), .B(n_385), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
O2A1O1Ixp33_ASAP7_75t_L g419 ( .A1(n_383), .A2(n_420), .B(n_421), .C(n_424), .Y(n_419) );
BUFx2_ASAP7_75t_L g400 ( .A(n_384), .Y(n_400) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_398), .B(n_410), .Y(n_397) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_407), .A2(n_413), .B1(n_414), .B2(n_417), .Y(n_412) );
OR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_409), .Y(n_407) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND4xp25_ASAP7_75t_L g418 ( .A(n_419), .B(n_427), .C(n_437), .D(n_443), .Y(n_418) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
AOI221xp5_ASAP7_75t_L g427 ( .A1(n_428), .A2(n_430), .B1(n_431), .B2(n_432), .C(n_434), .Y(n_427) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
CKINVDCx6p67_ASAP7_75t_R g444 ( .A(n_445), .Y(n_444) );
INVx3_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_446), .A2(n_745), .B1(n_746), .B2(n_747), .Y(n_744) );
CKINVDCx5p33_ASAP7_75t_R g446 ( .A(n_447), .Y(n_446) );
INVx3_ASAP7_75t_SL g747 ( .A(n_448), .Y(n_747) );
NOR2x2_ASAP7_75t_L g448 ( .A(n_449), .B(n_627), .Y(n_448) );
AO211x2_ASAP7_75t_L g449 ( .A1(n_450), .A2(n_472), .B(n_522), .C(n_595), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVxp67_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AND3x2_ASAP7_75t_L g676 ( .A(n_452), .B(n_557), .C(n_573), .Y(n_676) );
AND2x4_ASAP7_75t_L g679 ( .A(n_452), .B(n_680), .Y(n_679) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_462), .Y(n_452) );
NAND2x1p5_ASAP7_75t_L g535 ( .A(n_453), .B(n_536), .Y(n_535) );
INVx4_ASAP7_75t_L g588 ( .A(n_453), .Y(n_588) );
AND2x2_ASAP7_75t_SL g673 ( .A(n_453), .B(n_582), .Y(n_673) );
AND2x2_ASAP7_75t_L g716 ( .A(n_453), .B(n_537), .Y(n_716) );
INVx5_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx2_ASAP7_75t_L g565 ( .A(n_454), .Y(n_565) );
AND2x2_ASAP7_75t_L g584 ( .A(n_454), .B(n_528), .Y(n_584) );
AND2x2_ASAP7_75t_L g602 ( .A(n_454), .B(n_537), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_454), .B(n_536), .Y(n_662) );
NOR2x1_ASAP7_75t_SL g689 ( .A(n_454), .B(n_462), .Y(n_689) );
OR2x6_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_462), .B(n_528), .Y(n_527) );
AO21x2_ASAP7_75t_L g462 ( .A1(n_463), .A2(n_464), .B(n_470), .Y(n_462) );
NOR2xp33_ASAP7_75t_L g470 ( .A(n_463), .B(n_471), .Y(n_470) );
AO21x2_ASAP7_75t_L g561 ( .A1(n_463), .A2(n_464), .B(n_470), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_469), .Y(n_464) );
AO21x1_ASAP7_75t_L g472 ( .A1(n_473), .A2(n_504), .B(n_513), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
OAI22xp33_ASAP7_75t_L g570 ( .A1(n_474), .A2(n_571), .B1(n_575), .B2(n_576), .Y(n_570) );
OR2x2_ASAP7_75t_L g474 ( .A(n_475), .B(n_483), .Y(n_474) );
AND2x2_ASAP7_75t_L g631 ( .A(n_475), .B(n_519), .Y(n_631) );
BUFx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
AND2x4_ASAP7_75t_L g564 ( .A(n_476), .B(n_547), .Y(n_564) );
AND2x2_ASAP7_75t_L g636 ( .A(n_476), .B(n_521), .Y(n_636) );
AND2x2_ASAP7_75t_L g655 ( .A(n_476), .B(n_621), .Y(n_655) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx2_ASAP7_75t_L g514 ( .A(n_477), .Y(n_514) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_477), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_483), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_L g615 ( .A(n_484), .B(n_516), .Y(n_615) );
AND2x4_ASAP7_75t_L g484 ( .A(n_485), .B(n_496), .Y(n_484) );
AND2x2_ASAP7_75t_L g519 ( .A(n_485), .B(n_520), .Y(n_519) );
OR2x2_ASAP7_75t_L g552 ( .A(n_485), .B(n_553), .Y(n_552) );
AND2x2_ASAP7_75t_SL g612 ( .A(n_485), .B(n_548), .Y(n_612) );
INVx2_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
BUFx2_ASAP7_75t_L g705 ( .A(n_486), .Y(n_705) );
INVx2_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g547 ( .A(n_487), .Y(n_547) );
OAI21x1_ASAP7_75t_SL g487 ( .A1(n_488), .A2(n_490), .B(n_494), .Y(n_487) );
INVx1_ASAP7_75t_L g495 ( .A(n_489), .Y(n_495) );
INVx2_ASAP7_75t_L g553 ( .A(n_496), .Y(n_553) );
HB1xp67_ASAP7_75t_L g653 ( .A(n_496), .Y(n_653) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_498), .B(n_502), .Y(n_497) );
INVx2_ASAP7_75t_L g549 ( .A(n_504), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_504), .B(n_681), .Y(n_707) );
AND2x2_ASAP7_75t_L g726 ( .A(n_504), .B(n_716), .Y(n_726) );
BUFx2_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
AND2x4_ASAP7_75t_SL g594 ( .A(n_505), .B(n_553), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_507), .B(n_511), .Y(n_506) );
AND2x2_ASAP7_75t_SL g513 ( .A(n_514), .B(n_515), .Y(n_513) );
AND2x2_ASAP7_75t_L g593 ( .A(n_514), .B(n_594), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_514), .B(n_563), .Y(n_598) );
INVx1_ASAP7_75t_SL g725 ( .A(n_514), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_515), .B(n_676), .Y(n_675) );
AND2x2_ASAP7_75t_L g515 ( .A(n_516), .B(n_519), .Y(n_515) );
INVx1_ASAP7_75t_L g551 ( .A(n_516), .Y(n_551) );
AND2x2_ASAP7_75t_L g737 ( .A(n_516), .B(n_738), .Y(n_737) );
BUFx2_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g613 ( .A(n_517), .B(n_520), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_517), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g667 ( .A(n_517), .B(n_521), .Y(n_667) );
AND2x2_ASAP7_75t_L g698 ( .A(n_517), .B(n_699), .Y(n_698) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g563 ( .A(n_518), .B(n_521), .Y(n_563) );
INVxp67_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
BUFx3_ASAP7_75t_L g621 ( .A(n_518), .Y(n_621) );
AND2x2_ASAP7_75t_L g641 ( .A(n_519), .B(n_642), .Y(n_641) );
NAND2xp33_ASAP7_75t_L g654 ( .A(n_519), .B(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_520), .B(n_547), .Y(n_610) );
AND2x2_ASAP7_75t_L g699 ( .A(n_520), .B(n_548), .Y(n_699) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x2_ASAP7_75t_L g626 ( .A(n_521), .B(n_548), .Y(n_626) );
OR3x1_ASAP7_75t_L g522 ( .A(n_523), .B(n_570), .C(n_585), .Y(n_522) );
OAI321xp33_ASAP7_75t_L g523 ( .A1(n_524), .A2(n_535), .A3(n_545), .B1(n_550), .B2(n_554), .C(n_562), .Y(n_523) );
INVx1_ASAP7_75t_SL g524 ( .A(n_525), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_527), .Y(n_601) );
INVxp67_ASAP7_75t_SL g619 ( .A(n_527), .Y(n_619) );
OR2x2_ASAP7_75t_L g623 ( .A(n_527), .B(n_535), .Y(n_623) );
BUFx3_ASAP7_75t_L g557 ( .A(n_528), .Y(n_557) );
AND2x2_ASAP7_75t_L g574 ( .A(n_528), .B(n_560), .Y(n_574) );
INVx1_ASAP7_75t_L g591 ( .A(n_528), .Y(n_591) );
INVx2_ASAP7_75t_L g607 ( .A(n_528), .Y(n_607) );
OR2x2_ASAP7_75t_L g646 ( .A(n_528), .B(n_536), .Y(n_646) );
INVx2_ASAP7_75t_L g634 ( .A(n_535), .Y(n_634) );
AND2x2_ASAP7_75t_L g558 ( .A(n_536), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g573 ( .A(n_536), .Y(n_573) );
AND2x4_ASAP7_75t_L g582 ( .A(n_536), .B(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_536), .B(n_559), .Y(n_605) );
AND2x2_ASAP7_75t_L g712 ( .A(n_536), .B(n_607), .Y(n_712) );
INVx4_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_537), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_543), .Y(n_538) );
INVx1_ASAP7_75t_L g599 ( .A(n_545), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_546), .B(n_549), .Y(n_545) );
AND2x2_ASAP7_75t_L g686 ( .A(n_546), .B(n_613), .Y(n_686) );
INVx1_ASAP7_75t_SL g703 ( .A(n_546), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g732 ( .A(n_546), .B(n_679), .Y(n_732) );
AND2x4_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .Y(n_546) );
OR2x2_ASAP7_75t_L g575 ( .A(n_547), .B(n_548), .Y(n_575) );
AND2x2_ASAP7_75t_L g668 ( .A(n_549), .B(n_564), .Y(n_668) );
OR2x2_ASAP7_75t_L g550 ( .A(n_551), .B(n_552), .Y(n_550) );
NAND2xp5_ASAP7_75t_SL g691 ( .A(n_553), .B(n_564), .Y(n_691) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_555), .A2(n_704), .B1(n_709), .B2(n_711), .Y(n_708) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
AND2x2_ASAP7_75t_L g633 ( .A(n_556), .B(n_634), .Y(n_633) );
OR2x2_ASAP7_75t_L g728 ( .A(n_556), .B(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g684 ( .A(n_557), .B(n_602), .Y(n_684) );
AND2x4_ASAP7_75t_L g638 ( .A(n_558), .B(n_584), .Y(n_638) );
INVx1_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_560), .Y(n_736) );
INVx2_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
INVx1_ASAP7_75t_L g569 ( .A(n_561), .Y(n_569) );
INVx1_ASAP7_75t_L g583 ( .A(n_561), .Y(n_583) );
NAND4xp25_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .C(n_565), .D(n_566), .Y(n_562) );
AND2x2_ASAP7_75t_L g720 ( .A(n_563), .B(n_705), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_563), .B(n_731), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g639 ( .A(n_564), .B(n_640), .Y(n_639) );
OAI322xp33_ASAP7_75t_L g647 ( .A1(n_564), .A2(n_648), .A3(n_652), .B1(n_654), .B2(n_656), .C1(n_658), .C2(n_663), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_564), .B(n_613), .Y(n_663) );
INVx1_ASAP7_75t_L g731 ( .A(n_564), .Y(n_731) );
INVx2_ASAP7_75t_L g577 ( .A(n_565), .Y(n_577) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_568), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_569), .B(n_588), .Y(n_645) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_572), .B(n_615), .Y(n_614) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g618 ( .A(n_573), .Y(n_618) );
AND2x2_ASAP7_75t_L g690 ( .A(n_573), .B(n_601), .Y(n_690) );
AOI31xp33_ASAP7_75t_L g576 ( .A1(n_574), .A2(n_577), .A3(n_578), .B(n_581), .Y(n_576) );
AND2x2_ASAP7_75t_L g587 ( .A(n_574), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g715 ( .A(n_574), .B(n_716), .Y(n_715) );
AND2x2_ASAP7_75t_SL g722 ( .A(n_574), .B(n_602), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_574), .Y(n_723) );
INVx1_ASAP7_75t_SL g681 ( .A(n_575), .Y(n_681) );
NAND3xp33_ASAP7_75t_SL g709 ( .A(n_575), .B(n_703), .C(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g609 ( .A(n_580), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g590 ( .A(n_582), .B(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g651 ( .A(n_582), .Y(n_651) );
AOI322xp5_ASAP7_75t_L g733 ( .A1(n_582), .A2(n_612), .A3(n_615), .B1(n_734), .B2(n_735), .C1(n_737), .C2(n_739), .Y(n_733) );
AND2x2_ASAP7_75t_L g739 ( .A(n_582), .B(n_588), .Y(n_739) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_586), .A2(n_589), .B(n_592), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_588), .B(n_607), .Y(n_606) );
AND2x4_ASAP7_75t_L g734 ( .A(n_588), .B(n_621), .Y(n_734) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g660 ( .A(n_591), .Y(n_660) );
AND2x2_ASAP7_75t_L g688 ( .A(n_591), .B(n_689), .Y(n_688) );
AND2x2_ASAP7_75t_L g735 ( .A(n_591), .B(n_736), .Y(n_735) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx1_ASAP7_75t_L g640 ( .A(n_594), .Y(n_640) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
O2A1O1Ixp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_599), .B(n_600), .C(n_603), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g600 ( .A(n_601), .B(n_602), .Y(n_600) );
AND2x2_ASAP7_75t_L g657 ( .A(n_602), .B(n_607), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B(n_614), .C(n_616), .Y(n_603) );
OAI221xp5_ASAP7_75t_L g629 ( .A1(n_604), .A2(n_630), .B1(n_632), .B2(n_635), .C(n_637), .Y(n_629) );
OR2x2_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
INVx1_ASAP7_75t_L g649 ( .A(n_606), .Y(n_649) );
OR2x2_ASAP7_75t_L g669 ( .A(n_606), .B(n_670), .Y(n_669) );
AND2x2_ASAP7_75t_L g608 ( .A(n_609), .B(n_611), .Y(n_608) );
INVx1_ASAP7_75t_L g714 ( .A(n_609), .Y(n_714) );
INVx1_ASAP7_75t_L g738 ( .A(n_610), .Y(n_738) );
NAND2xp5_ASAP7_75t_SL g611 ( .A(n_612), .B(n_613), .Y(n_611) );
AND2x2_ASAP7_75t_L g620 ( .A(n_612), .B(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_612), .B(n_682), .Y(n_694) );
INVx1_ASAP7_75t_L g674 ( .A(n_613), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g616 ( .A1(n_617), .A2(n_620), .B1(n_622), .B2(n_624), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .Y(n_617) );
INVx1_ASAP7_75t_SL g682 ( .A(n_621), .Y(n_682) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
NAND4xp75_ASAP7_75t_L g627 ( .A(n_628), .B(n_664), .C(n_692), .D(n_717), .Y(n_627) );
NOR2xp67_ASAP7_75t_L g628 ( .A(n_629), .B(n_647), .Y(n_628) );
INVx1_ASAP7_75t_SL g630 ( .A(n_631), .Y(n_630) );
INVx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_SL g704 ( .A(n_636), .B(n_705), .Y(n_704) );
AOI22xp5_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_639), .B1(n_641), .B2(n_643), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_640), .B(n_703), .Y(n_702) );
INVx2_ASAP7_75t_SL g643 ( .A(n_644), .Y(n_643) );
OR2x2_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
INVx2_ASAP7_75t_L g680 ( .A(n_646), .Y(n_680) );
OR2x2_ASAP7_75t_L g695 ( .A(n_646), .B(n_696), .Y(n_695) );
NAND2xp5_ASAP7_75t_SL g648 ( .A(n_649), .B(n_650), .Y(n_648) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVx1_ASAP7_75t_L g710 ( .A(n_655), .Y(n_710) );
INVx1_ASAP7_75t_SL g656 ( .A(n_657), .Y(n_656) );
OAI21xp5_ASAP7_75t_SL g701 ( .A1(n_657), .A2(n_702), .B(n_704), .Y(n_701) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_665), .B(n_677), .Y(n_664) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_669), .B1(n_672), .B2(n_674), .C(n_675), .Y(n_665) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g713 ( .A1(n_667), .A2(n_714), .B(n_715), .Y(n_713) );
INVx3_ASAP7_75t_SL g672 ( .A(n_673), .Y(n_672) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_681), .A3(n_682), .B1(n_683), .B2(n_685), .C1(n_687), .C2(n_691), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_SL g685 ( .A(n_686), .Y(n_685) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_688), .B(n_690), .Y(n_687) );
INVx1_ASAP7_75t_L g700 ( .A(n_688), .Y(n_700) );
INVx1_ASAP7_75t_L g696 ( .A(n_689), .Y(n_696) );
AND2x2_ASAP7_75t_L g711 ( .A(n_689), .B(n_712), .Y(n_711) );
NOR2x1_ASAP7_75t_L g692 ( .A(n_693), .B(n_706), .Y(n_692) );
OAI221xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B1(n_697), .B2(n_700), .C(n_701), .Y(n_693) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g706 ( .A1(n_700), .A2(n_707), .B(n_708), .C(n_713), .Y(n_706) );
INVx2_ASAP7_75t_SL g729 ( .A(n_716), .Y(n_729) );
NOR2x1_ASAP7_75t_L g717 ( .A(n_718), .B(n_727), .Y(n_717) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_723), .B2(n_724), .Y(n_718) );
INVx1_ASAP7_75t_SL g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
OAI211xp5_ASAP7_75t_SL g727 ( .A1(n_728), .A2(n_730), .B(n_732), .C(n_733), .Y(n_727) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
INVx1_ASAP7_75t_SL g746 ( .A(n_741), .Y(n_746) );
CKINVDCx11_ASAP7_75t_R g741 ( .A(n_742), .Y(n_741) );
NOR2xp33_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
CKINVDCx5p33_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
CKINVDCx5p33_ASAP7_75t_R g753 ( .A(n_754), .Y(n_753) );
BUFx3_ASAP7_75t_L g754 ( .A(n_755), .Y(n_754) );
INVx1_ASAP7_75t_L g759 ( .A(n_755), .Y(n_759) );
CKINVDCx20_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
HB1xp67_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
CKINVDCx11_ASAP7_75t_R g763 ( .A(n_764), .Y(n_763) );
CKINVDCx20_ASAP7_75t_R g764 ( .A(n_765), .Y(n_764) );
CKINVDCx5p33_ASAP7_75t_R g766 ( .A(n_767), .Y(n_766) );
CKINVDCx5p33_ASAP7_75t_R g767 ( .A(n_768), .Y(n_767) );
BUFx8_ASAP7_75t_SL g768 ( .A(n_769), .Y(n_768) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_770), .Y(n_769) );
BUFx4f_ASAP7_75t_SL g779 ( .A(n_770), .Y(n_779) );
NAND2xp5_ASAP7_75t_SL g770 ( .A(n_771), .B(n_775), .Y(n_770) );
NOR2xp33_ASAP7_75t_L g776 ( .A(n_777), .B(n_778), .Y(n_776) );
INVx1_ASAP7_75t_SL g778 ( .A(n_779), .Y(n_778) );
endmodule