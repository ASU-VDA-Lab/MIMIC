module fake_netlist_1_7079_n_37 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_37);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_37;
wire n_20;
wire n_36;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx5p33_ASAP7_75t_R g11 ( .A(n_5), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_8), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_6), .Y(n_13) );
CKINVDCx5p33_ASAP7_75t_R g14 ( .A(n_3), .Y(n_14) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_4), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_0), .B(n_9), .Y(n_16) );
BUFx6f_ASAP7_75t_L g17 ( .A(n_1), .Y(n_17) );
AOI21xp33_ASAP7_75t_L g18 ( .A1(n_11), .A2(n_0), .B(n_1), .Y(n_18) );
NOR2xp33_ASAP7_75t_L g19 ( .A(n_15), .B(n_14), .Y(n_19) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_15), .B(n_2), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_13), .Y(n_21) );
INVx1_ASAP7_75t_SL g22 ( .A(n_12), .Y(n_22) );
AO31x2_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_13), .A3(n_17), .B(n_16), .Y(n_23) );
INVx3_ASAP7_75t_L g24 ( .A(n_21), .Y(n_24) );
OAI22xp5_ASAP7_75t_L g25 ( .A1(n_20), .A2(n_17), .B1(n_3), .B2(n_4), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_23), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
AND2x4_ASAP7_75t_L g28 ( .A(n_24), .B(n_19), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_27), .Y(n_29) );
OAI32xp33_ASAP7_75t_L g30 ( .A1(n_26), .A2(n_25), .A3(n_18), .B1(n_23), .B2(n_17), .Y(n_30) );
OAI21xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_26), .B(n_27), .Y(n_31) );
AOI221xp5_ASAP7_75t_L g32 ( .A1(n_30), .A2(n_28), .B1(n_22), .B2(n_25), .C(n_17), .Y(n_32) );
OAI22xp5_ASAP7_75t_L g33 ( .A1(n_32), .A2(n_28), .B1(n_17), .B2(n_30), .Y(n_33) );
XOR2xp5_ASAP7_75t_L g34 ( .A(n_31), .B(n_28), .Y(n_34) );
XOR2x2_ASAP7_75t_L g35 ( .A(n_34), .B(n_2), .Y(n_35) );
INVx2_ASAP7_75t_L g36 ( .A(n_33), .Y(n_36) );
AOI222xp33_ASAP7_75t_L g37 ( .A1(n_35), .A2(n_7), .B1(n_8), .B2(n_9), .C1(n_10), .C2(n_36), .Y(n_37) );
endmodule