module real_jpeg_4288_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_300;
wire n_221;
wire n_249;
wire n_292;
wire n_288;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_299;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_139;
wire n_188;
wire n_33;
wire n_65;
wire n_142;
wire n_175;
wire n_238;
wire n_76;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_259;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_187;
wire n_75;
wire n_97;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_216;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_127;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx8_ASAP7_75t_L g49 ( 
.A(n_0),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_1),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_1),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_2),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_2),
.A2(n_60),
.B1(n_68),
.B2(n_83),
.Y(n_82)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_2),
.A2(n_90),
.B(n_93),
.C(n_96),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_2),
.A2(n_60),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_2),
.A2(n_60),
.B1(n_139),
.B2(n_141),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_2),
.B(n_70),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_2),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_2),
.B(n_155),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_2),
.B(n_250),
.C(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_2),
.B(n_47),
.C(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_3),
.A2(n_183),
.B1(n_187),
.B2(n_188),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_3),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_4),
.A2(n_26),
.B1(n_66),
.B2(n_68),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_4),
.A2(n_26),
.B1(n_109),
.B2(n_111),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_4),
.A2(n_26),
.B1(n_154),
.B2(n_162),
.Y(n_161)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_5),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_5),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_5),
.Y(n_186)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_7),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_7),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_7),
.Y(n_126)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_7),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_8),
.Y(n_72)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_8),
.Y(n_78)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_8),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_8),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_10),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_10),
.Y(n_68)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_10),
.Y(n_77)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_10),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_11),
.Y(n_150)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_11),
.Y(n_152)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_11),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g250 ( 
.A(n_11),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_208),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_206),
.Y(n_13)
);

OR2x2_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_173),
.Y(n_14)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_15),
.B(n_173),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_122),
.C(n_166),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_17),
.B(n_211),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_88),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_64),
.B2(n_87),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_19),
.B(n_222),
.C(n_224),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_19),
.A2(n_20),
.B1(n_289),
.B2(n_290),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g19 ( 
.A(n_20),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_20),
.B(n_64),
.C(n_88),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_31),
.B1(n_45),
.B2(n_56),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g167 ( 
.A1(n_21),
.A2(n_31),
.B1(n_45),
.B2(n_56),
.Y(n_167)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_23),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_24),
.Y(n_63)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_30),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_31),
.B(n_45),
.Y(n_202)
);

NAND2x1_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_45),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_38),
.B1(n_40),
.B2(n_43),
.Y(n_32)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_36),
.Y(n_42)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_37),
.Y(n_51)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_42),
.Y(n_273)
);

BUFx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_45),
.Y(n_259)
);

AOI22x1_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_50),
.B1(n_52),
.B2(n_54),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_48),
.Y(n_140)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_49),
.Y(n_53)
);

INVx11_ASAP7_75t_L g143 ( 
.A(n_49),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g147 ( 
.A(n_49),
.Y(n_147)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_49),
.Y(n_248)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_51),
.Y(n_55)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_56),
.Y(n_201)
);

OAI21xp33_ASAP7_75t_L g93 ( 
.A1(n_57),
.A2(n_60),
.B(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g87 ( 
.A(n_64),
.Y(n_87)
);

OA22x2_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_69),
.B1(n_82),
.B2(n_86),
.Y(n_64)
);

OA22x2_ASAP7_75t_L g172 ( 
.A1(n_65),
.A2(n_69),
.B1(n_82),
.B2(n_86),
.Y(n_172)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g96 ( 
.A(n_68),
.Y(n_96)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_75),
.Y(n_69)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_70),
.Y(n_86)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_79),
.B2(n_80),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_97),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_89),
.A2(n_97),
.B1(n_98),
.B2(n_220),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_89),
.Y(n_220)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_95),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_97),
.A2(n_98),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_98),
.B(n_240),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_98),
.B(n_240),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_98),
.B(n_194),
.C(n_258),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_108),
.B1(n_115),
.B2(n_118),
.Y(n_98)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_99),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_99),
.A2(n_108),
.B1(n_118),
.B2(n_125),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_104),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_102),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_103),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_103),
.Y(n_130)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_107),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_107),
.Y(n_278)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_110),
.Y(n_119)
);

INVx4_ASAP7_75t_L g189 ( 
.A(n_110),
.Y(n_189)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_114),
.Y(n_121)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

INVx3_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_118),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_118),
.B(n_275),
.Y(n_274)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_122),
.B(n_166),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_135),
.B1(n_136),
.B2(n_165),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_123),
.Y(n_165)
);

NOR2xp67_ASAP7_75t_L g205 ( 
.A(n_123),
.B(n_136),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g123 ( 
.A1(n_124),
.A2(n_127),
.B(n_132),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_127),
.Y(n_180)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_131),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_133),
.A2(n_180),
.B1(n_181),
.B2(n_190),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_133),
.B(n_276),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_135),
.A2(n_136),
.B1(n_244),
.B2(n_252),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_135),
.B(n_252),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_135),
.A2(n_136),
.B1(n_167),
.B2(n_216),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_135),
.B(n_216),
.C(n_266),
.Y(n_292)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g136 ( 
.A(n_137),
.B(n_160),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_144),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_138),
.B(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_138),
.Y(n_196)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_140),
.Y(n_139)
);

INVx11_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_143),
.Y(n_154)
);

INVx5_ASAP7_75t_L g164 ( 
.A(n_143),
.Y(n_164)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_144),
.Y(n_171)
);

NOR2x1_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_155),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_148),
.B1(n_151),
.B2(n_153),
.Y(n_145)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AO22x1_ASAP7_75t_SL g155 ( 
.A1(n_151),
.A2(n_156),
.B1(n_157),
.B2(n_158),
.Y(n_155)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_155),
.B(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_155),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_161),
.Y(n_195)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_168),
.C(n_172),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_167),
.A2(n_168),
.B1(n_216),
.B2(n_217),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_167),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g194 ( 
.A1(n_170),
.A2(n_171),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_172),
.A2(n_200),
.B1(n_203),
.B2(n_204),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_172),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_172),
.A2(n_203),
.B1(n_214),
.B2(n_215),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_175),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B1(n_197),
.B2(n_198),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_179),
.B1(n_193),
.B2(n_194),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_188),
.Y(n_251)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_193),
.A2(n_194),
.B1(n_258),
.B2(n_260),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_193),
.A2(n_194),
.B1(n_285),
.B2(n_286),
.Y(n_284)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_194),
.B(n_285),
.C(n_287),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_198),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_205),
.Y(n_198)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_226),
.B(n_300),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_212),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_210),
.B(n_212),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_218),
.C(n_221),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_213),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_218),
.A2(n_219),
.B1(n_221),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_221),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_243),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_222),
.A2(n_223),
.B1(n_224),
.B2(n_225),
.Y(n_290)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_223),
.B(n_235),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_225),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_294),
.B(n_299),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_282),
.B(n_293),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_263),
.B(n_281),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_254),
.B(n_262),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_242),
.B(n_253),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_239),
.B(n_241),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_244),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_249),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

INVx4_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_261),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_261),
.Y(n_262)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_258),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_264),
.B(n_265),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_264),
.B(n_265),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_266),
.B(n_280),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_274),
.B2(n_279),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_267),
.B(n_279),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_272),
.Y(n_268)
);

INVx3_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_274),
.Y(n_279)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx8_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_283),
.B(n_292),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_292),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_284),
.A2(n_287),
.B1(n_288),
.B2(n_291),
.Y(n_283)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_284),
.Y(n_291)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);


endmodule