module fake_jpeg_18105_n_190 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_190);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_190;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_0),
.B(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_31),
.B(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_32),
.Y(n_58)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_29),
.Y(n_34)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_25),
.B(n_12),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_23),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_26),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_26),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_53),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_33),
.A2(n_18),
.B1(n_28),
.B2(n_27),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_59),
.B1(n_64),
.B2(n_45),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_33),
.A2(n_23),
.B1(n_28),
.B2(n_27),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_52),
.A2(n_24),
.B1(n_39),
.B2(n_42),
.Y(n_85)
);

AOI32xp33_ASAP7_75t_L g53 ( 
.A1(n_31),
.A2(n_16),
.A3(n_19),
.B1(n_14),
.B2(n_21),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_44),
.A2(n_45),
.B1(n_39),
.B2(n_43),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_20),
.C(n_26),
.Y(n_62)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_62),
.B(n_42),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_14),
.B1(n_24),
.B2(n_19),
.Y(n_64)
);

OA21x2_ASAP7_75t_L g66 ( 
.A1(n_49),
.A2(n_41),
.B(n_40),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_83),
.B1(n_2),
.B2(n_3),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_37),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_67),
.B(n_74),
.Y(n_96)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_16),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_69),
.B(n_12),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_55),
.B(n_38),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_70),
.B(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_72),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_50),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_78),
.C(n_2),
.Y(n_106)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_30),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_75),
.B(n_79),
.Y(n_97)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_76),
.Y(n_112)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_47),
.Y(n_77)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_55),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_55),
.B(n_38),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_50),
.B(n_36),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_82),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_51),
.B(n_36),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_84),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

AO22x2_ASAP7_75t_SL g87 ( 
.A1(n_63),
.A2(n_32),
.B1(n_34),
.B2(n_35),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_87),
.B(n_91),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_61),
.B(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_61),
.B(n_20),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_92),
.Y(n_107)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_20),
.Y(n_92)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_63),
.A2(n_35),
.B1(n_20),
.B2(n_17),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_93),
.A2(n_79),
.B1(n_83),
.B2(n_82),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_95),
.B(n_5),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_98),
.A2(n_99),
.B1(n_114),
.B2(n_115),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_66),
.A2(n_17),
.B1(n_3),
.B2(n_4),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_106),
.B(n_80),
.C(n_93),
.Y(n_125)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_71),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_72),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_65),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_116),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_106),
.B(n_78),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_117),
.B(n_123),
.Y(n_146)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_118),
.B(n_122),
.Y(n_139)
);

AO22x1_ASAP7_75t_SL g119 ( 
.A1(n_98),
.A2(n_66),
.B1(n_87),
.B2(n_73),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_131),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_100),
.A2(n_73),
.B1(n_68),
.B2(n_93),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_96),
.B(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_121),
.B(n_124),
.Y(n_144)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_102),
.B(n_70),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_130),
.C(n_117),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g126 ( 
.A(n_107),
.B(n_87),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_127),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_74),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_113),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_129),
.Y(n_134)
);

XNOR2x1_ASAP7_75t_SL g130 ( 
.A(n_102),
.B(n_93),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_100),
.A2(n_81),
.B1(n_90),
.B2(n_76),
.Y(n_131)
);

NAND2x1_ASAP7_75t_SL g132 ( 
.A(n_110),
.B(n_77),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_132),
.B(n_91),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_133),
.B(n_140),
.C(n_141),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_138),
.B(n_110),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_103),
.C(n_97),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_125),
.B(n_130),
.C(n_103),
.Y(n_141)
);

AOI322xp5_ASAP7_75t_SL g143 ( 
.A1(n_126),
.A2(n_115),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.C1(n_7),
.C2(n_101),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_143),
.B(n_7),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_145),
.A2(n_120),
.B(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_140),
.B(n_119),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_148),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_146),
.C(n_141),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_149),
.A2(n_154),
.B(n_156),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_150),
.B(n_155),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_131),
.C(n_128),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_151),
.C(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_139),
.Y(n_153)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_153),
.Y(n_161)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_137),
.B(n_119),
.C(n_128),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_142),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_137),
.A2(n_105),
.B(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_157),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_136),
.B(n_113),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

XOR2x1_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_145),
.Y(n_160)
);

AO21x1_ASAP7_75t_L g170 ( 
.A1(n_160),
.A2(n_148),
.B(n_156),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_163),
.B(n_167),
.C(n_165),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_136),
.C(n_134),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_167),
.B(n_112),
.C(n_109),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_144),
.Y(n_169)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_169),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_158),
.B1(n_154),
.B2(n_152),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_163),
.B(n_149),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_172),
.B(n_174),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_175),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_112),
.B1(n_111),
.B2(n_108),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_173),
.B(n_168),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_180),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_170),
.B(n_166),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_182),
.A2(n_183),
.B1(n_108),
.B2(n_176),
.Y(n_185)
);

AOI31xp67_ASAP7_75t_L g183 ( 
.A1(n_177),
.A2(n_164),
.A3(n_175),
.B(n_122),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_178),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_184),
.B(n_185),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_184),
.B(n_176),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_186),
.Y(n_188)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_188),
.A2(n_187),
.B(n_109),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_8),
.Y(n_190)
);


endmodule