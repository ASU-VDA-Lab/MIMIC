module fake_netlist_5_2179_n_1909 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1909);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1909;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_314;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_750;
wire n_742;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1735;
wire n_1697;
wire n_1575;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1835;
wire n_1726;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_SL g177 ( 
.A(n_18),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_93),
.Y(n_178)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_103),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_25),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_102),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_34),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_22),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_120),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_50),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_8),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_44),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_134),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_11),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_142),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_6),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_118),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_135),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_173),
.Y(n_195)
);

BUFx3_ASAP7_75t_L g196 ( 
.A(n_159),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_80),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_73),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_82),
.Y(n_199)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_149),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_139),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_78),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_169),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_12),
.Y(n_204)
);

INVx1_ASAP7_75t_SL g205 ( 
.A(n_46),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_147),
.Y(n_206)
);

BUFx10_ASAP7_75t_L g207 ( 
.A(n_130),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_17),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_112),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_156),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_152),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_79),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_51),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_53),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_33),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_175),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_100),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_35),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_19),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_110),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_128),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_7),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_17),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_23),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_146),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_123),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_121),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_106),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_95),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_71),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_7),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_66),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_124),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_167),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_0),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_42),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_34),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_157),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_46),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_92),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_163),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_53),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_36),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_55),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_23),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_165),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_32),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_168),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_75),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_151),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_18),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_98),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_2),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_24),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_166),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_11),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_61),
.Y(n_259)
);

BUFx10_ASAP7_75t_L g260 ( 
.A(n_35),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_43),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_99),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_69),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_10),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_114),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_87),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_83),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_138),
.Y(n_268)
);

INVx1_ASAP7_75t_SL g269 ( 
.A(n_150),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_77),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_72),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_59),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_117),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_116),
.Y(n_274)
);

BUFx10_ASAP7_75t_L g275 ( 
.A(n_113),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_58),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_70),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_21),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_70),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_59),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_69),
.Y(n_281)
);

BUFx10_ASAP7_75t_L g282 ( 
.A(n_96),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_52),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_47),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_109),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_43),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_104),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_140),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_91),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_41),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_164),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_45),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_148),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_36),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_171),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_174),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_162),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_86),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_76),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_28),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_65),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_37),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_160),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_32),
.Y(n_306)
);

BUFx2_ASAP7_75t_L g307 ( 
.A(n_132),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_126),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_119),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_60),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_136),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_12),
.Y(n_312)
);

BUFx10_ASAP7_75t_L g313 ( 
.A(n_153),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_45),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_28),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_60),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_55),
.Y(n_317)
);

INVx4_ASAP7_75t_R g318 ( 
.A(n_129),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_108),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_25),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_51),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_143),
.Y(n_322)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_144),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_127),
.Y(n_324)
);

INVx2_ASAP7_75t_SL g325 ( 
.A(n_170),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_19),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_5),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_89),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_13),
.Y(n_329)
);

INVx1_ASAP7_75t_SL g330 ( 
.A(n_90),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_15),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g332 ( 
.A(n_94),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_137),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_15),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_1),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_0),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_14),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_13),
.Y(n_338)
);

BUFx6f_ASAP7_75t_L g339 ( 
.A(n_133),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_88),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_68),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_154),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_8),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_10),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_54),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_48),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_42),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_66),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_97),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_115),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_24),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_14),
.Y(n_352)
);

INVx3_ASAP7_75t_L g353 ( 
.A(n_347),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_178),
.Y(n_354)
);

NOR2xp67_ASAP7_75t_L g355 ( 
.A(n_302),
.B(n_1),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_347),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_184),
.Y(n_357)
);

HB1xp67_ASAP7_75t_L g358 ( 
.A(n_225),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_347),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_347),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g362 ( 
.A(n_307),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_210),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_303),
.Y(n_364)
);

BUFx2_ASAP7_75t_L g365 ( 
.A(n_225),
.Y(n_365)
);

OR2x2_ASAP7_75t_L g366 ( 
.A(n_219),
.B(n_2),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_229),
.Y(n_367)
);

BUFx6f_ASAP7_75t_SL g368 ( 
.A(n_207),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_234),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_303),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_190),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_249),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_194),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_195),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_307),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g376 ( 
.A(n_191),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_200),
.B(n_3),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_219),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_224),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_198),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_200),
.B(n_3),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_232),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_199),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_232),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_248),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_202),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_248),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_252),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_252),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_258),
.Y(n_391)
);

INVxp33_ASAP7_75t_SL g392 ( 
.A(n_246),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_258),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_264),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_256),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_264),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_203),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_179),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g399 ( 
.A(n_246),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_272),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_319),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_272),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_277),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_228),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_277),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_283),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_180),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_283),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_206),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_182),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_R g411 ( 
.A(n_212),
.B(n_176),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_221),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_230),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_284),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_231),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_179),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_284),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_239),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_286),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_241),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_242),
.Y(n_421)
);

INVx4_ASAP7_75t_R g422 ( 
.A(n_196),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_209),
.B(n_4),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_286),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_295),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_247),
.Y(n_426)
);

INVxp67_ASAP7_75t_SL g427 ( 
.A(n_196),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g428 ( 
.A(n_209),
.B(n_4),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_306),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_306),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_310),
.Y(n_431)
);

INVxp33_ASAP7_75t_SL g432 ( 
.A(n_183),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_310),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_251),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_312),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_253),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_312),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_257),
.Y(n_438)
);

INVx1_ASAP7_75t_SL g439 ( 
.A(n_204),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_369),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_L g441 ( 
.A1(n_399),
.A2(n_301),
.B1(n_214),
.B2(n_223),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_362),
.B(n_325),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_369),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_356),
.Y(n_444)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_407),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_369),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_381),
.B(n_207),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_353),
.B(n_325),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_404),
.Y(n_452)
);

AND2x2_ASAP7_75t_L g453 ( 
.A(n_398),
.B(n_235),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_369),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_353),
.B(n_262),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_369),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_353),
.B(n_235),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_365),
.Y(n_458)
);

BUFx6f_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

AND2x6_ASAP7_75t_L g460 ( 
.A(n_377),
.B(n_234),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_416),
.B(n_265),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_427),
.B(n_266),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_423),
.B(n_428),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g464 ( 
.A(n_358),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_359),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_361),
.Y(n_466)
);

AND2x6_ASAP7_75t_L g467 ( 
.A(n_360),
.B(n_234),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_361),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_378),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_375),
.B(n_432),
.Y(n_470)
);

AND2x4_ASAP7_75t_L g471 ( 
.A(n_378),
.B(n_193),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_379),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

AND2x2_ASAP7_75t_L g474 ( 
.A(n_364),
.B(n_370),
.Y(n_474)
);

BUFx6f_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_370),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_365),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_355),
.Y(n_480)
);

INVxp33_ASAP7_75t_L g481 ( 
.A(n_366),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_383),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_383),
.B(n_351),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_385),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_385),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_439),
.Y(n_486)
);

BUFx2_ASAP7_75t_L g487 ( 
.A(n_354),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_386),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_386),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_388),
.B(n_267),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_388),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

INVx2_ASAP7_75t_L g493 ( 
.A(n_389),
.Y(n_493)
);

OR2x2_ASAP7_75t_L g494 ( 
.A(n_366),
.B(n_254),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_390),
.B(n_268),
.Y(n_495)
);

BUFx6f_ASAP7_75t_L g496 ( 
.A(n_390),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_391),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_391),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_393),
.Y(n_499)
);

OA21x2_ASAP7_75t_L g500 ( 
.A1(n_393),
.A2(n_341),
.B(n_334),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_L g501 ( 
.A(n_357),
.B(n_185),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_394),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_394),
.B(n_270),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_396),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_396),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_400),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_400),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_402),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_392),
.B(n_207),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_371),
.B(n_269),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_402),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_403),
.B(n_351),
.Y(n_512)
);

HB1xp67_ASAP7_75t_L g513 ( 
.A(n_403),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_405),
.Y(n_514)
);

HB1xp67_ASAP7_75t_L g515 ( 
.A(n_405),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_468),
.Y(n_517)
);

AO21x2_ASAP7_75t_L g518 ( 
.A1(n_463),
.A2(n_188),
.B(n_181),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_468),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_513),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_461),
.B(n_373),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_513),
.Y(n_522)
);

NAND3xp33_ASAP7_75t_L g523 ( 
.A(n_463),
.B(n_380),
.C(n_374),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_515),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_515),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_486),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_510),
.B(n_193),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_469),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_470),
.B(n_387),
.C(n_384),
.Y(n_529)
);

BUFx10_ASAP7_75t_L g530 ( 
.A(n_510),
.Y(n_530)
);

BUFx4f_ASAP7_75t_L g531 ( 
.A(n_500),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_486),
.Y(n_532)
);

BUFx2_ASAP7_75t_L g533 ( 
.A(n_452),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_469),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_448),
.B(n_509),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_452),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_472),
.Y(n_537)
);

OR2x2_ASAP7_75t_L g538 ( 
.A(n_458),
.B(n_376),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_460),
.A2(n_254),
.B1(n_334),
.B2(n_345),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_468),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_457),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_468),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_461),
.B(n_397),
.Y(n_543)
);

AND2x6_ASAP7_75t_L g544 ( 
.A(n_453),
.B(n_211),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_457),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_446),
.Y(n_546)
);

INVx6_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_444),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_472),
.Y(n_549)
);

BUFx3_ASAP7_75t_L g550 ( 
.A(n_457),
.Y(n_550)
);

OR2x6_ASAP7_75t_L g551 ( 
.A(n_487),
.B(n_341),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_473),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_473),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_444),
.Y(n_554)
);

BUFx10_ASAP7_75t_L g555 ( 
.A(n_442),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_460),
.A2(n_345),
.B1(n_344),
.B2(n_342),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_447),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_452),
.Y(n_558)
);

BUFx8_ASAP7_75t_SL g559 ( 
.A(n_458),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_448),
.B(n_211),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_458),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_487),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_447),
.Y(n_563)
);

AOI22xp33_ASAP7_75t_L g564 ( 
.A1(n_460),
.A2(n_344),
.B1(n_342),
.B2(n_323),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_488),
.Y(n_565)
);

INVx4_ASAP7_75t_L g566 ( 
.A(n_446),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_451),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_488),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_462),
.B(n_409),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_460),
.A2(n_226),
.B1(n_323),
.B2(n_368),
.Y(n_570)
);

INVxp67_ASAP7_75t_L g571 ( 
.A(n_480),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_489),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_509),
.B(n_226),
.Y(n_573)
);

BUFx3_ASAP7_75t_L g574 ( 
.A(n_457),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_470),
.B(n_234),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_489),
.Y(n_576)
);

INVx3_ASAP7_75t_L g577 ( 
.A(n_446),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_446),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_487),
.B(n_181),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_501),
.A2(n_438),
.B1(n_415),
.B2(n_434),
.Y(n_580)
);

OAI22xp33_ASAP7_75t_L g581 ( 
.A1(n_481),
.A2(n_205),
.B1(n_177),
.B2(n_317),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_491),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_460),
.A2(n_368),
.B1(n_197),
.B2(n_201),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_462),
.B(n_412),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_491),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_455),
.B(n_413),
.Y(n_586)
);

AND2x6_ASAP7_75t_L g587 ( 
.A(n_453),
.B(n_188),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_442),
.B(n_420),
.Y(n_588)
);

OR2x6_ASAP7_75t_L g589 ( 
.A(n_494),
.B(n_197),
.Y(n_589)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_441),
.Y(n_590)
);

BUFx3_ASAP7_75t_L g591 ( 
.A(n_500),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_446),
.Y(n_592)
);

BUFx2_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_455),
.B(n_234),
.Y(n_594)
);

BUFx10_ASAP7_75t_L g595 ( 
.A(n_445),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_497),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_480),
.Y(n_597)
);

INVx4_ASAP7_75t_L g598 ( 
.A(n_446),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_SL g599 ( 
.A(n_490),
.B(n_332),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_453),
.B(n_201),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_497),
.Y(n_601)
);

XNOR2xp5_ASAP7_75t_L g602 ( 
.A(n_441),
.B(n_363),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_451),
.Y(n_603)
);

NOR2x1p5_ASAP7_75t_L g604 ( 
.A(n_494),
.B(n_186),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_445),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_498),
.Y(n_606)
);

OAI21xp33_ASAP7_75t_SL g607 ( 
.A1(n_494),
.A2(n_217),
.B(n_216),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_450),
.A2(n_426),
.B1(n_418),
.B2(n_421),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_498),
.Y(n_609)
);

INVx4_ASAP7_75t_SL g610 ( 
.A(n_460),
.Y(n_610)
);

NOR2xp33_ASAP7_75t_L g611 ( 
.A(n_481),
.B(n_436),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_499),
.Y(n_612)
);

INVx4_ASAP7_75t_L g613 ( 
.A(n_446),
.Y(n_613)
);

INVxp67_ASAP7_75t_SL g614 ( 
.A(n_446),
.Y(n_614)
);

NAND2xp33_ASAP7_75t_SL g615 ( 
.A(n_450),
.B(n_233),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_465),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_465),
.Y(n_617)
);

INVx4_ASAP7_75t_L g618 ( 
.A(n_459),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_499),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_460),
.B(n_330),
.Y(n_620)
);

INVx3_ASAP7_75t_L g621 ( 
.A(n_459),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_479),
.B(n_406),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_460),
.B(n_271),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_SL g624 ( 
.A(n_490),
.B(n_332),
.Y(n_624)
);

NAND2xp5_ASAP7_75t_L g625 ( 
.A(n_460),
.B(n_285),
.Y(n_625)
);

INVx1_ASAP7_75t_SL g626 ( 
.A(n_483),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_466),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

BUFx8_ASAP7_75t_SL g629 ( 
.A(n_483),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_502),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_L g631 ( 
.A(n_495),
.B(n_503),
.Y(n_631)
);

AOI22xp5_ASAP7_75t_L g632 ( 
.A1(n_464),
.A2(n_368),
.B1(n_401),
.B2(n_395),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_460),
.B(n_287),
.Y(n_633)
);

AND2x2_ASAP7_75t_L g634 ( 
.A(n_474),
.B(n_408),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_477),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_483),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_495),
.B(n_503),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_SL g638 ( 
.A1(n_464),
.A2(n_281),
.B1(n_276),
.B2(n_335),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_506),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_506),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_508),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_508),
.Y(n_642)
);

INVx5_ASAP7_75t_L g643 ( 
.A(n_467),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_511),
.Y(n_644)
);

NOR2xp33_ASAP7_75t_SL g645 ( 
.A(n_512),
.B(n_367),
.Y(n_645)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_512),
.A2(n_372),
.B1(n_288),
.B2(n_289),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_511),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_512),
.B(n_189),
.C(n_187),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_500),
.Y(n_649)
);

AO21x2_ASAP7_75t_L g650 ( 
.A1(n_449),
.A2(n_217),
.B(n_216),
.Y(n_650)
);

AND2x6_ASAP7_75t_L g651 ( 
.A(n_471),
.B(n_220),
.Y(n_651)
);

INVx2_ASAP7_75t_SL g652 ( 
.A(n_500),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_466),
.B(n_292),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_474),
.B(n_408),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_500),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_459),
.Y(n_656)
);

OR2x2_ASAP7_75t_L g657 ( 
.A(n_514),
.B(n_414),
.Y(n_657)
);

INVx4_ASAP7_75t_L g658 ( 
.A(n_459),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_471),
.B(n_220),
.Y(n_659)
);

OR2x6_ASAP7_75t_L g660 ( 
.A(n_500),
.B(n_227),
.Y(n_660)
);

INVx1_ASAP7_75t_SL g661 ( 
.A(n_474),
.Y(n_661)
);

CKINVDCx20_ASAP7_75t_R g662 ( 
.A(n_449),
.Y(n_662)
);

NAND2xp33_ASAP7_75t_L g663 ( 
.A(n_467),
.B(n_332),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_471),
.B(n_332),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_471),
.B(n_332),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_514),
.Y(n_666)
);

AND2x6_ASAP7_75t_L g667 ( 
.A(n_471),
.B(n_227),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_485),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_477),
.Y(n_669)
);

AO22x2_ASAP7_75t_L g670 ( 
.A1(n_535),
.A2(n_309),
.B1(n_250),
.B2(n_273),
.Y(n_670)
);

NAND3xp33_ASAP7_75t_L g671 ( 
.A(n_527),
.B(n_208),
.C(n_192),
.Y(n_671)
);

O2A1O1Ixp5_ASAP7_75t_L g672 ( 
.A1(n_531),
.A2(n_485),
.B(n_340),
.C(n_273),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_543),
.B(n_631),
.Y(n_673)
);

AOI21xp5_ASAP7_75t_L g674 ( 
.A1(n_637),
.A2(n_443),
.B(n_440),
.Y(n_674)
);

BUFx6f_ASAP7_75t_SL g675 ( 
.A(n_595),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_591),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_521),
.B(n_485),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_531),
.B(n_339),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_626),
.B(n_661),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_591),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_532),
.B(n_240),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_569),
.B(n_485),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_584),
.B(n_485),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_611),
.B(n_588),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_541),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_655),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_SL g687 ( 
.A(n_531),
.B(n_339),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_541),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_545),
.Y(n_689)
);

INVxp33_ASAP7_75t_L g690 ( 
.A(n_629),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_L g691 ( 
.A1(n_535),
.A2(n_349),
.B1(n_300),
.B2(n_299),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_545),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_SL g693 ( 
.A(n_655),
.B(n_339),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_550),
.Y(n_694)
);

INVx1_ASAP7_75t_SL g695 ( 
.A(n_526),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_597),
.B(n_213),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_R g697 ( 
.A(n_562),
.B(n_296),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_518),
.A2(n_484),
.B1(n_477),
.B2(n_505),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_662),
.A2(n_600),
.B1(n_587),
.B2(n_636),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_636),
.B(n_477),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_548),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_586),
.B(n_477),
.Y(n_702)
);

BUFx6f_ASAP7_75t_L g703 ( 
.A(n_550),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_574),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_548),
.Y(n_705)
);

OAI22xp5_ASAP7_75t_L g706 ( 
.A1(n_523),
.A2(n_333),
.B1(n_311),
.B2(n_309),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_649),
.B(n_477),
.Y(n_707)
);

OR2x2_ASAP7_75t_L g708 ( 
.A(n_561),
.B(n_414),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_554),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_529),
.B(n_215),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_530),
.B(n_218),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_649),
.B(n_477),
.Y(n_712)
);

INVxp67_ASAP7_75t_SL g713 ( 
.A(n_652),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_574),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_662),
.A2(n_297),
.B1(n_305),
.B2(n_322),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_652),
.B(n_518),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_587),
.A2(n_328),
.B1(n_324),
.B2(n_350),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_570),
.B(n_339),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_634),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_634),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_654),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_654),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_518),
.B(n_477),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_528),
.B(n_484),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_534),
.B(n_484),
.Y(n_725)
);

AOI22xp33_ASAP7_75t_L g726 ( 
.A1(n_587),
.A2(n_484),
.B1(n_496),
.B2(n_505),
.Y(n_726)
);

BUFx2_ASAP7_75t_L g727 ( 
.A(n_526),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_530),
.B(n_222),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_635),
.Y(n_729)
);

AND2x4_ASAP7_75t_L g730 ( 
.A(n_659),
.B(n_250),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_537),
.B(n_484),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_659),
.B(n_274),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_549),
.B(n_484),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_657),
.Y(n_734)
);

INVx4_ASAP7_75t_L g735 ( 
.A(n_547),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_552),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_547),
.A2(n_274),
.B1(n_291),
.B2(n_294),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_553),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_565),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_568),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_572),
.B(n_484),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_576),
.B(n_484),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_582),
.Y(n_743)
);

AO221x1_ASAP7_75t_L g744 ( 
.A1(n_581),
.A2(n_339),
.B1(n_291),
.B2(n_294),
.C(n_298),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_585),
.B(n_496),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_L g746 ( 
.A(n_530),
.B(n_237),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_596),
.B(n_496),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_554),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_601),
.B(n_496),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_606),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_571),
.B(n_238),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_609),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_612),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_557),
.Y(n_754)
);

OAI22xp5_ASAP7_75t_SL g755 ( 
.A1(n_590),
.A2(n_236),
.B1(n_316),
.B2(n_327),
.Y(n_755)
);

AOI22xp5_ASAP7_75t_L g756 ( 
.A1(n_587),
.A2(n_298),
.B1(n_308),
.B2(n_311),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_SL g757 ( 
.A(n_620),
.B(n_496),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_559),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_593),
.B(n_244),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_619),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_SL g761 ( 
.A(n_610),
.B(n_496),
.Y(n_761)
);

A2O1A1Ixp33_ASAP7_75t_L g762 ( 
.A1(n_607),
.A2(n_340),
.B(n_333),
.C(n_308),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_SL g763 ( 
.A(n_605),
.B(n_331),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_557),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_610),
.B(n_496),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_587),
.A2(n_505),
.B1(n_496),
.B2(n_475),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_SL g767 ( 
.A(n_610),
.B(n_505),
.Y(n_767)
);

INVx2_ASAP7_75t_L g768 ( 
.A(n_563),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_628),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_583),
.B(n_505),
.Y(n_770)
);

NAND2xp33_ASAP7_75t_L g771 ( 
.A(n_544),
.B(n_467),
.Y(n_771)
);

AOI21xp5_ASAP7_75t_L g772 ( 
.A1(n_614),
.A2(n_443),
.B(n_440),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_630),
.B(n_505),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_639),
.B(n_505),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_668),
.B(n_505),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_563),
.Y(n_776)
);

INVx8_ASAP7_75t_L g777 ( 
.A(n_587),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_640),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_641),
.B(n_478),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_567),
.Y(n_780)
);

HB1xp67_ASAP7_75t_L g781 ( 
.A(n_629),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_547),
.Y(n_782)
);

BUFx3_ASAP7_75t_L g783 ( 
.A(n_520),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_567),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_538),
.B(n_245),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_642),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_600),
.A2(n_507),
.B1(n_504),
.B2(n_493),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_L g788 ( 
.A(n_644),
.B(n_478),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_647),
.Y(n_789)
);

AOI221xp5_ASAP7_75t_L g790 ( 
.A1(n_638),
.A2(n_338),
.B1(n_255),
.B2(n_343),
.C(n_259),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_SL g791 ( 
.A(n_659),
.B(n_475),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_527),
.B(n_475),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_666),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_603),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_595),
.B(n_240),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_603),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_600),
.A2(n_544),
.B1(n_573),
.B2(n_645),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_600),
.B(n_478),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_522),
.B(n_524),
.Y(n_799)
);

BUFx3_ASAP7_75t_L g800 ( 
.A(n_525),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_600),
.A2(n_476),
.B1(n_475),
.B2(n_504),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_SL g802 ( 
.A(n_623),
.B(n_475),
.Y(n_802)
);

BUFx5_ASAP7_75t_L g803 ( 
.A(n_544),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_625),
.B(n_475),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_600),
.B(n_478),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_633),
.B(n_475),
.Y(n_806)
);

NOR2xp33_ASAP7_75t_L g807 ( 
.A(n_555),
.B(n_261),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_544),
.B(n_482),
.Y(n_808)
);

OAI21xp5_ASAP7_75t_L g809 ( 
.A1(n_660),
.A2(n_456),
.B(n_454),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_555),
.B(n_263),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_580),
.B(n_482),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_544),
.B(n_575),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_555),
.B(n_475),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_544),
.B(n_482),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_646),
.B(n_278),
.Y(n_815)
);

INVx2_ASAP7_75t_SL g816 ( 
.A(n_595),
.Y(n_816)
);

AND2x2_ASAP7_75t_L g817 ( 
.A(n_622),
.B(n_240),
.Y(n_817)
);

OR2x6_ASAP7_75t_L g818 ( 
.A(n_579),
.B(n_417),
.Y(n_818)
);

INVx1_ASAP7_75t_L g819 ( 
.A(n_616),
.Y(n_819)
);

NAND2xp33_ASAP7_75t_L g820 ( 
.A(n_564),
.B(n_467),
.Y(n_820)
);

NOR2xp33_ASAP7_75t_L g821 ( 
.A(n_575),
.B(n_279),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_669),
.B(n_476),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_616),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_573),
.B(n_280),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_669),
.B(n_476),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_653),
.B(n_482),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_608),
.B(n_290),
.Y(n_827)
);

AOI22x1_ASAP7_75t_L g828 ( 
.A1(n_604),
.A2(n_456),
.B1(n_454),
.B2(n_443),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_617),
.B(n_492),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_617),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_627),
.B(n_492),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_627),
.Y(n_832)
);

AOI22xp33_ASAP7_75t_L g833 ( 
.A1(n_660),
.A2(n_476),
.B1(n_507),
.B2(n_504),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_560),
.B(n_492),
.Y(n_834)
);

NOR2xp33_ASAP7_75t_L g835 ( 
.A(n_579),
.B(n_293),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_560),
.B(n_492),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_599),
.B(n_493),
.Y(n_837)
);

OR2x6_ASAP7_75t_L g838 ( 
.A(n_579),
.B(n_417),
.Y(n_838)
);

NOR2xp67_ASAP7_75t_SL g839 ( 
.A(n_643),
.B(n_304),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_517),
.Y(n_840)
);

INVx2_ASAP7_75t_L g841 ( 
.A(n_517),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_673),
.B(n_589),
.Y(n_842)
);

BUFx2_ASAP7_75t_L g843 ( 
.A(n_727),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_701),
.Y(n_844)
);

NOR2xp33_ASAP7_75t_L g845 ( 
.A(n_684),
.B(n_562),
.Y(n_845)
);

BUFx4f_ASAP7_75t_L g846 ( 
.A(n_818),
.Y(n_846)
);

AOI21xp5_ASAP7_75t_L g847 ( 
.A1(n_702),
.A2(n_598),
.B(n_566),
.Y(n_847)
);

AOI21xp5_ASAP7_75t_L g848 ( 
.A1(n_713),
.A2(n_598),
.B(n_566),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_821),
.A2(n_648),
.B(n_624),
.C(n_599),
.Y(n_849)
);

AOI21xp5_ASAP7_75t_L g850 ( 
.A1(n_826),
.A2(n_598),
.B(n_566),
.Y(n_850)
);

OAI21xp5_ASAP7_75t_L g851 ( 
.A1(n_716),
.A2(n_660),
.B(n_624),
.Y(n_851)
);

AOI21x1_ASAP7_75t_L g852 ( 
.A1(n_678),
.A2(n_594),
.B(n_660),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_676),
.B(n_589),
.Y(n_853)
);

AOI21x1_ASAP7_75t_L g854 ( 
.A1(n_678),
.A2(n_594),
.B(n_665),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_676),
.B(n_589),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_811),
.A2(n_579),
.B1(n_551),
.B2(n_667),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_707),
.A2(n_613),
.B(n_658),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_680),
.B(n_589),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_758),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_712),
.A2(n_613),
.B(n_658),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_680),
.B(n_650),
.Y(n_861)
);

NOR2xp33_ASAP7_75t_L g862 ( 
.A(n_679),
.B(n_551),
.Y(n_862)
);

OR2x2_ASAP7_75t_L g863 ( 
.A(n_695),
.B(n_533),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_686),
.B(n_650),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_701),
.Y(n_865)
);

INVx3_ASAP7_75t_L g866 ( 
.A(n_703),
.Y(n_866)
);

BUFx4f_ASAP7_75t_L g867 ( 
.A(n_818),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_SL g868 ( 
.A(n_803),
.B(n_797),
.Y(n_868)
);

OAI22xp33_ASAP7_75t_L g869 ( 
.A1(n_719),
.A2(n_590),
.B1(n_551),
.B2(n_632),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_703),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_708),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_705),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_L g873 ( 
.A(n_686),
.B(n_650),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_699),
.B(n_536),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_687),
.A2(n_613),
.B(n_618),
.Y(n_875)
);

NOR2xp33_ASAP7_75t_L g876 ( 
.A(n_711),
.B(n_551),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_803),
.B(n_677),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_687),
.A2(n_618),
.B(n_658),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_803),
.B(n_643),
.Y(n_879)
);

INVxp67_ASAP7_75t_L g880 ( 
.A(n_681),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_703),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_817),
.B(n_602),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_693),
.A2(n_556),
.B(n_539),
.Y(n_883)
);

OAI21xp5_ASAP7_75t_L g884 ( 
.A1(n_693),
.A2(n_592),
.B(n_577),
.Y(n_884)
);

INVx4_ASAP7_75t_L g885 ( 
.A(n_703),
.Y(n_885)
);

AOI21x1_ASAP7_75t_L g886 ( 
.A1(n_802),
.A2(n_664),
.B(n_665),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_705),
.Y(n_887)
);

AOI21xp5_ASAP7_75t_L g888 ( 
.A1(n_812),
.A2(n_618),
.B(n_635),
.Y(n_888)
);

AOI21x1_ASAP7_75t_L g889 ( 
.A1(n_802),
.A2(n_664),
.B(n_542),
.Y(n_889)
);

NOR2xp33_ASAP7_75t_L g890 ( 
.A(n_728),
.B(n_615),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_709),
.Y(n_891)
);

AOI21xp5_ASAP7_75t_L g892 ( 
.A1(n_804),
.A2(n_635),
.B(n_643),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_682),
.B(n_651),
.Y(n_893)
);

NAND2x1p5_ASAP7_75t_L g894 ( 
.A(n_735),
.B(n_643),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_723),
.A2(n_546),
.B(n_577),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_688),
.Y(n_896)
);

OR2x2_ASAP7_75t_L g897 ( 
.A(n_734),
.B(n_536),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_804),
.A2(n_635),
.B(n_643),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_709),
.Y(n_899)
);

O2A1O1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_720),
.A2(n_663),
.B(n_507),
.C(n_493),
.Y(n_900)
);

BUFx6f_ASAP7_75t_L g901 ( 
.A(n_688),
.Y(n_901)
);

AOI21xp5_ASAP7_75t_L g902 ( 
.A1(n_806),
.A2(n_546),
.B(n_577),
.Y(n_902)
);

AOI21xp5_ASAP7_75t_L g903 ( 
.A1(n_806),
.A2(n_735),
.B(n_683),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_721),
.B(n_722),
.Y(n_904)
);

AOI21xp5_ASAP7_75t_L g905 ( 
.A1(n_735),
.A2(n_546),
.B(n_578),
.Y(n_905)
);

CKINVDCx8_ASAP7_75t_R g906 ( 
.A(n_758),
.Y(n_906)
);

AOI21xp5_ASAP7_75t_L g907 ( 
.A1(n_757),
.A2(n_578),
.B(n_592),
.Y(n_907)
);

OAI21xp5_ASAP7_75t_L g908 ( 
.A1(n_809),
.A2(n_578),
.B(n_592),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_736),
.B(n_651),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_738),
.B(n_651),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_757),
.A2(n_656),
.B(n_621),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_SL g912 ( 
.A(n_803),
.B(n_621),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_808),
.A2(n_656),
.B(n_621),
.Y(n_913)
);

O2A1O1Ixp33_ASAP7_75t_L g914 ( 
.A1(n_762),
.A2(n_663),
.B(n_493),
.C(n_504),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_814),
.A2(n_656),
.B(n_519),
.Y(n_915)
);

HB1xp67_ASAP7_75t_L g916 ( 
.A(n_783),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_700),
.A2(n_519),
.B(n_540),
.Y(n_917)
);

AND2x6_ASAP7_75t_L g918 ( 
.A(n_685),
.B(n_540),
.Y(n_918)
);

INVx3_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_748),
.Y(n_920)
);

INVx2_ASAP7_75t_L g921 ( 
.A(n_754),
.Y(n_921)
);

BUFx3_ASAP7_75t_L g922 ( 
.A(n_783),
.Y(n_922)
);

OAI321xp33_ASAP7_75t_L g923 ( 
.A1(n_706),
.A2(n_433),
.A3(n_431),
.B1(n_430),
.B2(n_429),
.C(n_425),
.Y(n_923)
);

A2O1A1Ixp33_ASAP7_75t_L g924 ( 
.A1(n_815),
.A2(n_615),
.B(n_558),
.C(n_542),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_754),
.Y(n_925)
);

NOR2xp33_ASAP7_75t_R g926 ( 
.A(n_816),
.B(n_558),
.Y(n_926)
);

AOI21xp5_ASAP7_75t_L g927 ( 
.A1(n_798),
.A2(n_440),
.B(n_443),
.Y(n_927)
);

AOI22xp5_ASAP7_75t_L g928 ( 
.A1(n_689),
.A2(n_667),
.B1(n_651),
.B2(n_516),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_777),
.Y(n_929)
);

O2A1O1Ixp33_ASAP7_75t_L g930 ( 
.A1(n_762),
.A2(n_507),
.B(n_516),
.C(n_419),
.Y(n_930)
);

OAI21xp33_ASAP7_75t_L g931 ( 
.A1(n_827),
.A2(n_321),
.B(n_326),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_739),
.B(n_651),
.Y(n_932)
);

AOI21x1_ASAP7_75t_L g933 ( 
.A1(n_813),
.A2(n_454),
.B(n_440),
.Y(n_933)
);

OAI21xp5_ASAP7_75t_L g934 ( 
.A1(n_672),
.A2(n_667),
.B(n_651),
.Y(n_934)
);

OAI21xp5_ASAP7_75t_L g935 ( 
.A1(n_805),
.A2(n_667),
.B(n_454),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_696),
.B(n_240),
.Y(n_936)
);

OAI21xp5_ASAP7_75t_L g937 ( 
.A1(n_674),
.A2(n_667),
.B(n_456),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_710),
.B(n_411),
.Y(n_938)
);

BUFx6f_ASAP7_75t_L g939 ( 
.A(n_777),
.Y(n_939)
);

INVx2_ASAP7_75t_L g940 ( 
.A(n_764),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_718),
.A2(n_516),
.B(n_431),
.C(n_430),
.Y(n_941)
);

INVx3_ASAP7_75t_L g942 ( 
.A(n_782),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_791),
.A2(n_456),
.B(n_516),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_799),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_764),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_746),
.B(n_559),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_692),
.A2(n_667),
.B1(n_476),
.B2(n_467),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_740),
.B(n_476),
.Y(n_948)
);

AOI21xp5_ASAP7_75t_L g949 ( 
.A1(n_791),
.A2(n_459),
.B(n_318),
.Y(n_949)
);

NOR2xp33_ASAP7_75t_L g950 ( 
.A(n_800),
.B(n_314),
.Y(n_950)
);

NOR2xp33_ASAP7_75t_L g951 ( 
.A(n_800),
.B(n_315),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_743),
.B(n_476),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_694),
.A2(n_352),
.B1(n_320),
.B2(n_329),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_729),
.A2(n_459),
.B(n_476),
.Y(n_954)
);

AND2x6_ASAP7_75t_L g955 ( 
.A(n_704),
.B(n_714),
.Y(n_955)
);

AND2x2_ASAP7_75t_L g956 ( 
.A(n_759),
.B(n_243),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

AND2x4_ASAP7_75t_L g958 ( 
.A(n_750),
.B(n_424),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_833),
.A2(n_771),
.B(n_777),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_768),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_776),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_752),
.B(n_459),
.Y(n_962)
);

AOI22xp5_ASAP7_75t_L g963 ( 
.A1(n_824),
.A2(n_467),
.B1(n_207),
.B2(n_275),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_771),
.A2(n_459),
.B(n_425),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_790),
.A2(n_835),
.B(n_785),
.C(n_671),
.Y(n_965)
);

AND2x2_ASAP7_75t_L g966 ( 
.A(n_795),
.B(n_243),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_753),
.B(n_760),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_776),
.Y(n_968)
);

BUFx2_ASAP7_75t_L g969 ( 
.A(n_818),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_777),
.A2(n_770),
.B(n_782),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_770),
.A2(n_437),
.B(n_435),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_834),
.A2(n_437),
.B(n_435),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_769),
.A2(n_778),
.B1(n_786),
.B2(n_789),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_793),
.B(n_337),
.Y(n_974)
);

AO21x1_ASAP7_75t_L g975 ( 
.A1(n_792),
.A2(n_433),
.B(n_429),
.Y(n_975)
);

NOR2x1p5_ASAP7_75t_SL g976 ( 
.A(n_803),
.B(n_422),
.Y(n_976)
);

O2A1O1Ixp33_ASAP7_75t_L g977 ( 
.A1(n_718),
.A2(n_313),
.B(n_275),
.C(n_282),
.Y(n_977)
);

AOI21xp5_ASAP7_75t_L g978 ( 
.A1(n_836),
.A2(n_348),
.B(n_346),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_837),
.A2(n_336),
.B(n_467),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_792),
.A2(n_467),
.B(n_131),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_779),
.A2(n_467),
.B(n_141),
.Y(n_981)
);

AOI21xp5_ASAP7_75t_L g982 ( 
.A1(n_788),
.A2(n_467),
.B(n_125),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_730),
.B(n_313),
.Y(n_983)
);

NOR2xp67_ASAP7_75t_L g984 ( 
.A(n_715),
.B(n_172),
.Y(n_984)
);

OAI22xp5_ASAP7_75t_L g985 ( 
.A1(n_818),
.A2(n_313),
.B1(n_282),
.B2(n_275),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_780),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_807),
.B(n_260),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_726),
.A2(n_122),
.B(n_81),
.Y(n_988)
);

OAI21xp5_ASAP7_75t_L g989 ( 
.A1(n_787),
.A2(n_313),
.B(n_282),
.Y(n_989)
);

AOI21x1_ASAP7_75t_L g990 ( 
.A1(n_775),
.A2(n_282),
.B(n_275),
.Y(n_990)
);

AOI21xp5_ASAP7_75t_L g991 ( 
.A1(n_724),
.A2(n_107),
.B(n_84),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_730),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_780),
.Y(n_993)
);

BUFx2_ASAP7_75t_L g994 ( 
.A(n_838),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_730),
.B(n_5),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_732),
.B(n_6),
.Y(n_996)
);

OAI22xp33_ASAP7_75t_L g997 ( 
.A1(n_838),
.A2(n_260),
.B1(n_243),
.B2(n_20),
.Y(n_997)
);

OAI22xp5_ASAP7_75t_L g998 ( 
.A1(n_838),
.A2(n_111),
.B1(n_101),
.B2(n_161),
.Y(n_998)
);

O2A1O1Ixp5_ASAP7_75t_L g999 ( 
.A1(n_784),
.A2(n_260),
.B(n_243),
.C(n_20),
.Y(n_999)
);

NOR2xp67_ASAP7_75t_L g1000 ( 
.A(n_691),
.B(n_155),
.Y(n_1000)
);

OAI22xp5_ASAP7_75t_L g1001 ( 
.A1(n_838),
.A2(n_105),
.B1(n_74),
.B2(n_260),
.Y(n_1001)
);

AO21x2_ASAP7_75t_L g1002 ( 
.A1(n_744),
.A2(n_773),
.B(n_725),
.Y(n_1002)
);

AOI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_732),
.A2(n_9),
.B1(n_16),
.B2(n_21),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_731),
.A2(n_9),
.B(n_16),
.Y(n_1004)
);

NOR2x1_ASAP7_75t_L g1005 ( 
.A(n_810),
.B(n_22),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_784),
.Y(n_1006)
);

OAI22xp5_ASAP7_75t_L g1007 ( 
.A1(n_670),
.A2(n_68),
.B1(n_27),
.B2(n_29),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_732),
.A2(n_26),
.B(n_27),
.C(n_29),
.Y(n_1008)
);

OAI21xp33_ASAP7_75t_L g1009 ( 
.A1(n_751),
.A2(n_26),
.B(n_30),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_733),
.A2(n_30),
.B(n_31),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_SL g1011 ( 
.A(n_763),
.B(n_31),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_670),
.B(n_33),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_741),
.A2(n_37),
.B(n_38),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_670),
.B(n_38),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_840),
.A2(n_39),
.B(n_40),
.Y(n_1015)
);

AND2x4_ASAP7_75t_L g1016 ( 
.A(n_794),
.B(n_39),
.Y(n_1016)
);

AO21x1_ASAP7_75t_L g1017 ( 
.A1(n_742),
.A2(n_40),
.B(n_41),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_840),
.A2(n_841),
.B(n_767),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_745),
.A2(n_747),
.B(n_774),
.Y(n_1019)
);

NOR2xp33_ASAP7_75t_L g1020 ( 
.A(n_819),
.B(n_44),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_749),
.A2(n_47),
.B(n_48),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_761),
.A2(n_50),
.B(n_52),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_830),
.B(n_54),
.Y(n_1023)
);

AND2x2_ASAP7_75t_L g1024 ( 
.A(n_697),
.B(n_67),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_822),
.A2(n_56),
.B(n_57),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_697),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_L g1027 ( 
.A(n_832),
.B(n_56),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_796),
.B(n_57),
.Y(n_1028)
);

NOR2xp33_ASAP7_75t_L g1029 ( 
.A(n_796),
.B(n_58),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_823),
.Y(n_1030)
);

INVx3_ASAP7_75t_L g1031 ( 
.A(n_823),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_841),
.Y(n_1032)
);

NOR2xp33_ASAP7_75t_L g1033 ( 
.A(n_845),
.B(n_755),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_959),
.A2(n_765),
.B(n_767),
.Y(n_1034)
);

O2A1O1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_965),
.A2(n_737),
.B(n_831),
.C(n_829),
.Y(n_1035)
);

AOI22xp5_ASAP7_75t_L g1036 ( 
.A1(n_890),
.A2(n_717),
.B1(n_803),
.B2(n_675),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_845),
.B(n_690),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_842),
.B(n_756),
.Y(n_1038)
);

INVx2_ASAP7_75t_SL g1039 ( 
.A(n_863),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_1031),
.Y(n_1040)
);

BUFx2_ASAP7_75t_L g1041 ( 
.A(n_843),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_944),
.B(n_803),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_1031),
.Y(n_1043)
);

OAI22xp5_ASAP7_75t_L g1044 ( 
.A1(n_876),
.A2(n_698),
.B1(n_828),
.B2(n_801),
.Y(n_1044)
);

OA22x2_ASAP7_75t_L g1045 ( 
.A1(n_944),
.A2(n_781),
.B1(n_675),
.B2(n_690),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_890),
.B(n_825),
.Y(n_1046)
);

HB1xp67_ASAP7_75t_L g1047 ( 
.A(n_916),
.Y(n_1047)
);

AND2x2_ASAP7_75t_L g1048 ( 
.A(n_882),
.B(n_822),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_868),
.A2(n_761),
.B(n_765),
.Y(n_1049)
);

NAND2xp5_ASAP7_75t_SL g1050 ( 
.A(n_992),
.B(n_766),
.Y(n_1050)
);

AOI21x1_ASAP7_75t_L g1051 ( 
.A1(n_877),
.A2(n_825),
.B(n_772),
.Y(n_1051)
);

AOI21x1_ASAP7_75t_L g1052 ( 
.A1(n_877),
.A2(n_839),
.B(n_820),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_891),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_SL g1054 ( 
.A(n_992),
.B(n_820),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_945),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_1015),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_1056)
);

OA22x2_ASAP7_75t_L g1057 ( 
.A1(n_880),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1057)
);

CKINVDCx14_ASAP7_75t_R g1058 ( 
.A(n_859),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_868),
.A2(n_64),
.B(n_65),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_876),
.B(n_67),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_987),
.B(n_967),
.Y(n_1061)
);

INVx2_ASAP7_75t_L g1062 ( 
.A(n_844),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_SL g1063 ( 
.A(n_992),
.B(n_853),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_903),
.A2(n_878),
.B(n_875),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_865),
.Y(n_1065)
);

AND2x4_ASAP7_75t_L g1066 ( 
.A(n_922),
.B(n_969),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_957),
.Y(n_1067)
);

HB1xp67_ASAP7_75t_L g1068 ( 
.A(n_916),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_960),
.Y(n_1069)
);

AND2x4_ASAP7_75t_L g1070 ( 
.A(n_994),
.B(n_896),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_871),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_848),
.A2(n_895),
.B(n_847),
.Y(n_1072)
);

OAI22xp5_ASAP7_75t_L g1073 ( 
.A1(n_855),
.A2(n_858),
.B1(n_856),
.B2(n_851),
.Y(n_1073)
);

OAI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_849),
.A2(n_864),
.B(n_861),
.Y(n_1074)
);

NOR3xp33_ASAP7_75t_SL g1075 ( 
.A(n_869),
.B(n_997),
.C(n_924),
.Y(n_1075)
);

A2O1A1Ixp33_ASAP7_75t_L g1076 ( 
.A1(n_1009),
.A2(n_883),
.B(n_862),
.C(n_1003),
.Y(n_1076)
);

NAND2x1p5_ASAP7_75t_L g1077 ( 
.A(n_929),
.B(n_939),
.Y(n_1077)
);

INVx3_ASAP7_75t_SL g1078 ( 
.A(n_897),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_961),
.Y(n_1079)
);

O2A1O1Ixp5_ASAP7_75t_L g1080 ( 
.A1(n_938),
.A2(n_934),
.B(n_949),
.C(n_937),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_872),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_887),
.Y(n_1082)
);

BUFx12f_ASAP7_75t_L g1083 ( 
.A(n_1026),
.Y(n_1083)
);

O2A1O1Ixp33_ASAP7_75t_L g1084 ( 
.A1(n_880),
.A2(n_997),
.B(n_931),
.C(n_1007),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_871),
.B(n_862),
.Y(n_1085)
);

OR2x6_ASAP7_75t_L g1086 ( 
.A(n_992),
.B(n_896),
.Y(n_1086)
);

BUFx3_ASAP7_75t_L g1087 ( 
.A(n_896),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_936),
.B(n_956),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_SL g1089 ( 
.A1(n_1029),
.A2(n_1020),
.B(n_935),
.C(n_900),
.Y(n_1089)
);

INVxp67_ASAP7_75t_L g1090 ( 
.A(n_950),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_869),
.B(n_874),
.Y(n_1091)
);

NAND3xp33_ASAP7_75t_SL g1092 ( 
.A(n_1011),
.B(n_946),
.C(n_926),
.Y(n_1092)
);

AOI22xp33_ASAP7_75t_L g1093 ( 
.A1(n_1012),
.A2(n_1014),
.B1(n_1017),
.B2(n_989),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_904),
.B(n_958),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_1016),
.Y(n_1095)
);

NOR2xp33_ASAP7_75t_L g1096 ( 
.A(n_950),
.B(n_951),
.Y(n_1096)
);

O2A1O1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_1008),
.A2(n_973),
.B(n_985),
.C(n_995),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_958),
.B(n_966),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_893),
.A2(n_850),
.B(n_888),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_899),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_996),
.A2(n_1027),
.B(n_1023),
.C(n_974),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_894),
.A2(n_857),
.B(n_860),
.Y(n_1102)
);

AND2x2_ASAP7_75t_L g1103 ( 
.A(n_951),
.B(n_1024),
.Y(n_1103)
);

A2O1A1Ixp33_ASAP7_75t_L g1104 ( 
.A1(n_1020),
.A2(n_1005),
.B(n_999),
.C(n_1029),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_866),
.B(n_881),
.Y(n_1105)
);

OAI22xp5_ASAP7_75t_L g1106 ( 
.A1(n_846),
.A2(n_867),
.B1(n_896),
.B2(n_901),
.Y(n_1106)
);

AND2x2_ASAP7_75t_L g1107 ( 
.A(n_946),
.B(n_1016),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_926),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_846),
.A2(n_867),
.B1(n_901),
.B2(n_873),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_901),
.B(n_983),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_866),
.B(n_881),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_SL g1112 ( 
.A(n_870),
.B(n_919),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_894),
.A2(n_970),
.B(n_908),
.Y(n_1113)
);

OAI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_901),
.A2(n_939),
.B1(n_929),
.B2(n_870),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_870),
.B(n_919),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_968),
.B(n_993),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_912),
.A2(n_879),
.B(n_1019),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_953),
.B(n_984),
.Y(n_1118)
);

AND2x2_ASAP7_75t_L g1119 ( 
.A(n_920),
.B(n_921),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_912),
.A2(n_879),
.B(n_884),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_1028),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_870),
.B(n_942),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_942),
.Y(n_1123)
);

INVxp67_ASAP7_75t_L g1124 ( 
.A(n_978),
.Y(n_1124)
);

AOI21xp5_ASAP7_75t_L g1125 ( 
.A1(n_913),
.A2(n_905),
.B(n_932),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_885),
.B(n_925),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_885),
.B(n_940),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_909),
.A2(n_910),
.B(n_915),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_R g1129 ( 
.A(n_906),
.B(n_929),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_998),
.A2(n_1001),
.B1(n_1000),
.B2(n_1021),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1032),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_986),
.B(n_1030),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_SL g1133 ( 
.A(n_929),
.B(n_939),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_892),
.A2(n_898),
.B(n_902),
.Y(n_1134)
);

BUFx2_ASAP7_75t_L g1135 ( 
.A(n_1006),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_911),
.A2(n_907),
.B(n_1018),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_939),
.B(n_928),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_962),
.Y(n_1138)
);

NOR2xp33_ASAP7_75t_L g1139 ( 
.A(n_948),
.B(n_952),
.Y(n_1139)
);

O2A1O1Ixp5_ASAP7_75t_SL g1140 ( 
.A1(n_977),
.A2(n_999),
.B(n_990),
.C(n_930),
.Y(n_1140)
);

CKINVDCx20_ASAP7_75t_R g1141 ( 
.A(n_963),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_SL g1142 ( 
.A(n_852),
.B(n_854),
.Y(n_1142)
);

O2A1O1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_977),
.A2(n_923),
.B(n_1010),
.C(n_1013),
.Y(n_1143)
);

INVx3_ASAP7_75t_L g1144 ( 
.A(n_918),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_889),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_971),
.A2(n_1022),
.B(n_1004),
.C(n_930),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_947),
.B(n_975),
.Y(n_1147)
);

AND2x2_ASAP7_75t_L g1148 ( 
.A(n_1002),
.B(n_972),
.Y(n_1148)
);

AOI22xp5_ASAP7_75t_L g1149 ( 
.A1(n_955),
.A2(n_918),
.B1(n_1002),
.B2(n_979),
.Y(n_1149)
);

AND2x2_ASAP7_75t_L g1150 ( 
.A(n_1025),
.B(n_941),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_976),
.A2(n_988),
.B(n_941),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_886),
.B(n_964),
.Y(n_1152)
);

NOR2xp33_ASAP7_75t_R g1153 ( 
.A(n_955),
.B(n_933),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_955),
.A2(n_918),
.B1(n_943),
.B2(n_927),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_900),
.B(n_917),
.Y(n_1155)
);

A2O1A1Ixp33_ASAP7_75t_L g1156 ( 
.A1(n_914),
.A2(n_991),
.B(n_980),
.C(n_981),
.Y(n_1156)
);

INVx6_ASAP7_75t_L g1157 ( 
.A(n_955),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_918),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_918),
.Y(n_1159)
);

A2O1A1Ixp33_ASAP7_75t_L g1160 ( 
.A1(n_914),
.A2(n_982),
.B(n_954),
.C(n_955),
.Y(n_1160)
);

A2O1A1Ixp33_ASAP7_75t_L g1161 ( 
.A1(n_890),
.A2(n_673),
.B(n_684),
.C(n_965),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_965),
.A2(n_673),
.B(n_684),
.C(n_842),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_842),
.A2(n_673),
.B1(n_684),
.B2(n_845),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_SL g1164 ( 
.A(n_842),
.B(n_673),
.Y(n_1164)
);

AND2x4_ASAP7_75t_L g1165 ( 
.A(n_922),
.B(n_969),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_842),
.B(n_673),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1031),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_916),
.Y(n_1168)
);

AOI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_959),
.A2(n_713),
.B(n_531),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_843),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_870),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_965),
.A2(n_673),
.B(n_684),
.C(n_842),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_870),
.Y(n_1173)
);

BUFx3_ASAP7_75t_L g1174 ( 
.A(n_843),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_L g1175 ( 
.A(n_845),
.B(n_673),
.Y(n_1175)
);

BUFx2_ASAP7_75t_L g1176 ( 
.A(n_843),
.Y(n_1176)
);

OAI22xp5_ASAP7_75t_L g1177 ( 
.A1(n_842),
.A2(n_673),
.B1(n_684),
.B2(n_845),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_959),
.A2(n_713),
.B(n_531),
.Y(n_1178)
);

CKINVDCx14_ASAP7_75t_R g1179 ( 
.A(n_859),
.Y(n_1179)
);

BUFx8_ASAP7_75t_SL g1180 ( 
.A(n_859),
.Y(n_1180)
);

NOR3xp33_ASAP7_75t_SL g1181 ( 
.A(n_869),
.B(n_558),
.C(n_536),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_891),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_L g1183 ( 
.A1(n_890),
.A2(n_673),
.B(n_684),
.C(n_965),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_842),
.B(n_673),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_870),
.Y(n_1185)
);

NOR2xp33_ASAP7_75t_L g1186 ( 
.A(n_845),
.B(n_673),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_842),
.B(n_673),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1031),
.Y(n_1188)
);

AND2x2_ASAP7_75t_L g1189 ( 
.A(n_882),
.B(n_679),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_891),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_959),
.A2(n_713),
.B(n_531),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_891),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1053),
.Y(n_1193)
);

O2A1O1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1175),
.A2(n_1186),
.B(n_1163),
.C(n_1177),
.Y(n_1194)
);

OAI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1175),
.A2(n_1186),
.B1(n_1033),
.B2(n_1096),
.Y(n_1195)
);

OAI21x1_ASAP7_75t_L g1196 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1196)
);

NOR2x1_ASAP7_75t_L g1197 ( 
.A(n_1042),
.B(n_1061),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1096),
.B(n_1090),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1199)
);

O2A1O1Ixp33_ASAP7_75t_L g1200 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_1033),
.C(n_1166),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1088),
.B(n_1103),
.Y(n_1201)
);

AND2x4_ASAP7_75t_L g1202 ( 
.A(n_1070),
.B(n_1095),
.Y(n_1202)
);

CKINVDCx20_ASAP7_75t_R g1203 ( 
.A(n_1180),
.Y(n_1203)
);

AO32x2_ASAP7_75t_L g1204 ( 
.A1(n_1073),
.A2(n_1044),
.A3(n_1109),
.B1(n_1106),
.B2(n_1093),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1064),
.A2(n_1134),
.B(n_1169),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_1058),
.Y(n_1206)
);

BUFx2_ASAP7_75t_L g1207 ( 
.A(n_1041),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1119),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1072),
.A2(n_1074),
.B(n_1113),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1184),
.B(n_1187),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1178),
.A2(n_1191),
.B(n_1172),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1162),
.A2(n_1080),
.B(n_1136),
.Y(n_1212)
);

BUFx2_ASAP7_75t_L g1213 ( 
.A(n_1176),
.Y(n_1213)
);

INVx2_ASAP7_75t_SL g1214 ( 
.A(n_1170),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1117),
.A2(n_1089),
.B(n_1035),
.Y(n_1215)
);

BUFx6f_ASAP7_75t_L g1216 ( 
.A(n_1185),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1051),
.A2(n_1128),
.B(n_1052),
.Y(n_1217)
);

NAND2x1_ASAP7_75t_L g1218 ( 
.A(n_1157),
.B(n_1086),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1089),
.A2(n_1137),
.B(n_1101),
.Y(n_1219)
);

OA21x2_ASAP7_75t_L g1220 ( 
.A1(n_1142),
.A2(n_1151),
.B(n_1160),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1091),
.A2(n_1097),
.B(n_1084),
.C(n_1076),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1091),
.A2(n_1076),
.B(n_1075),
.C(n_1143),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1137),
.A2(n_1164),
.B(n_1160),
.Y(n_1223)
);

AO32x2_ASAP7_75t_L g1224 ( 
.A1(n_1093),
.A2(n_1114),
.A3(n_1140),
.B1(n_1056),
.B2(n_1104),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_L g1225 ( 
.A(n_1164),
.B(n_1094),
.Y(n_1225)
);

OAI21x1_ASAP7_75t_L g1226 ( 
.A1(n_1034),
.A2(n_1142),
.B(n_1120),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1139),
.A2(n_1155),
.B(n_1046),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1139),
.A2(n_1124),
.B(n_1156),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1156),
.A2(n_1038),
.B(n_1050),
.Y(n_1229)
);

AND2x4_ASAP7_75t_L g1230 ( 
.A(n_1070),
.B(n_1066),
.Y(n_1230)
);

OAI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1049),
.A2(n_1060),
.B(n_1063),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1043),
.Y(n_1232)
);

NAND2xp5_ASAP7_75t_L g1233 ( 
.A(n_1189),
.B(n_1121),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1055),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1067),
.Y(n_1235)
);

AOI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1050),
.A2(n_1054),
.B(n_1130),
.Y(n_1236)
);

AOI21x1_ASAP7_75t_SL g1237 ( 
.A1(n_1118),
.A2(n_1148),
.B(n_1150),
.Y(n_1237)
);

NOR2xp33_ASAP7_75t_L g1238 ( 
.A(n_1085),
.B(n_1037),
.Y(n_1238)
);

NOR2x1_ASAP7_75t_L g1239 ( 
.A(n_1144),
.B(n_1063),
.Y(n_1239)
);

HB1xp67_ASAP7_75t_L g1240 ( 
.A(n_1071),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1039),
.B(n_1098),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1066),
.B(n_1165),
.Y(n_1242)
);

O2A1O1Ixp33_ASAP7_75t_SL g1243 ( 
.A1(n_1056),
.A2(n_1054),
.B(n_1147),
.C(n_1115),
.Y(n_1243)
);

AOI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1130),
.A2(n_1146),
.B(n_1147),
.Y(n_1244)
);

A2O1A1Ixp33_ASAP7_75t_L g1245 ( 
.A1(n_1110),
.A2(n_1059),
.B(n_1036),
.C(n_1181),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1146),
.A2(n_1110),
.B(n_1152),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1185),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1170),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1138),
.A2(n_1149),
.B(n_1133),
.Y(n_1249)
);

OAI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1048),
.A2(n_1116),
.B(n_1132),
.Y(n_1250)
);

AOI22xp5_ASAP7_75t_L g1251 ( 
.A1(n_1141),
.A2(n_1085),
.B1(n_1107),
.B2(n_1037),
.Y(n_1251)
);

CKINVDCx11_ASAP7_75t_R g1252 ( 
.A(n_1083),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1043),
.Y(n_1253)
);

A2O1A1Ixp33_ASAP7_75t_L g1254 ( 
.A1(n_1092),
.A2(n_1127),
.B(n_1126),
.C(n_1154),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_SL g1255 ( 
.A1(n_1159),
.A2(n_1105),
.B(n_1111),
.Y(n_1255)
);

AO31x2_ASAP7_75t_L g1256 ( 
.A1(n_1145),
.A2(n_1126),
.A3(n_1127),
.B(n_1192),
.Y(n_1256)
);

O2A1O1Ixp33_ASAP7_75t_L g1257 ( 
.A1(n_1078),
.A2(n_1068),
.B(n_1047),
.C(n_1168),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1135),
.B(n_1190),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1069),
.B(n_1182),
.Y(n_1259)
);

NAND3xp33_ASAP7_75t_SL g1260 ( 
.A(n_1129),
.B(n_1153),
.C(n_1131),
.Y(n_1260)
);

AOI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_1057),
.A2(n_1045),
.B1(n_1078),
.B2(n_1108),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1133),
.A2(n_1122),
.B(n_1112),
.Y(n_1262)
);

AO31x2_ASAP7_75t_L g1263 ( 
.A1(n_1079),
.A2(n_1040),
.A3(n_1167),
.B(n_1188),
.Y(n_1263)
);

AO31x2_ASAP7_75t_L g1264 ( 
.A1(n_1062),
.A2(n_1081),
.A3(n_1065),
.B(n_1100),
.Y(n_1264)
);

AOI21xp5_ASAP7_75t_L g1265 ( 
.A1(n_1112),
.A2(n_1122),
.B(n_1115),
.Y(n_1265)
);

O2A1O1Ixp33_ASAP7_75t_L g1266 ( 
.A1(n_1174),
.A2(n_1123),
.B(n_1165),
.C(n_1086),
.Y(n_1266)
);

A2O1A1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1144),
.A2(n_1087),
.B(n_1171),
.C(n_1173),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1087),
.B(n_1174),
.Y(n_1268)
);

AO22x2_ASAP7_75t_L g1269 ( 
.A1(n_1057),
.A2(n_1173),
.B1(n_1171),
.B2(n_1045),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1185),
.Y(n_1270)
);

NAND2xp33_ASAP7_75t_SL g1271 ( 
.A(n_1129),
.B(n_1153),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1086),
.B(n_1157),
.Y(n_1272)
);

BUFx2_ASAP7_75t_L g1273 ( 
.A(n_1179),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1157),
.B(n_1077),
.Y(n_1274)
);

BUFx2_ASAP7_75t_L g1275 ( 
.A(n_1077),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1189),
.B(n_532),
.Y(n_1276)
);

BUFx8_ASAP7_75t_L g1277 ( 
.A(n_1041),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1161),
.A2(n_673),
.B(n_1183),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_965),
.C(n_1056),
.Y(n_1279)
);

OAI22xp5_ASAP7_75t_L g1280 ( 
.A1(n_1175),
.A2(n_673),
.B1(n_1186),
.B2(n_1096),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1070),
.B(n_1095),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_SL g1283 ( 
.A(n_1096),
.B(n_673),
.Y(n_1283)
);

INVx1_ASAP7_75t_L g1284 ( 
.A(n_1053),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1175),
.B(n_673),
.Y(n_1286)
);

BUFx6f_ASAP7_75t_L g1287 ( 
.A(n_1185),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1288)
);

O2A1O1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_965),
.C(n_1056),
.Y(n_1289)
);

BUFx6f_ASAP7_75t_L g1290 ( 
.A(n_1185),
.Y(n_1290)
);

INVx6_ASAP7_75t_L g1291 ( 
.A(n_1170),
.Y(n_1291)
);

AO32x2_ASAP7_75t_L g1292 ( 
.A1(n_1163),
.A2(n_1177),
.A3(n_1007),
.B1(n_1073),
.B2(n_1044),
.Y(n_1292)
);

O2A1O1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1175),
.A2(n_673),
.B(n_1186),
.C(n_1177),
.Y(n_1293)
);

NOR2xp33_ASAP7_75t_L g1294 ( 
.A(n_1175),
.B(n_1186),
.Y(n_1294)
);

O2A1O1Ixp33_ASAP7_75t_L g1295 ( 
.A1(n_1175),
.A2(n_673),
.B(n_1186),
.C(n_1177),
.Y(n_1295)
);

AOI21xp5_ASAP7_75t_L g1296 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1175),
.B(n_673),
.Y(n_1297)
);

OAI21x1_ASAP7_75t_L g1298 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1298)
);

AOI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1157),
.Y(n_1300)
);

AND2x2_ASAP7_75t_L g1301 ( 
.A(n_1189),
.B(n_882),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1302)
);

BUFx10_ASAP7_75t_L g1303 ( 
.A(n_1066),
.Y(n_1303)
);

NOR3xp33_ASAP7_75t_L g1304 ( 
.A(n_1096),
.B(n_673),
.C(n_684),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_SL g1305 ( 
.A1(n_1097),
.A2(n_1059),
.B(n_1101),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1053),
.Y(n_1306)
);

AOI21xp5_ASAP7_75t_L g1307 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1307)
);

AOI21xp5_ASAP7_75t_L g1308 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1309)
);

AOI21xp33_ASAP7_75t_L g1310 ( 
.A1(n_1096),
.A2(n_673),
.B(n_684),
.Y(n_1310)
);

AND2x4_ASAP7_75t_L g1311 ( 
.A(n_1070),
.B(n_1095),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1313)
);

AO31x2_ASAP7_75t_L g1314 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1314)
);

AOI21xp5_ASAP7_75t_SL g1315 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_673),
.Y(n_1315)
);

A2O1A1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1175),
.A2(n_673),
.B(n_1186),
.C(n_1096),
.Y(n_1316)
);

AOI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1317)
);

CKINVDCx20_ASAP7_75t_R g1318 ( 
.A(n_1180),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1175),
.B(n_673),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1142),
.Y(n_1322)
);

CKINVDCx5p33_ASAP7_75t_R g1323 ( 
.A(n_1180),
.Y(n_1323)
);

NAND3xp33_ASAP7_75t_L g1324 ( 
.A(n_1175),
.B(n_673),
.C(n_684),
.Y(n_1324)
);

NOR2xp33_ASAP7_75t_SL g1325 ( 
.A(n_1180),
.B(n_532),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_965),
.C(n_1056),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1074),
.A2(n_1072),
.B(n_1142),
.Y(n_1327)
);

O2A1O1Ixp33_ASAP7_75t_SL g1328 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_965),
.C(n_1056),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_1144),
.B(n_1158),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1330)
);

INVx5_ASAP7_75t_L g1331 ( 
.A(n_1086),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1161),
.A2(n_1183),
.B(n_673),
.Y(n_1332)
);

INVx2_ASAP7_75t_SL g1333 ( 
.A(n_1170),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1053),
.Y(n_1334)
);

AO31x2_ASAP7_75t_L g1335 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1082),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1086),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1175),
.B(n_673),
.Y(n_1338)
);

AND2x4_ASAP7_75t_L g1339 ( 
.A(n_1070),
.B(n_1095),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1053),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1341)
);

A2O1A1Ixp33_ASAP7_75t_L g1342 ( 
.A1(n_1175),
.A2(n_673),
.B(n_1186),
.C(n_1096),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1053),
.Y(n_1343)
);

INVx2_ASAP7_75t_L g1344 ( 
.A(n_1082),
.Y(n_1344)
);

HB1xp67_ASAP7_75t_L g1345 ( 
.A(n_1071),
.Y(n_1345)
);

HB1xp67_ASAP7_75t_L g1346 ( 
.A(n_1071),
.Y(n_1346)
);

OAI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1102),
.A2(n_1099),
.B(n_1125),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1053),
.Y(n_1348)
);

AO31x2_ASAP7_75t_L g1349 ( 
.A1(n_1104),
.A2(n_1155),
.A3(n_1161),
.B(n_1183),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1072),
.A2(n_673),
.B(n_1074),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1047),
.Y(n_1351)
);

NAND2xp5_ASAP7_75t_L g1352 ( 
.A(n_1175),
.B(n_673),
.Y(n_1352)
);

OAI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1161),
.A2(n_673),
.B(n_1183),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1259),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1193),
.Y(n_1355)
);

BUFx2_ASAP7_75t_R g1356 ( 
.A(n_1323),
.Y(n_1356)
);

INVx4_ASAP7_75t_L g1357 ( 
.A(n_1331),
.Y(n_1357)
);

OAI22xp5_ASAP7_75t_L g1358 ( 
.A1(n_1324),
.A2(n_1195),
.B1(n_1342),
.B2(n_1316),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1304),
.A2(n_1310),
.B1(n_1280),
.B2(n_1324),
.Y(n_1359)
);

INVx6_ASAP7_75t_L g1360 ( 
.A(n_1277),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1294),
.A2(n_1283),
.B1(n_1352),
.B2(n_1286),
.Y(n_1361)
);

OAI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1297),
.A2(n_1338),
.B1(n_1319),
.B2(n_1251),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1234),
.Y(n_1363)
);

INVx4_ASAP7_75t_L g1364 ( 
.A(n_1331),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1235),
.Y(n_1365)
);

OAI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1251),
.A2(n_1261),
.B1(n_1238),
.B2(n_1210),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1284),
.Y(n_1367)
);

OAI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1261),
.A2(n_1353),
.B1(n_1278),
.B2(n_1244),
.Y(n_1368)
);

BUFx2_ASAP7_75t_L g1369 ( 
.A(n_1207),
.Y(n_1369)
);

INVx6_ASAP7_75t_L g1370 ( 
.A(n_1277),
.Y(n_1370)
);

INVx6_ASAP7_75t_L g1371 ( 
.A(n_1331),
.Y(n_1371)
);

OAI21xp5_ASAP7_75t_SL g1372 ( 
.A1(n_1293),
.A2(n_1295),
.B(n_1194),
.Y(n_1372)
);

CKINVDCx11_ASAP7_75t_R g1373 ( 
.A(n_1318),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1306),
.Y(n_1374)
);

INVx3_ASAP7_75t_L g1375 ( 
.A(n_1300),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1198),
.A2(n_1222),
.B1(n_1221),
.B2(n_1233),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1300),
.Y(n_1377)
);

BUFx5_ASAP7_75t_L g1378 ( 
.A(n_1329),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1334),
.Y(n_1379)
);

BUFx4_ASAP7_75t_SL g1380 ( 
.A(n_1206),
.Y(n_1380)
);

OAI22x1_ASAP7_75t_SL g1381 ( 
.A1(n_1214),
.A2(n_1333),
.B1(n_1325),
.B2(n_1252),
.Y(n_1381)
);

CKINVDCx11_ASAP7_75t_R g1382 ( 
.A(n_1273),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_L g1383 ( 
.A1(n_1201),
.A2(n_1305),
.B1(n_1301),
.B2(n_1350),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_L g1384 ( 
.A1(n_1282),
.A2(n_1302),
.B1(n_1312),
.B2(n_1317),
.Y(n_1384)
);

INVx8_ASAP7_75t_L g1385 ( 
.A(n_1329),
.Y(n_1385)
);

BUFx6f_ASAP7_75t_L g1386 ( 
.A(n_1291),
.Y(n_1386)
);

AOI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1241),
.A2(n_1225),
.B1(n_1276),
.B2(n_1260),
.Y(n_1387)
);

CKINVDCx20_ASAP7_75t_R g1388 ( 
.A(n_1213),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1296),
.A2(n_1308),
.B1(n_1313),
.B2(n_1299),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1340),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1343),
.Y(n_1391)
);

INVx8_ASAP7_75t_L g1392 ( 
.A(n_1329),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1348),
.Y(n_1393)
);

AOI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1307),
.A2(n_1341),
.B1(n_1197),
.B2(n_1219),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_SL g1395 ( 
.A1(n_1236),
.A2(n_1227),
.B1(n_1269),
.B2(n_1229),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1269),
.A2(n_1223),
.B1(n_1228),
.B2(n_1351),
.Y(n_1396)
);

INVx3_ASAP7_75t_SL g1397 ( 
.A(n_1291),
.Y(n_1397)
);

OAI22xp33_ASAP7_75t_L g1398 ( 
.A1(n_1258),
.A2(n_1208),
.B1(n_1250),
.B2(n_1346),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1336),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1254),
.A2(n_1245),
.B1(n_1315),
.B2(n_1332),
.Y(n_1400)
);

CKINVDCx6p67_ASAP7_75t_R g1401 ( 
.A(n_1303),
.Y(n_1401)
);

AND2x2_ASAP7_75t_L g1402 ( 
.A(n_1230),
.B(n_1242),
.Y(n_1402)
);

BUFx3_ASAP7_75t_L g1403 ( 
.A(n_1248),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1344),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1264),
.Y(n_1405)
);

INVx6_ASAP7_75t_L g1406 ( 
.A(n_1303),
.Y(n_1406)
);

BUFx4f_ASAP7_75t_L g1407 ( 
.A(n_1242),
.Y(n_1407)
);

CKINVDCx6p67_ASAP7_75t_R g1408 ( 
.A(n_1268),
.Y(n_1408)
);

BUFx12f_ASAP7_75t_L g1409 ( 
.A(n_1230),
.Y(n_1409)
);

BUFx2_ASAP7_75t_L g1410 ( 
.A(n_1240),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1232),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1253),
.Y(n_1412)
);

AOI22xp33_ASAP7_75t_SL g1413 ( 
.A1(n_1220),
.A2(n_1209),
.B1(n_1215),
.B2(n_1289),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1202),
.Y(n_1414)
);

AOI22xp33_ASAP7_75t_SL g1415 ( 
.A1(n_1220),
.A2(n_1328),
.B1(n_1326),
.B2(n_1279),
.Y(n_1415)
);

OAI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1200),
.A2(n_1345),
.B1(n_1257),
.B2(n_1218),
.Y(n_1416)
);

OAI21xp33_ASAP7_75t_L g1417 ( 
.A1(n_1197),
.A2(n_1231),
.B(n_1246),
.Y(n_1417)
);

AOI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1271),
.A2(n_1311),
.B1(n_1339),
.B2(n_1202),
.Y(n_1418)
);

CKINVDCx20_ASAP7_75t_R g1419 ( 
.A(n_1275),
.Y(n_1419)
);

BUFx10_ASAP7_75t_L g1420 ( 
.A(n_1281),
.Y(n_1420)
);

OAI21xp33_ASAP7_75t_L g1421 ( 
.A1(n_1212),
.A2(n_1249),
.B(n_1239),
.Y(n_1421)
);

CKINVDCx11_ASAP7_75t_R g1422 ( 
.A(n_1311),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1272),
.A2(n_1337),
.B1(n_1274),
.B2(n_1292),
.Y(n_1423)
);

BUFx10_ASAP7_75t_L g1424 ( 
.A(n_1216),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_SL g1425 ( 
.A1(n_1292),
.A2(n_1204),
.B1(n_1322),
.B2(n_1327),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_1263),
.Y(n_1426)
);

CKINVDCx5p33_ASAP7_75t_R g1427 ( 
.A(n_1247),
.Y(n_1427)
);

INVxp67_ASAP7_75t_SL g1428 ( 
.A(n_1266),
.Y(n_1428)
);

INVx1_ASAP7_75t_SL g1429 ( 
.A(n_1270),
.Y(n_1429)
);

INVx6_ASAP7_75t_L g1430 ( 
.A(n_1337),
.Y(n_1430)
);

INVx8_ASAP7_75t_L g1431 ( 
.A(n_1329),
.Y(n_1431)
);

AOI22xp33_ASAP7_75t_L g1432 ( 
.A1(n_1239),
.A2(n_1255),
.B1(n_1211),
.B2(n_1262),
.Y(n_1432)
);

INVxp67_ASAP7_75t_SL g1433 ( 
.A(n_1322),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1199),
.B(n_1349),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1199),
.B(n_1349),
.Y(n_1435)
);

OAI22xp33_ASAP7_75t_L g1436 ( 
.A1(n_1292),
.A2(n_1265),
.B1(n_1204),
.B2(n_1327),
.Y(n_1436)
);

AOI22xp33_ASAP7_75t_L g1437 ( 
.A1(n_1204),
.A2(n_1226),
.B1(n_1199),
.B2(n_1335),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1288),
.B(n_1349),
.Y(n_1438)
);

AOI22xp33_ASAP7_75t_L g1439 ( 
.A1(n_1247),
.A2(n_1290),
.B1(n_1287),
.B2(n_1217),
.Y(n_1439)
);

BUFx2_ASAP7_75t_L g1440 ( 
.A(n_1287),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1290),
.Y(n_1441)
);

CKINVDCx11_ASAP7_75t_R g1442 ( 
.A(n_1290),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1267),
.A2(n_1237),
.B1(n_1243),
.B2(n_1224),
.Y(n_1443)
);

CKINVDCx11_ASAP7_75t_R g1444 ( 
.A(n_1288),
.Y(n_1444)
);

INVx6_ASAP7_75t_L g1445 ( 
.A(n_1256),
.Y(n_1445)
);

AOI22xp33_ASAP7_75t_L g1446 ( 
.A1(n_1314),
.A2(n_1320),
.B1(n_1224),
.B2(n_1205),
.Y(n_1446)
);

AOI22xp33_ASAP7_75t_L g1447 ( 
.A1(n_1196),
.A2(n_1347),
.B1(n_1285),
.B2(n_1298),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_L g1448 ( 
.A1(n_1309),
.A2(n_673),
.B1(n_1186),
.B2(n_1175),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1321),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1330),
.A2(n_673),
.B1(n_1280),
.B2(n_1011),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_1203),
.Y(n_1453)
);

BUFx6f_ASAP7_75t_L g1454 ( 
.A(n_1291),
.Y(n_1454)
);

CKINVDCx11_ASAP7_75t_R g1455 ( 
.A(n_1203),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1291),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1259),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1458)
);

OAI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1324),
.A2(n_673),
.B1(n_1186),
.B2(n_1175),
.Y(n_1459)
);

BUFx4f_ASAP7_75t_SL g1460 ( 
.A(n_1203),
.Y(n_1460)
);

INVx5_ASAP7_75t_L g1461 ( 
.A(n_1331),
.Y(n_1461)
);

INVx6_ASAP7_75t_L g1462 ( 
.A(n_1277),
.Y(n_1462)
);

INVx8_ASAP7_75t_L g1463 ( 
.A(n_1331),
.Y(n_1463)
);

CKINVDCx11_ASAP7_75t_R g1464 ( 
.A(n_1203),
.Y(n_1464)
);

AOI22xp5_ASAP7_75t_L g1465 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1033),
.Y(n_1465)
);

AOI22xp33_ASAP7_75t_L g1466 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1466)
);

BUFx8_ASAP7_75t_L g1467 ( 
.A(n_1273),
.Y(n_1467)
);

AOI22xp33_ASAP7_75t_L g1468 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1468)
);

BUFx4f_ASAP7_75t_SL g1469 ( 
.A(n_1203),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1300),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1471)
);

INVx5_ASAP7_75t_L g1472 ( 
.A(n_1331),
.Y(n_1472)
);

OAI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1280),
.A2(n_673),
.B1(n_1324),
.B2(n_1195),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1259),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_SL g1475 ( 
.A1(n_1280),
.A2(n_673),
.B1(n_1011),
.B2(n_1033),
.Y(n_1475)
);

OAI22x1_ASAP7_75t_L g1476 ( 
.A1(n_1261),
.A2(n_1175),
.B1(n_1186),
.B2(n_1294),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1259),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1323),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1259),
.Y(n_1479)
);

AOI22xp33_ASAP7_75t_L g1480 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1096),
.B2(n_1175),
.Y(n_1480)
);

INVx6_ASAP7_75t_L g1481 ( 
.A(n_1277),
.Y(n_1481)
);

BUFx12f_ASAP7_75t_L g1482 ( 
.A(n_1252),
.Y(n_1482)
);

OAI22xp5_ASAP7_75t_L g1483 ( 
.A1(n_1324),
.A2(n_673),
.B1(n_1186),
.B2(n_1175),
.Y(n_1483)
);

AOI22xp33_ASAP7_75t_L g1484 ( 
.A1(n_1304),
.A2(n_673),
.B1(n_1280),
.B2(n_1310),
.Y(n_1484)
);

AND2x4_ASAP7_75t_L g1485 ( 
.A(n_1434),
.B(n_1435),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_1373),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1463),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_SL g1488 ( 
.A(n_1356),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1405),
.Y(n_1489)
);

OA21x2_ASAP7_75t_L g1490 ( 
.A1(n_1421),
.A2(n_1446),
.B(n_1389),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1426),
.Y(n_1491)
);

BUFx12f_ASAP7_75t_L g1492 ( 
.A(n_1455),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1447),
.A2(n_1449),
.B(n_1432),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1444),
.B(n_1434),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1475),
.A2(n_1400),
.B1(n_1465),
.B2(n_1480),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1435),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1410),
.Y(n_1497)
);

BUFx2_ASAP7_75t_L g1498 ( 
.A(n_1428),
.Y(n_1498)
);

OAI21x1_ASAP7_75t_L g1499 ( 
.A1(n_1447),
.A2(n_1449),
.B(n_1394),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1438),
.Y(n_1500)
);

OR2x6_ASAP7_75t_L g1501 ( 
.A(n_1417),
.B(n_1438),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1445),
.Y(n_1502)
);

OAI22xp5_ASAP7_75t_SL g1503 ( 
.A1(n_1475),
.A2(n_1452),
.B1(n_1451),
.B2(n_1458),
.Y(n_1503)
);

INVx1_ASAP7_75t_SL g1504 ( 
.A(n_1429),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1433),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1464),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1361),
.B(n_1362),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1433),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1354),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1436),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1355),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1436),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_1478),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1437),
.B(n_1372),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1362),
.B(n_1376),
.Y(n_1515)
);

INVx2_ASAP7_75t_L g1516 ( 
.A(n_1363),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1365),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1367),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1374),
.Y(n_1519)
);

AO31x2_ASAP7_75t_L g1520 ( 
.A1(n_1443),
.A2(n_1358),
.A3(n_1448),
.B(n_1483),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1379),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1390),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1391),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1437),
.B(n_1446),
.Y(n_1524)
);

INVx3_ASAP7_75t_L g1525 ( 
.A(n_1378),
.Y(n_1525)
);

OAI21x1_ASAP7_75t_L g1526 ( 
.A1(n_1384),
.A2(n_1439),
.B(n_1383),
.Y(n_1526)
);

OAI21x1_ASAP7_75t_L g1527 ( 
.A1(n_1416),
.A2(n_1393),
.B(n_1404),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_1453),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1459),
.A2(n_1468),
.B(n_1471),
.Y(n_1529)
);

OAI21x1_ASAP7_75t_L g1530 ( 
.A1(n_1399),
.A2(n_1411),
.B(n_1412),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1378),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1425),
.Y(n_1532)
);

OR2x6_ASAP7_75t_L g1533 ( 
.A(n_1463),
.B(n_1385),
.Y(n_1533)
);

OR2x2_ASAP7_75t_L g1534 ( 
.A(n_1423),
.B(n_1368),
.Y(n_1534)
);

OR2x2_ASAP7_75t_SL g1535 ( 
.A(n_1360),
.B(n_1370),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1466),
.A2(n_1484),
.B(n_1473),
.Y(n_1536)
);

CKINVDCx5p33_ASAP7_75t_R g1537 ( 
.A(n_1380),
.Y(n_1537)
);

INVx2_ASAP7_75t_L g1538 ( 
.A(n_1378),
.Y(n_1538)
);

CKINVDCx5p33_ASAP7_75t_R g1539 ( 
.A(n_1380),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1423),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1368),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1415),
.Y(n_1542)
);

BUFx2_ASAP7_75t_L g1543 ( 
.A(n_1428),
.Y(n_1543)
);

OAI21xp5_ASAP7_75t_L g1544 ( 
.A1(n_1450),
.A2(n_1484),
.B(n_1473),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1359),
.B(n_1457),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1474),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1415),
.Y(n_1547)
);

INVx2_ASAP7_75t_L g1548 ( 
.A(n_1477),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1395),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1479),
.Y(n_1550)
);

OR2x6_ASAP7_75t_L g1551 ( 
.A(n_1463),
.B(n_1431),
.Y(n_1551)
);

CKINVDCx11_ASAP7_75t_R g1552 ( 
.A(n_1482),
.Y(n_1552)
);

AND2x2_ASAP7_75t_L g1553 ( 
.A(n_1395),
.B(n_1396),
.Y(n_1553)
);

INVx4_ASAP7_75t_L g1554 ( 
.A(n_1461),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1369),
.Y(n_1555)
);

NAND4xp25_ASAP7_75t_L g1556 ( 
.A(n_1387),
.B(n_1450),
.C(n_1396),
.D(n_1413),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1413),
.B(n_1476),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1398),
.Y(n_1558)
);

OR2x6_ASAP7_75t_L g1559 ( 
.A(n_1392),
.B(n_1431),
.Y(n_1559)
);

OAI21x1_ASAP7_75t_L g1560 ( 
.A1(n_1418),
.A2(n_1377),
.B(n_1470),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1398),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_L g1562 ( 
.A(n_1366),
.B(n_1408),
.Y(n_1562)
);

HB1xp67_ASAP7_75t_SL g1563 ( 
.A(n_1356),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1375),
.A2(n_1470),
.B(n_1431),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_1472),
.Y(n_1565)
);

AO21x2_ASAP7_75t_L g1566 ( 
.A1(n_1366),
.A2(n_1402),
.B(n_1371),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_1357),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1364),
.Y(n_1568)
);

OA21x2_ASAP7_75t_L g1569 ( 
.A1(n_1440),
.A2(n_1441),
.B(n_1427),
.Y(n_1569)
);

OAI21x1_ASAP7_75t_L g1570 ( 
.A1(n_1375),
.A2(n_1364),
.B(n_1430),
.Y(n_1570)
);

AOI22xp33_ASAP7_75t_L g1571 ( 
.A1(n_1422),
.A2(n_1414),
.B1(n_1382),
.B2(n_1388),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_L g1572 ( 
.A(n_1403),
.B(n_1419),
.Y(n_1572)
);

CKINVDCx20_ASAP7_75t_R g1573 ( 
.A(n_1460),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_L g1574 ( 
.A(n_1407),
.B(n_1420),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1424),
.Y(n_1575)
);

OAI22xp5_ASAP7_75t_L g1576 ( 
.A1(n_1495),
.A2(n_1360),
.B1(n_1462),
.B2(n_1370),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1511),
.Y(n_1577)
);

A2O1A1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1536),
.A2(n_1407),
.B(n_1381),
.C(n_1456),
.Y(n_1578)
);

A2O1A1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1544),
.A2(n_1456),
.B(n_1454),
.C(n_1386),
.Y(n_1579)
);

OAI21xp5_ASAP7_75t_L g1580 ( 
.A1(n_1529),
.A2(n_1544),
.B(n_1515),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1509),
.B(n_1397),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1497),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1534),
.B(n_1397),
.Y(n_1583)
);

A2O1A1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1529),
.A2(n_1456),
.B(n_1386),
.C(n_1454),
.Y(n_1584)
);

NOR2x1p5_ASAP7_75t_L g1585 ( 
.A(n_1492),
.B(n_1401),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1532),
.B(n_1442),
.Y(n_1586)
);

OR2x6_ASAP7_75t_L g1587 ( 
.A(n_1501),
.B(n_1360),
.Y(n_1587)
);

OA21x2_ASAP7_75t_L g1588 ( 
.A1(n_1493),
.A2(n_1406),
.B(n_1409),
.Y(n_1588)
);

INVx3_ASAP7_75t_L g1589 ( 
.A(n_1564),
.Y(n_1589)
);

OAI21xp5_ASAP7_75t_SL g1590 ( 
.A1(n_1553),
.A2(n_1370),
.B(n_1462),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1524),
.B(n_1514),
.Y(n_1591)
);

AND2x2_ASAP7_75t_L g1592 ( 
.A(n_1524),
.B(n_1462),
.Y(n_1592)
);

NOR2x1_ASAP7_75t_SL g1593 ( 
.A(n_1501),
.B(n_1481),
.Y(n_1593)
);

A2O1A1Ixp33_ASAP7_75t_L g1594 ( 
.A1(n_1553),
.A2(n_1481),
.B(n_1467),
.C(n_1469),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1514),
.B(n_1481),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1494),
.B(n_1467),
.Y(n_1596)
);

NOR2xp33_ASAP7_75t_R g1597 ( 
.A(n_1537),
.B(n_1460),
.Y(n_1597)
);

NOR4xp25_ASAP7_75t_SL g1598 ( 
.A(n_1498),
.B(n_1469),
.C(n_1543),
.D(n_1539),
.Y(n_1598)
);

BUFx2_ASAP7_75t_L g1599 ( 
.A(n_1569),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1545),
.B(n_1546),
.Y(n_1600)
);

O2A1O1Ixp33_ASAP7_75t_SL g1601 ( 
.A1(n_1562),
.A2(n_1507),
.B(n_1542),
.C(n_1547),
.Y(n_1601)
);

OAI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1556),
.A2(n_1526),
.B(n_1541),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1556),
.A2(n_1549),
.B(n_1557),
.C(n_1541),
.Y(n_1603)
);

NAND2x1p5_ASAP7_75t_L g1604 ( 
.A(n_1498),
.B(n_1543),
.Y(n_1604)
);

AND2x4_ASAP7_75t_L g1605 ( 
.A(n_1531),
.B(n_1538),
.Y(n_1605)
);

OAI21xp5_ASAP7_75t_L g1606 ( 
.A1(n_1526),
.A2(n_1558),
.B(n_1561),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1538),
.B(n_1502),
.Y(n_1607)
);

OAI211xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1504),
.A2(n_1558),
.B(n_1561),
.C(n_1571),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1528),
.B(n_1572),
.Y(n_1609)
);

A2O1A1Ixp33_ASAP7_75t_L g1610 ( 
.A1(n_1540),
.A2(n_1542),
.B(n_1503),
.C(n_1510),
.Y(n_1610)
);

AND2x2_ASAP7_75t_L g1611 ( 
.A(n_1566),
.B(n_1555),
.Y(n_1611)
);

A2O1A1Ixp33_ASAP7_75t_L g1612 ( 
.A1(n_1540),
.A2(n_1503),
.B(n_1512),
.C(n_1527),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1511),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1564),
.Y(n_1614)
);

OAI21xp5_ASAP7_75t_L g1615 ( 
.A1(n_1560),
.A2(n_1499),
.B(n_1530),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1566),
.B(n_1511),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1485),
.B(n_1501),
.Y(n_1617)
);

OAI21xp5_ASAP7_75t_L g1618 ( 
.A1(n_1560),
.A2(n_1530),
.B(n_1570),
.Y(n_1618)
);

OR2x2_ASAP7_75t_L g1619 ( 
.A(n_1516),
.B(n_1521),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1569),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1538),
.B(n_1502),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_1492),
.Y(n_1622)
);

OR2x2_ASAP7_75t_L g1623 ( 
.A(n_1516),
.B(n_1521),
.Y(n_1623)
);

OR2x2_ASAP7_75t_L g1624 ( 
.A(n_1516),
.B(n_1521),
.Y(n_1624)
);

A2O1A1Ixp33_ASAP7_75t_L g1625 ( 
.A1(n_1548),
.A2(n_1550),
.B(n_1496),
.C(n_1500),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1485),
.B(n_1501),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1485),
.B(n_1517),
.Y(n_1627)
);

AOI22xp5_ASAP7_75t_L g1628 ( 
.A1(n_1566),
.A2(n_1573),
.B1(n_1574),
.B2(n_1506),
.Y(n_1628)
);

AOI22xp5_ASAP7_75t_L g1629 ( 
.A1(n_1492),
.A2(n_1506),
.B1(n_1559),
.B2(n_1533),
.Y(n_1629)
);

OA21x2_ASAP7_75t_L g1630 ( 
.A1(n_1491),
.A2(n_1489),
.B(n_1505),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1518),
.B(n_1519),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1491),
.A2(n_1489),
.B(n_1508),
.Y(n_1632)
);

INVx2_ASAP7_75t_L g1633 ( 
.A(n_1630),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1627),
.B(n_1490),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1600),
.B(n_1496),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1620),
.Y(n_1636)
);

NAND2x1_ASAP7_75t_L g1637 ( 
.A(n_1587),
.B(n_1554),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1580),
.A2(n_1506),
.B1(n_1550),
.B2(n_1552),
.Y(n_1638)
);

INVxp33_ASAP7_75t_L g1639 ( 
.A(n_1609),
.Y(n_1639)
);

HB1xp67_ASAP7_75t_L g1640 ( 
.A(n_1632),
.Y(n_1640)
);

AOI222xp33_ASAP7_75t_L g1641 ( 
.A1(n_1610),
.A2(n_1486),
.B1(n_1519),
.B2(n_1522),
.C1(n_1523),
.C2(n_1488),
.Y(n_1641)
);

BUFx2_ASAP7_75t_L g1642 ( 
.A(n_1618),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1617),
.B(n_1505),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1626),
.B(n_1508),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1616),
.B(n_1520),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1577),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1589),
.B(n_1525),
.Y(n_1647)
);

AND2x4_ASAP7_75t_L g1648 ( 
.A(n_1589),
.B(n_1614),
.Y(n_1648)
);

HB1xp67_ASAP7_75t_L g1649 ( 
.A(n_1599),
.Y(n_1649)
);

BUFx12f_ASAP7_75t_L g1650 ( 
.A(n_1622),
.Y(n_1650)
);

BUFx2_ASAP7_75t_L g1651 ( 
.A(n_1615),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1613),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1605),
.Y(n_1653)
);

AOI22xp5_ASAP7_75t_L g1654 ( 
.A1(n_1610),
.A2(n_1559),
.B1(n_1533),
.B2(n_1551),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1631),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1607),
.B(n_1621),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1606),
.B(n_1591),
.Y(n_1657)
);

INVx2_ASAP7_75t_SL g1658 ( 
.A(n_1648),
.Y(n_1658)
);

OAI221xp5_ASAP7_75t_L g1659 ( 
.A1(n_1638),
.A2(n_1578),
.B1(n_1603),
.B2(n_1608),
.C(n_1602),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1653),
.B(n_1611),
.Y(n_1660)
);

NOR3xp33_ASAP7_75t_L g1661 ( 
.A(n_1651),
.B(n_1576),
.C(n_1578),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1652),
.Y(n_1662)
);

NOR3xp33_ASAP7_75t_L g1663 ( 
.A(n_1651),
.B(n_1603),
.C(n_1584),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1645),
.B(n_1591),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1652),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1652),
.Y(n_1666)
);

INVx2_ASAP7_75t_L g1667 ( 
.A(n_1633),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1645),
.B(n_1619),
.Y(n_1668)
);

AND2x4_ASAP7_75t_L g1669 ( 
.A(n_1647),
.B(n_1593),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1656),
.B(n_1628),
.Y(n_1670)
);

AND2x2_ASAP7_75t_L g1671 ( 
.A(n_1656),
.B(n_1592),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1653),
.B(n_1592),
.Y(n_1672)
);

AOI221xp5_ASAP7_75t_L g1673 ( 
.A1(n_1657),
.A2(n_1601),
.B1(n_1612),
.B2(n_1582),
.C(n_1579),
.Y(n_1673)
);

AND2x4_ASAP7_75t_L g1674 ( 
.A(n_1647),
.B(n_1648),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1645),
.B(n_1623),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1646),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1646),
.Y(n_1677)
);

BUFx6f_ASAP7_75t_L g1678 ( 
.A(n_1650),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1633),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1657),
.B(n_1655),
.Y(n_1680)
);

OR2x2_ASAP7_75t_L g1681 ( 
.A(n_1657),
.B(n_1624),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1639),
.B(n_1622),
.Y(n_1682)
);

OAI22xp5_ASAP7_75t_L g1683 ( 
.A1(n_1638),
.A2(n_1579),
.B1(n_1584),
.B2(n_1612),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1635),
.B(n_1625),
.Y(n_1684)
);

HB1xp67_ASAP7_75t_L g1685 ( 
.A(n_1636),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1633),
.Y(n_1686)
);

INVx2_ASAP7_75t_SL g1687 ( 
.A(n_1648),
.Y(n_1687)
);

NOR3xp33_ASAP7_75t_SL g1688 ( 
.A(n_1635),
.B(n_1594),
.C(n_1590),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1633),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1634),
.B(n_1588),
.Y(n_1690)
);

NOR3xp33_ASAP7_75t_L g1691 ( 
.A(n_1651),
.B(n_1601),
.C(n_1594),
.Y(n_1691)
);

INVx3_ASAP7_75t_L g1692 ( 
.A(n_1674),
.Y(n_1692)
);

NAND2x1p5_ASAP7_75t_L g1693 ( 
.A(n_1678),
.B(n_1637),
.Y(n_1693)
);

NOR2xp33_ASAP7_75t_L g1694 ( 
.A(n_1682),
.B(n_1639),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1678),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1662),
.Y(n_1697)
);

NAND3xp33_ASAP7_75t_SL g1698 ( 
.A(n_1691),
.B(n_1641),
.C(n_1651),
.Y(n_1698)
);

NOR2xp67_ASAP7_75t_L g1699 ( 
.A(n_1658),
.B(n_1640),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1662),
.Y(n_1700)
);

OR2x2_ASAP7_75t_L g1701 ( 
.A(n_1680),
.B(n_1642),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1665),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1665),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1666),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1666),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1685),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1684),
.B(n_1643),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1685),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1678),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1664),
.B(n_1643),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1676),
.Y(n_1713)
);

AND2x4_ASAP7_75t_L g1714 ( 
.A(n_1669),
.B(n_1648),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1674),
.B(n_1642),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1676),
.Y(n_1716)
);

OR2x2_ASAP7_75t_L g1717 ( 
.A(n_1680),
.B(n_1655),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1672),
.B(n_1655),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1664),
.B(n_1643),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1667),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1668),
.B(n_1675),
.Y(n_1721)
);

NAND2xp5_ASAP7_75t_L g1722 ( 
.A(n_1681),
.B(n_1644),
.Y(n_1722)
);

OR2x2_ASAP7_75t_L g1723 ( 
.A(n_1668),
.B(n_1649),
.Y(n_1723)
);

INVx2_ASAP7_75t_L g1724 ( 
.A(n_1667),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1669),
.B(n_1648),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1677),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1677),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1695),
.B(n_1663),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1709),
.B(n_1663),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1696),
.B(n_1690),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1724),
.Y(n_1732)
);

NAND2xp33_ASAP7_75t_SL g1733 ( 
.A(n_1696),
.B(n_1688),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1692),
.B(n_1690),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1697),
.Y(n_1735)
);

NAND3xp33_ASAP7_75t_L g1736 ( 
.A(n_1694),
.B(n_1691),
.C(n_1661),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1706),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1711),
.B(n_1673),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1692),
.B(n_1690),
.Y(n_1739)
);

OR2x2_ASAP7_75t_L g1740 ( 
.A(n_1721),
.B(n_1675),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1724),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1721),
.B(n_1681),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1700),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1711),
.B(n_1673),
.Y(n_1744)
);

AOI32xp33_ASAP7_75t_L g1745 ( 
.A1(n_1698),
.A2(n_1661),
.A3(n_1659),
.B1(n_1683),
.B2(n_1670),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1700),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1702),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1702),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1724),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1703),
.Y(n_1750)
);

NOR2xp33_ASAP7_75t_L g1751 ( 
.A(n_1711),
.B(n_1650),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1692),
.B(n_1669),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1703),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1704),
.Y(n_1754)
);

AND2x4_ASAP7_75t_L g1755 ( 
.A(n_1699),
.B(n_1669),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1712),
.B(n_1670),
.Y(n_1756)
);

OR2x2_ASAP7_75t_L g1757 ( 
.A(n_1701),
.B(n_1649),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1692),
.B(n_1707),
.Y(n_1758)
);

AND2x2_ASAP7_75t_L g1759 ( 
.A(n_1707),
.B(n_1658),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1719),
.B(n_1671),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1704),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1708),
.B(n_1658),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1701),
.B(n_1723),
.Y(n_1763)
);

INVx3_ASAP7_75t_L g1764 ( 
.A(n_1714),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1705),
.Y(n_1765)
);

OR2x2_ASAP7_75t_L g1766 ( 
.A(n_1723),
.B(n_1649),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1693),
.A2(n_1659),
.B1(n_1654),
.B2(n_1688),
.Y(n_1767)
);

INVxp67_ASAP7_75t_L g1768 ( 
.A(n_1706),
.Y(n_1768)
);

OR2x2_ASAP7_75t_L g1769 ( 
.A(n_1710),
.B(n_1717),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1699),
.B(n_1678),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1735),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_SL g1772 ( 
.A(n_1745),
.B(n_1678),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1738),
.B(n_1744),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1734),
.Y(n_1774)
);

OR2x2_ASAP7_75t_L g1775 ( 
.A(n_1763),
.B(n_1710),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1770),
.B(n_1708),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1763),
.B(n_1742),
.Y(n_1777)
);

NAND2xp5_ASAP7_75t_L g1778 ( 
.A(n_1728),
.B(n_1671),
.Y(n_1778)
);

NOR2xp33_ASAP7_75t_L g1779 ( 
.A(n_1736),
.B(n_1650),
.Y(n_1779)
);

NOR2xp33_ASAP7_75t_L g1780 ( 
.A(n_1729),
.B(n_1650),
.Y(n_1780)
);

AND2x2_ASAP7_75t_L g1781 ( 
.A(n_1770),
.B(n_1715),
.Y(n_1781)
);

NOR2xp33_ASAP7_75t_L g1782 ( 
.A(n_1751),
.B(n_1650),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1768),
.B(n_1660),
.Y(n_1783)
);

INVxp67_ASAP7_75t_SL g1784 ( 
.A(n_1767),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1733),
.B(n_1660),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1733),
.B(n_1756),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1770),
.B(n_1715),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1735),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1737),
.B(n_1641),
.C(n_1683),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1764),
.B(n_1714),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1743),
.Y(n_1791)
);

AND3x2_ASAP7_75t_L g1792 ( 
.A(n_1730),
.B(n_1596),
.C(n_1595),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1743),
.Y(n_1793)
);

NOR2x1_ASAP7_75t_L g1794 ( 
.A(n_1755),
.B(n_1585),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1742),
.B(n_1660),
.Y(n_1795)
);

INVxp67_ASAP7_75t_L g1796 ( 
.A(n_1730),
.Y(n_1796)
);

NAND2x1p5_ASAP7_75t_L g1797 ( 
.A(n_1755),
.B(n_1678),
.Y(n_1797)
);

INVxp67_ASAP7_75t_L g1798 ( 
.A(n_1769),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1740),
.B(n_1718),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1746),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1732),
.Y(n_1801)
);

NAND2x1_ASAP7_75t_L g1802 ( 
.A(n_1755),
.B(n_1714),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1732),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1740),
.B(n_1718),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1764),
.B(n_1714),
.Y(n_1805)
);

AND2x2_ASAP7_75t_L g1806 ( 
.A(n_1764),
.B(n_1725),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1746),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1771),
.Y(n_1808)
);

AND2x4_ASAP7_75t_L g1809 ( 
.A(n_1794),
.B(n_1758),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1771),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1788),
.Y(n_1811)
);

OAI22xp5_ASAP7_75t_L g1812 ( 
.A1(n_1789),
.A2(n_1654),
.B1(n_1693),
.B2(n_1629),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1772),
.A2(n_1641),
.B(n_1693),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1788),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1773),
.B(n_1760),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1789),
.A2(n_1747),
.B(n_1731),
.Y(n_1816)
);

OAI22xp33_ASAP7_75t_L g1817 ( 
.A1(n_1784),
.A2(n_1654),
.B1(n_1583),
.B2(n_1604),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1769),
.C(n_1754),
.Y(n_1818)
);

AO22x1_ASAP7_75t_L g1819 ( 
.A1(n_1794),
.A2(n_1758),
.B1(n_1765),
.B2(n_1761),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1779),
.A2(n_1750),
.B(n_1748),
.Y(n_1820)
);

OAI21xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1785),
.A2(n_1752),
.B(n_1759),
.Y(n_1821)
);

AOI211x1_ASAP7_75t_SL g1822 ( 
.A1(n_1774),
.A2(n_1783),
.B(n_1778),
.C(n_1803),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1791),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1791),
.Y(n_1824)
);

HB1xp67_ASAP7_75t_L g1825 ( 
.A(n_1796),
.Y(n_1825)
);

AOI222xp33_ASAP7_75t_L g1826 ( 
.A1(n_1798),
.A2(n_1595),
.B1(n_1586),
.B2(n_1739),
.C1(n_1734),
.C2(n_1754),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1776),
.B(n_1759),
.Y(n_1827)
);

OAI22xp5_ASAP7_75t_L g1828 ( 
.A1(n_1802),
.A2(n_1780),
.B1(n_1797),
.B2(n_1777),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1777),
.B(n_1766),
.Y(n_1829)
);

NOR2xp33_ASAP7_75t_L g1830 ( 
.A(n_1782),
.B(n_1513),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1792),
.B(n_1766),
.Y(n_1831)
);

AND2x2_ASAP7_75t_SL g1832 ( 
.A(n_1776),
.B(n_1563),
.Y(n_1832)
);

NAND2xp33_ASAP7_75t_L g1833 ( 
.A(n_1797),
.B(n_1597),
.Y(n_1833)
);

OAI21xp5_ASAP7_75t_L g1834 ( 
.A1(n_1816),
.A2(n_1797),
.B(n_1775),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1825),
.B(n_1822),
.Y(n_1835)
);

OAI211xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1813),
.A2(n_1807),
.B(n_1800),
.C(n_1793),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1825),
.Y(n_1837)
);

AND2x2_ASAP7_75t_L g1838 ( 
.A(n_1832),
.B(n_1781),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1808),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1832),
.A2(n_1818),
.B1(n_1809),
.B2(n_1812),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1820),
.B(n_1781),
.Y(n_1841)
);

OAI22xp5_ASAP7_75t_L g1842 ( 
.A1(n_1809),
.A2(n_1831),
.B1(n_1828),
.B2(n_1802),
.Y(n_1842)
);

AOI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1833),
.A2(n_1787),
.B1(n_1774),
.B2(n_1805),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1810),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_L g1845 ( 
.A(n_1830),
.B(n_1787),
.Y(n_1845)
);

AOI22xp5_ASAP7_75t_L g1846 ( 
.A1(n_1821),
.A2(n_1826),
.B1(n_1827),
.B2(n_1817),
.Y(n_1846)
);

A2O1A1Ixp33_ASAP7_75t_L g1847 ( 
.A1(n_1815),
.A2(n_1775),
.B(n_1793),
.C(n_1807),
.Y(n_1847)
);

OAI22xp5_ASAP7_75t_L g1848 ( 
.A1(n_1829),
.A2(n_1804),
.B1(n_1799),
.B2(n_1795),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1811),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1814),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1817),
.A2(n_1830),
.B(n_1824),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1819),
.B(n_1800),
.Y(n_1852)
);

AND2x2_ASAP7_75t_L g1853 ( 
.A(n_1823),
.B(n_1790),
.Y(n_1853)
);

OAI211xp5_ASAP7_75t_L g1854 ( 
.A1(n_1835),
.A2(n_1803),
.B(n_1801),
.C(n_1806),
.Y(n_1854)
);

AOI22xp5_ASAP7_75t_L g1855 ( 
.A1(n_1840),
.A2(n_1806),
.B1(n_1805),
.B2(n_1790),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1838),
.B(n_1762),
.Y(n_1856)
);

INVxp67_ASAP7_75t_SL g1857 ( 
.A(n_1852),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1837),
.Y(n_1858)
);

OAI21xp5_ASAP7_75t_SL g1859 ( 
.A1(n_1834),
.A2(n_1586),
.B(n_1752),
.Y(n_1859)
);

AO22x1_ASAP7_75t_L g1860 ( 
.A1(n_1842),
.A2(n_1803),
.B1(n_1801),
.B2(n_1753),
.Y(n_1860)
);

XNOR2xp5_ASAP7_75t_L g1861 ( 
.A(n_1843),
.B(n_1535),
.Y(n_1861)
);

XNOR2x2_ASAP7_75t_SL g1862 ( 
.A(n_1846),
.B(n_1757),
.Y(n_1862)
);

INVx1_ASAP7_75t_L g1863 ( 
.A(n_1853),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1839),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1844),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_SL g1866 ( 
.A(n_1855),
.B(n_1845),
.Y(n_1866)
);

INVx1_ASAP7_75t_L g1867 ( 
.A(n_1863),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1858),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1856),
.B(n_1845),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1857),
.B(n_1841),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1864),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_L g1872 ( 
.A(n_1865),
.Y(n_1872)
);

INVxp33_ASAP7_75t_L g1873 ( 
.A(n_1861),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1862),
.A2(n_1847),
.B(n_1836),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_SL g1875 ( 
.A(n_1857),
.B(n_1851),
.Y(n_1875)
);

NAND3xp33_ASAP7_75t_L g1876 ( 
.A(n_1860),
.B(n_1836),
.C(n_1847),
.Y(n_1876)
);

OAI211xp5_ASAP7_75t_SL g1877 ( 
.A1(n_1875),
.A2(n_1859),
.B(n_1862),
.C(n_1854),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1872),
.Y(n_1878)
);

AOI211xp5_ASAP7_75t_SL g1879 ( 
.A1(n_1874),
.A2(n_1850),
.B(n_1849),
.C(n_1848),
.Y(n_1879)
);

NOR4xp75_ASAP7_75t_L g1880 ( 
.A(n_1866),
.B(n_1739),
.C(n_1581),
.D(n_1762),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_SL g1881 ( 
.A(n_1876),
.B(n_1801),
.Y(n_1881)
);

AOI31xp33_ASAP7_75t_L g1882 ( 
.A1(n_1873),
.A2(n_1757),
.A3(n_1535),
.B(n_1753),
.Y(n_1882)
);

O2A1O1Ixp33_ASAP7_75t_L g1883 ( 
.A1(n_1877),
.A2(n_1870),
.B(n_1868),
.C(n_1871),
.Y(n_1883)
);

NOR4xp75_ASAP7_75t_SL g1884 ( 
.A(n_1879),
.B(n_1869),
.C(n_1872),
.D(n_1867),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1878),
.Y(n_1885)
);

OAI22xp5_ASAP7_75t_SL g1886 ( 
.A1(n_1881),
.A2(n_1872),
.B1(n_1551),
.B2(n_1533),
.Y(n_1886)
);

NAND3xp33_ASAP7_75t_SL g1887 ( 
.A(n_1880),
.B(n_1598),
.C(n_1741),
.Y(n_1887)
);

AOI211xp5_ASAP7_75t_L g1888 ( 
.A1(n_1882),
.A2(n_1749),
.B(n_1741),
.C(n_1575),
.Y(n_1888)
);

OAI22x1_ASAP7_75t_L g1889 ( 
.A1(n_1885),
.A2(n_1749),
.B1(n_1725),
.B2(n_1687),
.Y(n_1889)
);

NAND4xp75_ASAP7_75t_L g1890 ( 
.A(n_1884),
.B(n_1883),
.C(n_1886),
.D(n_1888),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1887),
.Y(n_1891)
);

AND2x2_ASAP7_75t_L g1892 ( 
.A(n_1885),
.B(n_1725),
.Y(n_1892)
);

XOR2x1_ASAP7_75t_L g1893 ( 
.A(n_1885),
.B(n_1725),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1891),
.A2(n_1720),
.B(n_1722),
.Y(n_1894)
);

NOR2x1_ASAP7_75t_L g1895 ( 
.A(n_1890),
.B(n_1720),
.Y(n_1895)
);

AOI22x1_ASAP7_75t_L g1896 ( 
.A1(n_1891),
.A2(n_1554),
.B1(n_1565),
.B2(n_1575),
.Y(n_1896)
);

NOR2x1_ASAP7_75t_L g1897 ( 
.A(n_1895),
.B(n_1892),
.Y(n_1897)
);

OAI22xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1894),
.B1(n_1896),
.B2(n_1893),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1898),
.Y(n_1899)
);

NOR3xp33_ASAP7_75t_L g1900 ( 
.A(n_1898),
.B(n_1889),
.C(n_1487),
.Y(n_1900)
);

OAI22xp5_ASAP7_75t_SL g1901 ( 
.A1(n_1899),
.A2(n_1487),
.B1(n_1551),
.B2(n_1559),
.Y(n_1901)
);

NOR4xp25_ASAP7_75t_L g1902 ( 
.A(n_1900),
.B(n_1705),
.C(n_1726),
.D(n_1727),
.Y(n_1902)
);

OAI21xp5_ASAP7_75t_L g1903 ( 
.A1(n_1902),
.A2(n_1716),
.B(n_1713),
.Y(n_1903)
);

NAND2xp5_ASAP7_75t_L g1904 ( 
.A(n_1901),
.B(n_1713),
.Y(n_1904)
);

NAND2xp5_ASAP7_75t_L g1905 ( 
.A(n_1904),
.B(n_1716),
.Y(n_1905)
);

XNOR2xp5_ASAP7_75t_L g1906 ( 
.A(n_1905),
.B(n_1903),
.Y(n_1906)
);

OAI22xp33_ASAP7_75t_L g1907 ( 
.A1(n_1906),
.A2(n_1727),
.B1(n_1726),
.B2(n_1717),
.Y(n_1907)
);

OAI221xp5_ASAP7_75t_R g1908 ( 
.A1(n_1907),
.A2(n_1687),
.B1(n_1689),
.B2(n_1679),
.C(n_1686),
.Y(n_1908)
);

AOI211xp5_ASAP7_75t_L g1909 ( 
.A1(n_1908),
.A2(n_1487),
.B(n_1567),
.C(n_1568),
.Y(n_1909)
);


endmodule