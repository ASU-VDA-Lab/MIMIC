module real_aes_8967_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_725;
wire n_504;
wire n_119;
wire n_310;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_552;
wire n_402;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g482 ( .A1(n_0), .A2(n_143), .B(n_483), .C(n_486), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_1), .B(n_478), .Y(n_487) );
INVx1_ASAP7_75t_L g432 ( .A(n_2), .Y(n_432) );
INVx1_ASAP7_75t_L g141 ( .A(n_3), .Y(n_141) );
NAND2xp5_ASAP7_75t_SL g551 ( .A(n_4), .B(n_144), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_5), .A2(n_446), .B(n_522), .Y(n_521) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_6), .A2(n_151), .B(n_501), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_7), .A2(n_35), .B1(n_131), .B2(n_179), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_8), .B(n_151), .Y(n_159) );
AND2x6_ASAP7_75t_L g146 ( .A(n_9), .B(n_147), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g494 ( .A1(n_10), .A2(n_146), .B(n_451), .C(n_495), .Y(n_494) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_11), .B(n_36), .Y(n_433) );
INVx1_ASAP7_75t_L g122 ( .A(n_12), .Y(n_122) );
INVx1_ASAP7_75t_L g125 ( .A(n_13), .Y(n_125) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_14), .B(n_127), .Y(n_188) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_15), .B(n_144), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_16), .B(n_118), .Y(n_225) );
AO32x2_ASAP7_75t_L g195 ( .A1(n_17), .A2(n_117), .A3(n_151), .B1(n_170), .B2(n_196), .Y(n_195) );
AOI222xp33_ASAP7_75t_SL g101 ( .A1(n_18), .A2(n_39), .B1(n_102), .B2(n_724), .C1(n_725), .C2(n_727), .Y(n_101) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_19), .B(n_131), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_20), .B(n_118), .Y(n_148) );
AOI22xp33_ASAP7_75t_L g198 ( .A1(n_21), .A2(n_53), .B1(n_131), .B2(n_179), .Y(n_198) );
AOI22xp33_ASAP7_75t_SL g181 ( .A1(n_22), .A2(n_79), .B1(n_127), .B2(n_131), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_23), .B(n_131), .Y(n_211) );
A2O1A1Ixp33_ASAP7_75t_L g468 ( .A1(n_24), .A2(n_170), .B(n_451), .C(n_469), .Y(n_468) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_25), .A2(n_170), .B(n_451), .C(n_504), .Y(n_503) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_26), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_27), .B(n_172), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g479 ( .A1(n_28), .A2(n_446), .B(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_29), .B(n_172), .Y(n_213) );
INVx2_ASAP7_75t_L g129 ( .A(n_30), .Y(n_129) );
A2O1A1Ixp33_ASAP7_75t_L g448 ( .A1(n_31), .A2(n_449), .B(n_453), .C(n_459), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g163 ( .A(n_32), .B(n_131), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_33), .B(n_172), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_34), .B(n_190), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_37), .B(n_467), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g499 ( .A(n_38), .Y(n_499) );
INVx1_ASAP7_75t_L g724 ( .A(n_39), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_40), .B(n_144), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_41), .B(n_446), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g104 ( .A1(n_42), .A2(n_105), .B1(n_106), .B2(n_427), .Y(n_104) );
INVx1_ASAP7_75t_L g427 ( .A(n_42), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g744 ( .A1(n_42), .A2(n_44), .B1(n_427), .B2(n_745), .Y(n_744) );
A2O1A1Ixp33_ASAP7_75t_L g513 ( .A1(n_43), .A2(n_449), .B(n_459), .C(n_514), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g99 ( .A1(n_44), .A2(n_100), .B1(n_731), .B2(n_740), .C1(n_749), .C2(n_755), .Y(n_99) );
CKINVDCx20_ASAP7_75t_R g745 ( .A(n_44), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_45), .B(n_131), .Y(n_154) );
INVx1_ASAP7_75t_L g484 ( .A(n_46), .Y(n_484) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_47), .A2(n_87), .B1(n_179), .B2(n_180), .Y(n_178) );
INVx1_ASAP7_75t_L g515 ( .A(n_48), .Y(n_515) );
NAND2xp5_ASAP7_75t_SL g157 ( .A(n_49), .B(n_131), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g130 ( .A(n_50), .B(n_131), .Y(n_130) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_51), .B(n_446), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_52), .B(n_139), .Y(n_158) );
AOI22xp33_ASAP7_75t_SL g223 ( .A1(n_54), .A2(n_58), .B1(n_127), .B2(n_131), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g474 ( .A(n_55), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g167 ( .A(n_56), .B(n_131), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g187 ( .A(n_57), .B(n_131), .Y(n_187) );
INVx1_ASAP7_75t_L g147 ( .A(n_59), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_60), .B(n_446), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_61), .B(n_478), .Y(n_527) );
A2O1A1Ixp33_ASAP7_75t_L g524 ( .A1(n_62), .A2(n_133), .B(n_139), .C(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_63), .B(n_131), .Y(n_142) );
INVx1_ASAP7_75t_L g121 ( .A(n_64), .Y(n_121) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_65), .Y(n_736) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_66), .B(n_144), .Y(n_457) );
AO32x2_ASAP7_75t_L g176 ( .A1(n_67), .A2(n_151), .A3(n_170), .B1(n_177), .B2(n_182), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_68), .B(n_145), .Y(n_496) );
INVx1_ASAP7_75t_L g166 ( .A(n_69), .Y(n_166) );
INVx1_ASAP7_75t_L g208 ( .A(n_70), .Y(n_208) );
CKINVDCx16_ASAP7_75t_R g481 ( .A(n_71), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_72), .B(n_456), .Y(n_470) );
A2O1A1Ixp33_ASAP7_75t_L g548 ( .A1(n_73), .A2(n_451), .B(n_459), .C(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_SL g209 ( .A(n_74), .B(n_127), .Y(n_209) );
CKINVDCx16_ASAP7_75t_R g523 ( .A(n_75), .Y(n_523) );
INVx1_ASAP7_75t_L g735 ( .A(n_76), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_77), .Y(n_748) );
NAND2xp5_ASAP7_75t_SL g471 ( .A(n_78), .B(n_455), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_80), .B(n_179), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g462 ( .A(n_81), .Y(n_462) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_82), .B(n_127), .Y(n_212) );
INVx2_ASAP7_75t_L g119 ( .A(n_83), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g555 ( .A(n_84), .Y(n_555) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_85), .B(n_169), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_86), .B(n_127), .Y(n_155) );
OR2x2_ASAP7_75t_L g430 ( .A(n_88), .B(n_431), .Y(n_430) );
INVx2_ASAP7_75t_L g437 ( .A(n_88), .Y(n_437) );
OR2x2_ASAP7_75t_L g739 ( .A(n_88), .B(n_730), .Y(n_739) );
AOI22xp33_ASAP7_75t_L g222 ( .A1(n_89), .A2(n_98), .B1(n_127), .B2(n_128), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_90), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g454 ( .A(n_91), .Y(n_454) );
INVxp67_ASAP7_75t_L g526 ( .A(n_92), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_93), .B(n_127), .Y(n_164) );
INVx1_ASAP7_75t_L g492 ( .A(n_94), .Y(n_492) );
INVx1_ASAP7_75t_L g550 ( .A(n_95), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_96), .B(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g517 ( .A(n_97), .B(n_172), .Y(n_517) );
INVxp67_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
OAI22x1_ASAP7_75t_SL g102 ( .A1(n_103), .A2(n_428), .B1(n_434), .B2(n_438), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_104), .Y(n_103) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_104), .A2(n_428), .B1(n_436), .B2(n_726), .Y(n_725) );
OAI22xp5_ASAP7_75t_SL g742 ( .A1(n_105), .A2(n_106), .B1(n_743), .B2(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_393), .Y(n_106) );
NOR3xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_297), .C(n_381), .Y(n_107) );
NAND4xp25_ASAP7_75t_L g108 ( .A(n_109), .B(n_240), .C(n_262), .D(n_278), .Y(n_108) );
AOI221xp5_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_173), .B1(n_199), .B2(n_218), .C(n_226), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_112), .B(n_149), .Y(n_111) );
NAND2xp5_ASAP7_75t_SL g252 ( .A(n_112), .B(n_218), .Y(n_252) );
NAND4xp25_ASAP7_75t_L g292 ( .A(n_112), .B(n_280), .C(n_293), .D(n_295), .Y(n_292) );
INVxp67_ASAP7_75t_L g409 ( .A(n_112), .Y(n_409) );
INVx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g291 ( .A(n_113), .B(n_229), .Y(n_291) );
AND2x2_ASAP7_75t_L g315 ( .A(n_113), .B(n_149), .Y(n_315) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
AND2x2_ASAP7_75t_L g282 ( .A(n_114), .B(n_217), .Y(n_282) );
AND2x2_ASAP7_75t_L g322 ( .A(n_114), .B(n_303), .Y(n_322) );
AND2x2_ASAP7_75t_L g339 ( .A(n_114), .B(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_114), .B(n_150), .Y(n_363) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AND2x2_ASAP7_75t_L g216 ( .A(n_115), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g234 ( .A(n_115), .B(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g246 ( .A(n_115), .B(n_150), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_115), .B(n_160), .Y(n_268) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_123), .B(n_148), .Y(n_115) );
OA21x2_ASAP7_75t_L g160 ( .A1(n_116), .A2(n_161), .B(n_171), .Y(n_160) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
NOR2xp33_ASAP7_75t_L g498 ( .A(n_117), .B(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_118), .Y(n_151) );
AND2x2_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
AND2x2_ASAP7_75t_SL g172 ( .A(n_119), .B(n_120), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_121), .B(n_122), .Y(n_120) );
OAI21xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_137), .B(n_146), .Y(n_123) );
O2A1O1Ixp33_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B(n_130), .C(n_133), .Y(n_124) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_126), .A2(n_496), .B(n_497), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_126), .A2(n_505), .B(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_129), .Y(n_128) );
INVx2_ASAP7_75t_L g132 ( .A(n_129), .Y(n_132) );
INVx1_ASAP7_75t_L g140 ( .A(n_129), .Y(n_140) );
INVx3_ASAP7_75t_L g207 ( .A(n_131), .Y(n_207) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_131), .Y(n_552) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g179 ( .A(n_132), .Y(n_179) );
BUFx3_ASAP7_75t_L g180 ( .A(n_132), .Y(n_180) );
AND2x6_ASAP7_75t_L g451 ( .A(n_132), .B(n_452), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g549 ( .A1(n_133), .A2(n_550), .B(n_551), .C(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_134), .A2(n_211), .B(n_212), .Y(n_210) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g456 ( .A(n_135), .Y(n_456) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx3_ASAP7_75t_L g145 ( .A(n_136), .Y(n_145) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_136), .Y(n_169) );
INVx1_ASAP7_75t_L g190 ( .A(n_136), .Y(n_190) );
AND2x2_ASAP7_75t_L g447 ( .A(n_136), .B(n_140), .Y(n_447) );
INVx1_ASAP7_75t_L g452 ( .A(n_136), .Y(n_452) );
O2A1O1Ixp33_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_141), .B(n_142), .C(n_143), .Y(n_137) );
O2A1O1Ixp5_ASAP7_75t_L g165 ( .A1(n_138), .A2(n_166), .B(n_167), .C(n_168), .Y(n_165) );
AOI21xp5_ASAP7_75t_L g469 ( .A1(n_138), .A2(n_470), .B(n_471), .Y(n_469) );
INVx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
AOI21xp5_ASAP7_75t_L g156 ( .A1(n_143), .A2(n_157), .B(n_158), .Y(n_156) );
OAI22xp5_ASAP7_75t_L g196 ( .A1(n_143), .A2(n_169), .B1(n_197), .B2(n_198), .Y(n_196) );
OAI22xp5_ASAP7_75t_L g221 ( .A1(n_143), .A2(n_169), .B1(n_222), .B2(n_223), .Y(n_221) );
INVx2_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_144), .A2(n_154), .B(n_155), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_144), .A2(n_163), .B(n_164), .Y(n_162) );
O2A1O1Ixp5_ASAP7_75t_SL g206 ( .A1(n_144), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
NOR2xp33_ASAP7_75t_L g525 ( .A(n_144), .B(n_526), .Y(n_525) );
INVx5_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
OAI22xp5_ASAP7_75t_SL g177 ( .A1(n_145), .A2(n_169), .B1(n_178), .B2(n_181), .Y(n_177) );
OAI21xp5_ASAP7_75t_L g152 ( .A1(n_146), .A2(n_153), .B(n_156), .Y(n_152) );
BUFx3_ASAP7_75t_L g170 ( .A(n_146), .Y(n_170) );
OAI21xp5_ASAP7_75t_L g185 ( .A1(n_146), .A2(n_186), .B(n_191), .Y(n_185) );
OAI21xp5_ASAP7_75t_L g205 ( .A1(n_146), .A2(n_206), .B(n_210), .Y(n_205) );
AND2x4_ASAP7_75t_L g446 ( .A(n_146), .B(n_447), .Y(n_446) );
INVx4_ASAP7_75t_SL g460 ( .A(n_146), .Y(n_460) );
NAND2x1p5_ASAP7_75t_L g493 ( .A(n_146), .B(n_447), .Y(n_493) );
AND2x2_ASAP7_75t_L g249 ( .A(n_149), .B(n_250), .Y(n_249) );
AOI221xp5_ASAP7_75t_L g298 ( .A1(n_149), .A2(n_299), .B1(n_302), .B2(n_304), .C(n_308), .Y(n_298) );
AND2x2_ASAP7_75t_L g357 ( .A(n_149), .B(n_322), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_149), .B(n_339), .Y(n_391) );
AND2x2_ASAP7_75t_L g149 ( .A(n_150), .B(n_160), .Y(n_149) );
INVx3_ASAP7_75t_L g217 ( .A(n_150), .Y(n_217) );
AND2x2_ASAP7_75t_L g266 ( .A(n_150), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g320 ( .A(n_150), .B(n_235), .Y(n_320) );
AND2x2_ASAP7_75t_L g378 ( .A(n_150), .B(n_379), .Y(n_378) );
OA21x2_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_152), .B(n_159), .Y(n_150) );
INVx4_ASAP7_75t_L g220 ( .A(n_151), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_151), .A2(n_502), .B(n_503), .Y(n_501) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_151), .Y(n_520) );
AND2x2_ASAP7_75t_L g218 ( .A(n_160), .B(n_219), .Y(n_218) );
INVx2_ASAP7_75t_L g235 ( .A(n_160), .Y(n_235) );
INVx1_ASAP7_75t_L g290 ( .A(n_160), .Y(n_290) );
HB1xp67_ASAP7_75t_L g296 ( .A(n_160), .Y(n_296) );
AND2x2_ASAP7_75t_L g341 ( .A(n_160), .B(n_217), .Y(n_341) );
OR2x2_ASAP7_75t_L g380 ( .A(n_160), .B(n_219), .Y(n_380) );
OAI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_165), .B(n_170), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_168), .A2(n_192), .B(n_193), .Y(n_191) );
INVx2_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx4_ASAP7_75t_L g485 ( .A(n_169), .Y(n_485) );
NAND3xp33_ASAP7_75t_L g239 ( .A(n_170), .B(n_220), .C(n_221), .Y(n_239) );
INVx2_ASAP7_75t_L g182 ( .A(n_172), .Y(n_182) );
OA21x2_ASAP7_75t_L g184 ( .A1(n_172), .A2(n_185), .B(n_194), .Y(n_184) );
OA21x2_ASAP7_75t_L g204 ( .A1(n_172), .A2(n_205), .B(n_213), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g444 ( .A1(n_172), .A2(n_445), .B(n_448), .Y(n_444) );
INVx1_ASAP7_75t_L g475 ( .A(n_172), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_172), .A2(n_512), .B(n_513), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_173), .B(n_260), .Y(n_259) );
AND2x2_ASAP7_75t_L g173 ( .A(n_174), .B(n_183), .Y(n_173) );
AND2x2_ASAP7_75t_L g376 ( .A(n_174), .B(n_373), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_174), .B(n_358), .Y(n_408) );
BUFx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
AND2x2_ASAP7_75t_L g307 ( .A(n_175), .B(n_231), .Y(n_307) );
AND2x2_ASAP7_75t_L g356 ( .A(n_175), .B(n_202), .Y(n_356) );
INVx1_ASAP7_75t_L g402 ( .A(n_175), .Y(n_402) );
INVx1_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_176), .Y(n_215) );
AND2x2_ASAP7_75t_L g257 ( .A(n_176), .B(n_231), .Y(n_257) );
INVx1_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
AND2x2_ASAP7_75t_L g280 ( .A(n_176), .B(n_195), .Y(n_280) );
HB1xp67_ASAP7_75t_L g458 ( .A(n_180), .Y(n_458) );
INVx2_ASAP7_75t_L g486 ( .A(n_180), .Y(n_486) );
INVx1_ASAP7_75t_L g472 ( .A(n_182), .Y(n_472) );
AND2x2_ASAP7_75t_L g348 ( .A(n_183), .B(n_256), .Y(n_348) );
INVx2_ASAP7_75t_L g413 ( .A(n_183), .Y(n_413) );
AND2x2_ASAP7_75t_L g183 ( .A(n_184), .B(n_195), .Y(n_183) );
AND2x2_ASAP7_75t_L g230 ( .A(n_184), .B(n_231), .Y(n_230) );
OR2x2_ASAP7_75t_L g243 ( .A(n_184), .B(n_203), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_184), .B(n_202), .Y(n_271) );
INVx1_ASAP7_75t_L g277 ( .A(n_184), .Y(n_277) );
INVx1_ASAP7_75t_L g294 ( .A(n_184), .Y(n_294) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_184), .Y(n_306) );
INVx2_ASAP7_75t_L g374 ( .A(n_184), .Y(n_374) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_187), .A2(n_188), .B(n_189), .Y(n_186) );
INVx1_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g231 ( .A(n_195), .Y(n_231) );
BUFx2_ASAP7_75t_L g328 ( .A(n_195), .Y(n_328) );
AND2x2_ASAP7_75t_L g373 ( .A(n_195), .B(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_214), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_201), .B(n_310), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_201), .A2(n_372), .B(n_386), .Y(n_396) );
AND2x2_ASAP7_75t_L g421 ( .A(n_201), .B(n_307), .Y(n_421) );
BUFx2_ASAP7_75t_L g201 ( .A(n_202), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_203), .Y(n_202) );
INVx1_ASAP7_75t_L g343 ( .A(n_203), .Y(n_343) );
AND2x2_ASAP7_75t_L g372 ( .A(n_203), .B(n_373), .Y(n_372) );
INVx2_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_204), .Y(n_256) );
INVx2_ASAP7_75t_L g275 ( .A(n_204), .Y(n_275) );
OR2x2_ASAP7_75t_L g276 ( .A(n_204), .B(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
INVx2_ASAP7_75t_L g229 ( .A(n_215), .Y(n_229) );
OR2x2_ASAP7_75t_L g242 ( .A(n_215), .B(n_243), .Y(n_242) );
AND2x2_ASAP7_75t_L g310 ( .A(n_215), .B(n_306), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_215), .B(n_406), .Y(n_405) );
OR2x2_ASAP7_75t_L g411 ( .A(n_215), .B(n_412), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_215), .B(n_348), .Y(n_423) );
AND2x2_ASAP7_75t_L g302 ( .A(n_216), .B(n_303), .Y(n_302) );
AND2x2_ASAP7_75t_L g325 ( .A(n_216), .B(n_218), .Y(n_325) );
INVx2_ASAP7_75t_L g237 ( .A(n_217), .Y(n_237) );
AND2x2_ASAP7_75t_L g265 ( .A(n_217), .B(n_238), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_217), .B(n_290), .Y(n_346) );
AND2x2_ASAP7_75t_L g260 ( .A(n_218), .B(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g407 ( .A(n_218), .Y(n_407) );
AND2x2_ASAP7_75t_L g419 ( .A(n_218), .B(n_282), .Y(n_419) );
AND2x2_ASAP7_75t_L g245 ( .A(n_219), .B(n_235), .Y(n_245) );
INVx1_ASAP7_75t_L g340 ( .A(n_219), .Y(n_340) );
AO21x1_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B(n_224), .Y(n_219) );
NOR2xp33_ASAP7_75t_L g461 ( .A(n_220), .B(n_462), .Y(n_461) );
INVx3_ASAP7_75t_L g478 ( .A(n_220), .Y(n_478) );
AO21x2_ASAP7_75t_L g490 ( .A1(n_220), .A2(n_491), .B(n_498), .Y(n_490) );
AO21x2_ASAP7_75t_L g546 ( .A1(n_220), .A2(n_547), .B(n_554), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_220), .B(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x4_ASAP7_75t_L g238 ( .A(n_225), .B(n_239), .Y(n_238) );
INVxp67_ASAP7_75t_L g226 ( .A(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_232), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g285 ( .A(n_229), .B(n_276), .Y(n_285) );
OR2x2_ASAP7_75t_L g417 ( .A(n_229), .B(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g334 ( .A(n_230), .B(n_275), .Y(n_334) );
AND2x2_ASAP7_75t_L g342 ( .A(n_230), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g401 ( .A(n_230), .B(n_402), .Y(n_401) );
AND2x2_ASAP7_75t_L g425 ( .A(n_230), .B(n_272), .Y(n_425) );
NOR2xp67_ASAP7_75t_L g383 ( .A(n_231), .B(n_384), .Y(n_383) );
OR2x2_ASAP7_75t_L g412 ( .A(n_231), .B(n_275), .Y(n_412) );
INVx1_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
NAND2x1p5_ASAP7_75t_L g233 ( .A(n_234), .B(n_236), .Y(n_233) );
AND2x2_ASAP7_75t_L g264 ( .A(n_234), .B(n_265), .Y(n_264) );
INVxp67_ASAP7_75t_L g426 ( .A(n_234), .Y(n_426) );
NOR2x1_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
INVx1_ASAP7_75t_L g261 ( .A(n_237), .Y(n_261) );
AND2x2_ASAP7_75t_L g312 ( .A(n_237), .B(n_245), .Y(n_312) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_237), .B(n_380), .Y(n_406) );
INVx2_ASAP7_75t_L g251 ( .A(n_238), .Y(n_251) );
INVx3_ASAP7_75t_L g303 ( .A(n_238), .Y(n_303) );
OR2x2_ASAP7_75t_L g331 ( .A(n_238), .B(n_332), .Y(n_331) );
AOI311xp33_ASAP7_75t_L g240 ( .A1(n_241), .A2(n_244), .A3(n_246), .B(n_247), .C(n_258), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g278 ( .A1(n_241), .A2(n_279), .B(n_281), .C(n_283), .Y(n_278) );
INVx2_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx2_ASAP7_75t_SL g263 ( .A(n_243), .Y(n_263) );
INVx2_ASAP7_75t_L g244 ( .A(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g281 ( .A(n_245), .B(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_245), .B(n_261), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_245), .B(n_246), .Y(n_414) );
AND2x2_ASAP7_75t_L g336 ( .A(n_246), .B(n_250), .Y(n_336) );
AOI21xp33_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_252), .B(n_253), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g394 ( .A(n_250), .B(n_282), .Y(n_394) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g267 ( .A(n_251), .B(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g288 ( .A(n_251), .Y(n_288) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_257), .Y(n_254) );
AND2x2_ASAP7_75t_L g279 ( .A(n_255), .B(n_280), .Y(n_279) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
INVx1_ASAP7_75t_L g324 ( .A(n_257), .Y(n_324) );
AND2x4_ASAP7_75t_L g386 ( .A(n_257), .B(n_355), .Y(n_386) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AOI222xp33_ASAP7_75t_L g337 ( .A1(n_260), .A2(n_326), .B1(n_338), .B2(n_342), .C1(n_344), .C2(n_348), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_264), .B(n_266), .C(n_269), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_263), .B(n_307), .Y(n_330) );
INVx1_ASAP7_75t_L g352 ( .A(n_265), .Y(n_352) );
INVx1_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
OR2x2_ASAP7_75t_L g351 ( .A(n_268), .B(n_352), .Y(n_351) );
OAI21xp33_ASAP7_75t_SL g269 ( .A1(n_270), .A2(n_272), .B(n_276), .Y(n_269) );
NAND3xp33_ASAP7_75t_L g287 ( .A(n_270), .B(n_288), .C(n_289), .Y(n_287) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_270), .A2(n_307), .B(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
INVx1_ASAP7_75t_SL g272 ( .A(n_273), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_275), .Y(n_273) );
HB1xp67_ASAP7_75t_L g327 ( .A(n_274), .Y(n_327) );
AND2x2_ASAP7_75t_SL g293 ( .A(n_275), .B(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g384 ( .A(n_275), .Y(n_384) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_275), .Y(n_400) );
INVx2_ASAP7_75t_L g358 ( .A(n_276), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_280), .B(n_301), .Y(n_300) );
INVx2_ASAP7_75t_L g332 ( .A(n_282), .Y(n_332) );
OAI221xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_286), .B1(n_287), .B2(n_291), .C(n_292), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_286), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_SL g420 ( .A(n_286), .Y(n_420) );
INVx1_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g301 ( .A(n_293), .Y(n_301) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_293), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g359 ( .A(n_293), .B(n_307), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_293), .B(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g392 ( .A(n_293), .B(n_327), .Y(n_392) );
BUFx3_ASAP7_75t_L g355 ( .A(n_294), .Y(n_355) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
NAND5xp2_ASAP7_75t_L g297 ( .A(n_298), .B(n_316), .C(n_337), .D(n_349), .E(n_364), .Y(n_297) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AOI32xp33_ASAP7_75t_L g389 ( .A1(n_301), .A2(n_328), .A3(n_344), .B1(n_390), .B2(n_392), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_303), .B(n_362), .Y(n_361) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
INVx1_ASAP7_75t_SL g313 ( .A(n_307), .Y(n_313) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_309), .A2(n_311), .B1(n_313), .B2(n_314), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx1_ASAP7_75t_SL g314 ( .A(n_315), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_323), .B1(n_325), .B2(n_326), .C(n_329), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g388 ( .A(n_320), .B(n_339), .Y(n_388) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g403 ( .A1(n_325), .A2(n_386), .B1(n_404), .B2(n_409), .C(n_410), .Y(n_403) );
AND2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx2_ASAP7_75t_L g369 ( .A(n_328), .Y(n_369) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_330), .A2(n_331), .B1(n_333), .B2(n_335), .Y(n_329) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_SL g335 ( .A(n_336), .Y(n_335) );
AND2x2_ASAP7_75t_L g338 ( .A(n_339), .B(n_341), .Y(n_338) );
INVx1_ASAP7_75t_L g347 ( .A(n_339), .Y(n_347) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B1(n_357), .B2(n_358), .C1(n_359), .C2(n_360), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
OAI22xp33_ASAP7_75t_L g404 ( .A1(n_358), .A2(n_405), .B1(n_407), .B2(n_408), .Y(n_404) );
INVx1_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
AOI21xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_367), .B(n_370), .Y(n_364) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
AOI21xp33_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B(n_377), .Y(n_370) );
INVx2_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
INVx1_ASAP7_75t_L g418 ( .A(n_373), .Y(n_418) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g381 ( .A1(n_382), .A2(n_385), .B(n_387), .C(n_389), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
AOI211xp5_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_395), .B(n_397), .C(n_422), .Y(n_393) );
CKINVDCx16_ASAP7_75t_R g398 ( .A(n_394), .Y(n_398) );
INVxp67_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OAI211xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_399), .B(n_403), .C(n_415), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AOI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_413), .B(n_414), .Y(n_410) );
AOI22xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_419), .B1(n_420), .B2(n_421), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
AOI21xp33_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_426), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx2_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
OR2x2_ASAP7_75t_L g436 ( .A(n_431), .B(n_437), .Y(n_436) );
INVx2_ASAP7_75t_L g730 ( .A(n_431), .Y(n_730) );
AND2x2_ASAP7_75t_L g431 ( .A(n_432), .B(n_433), .Y(n_431) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
NOR2x2_ASAP7_75t_L g729 ( .A(n_437), .B(n_730), .Y(n_729) );
INVx2_ASAP7_75t_L g726 ( .A(n_438), .Y(n_726) );
OR3x2_ASAP7_75t_L g438 ( .A(n_439), .B(n_638), .C(n_681), .Y(n_438) );
NAND5xp2_ASAP7_75t_L g439 ( .A(n_440), .B(n_565), .C(n_595), .D(n_612), .E(n_627), .Y(n_439) );
AOI221xp5_ASAP7_75t_SL g440 ( .A1(n_441), .A2(n_488), .B1(n_528), .B2(n_534), .C(n_538), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_442), .B(n_463), .Y(n_441) );
OR2x2_ASAP7_75t_L g543 ( .A(n_442), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g582 ( .A(n_442), .B(n_583), .Y(n_582) );
AND2x2_ASAP7_75t_L g600 ( .A(n_442), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_442), .B(n_536), .Y(n_617) );
OR2x2_ASAP7_75t_L g629 ( .A(n_442), .B(n_630), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_442), .B(n_588), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g661 ( .A(n_442), .B(n_662), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_442), .B(n_566), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_442), .B(n_574), .Y(n_680) );
AND2x2_ASAP7_75t_L g712 ( .A(n_442), .B(n_476), .Y(n_712) );
HB1xp67_ASAP7_75t_L g720 ( .A(n_442), .Y(n_720) );
INVx5_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_443), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g540 ( .A(n_443), .B(n_518), .Y(n_540) );
BUFx2_ASAP7_75t_L g562 ( .A(n_443), .Y(n_562) );
AND2x2_ASAP7_75t_L g591 ( .A(n_443), .B(n_464), .Y(n_591) );
AND2x2_ASAP7_75t_L g646 ( .A(n_443), .B(n_544), .Y(n_646) );
OR2x6_ASAP7_75t_L g443 ( .A(n_444), .B(n_461), .Y(n_443) );
BUFx2_ASAP7_75t_L g467 ( .A(n_446), .Y(n_467) );
INVx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
O2A1O1Ixp33_ASAP7_75t_SL g480 ( .A1(n_450), .A2(n_460), .B(n_481), .C(n_482), .Y(n_480) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_450), .A2(n_460), .B(n_523), .C(n_524), .Y(n_522) );
INVx5_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
O2A1O1Ixp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_455), .B(n_457), .C(n_458), .Y(n_453) );
O2A1O1Ixp33_ASAP7_75t_L g514 ( .A1(n_455), .A2(n_458), .B(n_515), .C(n_516), .Y(n_514) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_463), .B(n_600), .Y(n_609) );
OAI32xp33_ASAP7_75t_L g623 ( .A1(n_463), .A2(n_559), .A3(n_624), .B1(n_625), .B2(n_626), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_463), .B(n_625), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_463), .B(n_543), .Y(n_666) );
INVx1_ASAP7_75t_SL g695 ( .A(n_463), .Y(n_695) );
NAND4xp25_ASAP7_75t_L g704 ( .A(n_463), .B(n_490), .C(n_646), .D(n_705), .Y(n_704) );
AND2x4_ASAP7_75t_L g463 ( .A(n_464), .B(n_476), .Y(n_463) );
INVx5_ASAP7_75t_L g537 ( .A(n_464), .Y(n_537) );
AND2x2_ASAP7_75t_L g566 ( .A(n_464), .B(n_477), .Y(n_566) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_464), .Y(n_645) );
AND2x2_ASAP7_75t_L g715 ( .A(n_464), .B(n_662), .Y(n_715) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_473), .Y(n_464) );
AOI21xp5_ASAP7_75t_SL g465 ( .A1(n_466), .A2(n_468), .B(n_472), .Y(n_465) );
NOR2xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_475), .Y(n_473) );
AND2x4_ASAP7_75t_L g588 ( .A(n_476), .B(n_537), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g597 ( .A(n_476), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g622 ( .A(n_476), .B(n_544), .Y(n_622) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
AND2x2_ASAP7_75t_L g536 ( .A(n_477), .B(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g574 ( .A(n_477), .B(n_546), .Y(n_574) );
AND2x2_ASAP7_75t_L g583 ( .A(n_477), .B(n_545), .Y(n_583) );
OA21x2_ASAP7_75t_L g477 ( .A1(n_478), .A2(n_479), .B(n_487), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
AOI222xp33_ASAP7_75t_L g651 ( .A1(n_488), .A2(n_652), .B1(n_654), .B2(n_656), .C1(n_659), .C2(n_660), .Y(n_651) );
AND2x4_ASAP7_75t_L g488 ( .A(n_489), .B(n_507), .Y(n_488) );
AND2x2_ASAP7_75t_L g584 ( .A(n_489), .B(n_585), .Y(n_584) );
NAND3xp33_ASAP7_75t_L g701 ( .A(n_489), .B(n_562), .C(n_702), .Y(n_701) );
AND2x2_ASAP7_75t_L g489 ( .A(n_490), .B(n_500), .Y(n_489) );
INVx5_ASAP7_75t_SL g533 ( .A(n_490), .Y(n_533) );
OAI322xp33_ASAP7_75t_L g538 ( .A1(n_490), .A2(n_539), .A3(n_541), .B1(n_542), .B2(n_556), .C1(n_559), .C2(n_561), .Y(n_538) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_490), .B(n_531), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_490), .B(n_519), .Y(n_710) );
OAI21xp5_ASAP7_75t_L g491 ( .A1(n_492), .A2(n_493), .B(n_494), .Y(n_491) );
INVx2_ASAP7_75t_L g531 ( .A(n_500), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_500), .B(n_509), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_507), .B(n_569), .Y(n_624) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g603 ( .A(n_508), .B(n_604), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_518), .Y(n_508) );
OR2x2_ASAP7_75t_L g532 ( .A(n_509), .B(n_533), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_509), .B(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g571 ( .A(n_509), .B(n_519), .Y(n_571) );
AND2x2_ASAP7_75t_L g594 ( .A(n_509), .B(n_531), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g605 ( .A(n_509), .B(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g610 ( .A(n_509), .B(n_569), .Y(n_610) );
AND2x2_ASAP7_75t_L g618 ( .A(n_509), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_509), .B(n_578), .Y(n_668) );
INVx5_ASAP7_75t_SL g509 ( .A(n_510), .Y(n_509) );
AND2x2_ASAP7_75t_L g558 ( .A(n_510), .B(n_533), .Y(n_558) );
OR2x2_ASAP7_75t_L g559 ( .A(n_510), .B(n_560), .Y(n_559) );
AND2x2_ASAP7_75t_L g585 ( .A(n_510), .B(n_519), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_510), .B(n_632), .Y(n_673) );
OR2x2_ASAP7_75t_L g689 ( .A(n_510), .B(n_633), .Y(n_689) );
AND2x2_ASAP7_75t_SL g696 ( .A(n_510), .B(n_650), .Y(n_696) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_510), .Y(n_703) );
OR2x6_ASAP7_75t_L g510 ( .A(n_511), .B(n_517), .Y(n_510) );
AND2x2_ASAP7_75t_L g557 ( .A(n_518), .B(n_558), .Y(n_557) );
AND2x2_ASAP7_75t_L g607 ( .A(n_518), .B(n_531), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_518), .B(n_533), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_518), .B(n_569), .Y(n_691) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_519), .B(n_533), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_519), .B(n_531), .Y(n_579) );
OR2x2_ASAP7_75t_L g633 ( .A(n_519), .B(n_531), .Y(n_633) );
AND2x2_ASAP7_75t_L g650 ( .A(n_519), .B(n_530), .Y(n_650) );
INVxp67_ASAP7_75t_L g672 ( .A(n_519), .Y(n_672) );
AND2x2_ASAP7_75t_L g699 ( .A(n_519), .B(n_569), .Y(n_699) );
HB1xp67_ASAP7_75t_L g706 ( .A(n_519), .Y(n_706) );
OA21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_519) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_530), .B(n_580), .Y(n_653) );
INVx1_ASAP7_75t_SL g530 ( .A(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g569 ( .A(n_531), .B(n_533), .Y(n_569) );
OR2x2_ASAP7_75t_L g636 ( .A(n_531), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g580 ( .A(n_532), .Y(n_580) );
OR2x2_ASAP7_75t_L g641 ( .A(n_532), .B(n_633), .Y(n_641) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
INVx1_ASAP7_75t_L g541 ( .A(n_536), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_536), .B(n_600), .Y(n_599) );
OR2x2_ASAP7_75t_L g542 ( .A(n_537), .B(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_537), .B(n_564), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_537), .B(n_544), .Y(n_576) );
INVx2_ASAP7_75t_L g621 ( .A(n_537), .Y(n_621) );
AND2x2_ASAP7_75t_L g634 ( .A(n_537), .B(n_574), .Y(n_634) );
AND2x2_ASAP7_75t_L g659 ( .A(n_537), .B(n_583), .Y(n_659) );
INVx1_ASAP7_75t_L g611 ( .A(n_542), .Y(n_611) );
INVx2_ASAP7_75t_SL g598 ( .A(n_543), .Y(n_598) );
INVx1_ASAP7_75t_L g601 ( .A(n_544), .Y(n_601) );
INVx2_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g564 ( .A(n_545), .Y(n_564) );
INVx2_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
BUFx2_ASAP7_75t_L g662 ( .A(n_546), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_548), .B(n_553), .Y(n_547) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g631 ( .A(n_558), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
AOI22xp5_ASAP7_75t_L g639 ( .A1(n_558), .A2(n_640), .B1(n_642), .B2(n_647), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_558), .B(n_650), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_559), .B(n_653), .Y(n_652) );
INVx1_ASAP7_75t_SL g593 ( .A(n_560), .Y(n_593) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OR2x2_ASAP7_75t_L g575 ( .A(n_562), .B(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_562), .B(n_566), .Y(n_626) );
AND2x2_ASAP7_75t_L g649 ( .A(n_562), .B(n_650), .Y(n_649) );
BUFx2_ASAP7_75t_L g625 ( .A(n_564), .Y(n_625) );
AOI211xp5_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_567), .B(n_572), .C(n_586), .Y(n_565) );
INVx1_ASAP7_75t_L g589 ( .A(n_566), .Y(n_589) );
OAI221xp5_ASAP7_75t_SL g697 ( .A1(n_566), .A2(n_698), .B1(n_700), .B2(n_701), .C(n_704), .Y(n_697) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
INVx1_ASAP7_75t_L g716 ( .A(n_569), .Y(n_716) );
INVx1_ASAP7_75t_L g570 ( .A(n_571), .Y(n_570) );
OR2x2_ASAP7_75t_L g665 ( .A(n_571), .B(n_604), .Y(n_665) );
A2O1A1Ixp33_ASAP7_75t_L g572 ( .A1(n_573), .A2(n_575), .B(n_577), .C(n_581), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_578), .B(n_580), .Y(n_577) );
INVx1_ASAP7_75t_SL g578 ( .A(n_579), .Y(n_578) );
OAI32xp33_ASAP7_75t_L g690 ( .A1(n_579), .A2(n_580), .A3(n_643), .B1(n_680), .B2(n_691), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_584), .Y(n_581) );
AND2x2_ASAP7_75t_L g722 ( .A(n_582), .B(n_621), .Y(n_722) );
AND2x2_ASAP7_75t_L g669 ( .A(n_583), .B(n_621), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_583), .B(n_591), .Y(n_687) );
AOI31xp33_ASAP7_75t_SL g586 ( .A1(n_587), .A2(n_589), .A3(n_590), .B(n_592), .Y(n_586) );
INVxp67_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_588), .B(n_600), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_588), .B(n_598), .Y(n_685) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_588), .A2(n_618), .B1(n_708), .B2(n_711), .C(n_713), .Y(n_707) );
CKINVDCx16_ASAP7_75t_R g590 ( .A(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g613 ( .A(n_593), .B(n_614), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_602), .B1(n_605), .B2(n_608), .C1(n_610), .C2(n_611), .Y(n_595) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx1_ASAP7_75t_L g678 ( .A(n_597), .Y(n_678) );
INVx1_ASAP7_75t_L g700 ( .A(n_600), .Y(n_700) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_603), .A2(n_714), .B1(n_716), .B2(n_717), .Y(n_713) );
INVx1_ASAP7_75t_L g619 ( .A(n_604), .Y(n_619) );
INVx1_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_616), .B1(n_618), .B2(n_620), .C(n_623), .Y(n_612) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
OR2x2_ASAP7_75t_L g657 ( .A(n_615), .B(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g709 ( .A(n_615), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
INVx1_ASAP7_75t_L g684 ( .A(n_620), .Y(n_684) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g648 ( .A(n_621), .Y(n_648) );
INVx1_ASAP7_75t_L g630 ( .A(n_622), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_625), .B(n_712), .Y(n_717) );
AOI22xp33_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_631), .B1(n_634), .B2(n_635), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_SL g721 ( .A(n_634), .Y(n_721) );
INVxp33_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_636), .B(n_680), .Y(n_679) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_637), .A2(n_671), .A3(n_672), .B1(n_673), .B2(n_674), .Y(n_670) );
NAND4xp25_ASAP7_75t_L g638 ( .A(n_639), .B(n_651), .C(n_663), .D(n_675), .Y(n_638) );
INVx1_ASAP7_75t_SL g640 ( .A(n_641), .Y(n_640) );
NAND2xp33_ASAP7_75t_SL g642 ( .A(n_643), .B(n_644), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_645), .B(n_646), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_646), .B(n_695), .Y(n_694) );
AND2x2_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
CKINVDCx16_ASAP7_75t_R g656 ( .A(n_657), .Y(n_656) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_660), .A2(n_676), .B1(n_693), .B2(n_696), .C(n_697), .Y(n_692) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AND2x2_ASAP7_75t_L g711 ( .A(n_662), .B(n_712), .Y(n_711) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B1(n_667), .B2(n_669), .C(n_670), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g702 ( .A(n_672), .B(n_703), .Y(n_702) );
AOI21xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .B(n_679), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g681 ( .A(n_682), .B(n_692), .C(n_707), .D(n_718), .Y(n_681) );
O2A1O1Ixp33_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_686), .B(n_688), .C(n_690), .Y(n_682) );
NAND2xp5_ASAP7_75t_SL g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVxp67_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g723 ( .A(n_710), .Y(n_723) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
OAI21xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B(n_723), .Y(n_718) );
NOR2xp33_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NAND2xp33_ASAP7_75t_L g732 ( .A(n_733), .B(n_737), .Y(n_732) );
NOR2xp33_ASAP7_75t_SL g733 ( .A(n_734), .B(n_736), .Y(n_733) );
INVx1_ASAP7_75t_SL g754 ( .A(n_734), .Y(n_754) );
INVx1_ASAP7_75t_L g753 ( .A(n_736), .Y(n_753) );
OA21x2_ASAP7_75t_L g756 ( .A1(n_736), .A2(n_754), .B(n_757), .Y(n_756) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_SL g738 ( .A(n_739), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g741 ( .A1(n_739), .A2(n_742), .B(n_746), .Y(n_741) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_739), .Y(n_747) );
BUFx2_ASAP7_75t_L g757 ( .A(n_739), .Y(n_757) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
CKINVDCx20_ASAP7_75t_R g743 ( .A(n_744), .Y(n_743) );
NOR2xp33_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_750), .Y(n_749) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_752), .B(n_754), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
endmodule