module fake_jpeg_24333_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g7 ( 
.A(n_2),
.Y(n_7)
);

BUFx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

BUFx3_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

INVx8_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_5),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

OA22x2_ASAP7_75t_L g15 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_15)
);

XNOR2xp5_ASAP7_75t_L g27 ( 
.A(n_15),
.B(n_19),
.Y(n_27)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx10_ASAP7_75t_R g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx10_ASAP7_75t_R g24 ( 
.A(n_17),
.Y(n_24)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_18),
.A2(n_20),
.B(n_11),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_10),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_14),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_21),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_18),
.B(n_13),
.C(n_11),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_20),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_26),
.B(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_28),
.A2(n_31),
.B1(n_10),
.B2(n_16),
.Y(n_33)
);

NOR3xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_32),
.C(n_12),
.Y(n_35)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_15),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_14),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.C(n_19),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_21),
.B1(n_22),
.B2(n_15),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_35),
.A2(n_12),
.B(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_38),
.Y(n_41)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_40),
.B1(n_15),
.B2(n_10),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_35),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_34),
.C(n_17),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_43),
.Y(n_45)
);

AOI322xp5_ASAP7_75t_L g44 ( 
.A1(n_42),
.A2(n_8),
.A3(n_13),
.B1(n_7),
.B2(n_6),
.C1(n_5),
.C2(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_44),
.B(n_41),
.Y(n_46)
);

AOI322xp5_ASAP7_75t_L g47 ( 
.A1(n_46),
.A2(n_1),
.A3(n_7),
.B1(n_8),
.B2(n_45),
.C1(n_41),
.C2(n_33),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g48 ( 
.A(n_47),
.B(n_8),
.Y(n_48)
);


endmodule