module fake_ariane_257_n_5709 (n_295, n_356, n_556, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_386, n_307, n_516, n_589, n_332, n_581, n_294, n_646, n_197, n_640, n_463, n_176, n_34, n_404, n_172, n_678, n_651, n_347, n_423, n_183, n_469, n_479, n_603, n_373, n_299, n_541, n_499, n_12, n_564, n_133, n_610, n_66, n_205, n_341, n_71, n_109, n_245, n_421, n_96, n_549, n_522, n_319, n_49, n_591, n_20, n_690, n_416, n_283, n_50, n_187, n_525, n_367, n_649, n_598, n_345, n_374, n_318, n_103, n_244, n_643, n_679, n_226, n_220, n_261, n_682, n_36, n_663, n_370, n_189, n_72, n_286, n_443, n_586, n_57, n_686, n_605, n_424, n_528, n_584, n_387, n_406, n_117, n_139, n_524, n_85, n_130, n_349, n_391, n_634, n_466, n_346, n_214, n_348, n_552, n_2, n_462, n_607, n_670, n_32, n_410, n_379, n_445, n_515, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_441, n_568, n_385, n_637, n_73, n_327, n_77, n_372, n_377, n_15, n_396, n_631, n_23, n_399, n_554, n_520, n_87, n_279, n_207, n_363, n_354, n_41, n_140, n_419, n_151, n_28, n_146, n_230, n_270, n_194, n_633, n_154, n_338, n_142, n_285, n_473, n_186, n_202, n_145, n_193, n_500, n_665, n_59, n_336, n_315, n_594, n_311, n_239, n_402, n_35, n_272, n_54, n_8, n_668, n_339, n_672, n_487, n_167, n_90, n_38, n_422, n_47, n_153, n_18, n_648, n_269, n_597, n_75, n_158, n_69, n_259, n_95, n_446, n_553, n_143, n_566, n_578, n_625, n_152, n_405, n_557, n_120, n_169, n_106, n_173, n_242, n_645, n_309, n_320, n_115, n_331, n_559, n_401, n_485, n_267, n_495, n_504, n_647, n_483, n_335, n_435, n_350, n_291, n_344, n_381, n_426, n_433, n_481, n_600, n_398, n_62, n_210, n_200, n_529, n_502, n_166, n_253, n_561, n_218, n_79, n_3, n_271, n_465, n_486, n_507, n_247, n_569, n_567, n_91, n_240, n_369, n_128, n_224, n_44, n_82, n_31, n_547, n_420, n_562, n_518, n_439, n_604, n_614, n_677, n_222, n_478, n_510, n_256, n_326, n_681, n_227, n_48, n_188, n_323, n_550, n_635, n_330, n_400, n_689, n_11, n_129, n_126, n_282, n_328, n_368, n_590, n_277, n_248, n_301, n_467, n_432, n_545, n_536, n_644, n_293, n_620, n_228, n_325, n_276, n_93, n_688, n_636, n_427, n_108, n_587, n_497, n_303, n_671, n_442, n_168, n_81, n_1, n_206, n_352, n_538, n_576, n_511, n_611, n_238, n_365, n_429, n_455, n_654, n_588, n_638, n_136, n_334, n_192, n_661, n_488, n_667, n_300, n_533, n_505, n_14, n_163, n_88, n_141, n_390, n_498, n_104, n_501, n_438, n_314, n_684, n_16, n_440, n_627, n_273, n_305, n_539, n_312, n_233, n_56, n_60, n_388, n_333, n_449, n_612, n_413, n_392, n_376, n_512, n_579, n_459, n_685, n_221, n_321, n_86, n_361, n_458, n_89, n_149, n_383, n_623, n_237, n_175, n_453, n_74, n_491, n_19, n_40, n_181, n_616, n_617, n_658, n_630, n_570, n_53, n_260, n_362, n_543, n_310, n_236, n_601, n_683, n_565, n_281, n_24, n_7, n_628, n_461, n_209, n_262, n_490, n_17, n_225, n_235, n_660, n_464, n_575, n_546, n_297, n_662, n_641, n_503, n_290, n_527, n_46, n_84, n_371, n_199, n_107, n_639, n_217, n_452, n_673, n_676, n_178, n_42, n_551, n_308, n_417, n_201, n_70, n_572, n_343, n_10, n_414, n_571, n_680, n_287, n_302, n_380, n_6, n_582, n_94, n_284, n_4, n_448, n_593, n_249, n_534, n_37, n_58, n_65, n_123, n_212, n_355, n_444, n_609, n_278, n_255, n_560, n_450, n_257, n_148, n_652, n_451, n_613, n_475, n_135, n_409, n_171, n_519, n_384, n_468, n_61, n_526, n_102, n_182, n_674, n_482, n_316, n_196, n_125, n_43, n_577, n_407, n_13, n_27, n_254, n_596, n_476, n_460, n_219, n_55, n_535, n_231, n_366, n_656, n_555, n_234, n_492, n_574, n_280, n_215, n_252, n_629, n_664, n_161, n_454, n_298, n_532, n_68, n_415, n_78, n_63, n_655, n_99, n_540, n_216, n_544, n_5, n_599, n_514, n_418, n_537, n_223, n_403, n_25, n_83, n_389, n_657, n_513, n_288, n_179, n_395, n_621, n_195, n_606, n_213, n_110, n_304, n_659, n_67, n_509, n_583, n_306, n_666, n_313, n_92, n_430, n_626, n_493, n_203, n_378, n_436, n_150, n_98, n_375, n_113, n_114, n_33, n_324, n_585, n_669, n_619, n_337, n_437, n_111, n_21, n_274, n_622, n_472, n_296, n_265, n_208, n_456, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_615, n_521, n_51, n_496, n_76, n_342, n_26, n_246, n_517, n_530, n_0, n_428, n_159, n_358, n_105, n_580, n_608, n_30, n_494, n_131, n_263, n_434, n_360, n_563, n_229, n_394, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_329, n_185, n_340, n_289, n_9, n_112, n_45, n_542, n_548, n_523, n_268, n_266, n_470, n_457, n_164, n_157, n_632, n_184, n_177, n_477, n_364, n_258, n_650, n_425, n_431, n_508, n_624, n_118, n_121, n_618, n_411, n_484, n_353, n_22, n_241, n_29, n_357, n_412, n_687, n_447, n_191, n_382, n_489, n_80, n_480, n_211, n_642, n_97, n_408, n_595, n_322, n_251, n_506, n_602, n_558, n_592, n_116, n_397, n_471, n_351, n_39, n_393, n_474, n_653, n_359, n_155, n_573, n_127, n_531, n_675, n_5709);

input n_295;
input n_356;
input n_556;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_386;
input n_307;
input n_516;
input n_589;
input n_332;
input n_581;
input n_294;
input n_646;
input n_197;
input n_640;
input n_463;
input n_176;
input n_34;
input n_404;
input n_172;
input n_678;
input n_651;
input n_347;
input n_423;
input n_183;
input n_469;
input n_479;
input n_603;
input n_373;
input n_299;
input n_541;
input n_499;
input n_12;
input n_564;
input n_133;
input n_610;
input n_66;
input n_205;
input n_341;
input n_71;
input n_109;
input n_245;
input n_421;
input n_96;
input n_549;
input n_522;
input n_319;
input n_49;
input n_591;
input n_20;
input n_690;
input n_416;
input n_283;
input n_50;
input n_187;
input n_525;
input n_367;
input n_649;
input n_598;
input n_345;
input n_374;
input n_318;
input n_103;
input n_244;
input n_643;
input n_679;
input n_226;
input n_220;
input n_261;
input n_682;
input n_36;
input n_663;
input n_370;
input n_189;
input n_72;
input n_286;
input n_443;
input n_586;
input n_57;
input n_686;
input n_605;
input n_424;
input n_528;
input n_584;
input n_387;
input n_406;
input n_117;
input n_139;
input n_524;
input n_85;
input n_130;
input n_349;
input n_391;
input n_634;
input n_466;
input n_346;
input n_214;
input n_348;
input n_552;
input n_2;
input n_462;
input n_607;
input n_670;
input n_32;
input n_410;
input n_379;
input n_445;
input n_515;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_441;
input n_568;
input n_385;
input n_637;
input n_73;
input n_327;
input n_77;
input n_372;
input n_377;
input n_15;
input n_396;
input n_631;
input n_23;
input n_399;
input n_554;
input n_520;
input n_87;
input n_279;
input n_207;
input n_363;
input n_354;
input n_41;
input n_140;
input n_419;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_633;
input n_154;
input n_338;
input n_142;
input n_285;
input n_473;
input n_186;
input n_202;
input n_145;
input n_193;
input n_500;
input n_665;
input n_59;
input n_336;
input n_315;
input n_594;
input n_311;
input n_239;
input n_402;
input n_35;
input n_272;
input n_54;
input n_8;
input n_668;
input n_339;
input n_672;
input n_487;
input n_167;
input n_90;
input n_38;
input n_422;
input n_47;
input n_153;
input n_18;
input n_648;
input n_269;
input n_597;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_446;
input n_553;
input n_143;
input n_566;
input n_578;
input n_625;
input n_152;
input n_405;
input n_557;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_645;
input n_309;
input n_320;
input n_115;
input n_331;
input n_559;
input n_401;
input n_485;
input n_267;
input n_495;
input n_504;
input n_647;
input n_483;
input n_335;
input n_435;
input n_350;
input n_291;
input n_344;
input n_381;
input n_426;
input n_433;
input n_481;
input n_600;
input n_398;
input n_62;
input n_210;
input n_200;
input n_529;
input n_502;
input n_166;
input n_253;
input n_561;
input n_218;
input n_79;
input n_3;
input n_271;
input n_465;
input n_486;
input n_507;
input n_247;
input n_569;
input n_567;
input n_91;
input n_240;
input n_369;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_547;
input n_420;
input n_562;
input n_518;
input n_439;
input n_604;
input n_614;
input n_677;
input n_222;
input n_478;
input n_510;
input n_256;
input n_326;
input n_681;
input n_227;
input n_48;
input n_188;
input n_323;
input n_550;
input n_635;
input n_330;
input n_400;
input n_689;
input n_11;
input n_129;
input n_126;
input n_282;
input n_328;
input n_368;
input n_590;
input n_277;
input n_248;
input n_301;
input n_467;
input n_432;
input n_545;
input n_536;
input n_644;
input n_293;
input n_620;
input n_228;
input n_325;
input n_276;
input n_93;
input n_688;
input n_636;
input n_427;
input n_108;
input n_587;
input n_497;
input n_303;
input n_671;
input n_442;
input n_168;
input n_81;
input n_1;
input n_206;
input n_352;
input n_538;
input n_576;
input n_511;
input n_611;
input n_238;
input n_365;
input n_429;
input n_455;
input n_654;
input n_588;
input n_638;
input n_136;
input n_334;
input n_192;
input n_661;
input n_488;
input n_667;
input n_300;
input n_533;
input n_505;
input n_14;
input n_163;
input n_88;
input n_141;
input n_390;
input n_498;
input n_104;
input n_501;
input n_438;
input n_314;
input n_684;
input n_16;
input n_440;
input n_627;
input n_273;
input n_305;
input n_539;
input n_312;
input n_233;
input n_56;
input n_60;
input n_388;
input n_333;
input n_449;
input n_612;
input n_413;
input n_392;
input n_376;
input n_512;
input n_579;
input n_459;
input n_685;
input n_221;
input n_321;
input n_86;
input n_361;
input n_458;
input n_89;
input n_149;
input n_383;
input n_623;
input n_237;
input n_175;
input n_453;
input n_74;
input n_491;
input n_19;
input n_40;
input n_181;
input n_616;
input n_617;
input n_658;
input n_630;
input n_570;
input n_53;
input n_260;
input n_362;
input n_543;
input n_310;
input n_236;
input n_601;
input n_683;
input n_565;
input n_281;
input n_24;
input n_7;
input n_628;
input n_461;
input n_209;
input n_262;
input n_490;
input n_17;
input n_225;
input n_235;
input n_660;
input n_464;
input n_575;
input n_546;
input n_297;
input n_662;
input n_641;
input n_503;
input n_290;
input n_527;
input n_46;
input n_84;
input n_371;
input n_199;
input n_107;
input n_639;
input n_217;
input n_452;
input n_673;
input n_676;
input n_178;
input n_42;
input n_551;
input n_308;
input n_417;
input n_201;
input n_70;
input n_572;
input n_343;
input n_10;
input n_414;
input n_571;
input n_680;
input n_287;
input n_302;
input n_380;
input n_6;
input n_582;
input n_94;
input n_284;
input n_4;
input n_448;
input n_593;
input n_249;
input n_534;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_355;
input n_444;
input n_609;
input n_278;
input n_255;
input n_560;
input n_450;
input n_257;
input n_148;
input n_652;
input n_451;
input n_613;
input n_475;
input n_135;
input n_409;
input n_171;
input n_519;
input n_384;
input n_468;
input n_61;
input n_526;
input n_102;
input n_182;
input n_674;
input n_482;
input n_316;
input n_196;
input n_125;
input n_43;
input n_577;
input n_407;
input n_13;
input n_27;
input n_254;
input n_596;
input n_476;
input n_460;
input n_219;
input n_55;
input n_535;
input n_231;
input n_366;
input n_656;
input n_555;
input n_234;
input n_492;
input n_574;
input n_280;
input n_215;
input n_252;
input n_629;
input n_664;
input n_161;
input n_454;
input n_298;
input n_532;
input n_68;
input n_415;
input n_78;
input n_63;
input n_655;
input n_99;
input n_540;
input n_216;
input n_544;
input n_5;
input n_599;
input n_514;
input n_418;
input n_537;
input n_223;
input n_403;
input n_25;
input n_83;
input n_389;
input n_657;
input n_513;
input n_288;
input n_179;
input n_395;
input n_621;
input n_195;
input n_606;
input n_213;
input n_110;
input n_304;
input n_659;
input n_67;
input n_509;
input n_583;
input n_306;
input n_666;
input n_313;
input n_92;
input n_430;
input n_626;
input n_493;
input n_203;
input n_378;
input n_436;
input n_150;
input n_98;
input n_375;
input n_113;
input n_114;
input n_33;
input n_324;
input n_585;
input n_669;
input n_619;
input n_337;
input n_437;
input n_111;
input n_21;
input n_274;
input n_622;
input n_472;
input n_296;
input n_265;
input n_208;
input n_456;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_615;
input n_521;
input n_51;
input n_496;
input n_76;
input n_342;
input n_26;
input n_246;
input n_517;
input n_530;
input n_0;
input n_428;
input n_159;
input n_358;
input n_105;
input n_580;
input n_608;
input n_30;
input n_494;
input n_131;
input n_263;
input n_434;
input n_360;
input n_563;
input n_229;
input n_394;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_329;
input n_185;
input n_340;
input n_289;
input n_9;
input n_112;
input n_45;
input n_542;
input n_548;
input n_523;
input n_268;
input n_266;
input n_470;
input n_457;
input n_164;
input n_157;
input n_632;
input n_184;
input n_177;
input n_477;
input n_364;
input n_258;
input n_650;
input n_425;
input n_431;
input n_508;
input n_624;
input n_118;
input n_121;
input n_618;
input n_411;
input n_484;
input n_353;
input n_22;
input n_241;
input n_29;
input n_357;
input n_412;
input n_687;
input n_447;
input n_191;
input n_382;
input n_489;
input n_80;
input n_480;
input n_211;
input n_642;
input n_97;
input n_408;
input n_595;
input n_322;
input n_251;
input n_506;
input n_602;
input n_558;
input n_592;
input n_116;
input n_397;
input n_471;
input n_351;
input n_39;
input n_393;
input n_474;
input n_653;
input n_359;
input n_155;
input n_573;
input n_127;
input n_531;
input n_675;

output n_5709;

wire n_2752;
wire n_3527;
wire n_4474;
wire n_4030;
wire n_4770;
wire n_5093;
wire n_3152;
wire n_4586;
wire n_3056;
wire n_3500;
wire n_2679;
wire n_5402;
wire n_2182;
wire n_5553;
wire n_2680;
wire n_3264;
wire n_1250;
wire n_2993;
wire n_4283;
wire n_2879;
wire n_4403;
wire n_4962;
wire n_1430;
wire n_2002;
wire n_1238;
wire n_2729;
wire n_4302;
wire n_4547;
wire n_5090;
wire n_3765;
wire n_864;
wire n_5302;
wire n_1096;
wire n_1379;
wire n_2376;
wire n_2790;
wire n_2207;
wire n_3954;
wire n_4982;
wire n_2042;
wire n_1131;
wire n_5479;
wire n_2646;
wire n_737;
wire n_2653;
wire n_4610;
wire n_3115;
wire n_4028;
wire n_5263;
wire n_5565;
wire n_2482;
wire n_1682;
wire n_958;
wire n_2554;
wire n_4321;
wire n_1985;
wire n_5590;
wire n_2621;
wire n_4853;
wire n_1909;
wire n_5229;
wire n_4260;
wire n_903;
wire n_3348;
wire n_3261;
wire n_1761;
wire n_1690;
wire n_2807;
wire n_1018;
wire n_4512;
wire n_4132;
wire n_1364;
wire n_2390;
wire n_4500;
wire n_2322;
wire n_1107;
wire n_2663;
wire n_5481;
wire n_4824;
wire n_5340;
wire n_3545;
wire n_1428;
wire n_1284;
wire n_4741;
wire n_1241;
wire n_4143;
wire n_4273;
wire n_901;
wire n_4136;
wire n_3144;
wire n_2359;
wire n_1519;
wire n_4567;
wire n_786;
wire n_3552;
wire n_2950;
wire n_3639;
wire n_3254;
wire n_2227;
wire n_2301;
wire n_3121;
wire n_2847;
wire n_5589;
wire n_3015;
wire n_3870;
wire n_3749;
wire n_1676;
wire n_1085;
wire n_5691;
wire n_3482;
wire n_5403;
wire n_823;
wire n_1900;
wire n_4268;
wire n_863;
wire n_3960;
wire n_2433;
wire n_3975;
wire n_899;
wire n_2004;
wire n_4018;
wire n_1495;
wire n_3325;
wire n_4227;
wire n_5158;
wire n_5152;
wire n_1917;
wire n_2456;
wire n_5092;
wire n_1924;
wire n_1811;
wire n_3612;
wire n_4505;
wire n_1840;
wire n_5247;
wire n_5464;
wire n_4476;
wire n_844;
wire n_1267;
wire n_2956;
wire n_5210;
wire n_1213;
wire n_2382;
wire n_780;
wire n_5292;
wire n_1918;
wire n_4119;
wire n_4443;
wire n_4000;
wire n_2686;
wire n_5086;
wire n_1949;
wire n_1140;
wire n_3458;
wire n_3511;
wire n_2077;
wire n_1121;
wire n_3012;
wire n_1947;
wire n_4529;
wire n_3850;
wire n_1216;
wire n_4908;
wire n_3754;
wire n_5060;
wire n_4432;
wire n_2263;
wire n_3518;
wire n_2800;
wire n_2116;
wire n_4530;
wire n_1432;
wire n_2245;
wire n_5614;
wire n_5391;
wire n_5452;
wire n_3359;
wire n_3841;
wire n_5249;
wire n_851;
wire n_3900;
wire n_3413;
wire n_5076;
wire n_3539;
wire n_5062;
wire n_2134;
wire n_3862;
wire n_930;
wire n_4912;
wire n_4226;
wire n_4311;
wire n_3284;
wire n_5046;
wire n_1386;
wire n_3506;
wire n_4827;
wire n_1842;
wire n_4993;
wire n_3678;
wire n_2791;
wire n_1661;
wire n_3212;
wire n_4871;
wire n_3529;
wire n_4405;
wire n_966;
wire n_992;
wire n_3549;
wire n_3914;
wire n_5586;
wire n_1692;
wire n_2611;
wire n_5468;
wire n_3029;
wire n_4745;
wire n_2398;
wire n_4233;
wire n_4791;
wire n_5056;
wire n_1178;
wire n_2015;
wire n_5204;
wire n_2877;
wire n_4951;
wire n_4959;
wire n_3000;
wire n_2930;
wire n_2745;
wire n_2087;
wire n_2161;
wire n_746;
wire n_1357;
wire n_1787;
wire n_1389;
wire n_3172;
wire n_2659;
wire n_4033;
wire n_3747;
wire n_4905;
wire n_4508;
wire n_4045;
wire n_4894;
wire n_3651;
wire n_1812;
wire n_3614;
wire n_959;
wire n_2257;
wire n_1101;
wire n_1343;
wire n_3116;
wire n_4141;
wire n_3784;
wire n_3372;
wire n_3891;
wire n_4422;
wire n_1623;
wire n_3559;
wire n_5179;
wire n_2435;
wire n_5680;
wire n_1932;
wire n_1780;
wire n_2825;
wire n_5685;
wire n_5549;
wire n_1087;
wire n_2388;
wire n_2273;
wire n_1911;
wire n_3496;
wire n_4364;
wire n_3493;
wire n_3700;
wire n_4307;
wire n_2795;
wire n_1841;
wire n_1680;
wire n_2954;
wire n_4438;
wire n_974;
wire n_3814;
wire n_4367;
wire n_5134;
wire n_2467;
wire n_4195;
wire n_5091;
wire n_4866;
wire n_1447;
wire n_1220;
wire n_2019;
wire n_5708;
wire n_698;
wire n_3010;
wire n_2160;
wire n_1992;
wire n_5454;
wire n_1209;
wire n_4254;
wire n_3438;
wire n_2625;
wire n_5373;
wire n_1578;
wire n_3147;
wire n_3661;
wire n_3320;
wire n_4179;
wire n_2144;
wire n_1029;
wire n_2649;
wire n_1247;
wire n_1568;
wire n_2919;
wire n_3108;
wire n_2632;
wire n_5557;
wire n_4314;
wire n_2980;
wire n_1728;
wire n_4315;
wire n_5647;
wire n_3239;
wire n_2631;
wire n_3311;
wire n_3516;
wire n_4442;
wire n_4857;
wire n_1651;
wire n_3087;
wire n_4637;
wire n_5523;
wire n_2697;
wire n_1263;
wire n_1817;
wire n_3704;
wire n_2677;
wire n_4296;
wire n_2483;
wire n_5088;
wire n_1032;
wire n_1592;
wire n_5392;
wire n_4714;
wire n_3074;
wire n_2655;
wire n_3589;
wire n_1743;
wire n_720;
wire n_1943;
wire n_5138;
wire n_4588;
wire n_5149;
wire n_1163;
wire n_3054;
wire n_4970;
wire n_5280;
wire n_4153;
wire n_1868;
wire n_5052;
wire n_3601;
wire n_5137;
wire n_2373;
wire n_3881;
wire n_5089;
wire n_2099;
wire n_3759;
wire n_3323;
wire n_4643;
wire n_2617;
wire n_808;
wire n_2476;
wire n_2814;
wire n_4133;
wire n_2636;
wire n_1439;
wire n_3466;
wire n_2074;
wire n_5031;
wire n_1665;
wire n_2122;
wire n_4543;
wire n_4337;
wire n_5082;
wire n_4788;
wire n_1414;
wire n_2067;
wire n_4555;
wire n_5230;
wire n_1901;
wire n_4486;
wire n_3465;
wire n_2117;
wire n_1053;
wire n_5296;
wire n_5398;
wire n_1906;
wire n_2194;
wire n_4780;
wire n_4640;
wire n_1828;
wire n_1304;
wire n_3335;
wire n_3007;
wire n_2267;
wire n_1349;
wire n_1061;
wire n_2102;
wire n_4157;
wire n_3477;
wire n_3370;
wire n_874;
wire n_3949;
wire n_2286;
wire n_5192;
wire n_4247;
wire n_707;
wire n_5051;
wire n_5336;
wire n_3036;
wire n_2783;
wire n_4583;
wire n_1015;
wire n_1162;
wire n_4292;
wire n_2118;
wire n_1490;
wire n_5552;
wire n_3764;
wire n_1553;
wire n_4773;
wire n_1760;
wire n_5028;
wire n_1086;
wire n_3025;
wire n_3051;
wire n_2802;
wire n_986;
wire n_1104;
wire n_887;
wire n_2125;
wire n_1156;
wire n_4974;
wire n_5123;
wire n_2861;
wire n_4344;
wire n_5242;
wire n_3130;
wire n_1188;
wire n_1498;
wire n_4856;
wire n_2618;
wire n_4216;
wire n_957;
wire n_1242;
wire n_2707;
wire n_5596;
wire n_2849;
wire n_1489;
wire n_2756;
wire n_3781;
wire n_2217;
wire n_4864;
wire n_2226;
wire n_5127;
wire n_4313;
wire n_5255;
wire n_4460;
wire n_4670;
wire n_1119;
wire n_3713;
wire n_1863;
wire n_5536;
wire n_4798;
wire n_1500;
wire n_4946;
wire n_4848;
wire n_4297;
wire n_4941;
wire n_4229;
wire n_5071;
wire n_3337;
wire n_1189;
wire n_3750;
wire n_3424;
wire n_3356;
wire n_1523;
wire n_2190;
wire n_3931;
wire n_2516;
wire n_4991;
wire n_3070;
wire n_1005;
wire n_3275;
wire n_5198;
wire n_3245;
wire n_2894;
wire n_2452;
wire n_4182;
wire n_2827;
wire n_3214;
wire n_3085;
wire n_3373;
wire n_4252;
wire n_5539;
wire n_5009;
wire n_3710;
wire n_1844;
wire n_1957;
wire n_1953;
wire n_1219;
wire n_710;
wire n_3944;
wire n_5632;
wire n_4729;
wire n_1793;
wire n_4446;
wire n_4662;
wire n_5613;
wire n_4800;
wire n_1373;
wire n_1540;
wire n_5427;
wire n_4440;
wire n_1797;
wire n_4425;
wire n_5450;
wire n_832;
wire n_744;
wire n_2821;
wire n_3696;
wire n_1331;
wire n_4781;
wire n_1529;
wire n_3531;
wire n_5124;
wire n_4237;
wire n_5297;
wire n_4828;
wire n_3333;
wire n_4652;
wire n_4114;
wire n_1007;
wire n_1580;
wire n_3135;
wire n_4925;
wire n_2448;
wire n_2211;
wire n_951;
wire n_5318;
wire n_5374;
wire n_2424;
wire n_4697;
wire n_4765;
wire n_5108;
wire n_722;
wire n_3277;
wire n_4863;
wire n_1766;
wire n_5463;
wire n_1338;
wire n_2978;
wire n_4859;
wire n_4568;
wire n_3617;
wire n_704;
wire n_2958;
wire n_1714;
wire n_1044;
wire n_4429;
wire n_5435;
wire n_3340;
wire n_5053;
wire n_5476;
wire n_5483;
wire n_1243;
wire n_5511;
wire n_3486;
wire n_2457;
wire n_2992;
wire n_3197;
wire n_3256;
wire n_1878;
wire n_3646;
wire n_2520;
wire n_811;
wire n_791;
wire n_3864;
wire n_4694;
wire n_1025;
wire n_4664;
wire n_3450;
wire n_4633;
wire n_2026;
wire n_4050;
wire n_3173;
wire n_1406;
wire n_5073;
wire n_4306;
wire n_2684;
wire n_2726;
wire n_4006;
wire n_3266;
wire n_3102;
wire n_1499;
wire n_4288;
wire n_3452;
wire n_4098;
wire n_2691;
wire n_4511;
wire n_3422;
wire n_4675;
wire n_695;
wire n_2991;
wire n_5419;
wire n_1596;
wire n_4289;
wire n_4972;
wire n_2723;
wire n_1476;
wire n_2016;
wire n_3925;
wire n_4689;
wire n_5165;
wire n_2850;
wire n_1874;
wire n_5077;
wire n_3780;
wire n_1657;
wire n_3753;
wire n_1488;
wire n_4846;
wire n_1330;
wire n_906;
wire n_2295;
wire n_5225;
wire n_4076;
wire n_3142;
wire n_3129;
wire n_3495;
wire n_3843;
wire n_4805;
wire n_2606;
wire n_2386;
wire n_4822;
wire n_1829;
wire n_4635;
wire n_1450;
wire n_5532;
wire n_3740;
wire n_5441;
wire n_2417;
wire n_1815;
wire n_1493;
wire n_2911;
wire n_3313;
wire n_2354;
wire n_4281;
wire n_3945;
wire n_3726;
wire n_4419;
wire n_5405;
wire n_1256;
wire n_5365;
wire n_3560;
wire n_3345;
wire n_3421;
wire n_1448;
wire n_1009;
wire n_3548;
wire n_4906;
wire n_4630;
wire n_4829;
wire n_2612;
wire n_5259;
wire n_3236;
wire n_1995;
wire n_1397;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_4966;
wire n_2250;
wire n_1117;
wire n_3321;
wire n_1303;
wire n_4188;
wire n_2001;
wire n_2506;
wire n_2413;
wire n_4825;
wire n_2610;
wire n_3715;
wire n_1593;
wire n_2626;
wire n_2892;
wire n_2605;
wire n_2804;
wire n_5006;
wire n_4882;
wire n_3206;
wire n_1035;
wire n_3475;
wire n_4878;
wire n_2070;
wire n_3842;
wire n_1367;
wire n_4202;
wire n_2044;
wire n_5679;
wire n_3886;
wire n_825;
wire n_732;
wire n_2619;
wire n_1192;
wire n_5141;
wire n_3098;
wire n_4503;
wire n_1291;
wire n_5208;
wire n_5113;
wire n_3987;
wire n_5205;
wire n_4249;
wire n_3160;
wire n_1160;
wire n_2968;
wire n_1882;
wire n_1976;
wire n_2711;
wire n_3223;
wire n_3386;
wire n_3921;
wire n_2177;
wire n_2766;
wire n_4196;
wire n_1197;
wire n_2613;
wire n_5667;
wire n_1517;
wire n_2647;
wire n_5508;
wire n_5105;
wire n_3920;
wire n_3444;
wire n_3851;
wire n_1671;
wire n_5027;
wire n_2343;
wire n_1048;
wire n_775;
wire n_3380;
wire n_5688;
wire n_2826;
wire n_869;
wire n_846;
wire n_1398;
wire n_1921;
wire n_5629;
wire n_2411;
wire n_4631;
wire n_1504;
wire n_2110;
wire n_5377;
wire n_3822;
wire n_889;
wire n_4355;
wire n_3818;
wire n_5599;
wire n_3587;
wire n_2608;
wire n_1948;
wire n_4155;
wire n_810;
wire n_4278;
wire n_4710;
wire n_1959;
wire n_3497;
wire n_4542;
wire n_5451;
wire n_3243;
wire n_4326;
wire n_2121;
wire n_3865;
wire n_5460;
wire n_4685;
wire n_3927;
wire n_2068;
wire n_3595;
wire n_1194;
wire n_4060;
wire n_1647;
wire n_1454;
wire n_2459;
wire n_941;
wire n_3396;
wire n_5517;
wire n_5426;
wire n_4093;
wire n_5693;
wire n_5695;
wire n_4123;
wire n_4294;
wire n_1521;
wire n_1940;
wire n_3683;
wire n_4452;
wire n_3887;
wire n_3195;
wire n_5587;
wire n_4722;
wire n_3048;
wire n_3339;
wire n_4126;
wire n_4164;
wire n_5030;
wire n_2963;
wire n_5674;
wire n_2561;
wire n_1056;
wire n_5584;
wire n_3168;
wire n_5320;
wire n_4079;
wire n_1749;
wire n_1653;
wire n_4088;
wire n_2669;
wire n_3911;
wire n_3802;
wire n_4366;
wire n_1584;
wire n_848;
wire n_5125;
wire n_4922;
wire n_4733;
wire n_1814;
wire n_2441;
wire n_4041;
wire n_2688;
wire n_4208;
wire n_4623;
wire n_4935;
wire n_4509;
wire n_2073;
wire n_4004;
wire n_5238;
wire n_750;
wire n_834;
wire n_3630;
wire n_1612;
wire n_800;
wire n_1910;
wire n_2189;
wire n_4194;
wire n_2018;
wire n_2672;
wire n_2602;
wire n_724;
wire n_2931;
wire n_3433;
wire n_5556;
wire n_3597;
wire n_1956;
wire n_1589;
wire n_4111;
wire n_5633;
wire n_3786;
wire n_875;
wire n_2828;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_4204;
wire n_3553;
wire n_5323;
wire n_3645;
wire n_793;
wire n_5705;
wire n_4996;
wire n_1485;
wire n_2883;
wire n_4411;
wire n_4317;
wire n_3550;
wire n_5510;
wire n_4785;
wire n_2870;
wire n_1494;
wire n_1893;
wire n_1805;
wire n_4068;
wire n_5440;
wire n_2270;
wire n_4163;
wire n_3294;
wire n_2443;
wire n_3610;
wire n_5011;
wire n_1554;
wire n_3279;
wire n_5513;
wire n_972;
wire n_4262;
wire n_2923;
wire n_2843;
wire n_3714;
wire n_4832;
wire n_3676;
wire n_2010;
wire n_5197;
wire n_1679;
wire n_3109;
wire n_1952;
wire n_2394;
wire n_3125;
wire n_5128;
wire n_2356;
wire n_5618;
wire n_4672;
wire n_2564;
wire n_3558;
wire n_3034;
wire n_3502;
wire n_783;
wire n_4053;
wire n_1127;
wire n_1008;
wire n_3963;
wire n_3091;
wire n_1024;
wire n_5157;
wire n_4496;
wire n_2518;
wire n_936;
wire n_4596;
wire n_5178;
wire n_3105;
wire n_1525;
wire n_4628;
wire n_1775;
wire n_908;
wire n_1036;
wire n_4083;
wire n_1270;
wire n_1272;
wire n_2794;
wire n_2901;
wire n_3940;
wire n_3225;
wire n_3621;
wire n_5529;
wire n_3473;
wire n_3680;
wire n_3565;
wire n_5388;
wire n_5354;
wire n_2453;
wire n_3331;
wire n_1788;
wire n_2138;
wire n_3040;
wire n_4230;
wire n_3360;
wire n_1930;
wire n_1809;
wire n_3585;
wire n_1843;
wire n_2000;
wire n_5276;
wire n_4037;
wire n_3804;
wire n_4659;
wire n_3211;
wire n_917;
wire n_5196;
wire n_2096;
wire n_2440;
wire n_2556;
wire n_2215;
wire n_3847;
wire n_4073;
wire n_1261;
wire n_3633;
wire n_857;
wire n_1235;
wire n_2584;
wire n_4001;
wire n_1462;
wire n_5701;
wire n_1064;
wire n_1446;
wire n_1701;
wire n_3111;
wire n_731;
wire n_1813;
wire n_2997;
wire n_1573;
wire n_3258;
wire n_758;
wire n_3691;
wire n_2252;
wire n_1996;
wire n_1106;
wire n_2009;
wire n_784;
wire n_4339;
wire n_4690;
wire n_2987;
wire n_1473;
wire n_1076;
wire n_1348;
wire n_2651;
wire n_753;
wire n_2733;
wire n_2445;
wire n_2103;
wire n_4024;
wire n_4169;
wire n_3316;
wire n_4023;
wire n_4253;
wire n_2522;
wire n_3632;
wire n_1344;
wire n_4064;
wire n_3351;
wire n_5478;
wire n_1141;
wire n_3457;
wire n_5384;
wire n_840;
wire n_2324;
wire n_5283;
wire n_3454;
wire n_2139;
wire n_2521;
wire n_5686;
wire n_2740;
wire n_1991;
wire n_4066;
wire n_4681;
wire n_3303;
wire n_4414;
wire n_2541;
wire n_5094;
wire n_3232;
wire n_1113;
wire n_3768;
wire n_4295;
wire n_1615;
wire n_4100;
wire n_1265;
wire n_2372;
wire n_2105;
wire n_3445;
wire n_1806;
wire n_4087;
wire n_1409;
wire n_1684;
wire n_1588;
wire n_1148;
wire n_1673;
wire n_4473;
wire n_4619;
wire n_5371;
wire n_2290;
wire n_4398;
wire n_5026;
wire n_2856;
wire n_3235;
wire n_5350;
wire n_3265;
wire n_3018;
wire n_1875;
wire n_2429;
wire n_5286;
wire n_4449;
wire n_3285;
wire n_4607;
wire n_1039;
wire n_5676;
wire n_5040;
wire n_1150;
wire n_4266;
wire n_1628;
wire n_2971;
wire n_4407;
wire n_4695;
wire n_1136;
wire n_1190;
wire n_3628;
wire n_4777;
wire n_5243;
wire n_3941;
wire n_1915;
wire n_5399;
wire n_2846;
wire n_3371;
wire n_4918;
wire n_3872;
wire n_4415;
wire n_5110;
wire n_1964;
wire n_3659;
wire n_3928;
wire n_1777;
wire n_3366;
wire n_3441;
wire n_3020;
wire n_4146;
wire n_4947;
wire n_708;
wire n_2545;
wire n_2513;
wire n_4408;
wire n_2115;
wire n_2017;
wire n_1810;
wire n_1347;
wire n_4976;
wire n_860;
wire n_3555;
wire n_3534;
wire n_4548;
wire n_2670;
wire n_3556;
wire n_896;
wire n_4574;
wire n_2644;
wire n_4557;
wire n_3071;
wire n_1698;
wire n_1337;
wire n_774;
wire n_2148;
wire n_5548;
wire n_1168;
wire n_4663;
wire n_3296;
wire n_3794;
wire n_3762;
wire n_4624;
wire n_4963;
wire n_5136;
wire n_4205;
wire n_3293;
wire n_4902;
wire n_1683;
wire n_4686;
wire n_2384;
wire n_1705;
wire n_768;
wire n_3707;
wire n_3895;
wire n_1091;
wire n_3149;
wire n_3934;
wire n_4338;
wire n_2058;
wire n_3231;
wire n_1846;
wire n_4161;
wire n_5304;
wire n_5437;
wire n_1581;
wire n_946;
wire n_757;
wire n_2047;
wire n_3058;
wire n_1655;
wire n_3398;
wire n_3709;
wire n_1146;
wire n_5355;
wire n_998;
wire n_3592;
wire n_5321;
wire n_2536;
wire n_1604;
wire n_3399;
wire n_4772;
wire n_1368;
wire n_963;
wire n_4120;
wire n_925;
wire n_2880;
wire n_1313;
wire n_1001;
wire n_3722;
wire n_4716;
wire n_4654;
wire n_1115;
wire n_1339;
wire n_1051;
wire n_5116;
wire n_3771;
wire n_719;
wire n_3158;
wire n_3221;
wire n_2316;
wire n_1010;
wire n_2830;
wire n_5500;
wire n_4622;
wire n_4757;
wire n_803;
wire n_1871;
wire n_5669;
wire n_5672;
wire n_4016;
wire n_3334;
wire n_5621;
wire n_2940;
wire n_3427;
wire n_3162;
wire n_5569;
wire n_4591;
wire n_5515;
wire n_3083;
wire n_4570;
wire n_2491;
wire n_1931;
wire n_5559;
wire n_2259;
wire n_5337;
wire n_849;
wire n_5059;
wire n_4655;
wire n_1820;
wire n_1233;
wire n_4493;
wire n_1808;
wire n_1635;
wire n_1704;
wire n_4896;
wire n_4851;
wire n_2479;
wire n_886;
wire n_1308;
wire n_1451;
wire n_1487;
wire n_5528;
wire n_5605;
wire n_3432;
wire n_2163;
wire n_1938;
wire n_2484;
wire n_5358;
wire n_1469;
wire n_4901;
wire n_3480;
wire n_1355;
wire n_4213;
wire n_4127;
wire n_2500;
wire n_2334;
wire n_5467;
wire n_1169;
wire n_789;
wire n_3181;
wire n_5493;
wire n_1916;
wire n_4602;
wire n_1713;
wire n_1436;
wire n_2818;
wire n_4900;
wire n_3578;
wire n_1109;
wire n_2537;
wire n_3745;
wire n_3487;
wire n_3668;
wire n_2011;
wire n_1515;
wire n_817;
wire n_1566;
wire n_2837;
wire n_717;
wire n_952;
wire n_2446;
wire n_4116;
wire n_5360;
wire n_2671;
wire n_2702;
wire n_4363;
wire n_3561;
wire n_1839;
wire n_1138;
wire n_4103;
wire n_2529;
wire n_2374;
wire n_5439;
wire n_1225;
wire n_3154;
wire n_1366;
wire n_3938;
wire n_2278;
wire n_1424;
wire n_4736;
wire n_2976;
wire n_4842;
wire n_5250;
wire n_4416;
wire n_4439;
wire n_870;
wire n_4985;
wire n_3382;
wire n_3930;
wire n_3808;
wire n_5471;
wire n_2248;
wire n_813;
wire n_4660;
wire n_3081;
wire n_5497;
wire n_5519;
wire n_995;
wire n_2579;
wire n_1961;
wire n_1535;
wire n_2960;
wire n_3270;
wire n_871;
wire n_2844;
wire n_1979;
wire n_829;
wire n_4814;
wire n_2221;
wire n_5502;
wire n_1283;
wire n_2317;
wire n_2838;
wire n_1736;
wire n_2200;
wire n_2781;
wire n_2442;
wire n_3657;
wire n_5706;
wire n_2634;
wire n_2746;
wire n_5098;
wire n_721;
wire n_1084;
wire n_1276;
wire n_5145;
wire n_2878;
wire n_3830;
wire n_3252;
wire n_5466;
wire n_1528;
wire n_3315;
wire n_3523;
wire n_3999;
wire n_3420;
wire n_3859;
wire n_868;
wire n_5213;
wire n_3474;
wire n_2458;
wire n_5592;
wire n_5620;
wire n_3150;
wire n_5491;
wire n_1542;
wire n_4831;
wire n_4782;
wire n_1539;
wire n_2859;
wire n_5216;
wire n_3412;
wire n_1851;
wire n_2162;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_5703;
wire n_1636;
wire n_4597;
wire n_4546;
wire n_5187;
wire n_4031;
wire n_5119;
wire n_1254;
wire n_4147;
wire n_1703;
wire n_3073;
wire n_3571;
wire n_4576;
wire n_3297;
wire n_5148;
wire n_3003;
wire n_4340;
wire n_3136;
wire n_2867;
wire n_5330;
wire n_2899;
wire n_1560;
wire n_4284;
wire n_3274;
wire n_3877;
wire n_5526;
wire n_5202;
wire n_3817;
wire n_2722;
wire n_3728;
wire n_5107;
wire n_4680;
wire n_5067;
wire n_1012;
wire n_2061;
wire n_2685;
wire n_2512;
wire n_1790;
wire n_2788;
wire n_1443;
wire n_5264;
wire n_2595;
wire n_1465;
wire n_3084;
wire n_705;
wire n_4593;
wire n_4562;
wire n_3860;
wire n_2909;
wire n_3554;
wire n_2717;
wire n_1391;
wire n_2981;
wire n_1006;
wire n_4995;
wire n_1159;
wire n_4498;
wire n_772;
wire n_1245;
wire n_2743;
wire n_1669;
wire n_2969;
wire n_3429;
wire n_1675;
wire n_2466;
wire n_3758;
wire n_5423;
wire n_2568;
wire n_2271;
wire n_2326;
wire n_3485;
wire n_1594;
wire n_4109;
wire n_1935;
wire n_3777;
wire n_1872;
wire n_1585;
wire n_3767;
wire n_3692;
wire n_1351;
wire n_3234;
wire n_2216;
wire n_2426;
wire n_4850;
wire n_1260;
wire n_3716;
wire n_2926;
wire n_4937;
wire n_798;
wire n_5574;
wire n_3391;
wire n_912;
wire n_4786;
wire n_5203;
wire n_4354;
wire n_4235;
wire n_3159;
wire n_2855;
wire n_794;
wire n_2848;
wire n_3306;
wire n_2185;
wire n_4345;
wire n_1292;
wire n_1026;
wire n_3460;
wire n_1610;
wire n_5155;
wire n_2202;
wire n_2952;
wire n_3530;
wire n_2693;
wire n_5408;
wire n_5540;
wire n_3240;
wire n_5066;
wire n_931;
wire n_3362;
wire n_4992;
wire n_4130;
wire n_967;
wire n_5130;
wire n_4175;
wire n_1079;
wire n_5200;
wire n_3393;
wire n_2836;
wire n_2864;
wire n_4456;
wire n_1717;
wire n_2172;
wire n_2601;
wire n_1880;
wire n_2365;
wire n_5684;
wire n_1399;
wire n_1855;
wire n_2333;
wire n_3629;
wire n_4948;
wire n_5413;
wire n_1903;
wire n_2147;
wire n_4020;
wire n_5111;
wire n_5150;
wire n_1226;
wire n_2224;
wire n_1970;
wire n_3724;
wire n_3287;
wire n_2167;
wire n_2293;
wire n_3046;
wire n_2921;
wire n_1240;
wire n_4984;
wire n_4055;
wire n_4410;
wire n_3980;
wire n_5444;
wire n_3257;
wire n_3730;
wire n_5615;
wire n_3979;
wire n_5097;
wire n_2695;
wire n_2598;
wire n_3727;
wire n_976;
wire n_4003;
wire n_1832;
wire n_767;
wire n_2302;
wire n_3014;
wire n_2294;
wire n_2274;
wire n_5640;
wire n_3342;
wire n_2895;
wire n_3796;
wire n_3884;
wire n_4492;
wire n_3625;
wire n_5550;
wire n_3375;
wire n_2768;
wire n_3760;
wire n_5661;
wire n_4975;
wire n_3515;
wire n_2363;
wire n_5306;
wire n_2728;
wire n_2025;
wire n_3744;
wire n_5457;
wire n_5159;
wire n_4022;
wire n_1020;
wire n_2495;
wire n_1058;
wire n_4336;
wire n_5314;
wire n_5231;
wire n_5064;
wire n_2223;
wire n_1279;
wire n_2511;
wire n_3981;
wire n_2681;
wire n_1689;
wire n_2535;
wire n_1255;
wire n_3031;
wire n_2335;
wire n_5482;
wire n_3215;
wire n_1401;
wire n_3138;
wire n_776;
wire n_2860;
wire n_2041;
wire n_1933;
wire n_4494;
wire n_4201;
wire n_5287;
wire n_4719;
wire n_5651;
wire n_3577;
wire n_4074;
wire n_3994;
wire n_4636;
wire n_4983;
wire n_3185;
wire n_1217;
wire n_2662;
wire n_4386;
wire n_3917;
wire n_1231;
wire n_5623;
wire n_5041;
wire n_4275;
wire n_3774;
wire n_5023;
wire n_5524;
wire n_926;
wire n_2296;
wire n_2178;
wire n_4243;
wire n_2765;
wire n_4225;
wire n_4658;
wire n_4186;
wire n_1501;
wire n_2241;
wire n_4699;
wire n_5139;
wire n_4096;
wire n_2531;
wire n_1570;
wire n_3377;
wire n_1518;
wire n_4907;
wire n_3961;
wire n_5153;
wire n_855;
wire n_2059;
wire n_4713;
wire n_1287;
wire n_1611;
wire n_3374;
wire n_4870;
wire n_4818;
wire n_4916;
wire n_4323;
wire n_1899;
wire n_5376;
wire n_3508;
wire n_4129;
wire n_5488;
wire n_1105;
wire n_3599;
wire n_5646;
wire n_4480;
wire n_3734;
wire n_3401;
wire n_983;
wire n_699;
wire n_3542;
wire n_3263;
wire n_2523;
wire n_1945;
wire n_2418;
wire n_1377;
wire n_1614;
wire n_5328;
wire n_3819;
wire n_3222;
wire n_1740;
wire n_4616;
wire n_5016;
wire n_5470;
wire n_1092;
wire n_3205;
wire n_4374;
wire n_2225;
wire n_1963;
wire n_3868;
wire n_729;
wire n_2218;
wire n_1122;
wire n_1408;
wire n_2593;
wire n_1693;
wire n_2741;
wire n_2184;
wire n_2714;
wire n_5362;
wire n_2754;
wire n_4580;
wire n_1218;
wire n_3611;
wire n_5147;
wire n_4826;
wire n_3959;
wire n_3338;
wire n_2962;
wire n_4514;
wire n_1543;
wire n_877;
wire n_3995;
wire n_3908;
wire n_1055;
wire n_1395;
wire n_3892;
wire n_1346;
wire n_1089;
wire n_1502;
wire n_3501;
wire n_1478;
wire n_2555;
wire n_3216;
wire n_3568;
wire n_2708;
wire n_735;
wire n_4844;
wire n_1294;
wire n_4049;
wire n_2661;
wire n_845;
wire n_1649;
wire n_2470;
wire n_1297;
wire n_3551;
wire n_1708;
wire n_5037;
wire n_5650;
wire n_5581;
wire n_4677;
wire n_5189;
wire n_4525;
wire n_3364;
wire n_2643;
wire n_755;
wire n_3766;
wire n_3985;
wire n_5055;
wire n_4369;
wire n_3826;
wire n_5648;
wire n_2266;
wire n_4324;
wire n_842;
wire n_1898;
wire n_1741;
wire n_1907;
wire n_742;
wire n_5160;
wire n_1719;
wire n_2742;
wire n_769;
wire n_3671;
wire n_2366;
wire n_1753;
wire n_5484;
wire n_1372;
wire n_1895;
wire n_4104;
wire n_982;
wire n_3791;
wire n_915;
wire n_2008;
wire n_4989;
wire n_3064;
wire n_3199;
wire n_2127;
wire n_3151;
wire n_3016;
wire n_2460;
wire n_1319;
wire n_3367;
wire n_3669;
wire n_3956;
wire n_4898;
wire n_4081;
wire n_2292;
wire n_2480;
wire n_4528;
wire n_2772;
wire n_1700;
wire n_1332;
wire n_5385;
wire n_1747;
wire n_3990;
wire n_5622;
wire n_1171;
wire n_5635;
wire n_4069;
wire n_3582;
wire n_4280;
wire n_1867;
wire n_5609;
wire n_3993;
wire n_2576;
wire n_3459;
wire n_4811;
wire n_2696;
wire n_5595;
wire n_5256;
wire n_4779;
wire n_2140;
wire n_2157;
wire n_1966;
wire n_5380;
wire n_1400;
wire n_3735;
wire n_1527;
wire n_1513;
wire n_3656;
wire n_4524;
wire n_2831;
wire n_3069;
wire n_4657;
wire n_5568;
wire n_4891;
wire n_2629;
wire n_3369;
wire n_1257;
wire n_1954;
wire n_3964;
wire n_5364;
wire n_3302;
wire n_5597;
wire n_2486;
wire n_1897;
wire n_5469;
wire n_2137;
wire n_3685;
wire n_4977;
wire n_2492;
wire n_2939;
wire n_3425;
wire n_4876;
wire n_5021;
wire n_1449;
wire n_2900;
wire n_797;
wire n_2912;
wire n_1405;
wire n_3813;
wire n_5312;
wire n_2622;
wire n_3447;
wire n_1757;
wire n_1950;
wire n_2264;
wire n_805;
wire n_2032;
wire n_2090;
wire n_3124;
wire n_3811;
wire n_4200;
wire n_2249;
wire n_3411;
wire n_5222;
wire n_3463;
wire n_2785;
wire n_730;
wire n_4938;
wire n_1281;
wire n_2574;
wire n_2364;
wire n_1856;
wire n_1524;
wire n_2928;
wire n_5505;
wire n_1118;
wire n_4604;
wire n_2905;
wire n_2884;
wire n_3408;
wire n_1293;
wire n_961;
wire n_726;
wire n_5504;
wire n_878;
wire n_4118;
wire n_3857;
wire n_3110;
wire n_4239;
wire n_3157;
wire n_1180;
wire n_1697;
wire n_2730;
wire n_5129;
wire n_806;
wire n_1350;
wire n_4704;
wire n_2720;
wire n_1561;
wire n_5494;
wire n_2405;
wire n_2700;
wire n_1616;
wire n_2416;
wire n_2064;
wire n_3640;
wire n_5663;
wire n_5161;
wire n_1557;
wire n_4744;
wire n_5378;
wire n_5626;
wire n_4706;
wire n_2022;
wire n_3879;
wire n_4343;
wire n_1505;
wire n_2408;
wire n_4764;
wire n_5389;
wire n_4990;
wire n_2986;
wire n_949;
wire n_2454;
wire n_3591;
wire n_2760;
wire n_4919;
wire n_1208;
wire n_3317;
wire n_5653;
wire n_4835;
wire n_1151;
wire n_4420;
wire n_2244;
wire n_2143;
wire n_2393;
wire n_4251;
wire n_5266;
wire n_4559;
wire n_4742;
wire n_5038;
wire n_3566;
wire n_1133;
wire n_883;
wire n_4372;
wire n_5396;
wire n_4097;
wire n_4162;
wire n_5293;
wire n_779;
wire n_4790;
wire n_4173;
wire n_5309;
wire n_3573;
wire n_2943;
wire n_3319;
wire n_2247;
wire n_2230;
wire n_1269;
wire n_4727;
wire n_1547;
wire n_1438;
wire n_3654;
wire n_5627;
wire n_1047;
wire n_3783;
wire n_4008;
wire n_2158;
wire n_3643;
wire n_2285;
wire n_3184;
wire n_1288;
wire n_2173;
wire n_3982;
wire n_3647;
wire n_1143;
wire n_3973;
wire n_4799;
wire n_4534;
wire n_5636;
wire n_4960;
wire n_1153;
wire n_1103;
wire n_5707;
wire n_5594;
wire n_3738;
wire n_894;
wire n_5697;
wire n_1380;
wire n_2020;
wire n_5606;
wire n_2310;
wire n_3600;
wire n_1023;
wire n_914;
wire n_5382;
wire n_4327;
wire n_3190;
wire n_3027;
wire n_4011;
wire n_3695;
wire n_3800;
wire n_3462;
wire n_3906;
wire n_3011;
wire n_3395;
wire n_2820;
wire n_3733;
wire n_1165;
wire n_3967;
wire n_4370;
wire n_5638;
wire n_4816;
wire n_4091;
wire n_5058;
wire n_1417;
wire n_3096;
wire n_4166;
wire n_2777;
wire n_5356;
wire n_2234;
wire n_1341;
wire n_3233;
wire n_2431;
wire n_3322;
wire n_1603;
wire n_4478;
wire n_2935;
wire n_4246;
wire n_715;
wire n_1066;
wire n_2863;
wire n_2331;
wire n_4632;
wire n_4061;
wire n_2920;
wire n_1712;
wire n_3344;
wire n_4754;
wire n_1534;
wire n_1290;
wire n_4375;
wire n_2396;
wire n_3368;
wire n_1559;
wire n_3117;
wire n_4684;
wire n_743;
wire n_1546;
wire n_3384;
wire n_5279;
wire n_2592;
wire n_3490;
wire n_962;
wire n_5043;
wire n_4241;
wire n_1622;
wire n_2751;
wire n_3113;
wire n_4183;
wire n_918;
wire n_1968;
wire n_5645;
wire n_5020;
wire n_2842;
wire n_2196;
wire n_3603;
wire n_2371;
wire n_1978;
wire n_3720;
wire n_5232;
wire n_2560;
wire n_4256;
wire n_1164;
wire n_1193;
wire n_1345;
wire n_5035;
wire n_3037;
wire n_1336;
wire n_1033;
wire n_5453;
wire n_4333;
wire n_5339;
wire n_5443;
wire n_1166;
wire n_2007;
wire n_3363;
wire n_1158;
wire n_1803;
wire n_872;
wire n_3522;
wire n_4455;
wire n_3241;
wire n_3899;
wire n_5631;
wire n_3481;
wire n_5101;
wire n_2236;
wire n_692;
wire n_4457;
wire n_2150;
wire n_1816;
wire n_2803;
wire n_2887;
wire n_2648;
wire n_4735;
wire n_3305;
wire n_3810;
wire n_5170;
wire n_4062;
wire n_2093;
wire n_3354;
wire n_5608;
wire n_2204;
wire n_1481;
wire n_2040;
wire n_2151;
wire n_2455;
wire n_827;
wire n_3437;
wire n_2231;
wire n_4212;
wire n_4584;
wire n_5702;
wire n_3574;
wire n_2530;
wire n_2289;
wire n_2299;
wire n_751;
wire n_1027;
wire n_1070;
wire n_2406;
wire n_4477;
wire n_4110;
wire n_5182;
wire n_1221;
wire n_4217;
wire n_5277;
wire n_792;
wire n_1262;
wire n_1942;
wire n_2951;
wire n_3807;
wire n_4048;
wire n_1579;
wire n_4949;
wire n_2181;
wire n_2014;
wire n_2974;
wire n_923;
wire n_1124;
wire n_1326;
wire n_3969;
wire n_2282;
wire n_4605;
wire n_981;
wire n_3873;
wire n_4649;
wire n_1204;
wire n_2428;
wire n_994;
wire n_1360;
wire n_2858;
wire n_3076;
wire n_3410;
wire n_5415;
wire n_856;
wire n_4592;
wire n_4999;
wire n_1564;
wire n_2872;
wire n_3701;
wire n_3706;
wire n_4820;
wire n_1858;
wire n_1678;
wire n_2589;
wire n_4086;
wire n_1482;
wire n_1361;
wire n_4656;
wire n_1520;
wire n_4862;
wire n_5687;
wire n_1411;
wire n_1359;
wire n_3536;
wire n_1721;
wire n_3782;
wire n_1317;
wire n_3594;
wire n_5383;
wire n_2385;
wire n_5690;
wire n_1980;
wire n_4177;
wire n_2501;
wire n_1385;
wire n_1998;
wire n_5029;
wire n_2675;
wire n_2604;
wire n_3521;
wire n_3855;
wire n_2985;
wire n_5218;
wire n_2630;
wire n_2028;
wire n_919;
wire n_3114;
wire n_2092;
wire n_3622;
wire n_2773;
wire n_2817;
wire n_2402;
wire n_1458;
wire n_3047;
wire n_3163;
wire n_5361;
wire n_1550;
wire n_1358;
wire n_1200;
wire n_826;
wire n_5512;
wire n_2808;
wire n_2344;
wire n_3520;
wire n_2392;
wire n_3272;
wire n_3122;
wire n_3687;
wire n_2787;
wire n_5617;
wire n_3799;
wire n_3133;
wire n_2805;
wire n_1268;
wire n_2676;
wire n_2770;
wire n_4550;
wire n_4347;
wire n_702;
wire n_5193;
wire n_4933;
wire n_968;
wire n_4144;
wire n_5514;
wire n_5611;
wire n_2375;
wire n_3278;
wire n_5579;
wire n_4167;
wire n_3608;
wire n_4895;
wire n_1282;
wire n_4726;
wire n_5573;
wire n_5143;
wire n_1755;
wire n_5188;
wire n_5049;
wire n_2212;
wire n_5308;
wire n_4434;
wire n_5068;
wire n_2569;
wire n_4019;
wire n_4199;
wire n_816;
wire n_1322;
wire n_3829;
wire n_4510;
wire n_5057;
wire n_5425;
wire n_5273;
wire n_2469;
wire n_1125;
wire n_2358;
wire n_1710;
wire n_3546;
wire n_2355;
wire n_1390;
wire n_3068;
wire n_1629;
wire n_1094;
wire n_5683;
wire n_1510;
wire n_3002;
wire n_1099;
wire n_5248;
wire n_4899;
wire n_3146;
wire n_3038;
wire n_759;
wire n_4156;
wire n_1727;
wire n_3693;
wire n_3132;
wire n_5002;
wire n_5487;
wire n_5649;
wire n_5531;
wire n_831;
wire n_3681;
wire n_5666;
wire n_3970;
wire n_778;
wire n_2351;
wire n_1619;
wire n_3188;
wire n_4448;
wire n_3218;
wire n_1152;
wire n_2447;
wire n_2101;
wire n_4193;
wire n_1236;
wire n_4579;
wire n_4776;
wire n_2704;
wire n_1334;
wire n_3729;
wire n_4471;
wire n_4392;
wire n_3103;
wire n_2048;
wire n_3028;
wire n_4691;
wire n_3148;
wire n_3775;
wire n_5682;
wire n_5461;
wire n_3966;
wire n_4397;
wire n_3616;
wire n_4753;
wire n_4803;
wire n_1289;
wire n_1831;
wire n_3874;
wire n_2191;
wire n_4165;
wire n_2056;
wire n_2852;
wire n_2515;
wire n_1600;
wire n_1144;
wire n_838;
wire n_1941;
wire n_3637;
wire n_1017;
wire n_734;
wire n_4893;
wire n_2240;
wire n_4258;
wire n_709;
wire n_2917;
wire n_3194;
wire n_2432;
wire n_2085;
wire n_5033;
wire n_1686;
wire n_4232;
wire n_5075;
wire n_2097;
wire n_3461;
wire n_1410;
wire n_939;
wire n_2297;
wire n_4203;
wire n_5400;
wire n_1325;
wire n_1223;
wire n_5347;
wire n_2957;
wire n_1983;
wire n_4767;
wire n_4569;
wire n_948;
wire n_3820;
wire n_5144;
wire n_3072;
wire n_2961;
wire n_4468;
wire n_5509;
wire n_1923;
wire n_3848;
wire n_3631;
wire n_5169;
wire n_4885;
wire n_1479;
wire n_4698;
wire n_1031;
wire n_3674;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_5349;
wire n_3763;
wire n_933;
wire n_3499;
wire n_5534;
wire n_1821;
wire n_3910;
wire n_3947;
wire n_2585;
wire n_5183;
wire n_3361;
wire n_2995;
wire n_4533;
wire n_4287;
wire n_3228;
wire n_2164;
wire n_1732;
wire n_2678;
wire n_1186;
wire n_2052;
wire n_4761;
wire n_4627;
wire n_4556;
wire n_2205;
wire n_2183;
wire n_1724;
wire n_3088;
wire n_1707;
wire n_2080;
wire n_5254;
wire n_3590;
wire n_1126;
wire n_5079;
wire n_2761;
wire n_2357;
wire n_4520;
wire n_895;
wire n_1639;
wire n_2421;
wire n_1302;
wire n_3295;
wire n_3849;
wire n_4263;
wire n_4444;
wire n_5039;
wire n_1818;
wire n_4265;
wire n_3557;
wire n_1598;
wire n_2269;
wire n_1583;
wire n_4612;
wire n_5375;
wire n_5438;
wire n_1264;
wire n_4149;
wire n_1827;
wire n_4958;
wire n_1752;
wire n_2361;
wire n_4538;
wire n_3030;
wire n_3505;
wire n_5563;
wire n_3075;
wire n_1102;
wire n_2239;
wire n_1296;
wire n_4730;
wire n_4421;
wire n_2464;
wire n_3697;
wire n_882;
wire n_2304;
wire n_2514;
wire n_1299;
wire n_3430;
wire n_2063;
wire n_3489;
wire n_5012;
wire n_2079;
wire n_2152;
wire n_4967;
wire n_2517;
wire n_4696;
wire n_3484;
wire n_4971;
wire n_2095;
wire n_5664;
wire n_2738;
wire n_2590;
wire n_4661;
wire n_2797;
wire n_3041;
wire n_1421;
wire n_2208;
wire n_2423;
wire n_5422;
wire n_5246;
wire n_4376;
wire n_3832;
wire n_3525;
wire n_3712;
wire n_4305;
wire n_1069;
wire n_2037;
wire n_2953;
wire n_2823;
wire n_3684;
wire n_5404;
wire n_913;
wire n_1681;
wire n_4834;
wire n_1507;
wire n_5332;
wire n_2866;
wire n_3153;
wire n_1174;
wire n_2346;
wire n_4692;
wire n_1353;
wire n_3268;
wire n_2559;
wire n_5616;
wire n_1383;
wire n_4259;
wire n_2030;
wire n_850;
wire n_4299;
wire n_5625;
wire n_2407;
wire n_5367;
wire n_2243;
wire n_5288;
wire n_2694;
wire n_5601;
wire n_3742;
wire n_4965;
wire n_1837;
wire n_4178;
wire n_2006;
wire n_4953;
wire n_4813;
wire n_3352;
wire n_2367;
wire n_5294;
wire n_5570;
wire n_2731;
wire n_3703;
wire n_5411;
wire n_5670;
wire n_1246;
wire n_5265;
wire n_2123;
wire n_2238;
wire n_4793;
wire n_4802;
wire n_1196;
wire n_3435;
wire n_2380;
wire n_1187;
wire n_4897;
wire n_1298;
wire n_1745;
wire n_4674;
wire n_4796;
wire n_1088;
wire n_766;
wire n_5184;
wire n_2750;
wire n_2547;
wire n_945;
wire n_4575;
wire n_3665;
wire n_3063;
wire n_3281;
wire n_3535;
wire n_5061;
wire n_2288;
wire n_3858;
wire n_4653;
wire n_4589;
wire n_3220;
wire n_4581;
wire n_4625;
wire n_2107;
wire n_5070;
wire n_4845;
wire n_4148;
wire n_3679;
wire n_738;
wire n_5575;
wire n_4968;
wire n_2342;
wire n_4590;
wire n_5177;
wire n_4038;
wire n_3856;
wire n_5316;
wire n_2735;
wire n_953;
wire n_4214;
wire n_1888;
wire n_5290;
wire n_1224;
wire n_2109;
wire n_1425;
wire n_2709;
wire n_3419;
wire n_989;
wire n_5048;
wire n_2233;
wire n_5363;
wire n_5665;
wire n_795;
wire n_4892;
wire n_1936;
wire n_3890;
wire n_821;
wire n_770;
wire n_5607;
wire n_1514;
wire n_2782;
wire n_3929;
wire n_971;
wire n_4353;
wire n_2201;
wire n_4950;
wire n_1650;
wire n_4176;
wire n_4124;
wire n_4431;
wire n_1404;
wire n_3347;
wire n_4797;
wire n_4823;
wire n_5462;
wire n_4488;
wire n_5278;
wire n_2779;
wire n_3627;
wire n_3596;
wire n_5214;
wire n_3756;
wire n_4077;
wire n_3209;
wire n_5220;
wire n_4608;
wire n_3948;
wire n_4839;
wire n_1074;
wire n_1765;
wire n_1977;
wire n_2650;
wire n_4454;
wire n_4184;
wire n_2332;
wire n_2391;
wire n_1295;
wire n_2060;
wire n_3883;
wire n_1013;
wire n_4032;
wire n_2571;
wire n_4929;
wire n_2874;
wire n_4117;
wire n_3049;
wire n_3634;
wire n_5436;
wire n_2341;
wire n_1654;
wire n_3066;
wire n_2045;
wire n_3913;
wire n_5341;
wire n_2575;
wire n_3739;
wire n_1230;
wire n_5140;
wire n_1597;
wire n_2942;
wire n_1771;
wire n_4541;
wire n_3271;
wire n_3164;
wire n_3861;
wire n_5096;
wire n_2043;
wire n_4171;
wire n_4815;
wire n_4665;
wire n_5639;
wire n_4884;
wire n_3580;
wire n_1437;
wire n_4276;
wire n_1378;
wire n_5268;
wire n_5050;
wire n_5240;
wire n_5503;
wire n_1461;
wire n_1876;
wire n_1830;
wire n_5001;
wire n_5658;
wire n_1112;
wire n_700;
wire n_4174;
wire n_5131;
wire n_5546;
wire n_5174;
wire n_2145;
wire n_4801;
wire n_4582;
wire n_4774;
wire n_4108;
wire n_5289;
wire n_3119;
wire n_4740;
wire n_1108;
wire n_1274;
wire n_4394;
wire n_5544;
wire n_5660;
wire n_4920;
wire n_3909;
wire n_4220;
wire n_2703;
wire n_5069;
wire n_5541;
wire n_5610;
wire n_916;
wire n_2810;
wire n_1884;
wire n_1555;
wire n_762;
wire n_1253;
wire n_1468;
wire n_4378;
wire n_5166;
wire n_2683;
wire n_4180;
wire n_4459;
wire n_3624;
wire n_1182;
wire n_4594;
wire n_2748;
wire n_4642;
wire n_1376;
wire n_2925;
wire n_1435;
wire n_1750;
wire n_1506;
wire n_3544;
wire n_5300;
wire n_2072;
wire n_3852;
wire n_5233;
wire n_5381;
wire n_1491;
wire n_2628;
wire n_3219;
wire n_1083;
wire n_5333;
wire n_4914;
wire n_3510;
wire n_4587;
wire n_1139;
wire n_3688;
wire n_5008;
wire n_1312;
wire n_3871;
wire n_892;
wire n_3757;
wire n_1567;
wire n_2219;
wire n_2100;
wire n_3666;
wire n_5538;
wire n_990;
wire n_867;
wire n_3479;
wire n_944;
wire n_5499;
wire n_749;
wire n_2888;
wire n_3998;
wire n_4150;
wire n_1920;
wire n_4285;
wire n_2668;
wire n_2701;
wire n_2400;
wire n_3741;
wire n_5582;
wire n_2567;
wire n_2557;
wire n_1908;
wire n_5675;
wire n_1155;
wire n_2755;
wire n_1071;
wire n_5109;
wire n_712;
wire n_909;
wire n_1392;
wire n_2066;
wire n_5281;
wire n_2762;
wire n_964;
wire n_2220;
wire n_4433;
wire n_2829;
wire n_1914;
wire n_2253;
wire n_2130;
wire n_4861;
wire n_2021;
wire n_1563;
wire n_3673;
wire n_3052;
wire n_2507;
wire n_1633;
wire n_4621;
wire n_3187;
wire n_4451;
wire n_5285;
wire n_2328;
wire n_2434;
wire n_1234;
wire n_3936;
wire n_5564;
wire n_2261;
wire n_3082;
wire n_5162;
wire n_5442;
wire n_2473;
wire n_4784;
wire n_2438;
wire n_3210;
wire n_3867;
wire n_3397;
wire n_1646;
wire n_2262;
wire n_4613;
wire n_2565;
wire n_1237;
wire n_1095;
wire n_3078;
wire n_3971;
wire n_5630;
wire n_5117;
wire n_4979;
wire n_3869;
wire n_1531;
wire n_2113;
wire n_1387;
wire n_3711;
wire n_5054;
wire n_3171;
wire n_5394;
wire n_4751;
wire n_4242;
wire n_1951;
wire n_2490;
wire n_2558;
wire n_1496;
wire n_2812;
wire n_3300;
wire n_5496;
wire n_3104;
wire n_4122;
wire n_2132;
wire n_4522;
wire n_4952;
wire n_4426;
wire n_5699;
wire n_4362;
wire n_3267;
wire n_3946;
wire n_2112;
wire n_2640;
wire n_5000;
wire n_4634;
wire n_4932;
wire n_1795;
wire n_1384;
wire n_2237;
wire n_2983;
wire n_5211;
wire n_4089;
wire n_3513;
wire n_1173;
wire n_3498;
wire n_5132;
wire n_2350;
wire n_5535;
wire n_1068;
wire n_1198;
wire n_4506;
wire n_4728;
wire n_1886;
wire n_4346;
wire n_1648;
wire n_2187;
wire n_1413;
wire n_2481;
wire n_3863;
wire n_2327;
wire n_3882;
wire n_3916;
wire n_1365;
wire n_3968;
wire n_3675;
wire n_2437;
wire n_2841;
wire n_3332;
wire n_2055;
wire n_2998;
wire n_1423;
wire n_4359;
wire n_1609;
wire n_2822;
wire n_1939;
wire n_2308;
wire n_2242;
wire n_4447;
wire n_2937;
wire n_4293;
wire n_5176;
wire n_4039;
wire n_1798;
wire n_3057;
wire n_1608;
wire n_3983;
wire n_703;
wire n_3318;
wire n_3385;
wire n_3773;
wire n_3494;
wire n_1278;
wire n_5074;
wire n_3788;
wire n_3939;
wire n_727;
wire n_3569;
wire n_3837;
wire n_4942;
wire n_3835;
wire n_2496;
wire n_3260;
wire n_3349;
wire n_4348;
wire n_1602;
wire n_3139;
wire n_3801;
wire n_5681;
wire n_2338;
wire n_5261;
wire n_1080;
wire n_3636;
wire n_3653;
wire n_3823;
wire n_3403;
wire n_2057;
wire n_1205;
wire n_2716;
wire n_2944;
wire n_2780;
wire n_3439;
wire n_1120;
wire n_1202;
wire n_4084;
wire n_1371;
wire n_4240;
wire n_2033;
wire n_4121;
wire n_3602;
wire n_2774;
wire n_2799;
wire n_4393;
wire n_3984;
wire n_1586;
wire n_1431;
wire n_4389;
wire n_1763;
wire n_5641;
wire n_4461;
wire n_2763;
wire n_3156;
wire n_1859;
wire n_2660;
wire n_3426;
wire n_4615;
wire n_3044;
wire n_3492;
wire n_3737;
wire n_5657;
wire n_2379;
wire n_3579;
wire n_1667;
wire n_888;
wire n_3896;
wire n_2300;
wire n_4067;
wire n_1677;
wire n_5244;
wire n_5114;
wire n_4551;
wire n_4521;
wire n_2284;
wire n_3005;
wire n_5420;
wire n_2283;
wire n_5206;
wire n_2526;
wire n_1097;
wire n_1711;
wire n_4387;
wire n_2508;
wire n_3186;
wire n_2594;
wire n_1239;
wire n_5298;
wire n_3417;
wire n_890;
wire n_3626;
wire n_4598;
wire n_4464;
wire n_5106;
wire n_4789;
wire n_3180;
wire n_3423;
wire n_1081;
wire n_2119;
wire n_2493;
wire n_5080;
wire n_4565;
wire n_3392;
wire n_1800;
wire n_5081;
wire n_2904;
wire n_3353;
wire n_2946;
wire n_3512;
wire n_1860;
wire n_1734;
wire n_4552;
wire n_2840;
wire n_4482;
wire n_837;
wire n_812;
wire n_4172;
wire n_4040;
wire n_3024;
wire n_5567;
wire n_5406;
wire n_4328;
wire n_1854;
wire n_5191;
wire n_1206;
wire n_1729;
wire n_1508;
wire n_2893;
wire n_4940;
wire n_785;
wire n_3161;
wire n_2389;
wire n_1309;
wire n_999;
wire n_2280;
wire n_1394;
wire n_5085;
wire n_3365;
wire n_4113;
wire n_873;
wire n_3977;
wire n_2468;
wire n_2171;
wire n_4112;
wire n_5602;
wire n_2035;
wire n_4928;
wire n_2614;
wire n_5428;
wire n_2494;
wire n_1538;
wire n_4865;
wire n_2128;
wire n_4071;
wire n_4436;
wire n_3586;
wire n_4160;
wire n_1668;
wire n_4137;
wire n_1078;
wire n_5417;
wire n_4545;
wire n_4758;
wire n_1161;
wire n_4840;
wire n_3097;
wire n_4395;
wire n_4873;
wire n_3507;
wire n_1191;
wire n_4535;
wire n_4385;
wire n_1215;
wire n_3748;
wire n_4731;
wire n_2337;
wire n_1786;
wire n_3732;
wire n_1804;
wire n_4671;
wire n_2272;
wire n_5571;
wire n_4766;
wire n_4558;
wire n_1318;
wire n_1632;
wire n_1769;
wire n_1929;
wire n_4319;
wire n_2929;
wire n_4358;
wire n_1526;
wire n_4874;
wire n_2656;
wire n_4904;
wire n_1997;
wire n_1137;
wire n_1258;
wire n_1733;
wire n_4651;
wire n_943;
wire n_3167;
wire n_4748;
wire n_1807;
wire n_1123;
wire n_2857;
wire n_1784;
wire n_4618;
wire n_3787;
wire n_4025;
wire n_1321;
wire n_3050;
wire n_3919;
wire n_752;
wire n_985;
wire n_5506;
wire n_5475;
wire n_2412;
wire n_3298;
wire n_3107;
wire n_1352;
wire n_5431;
wire n_5100;
wire n_2383;
wire n_2764;
wire n_1822;
wire n_1441;
wire n_5315;
wire n_2633;
wire n_3708;
wire n_2907;
wire n_1429;
wire n_2353;
wire n_2528;
wire n_1778;
wire n_1154;
wire n_4910;
wire n_1759;
wire n_2325;
wire n_4724;
wire n_1130;
wire n_3718;
wire n_756;
wire n_3390;
wire n_2298;
wire n_1016;
wire n_1149;
wire n_4666;
wire n_3140;
wire n_2320;
wire n_4082;
wire n_979;
wire n_3976;
wire n_2813;
wire n_897;
wire n_2546;
wire n_3381;
wire n_3736;
wire n_4466;
wire n_891;
wire n_885;
wire n_1659;
wire n_3955;
wire n_5366;
wire n_5322;
wire n_1864;
wire n_5414;
wire n_3086;
wire n_1887;
wire n_3165;
wire n_3336;
wire n_3635;
wire n_3541;
wire n_2502;
wire n_5151;
wire n_714;
wire n_3605;
wire n_5307;
wire n_2170;
wire n_4721;
wire n_725;
wire n_1577;
wire n_5003;
wire n_3840;
wire n_2198;
wire n_5369;
wire n_3067;
wire n_3809;
wire n_4921;
wire n_1852;
wire n_801;
wire n_4377;
wire n_818;
wire n_2410;
wire n_2314;
wire n_5156;
wire n_5593;
wire n_5270;
wire n_3468;
wire n_1877;
wire n_4301;
wire n_5313;
wire n_2133;
wire n_2497;
wire n_879;
wire n_5446;
wire n_4561;
wire n_3291;
wire n_1541;
wire n_1472;
wire n_1050;
wire n_2578;
wire n_1201;
wire n_2475;
wire n_1185;
wire n_4715;
wire n_2715;
wire n_2665;
wire n_4879;
wire n_5044;
wire n_3755;
wire n_1090;
wire n_4536;
wire n_4304;
wire n_4927;
wire n_4078;
wire n_5459;
wire n_1624;
wire n_1801;
wire n_2854;
wire n_4418;
wire n_3341;
wire n_4125;
wire n_5390;
wire n_5351;
wire n_5267;
wire n_1116;
wire n_5024;
wire n_3043;
wire n_2747;
wire n_1511;
wire n_5275;
wire n_3226;
wire n_3378;
wire n_1641;
wire n_3731;
wire n_4527;
wire n_4291;
wire n_4151;
wire n_2845;
wire n_4412;
wire n_2036;
wire n_843;
wire n_3358;
wire n_2003;
wire n_2533;
wire n_1307;
wire n_4682;
wire n_1128;
wire n_2419;
wire n_2330;
wire n_5078;
wire n_4810;
wire n_3189;
wire n_2309;
wire n_4957;
wire n_4855;
wire n_1955;
wire n_3289;
wire n_1440;
wire n_1370;
wire n_5005;
wire n_1549;
wire n_5207;
wire n_2658;
wire n_5624;
wire n_3620;
wire n_4601;
wire n_1065;
wire n_4518;
wire n_2767;
wire n_5474;
wire n_3376;
wire n_1362;
wire n_3123;
wire n_5447;
wire n_2692;
wire n_1300;
wire n_1960;
wire n_4102;
wire n_4308;
wire n_5700;
wire n_2862;
wire n_4325;
wire n_1420;
wire n_2645;
wire n_2553;
wire n_4711;
wire n_2749;
wire n_4413;
wire n_1210;
wire n_3307;
wire n_1885;
wire n_3251;
wire n_3288;
wire n_2833;
wire n_1038;
wire n_3723;
wire n_4135;
wire n_5223;
wire n_5662;
wire n_3880;
wire n_3904;
wire n_3008;
wire n_4821;
wire n_3242;
wire n_3405;
wire n_2313;
wire n_1022;
wire n_5465;
wire n_3532;
wire n_5154;
wire n_2609;
wire n_1767;
wire n_4138;
wire n_1040;
wire n_3131;
wire n_1973;
wire n_1444;
wire n_820;
wire n_2882;
wire n_2303;
wire n_4384;
wire n_4639;
wire n_1664;
wire n_4577;
wire n_2154;
wire n_1986;
wire n_2624;
wire n_2054;
wire n_1857;
wire n_3926;
wire n_4481;
wire n_984;
wire n_5087;
wire n_1552;
wire n_2938;
wire n_2498;
wire n_3992;
wire n_1772;
wire n_1311;
wire n_3106;
wire n_2881;
wire n_3092;
wire n_4270;
wire n_697;
wire n_4620;
wire n_5397;
wire n_4924;
wire n_4044;
wire n_2305;
wire n_880;
wire n_5566;
wire n_3304;
wire n_4388;
wire n_3247;
wire n_739;
wire n_1028;
wire n_4271;
wire n_2180;
wire n_4406;
wire n_2809;
wire n_5652;
wire n_975;
wire n_1645;
wire n_932;
wire n_2276;
wire n_3301;
wire n_2910;
wire n_2503;
wire n_3785;
wire n_5492;
wire n_2465;
wire n_5501;
wire n_2972;
wire n_4401;
wire n_2586;
wire n_2989;
wire n_3178;
wire n_2251;
wire n_3100;
wire n_3721;
wire n_3389;
wire n_2126;
wire n_2425;
wire n_5692;
wire n_4973;
wire n_4792;
wire n_1601;
wire n_3537;
wire n_4402;
wire n_2487;
wire n_5473;
wire n_1834;
wire n_1011;
wire n_2534;
wire n_2941;
wire n_4286;
wire n_3638;
wire n_3576;
wire n_5562;
wire n_4858;
wire n_1445;
wire n_5370;
wire n_4435;
wire n_3248;
wire n_5317;
wire n_5458;
wire n_2387;
wire n_4318;
wire n_5227;
wire n_830;
wire n_987;
wire n_2510;
wire n_3570;
wire n_3227;
wire n_5359;
wire n_4673;
wire n_2793;
wire n_5282;
wire n_2639;
wire n_4738;
wire n_2603;
wire n_5386;
wire n_1167;
wire n_4554;
wire n_4526;
wire n_4105;
wire n_969;
wire n_3663;
wire n_1663;
wire n_2086;
wire n_1926;
wire n_1630;
wire n_1720;
wire n_2409;
wire n_2966;
wire n_3431;
wire n_3355;
wire n_1738;
wire n_3897;
wire n_1735;
wire n_4005;
wire n_4181;
wire n_2543;
wire n_2321;
wire n_1077;
wire n_2597;
wire n_956;
wire n_765;
wire n_4092;
wire n_4875;
wire n_4255;
wire n_2758;
wire n_5036;
wire n_1271;
wire n_2186;
wire n_4647;
wire n_3575;
wire n_2471;
wire n_3042;
wire n_1067;
wire n_1323;
wire n_1937;
wire n_4142;
wire n_5118;
wire n_900;
wire n_5485;
wire n_5525;
wire n_3004;
wire n_1551;
wire n_4849;
wire n_5271;
wire n_2039;
wire n_1285;
wire n_733;
wire n_761;
wire n_3838;
wire n_4059;
wire n_5194;
wire n_5445;
wire n_2734;
wire n_4499;
wire n_4504;
wire n_3598;
wire n_4917;
wire n_2420;
wire n_3273;
wire n_2918;
wire n_835;
wire n_1865;
wire n_2641;
wire n_2463;
wire n_2580;
wire n_1792;
wire n_5628;
wire n_5245;
wire n_2062;
wire n_4489;
wire n_822;
wire n_1459;
wire n_2153;
wire n_5329;
wire n_5472;
wire n_839;
wire n_1754;
wire n_4833;
wire n_3394;
wire n_2235;
wire n_1575;
wire n_4564;
wire n_1848;
wire n_1172;
wire n_3776;
wire n_2775;
wire n_3903;
wire n_3581;
wire n_5072;
wire n_3778;
wire n_4322;
wire n_2260;
wire n_1660;
wire n_1315;
wire n_4080;
wire n_2206;
wire n_997;
wire n_1643;
wire n_4185;
wire n_1320;
wire n_3001;
wire n_5260;
wire n_4981;
wire n_2347;
wire n_4676;
wire n_2657;
wire n_2990;
wire n_2538;
wire n_2034;
wire n_3932;
wire n_1934;
wire n_2577;
wire n_2362;
wire n_5372;
wire n_4507;
wire n_4756;
wire n_1576;
wire n_2422;
wire n_2933;
wire n_3387;
wire n_3952;
wire n_4365;
wire n_3584;
wire n_4349;
wire n_3446;
wire n_1059;
wire n_2736;
wire n_3825;
wire n_4198;
wire n_977;
wire n_2339;
wire n_2532;
wire n_4373;
wire n_1866;
wire n_2664;
wire n_4154;
wire n_4390;
wire n_1782;
wire n_1558;
wire n_4107;
wire n_2519;
wire n_4380;
wire n_4361;
wire n_4609;
wire n_2360;
wire n_4453;
wire n_723;
wire n_1393;
wire n_4571;
wire n_3137;
wire n_2544;
wire n_809;
wire n_3032;
wire n_5612;
wire n_4886;
wire n_5172;
wire n_881;
wire n_1477;
wire n_1019;
wire n_1982;
wire n_5311;
wire n_910;
wire n_5164;
wire n_4964;
wire n_4700;
wire n_4002;
wire n_1114;
wire n_1742;
wire n_4679;
wire n_3815;
wire n_1768;
wire n_2193;
wire n_2369;
wire n_1199;
wire n_1273;
wire n_2982;
wire n_5495;
wire n_4483;
wire n_3061;
wire n_2587;
wire n_3504;
wire n_5547;
wire n_4693;
wire n_1043;
wire n_5121;
wire n_4956;
wire n_2869;
wire n_5379;
wire n_4487;
wire n_2674;
wire n_1737;
wire n_1613;
wire n_3026;
wire n_2979;
wire n_4329;
wire n_5291;
wire n_4010;
wire n_4501;
wire n_4808;
wire n_3902;
wire n_3244;
wire n_1779;
wire n_2562;
wire n_3112;
wire n_954;
wire n_2051;
wire n_3196;
wire n_2673;
wire n_4678;
wire n_1591;
wire n_5301;
wire n_5126;
wire n_2548;
wire n_3488;
wire n_2381;
wire n_2744;
wire n_1967;
wire n_2179;
wire n_1280;
wire n_3779;
wire n_1063;
wire n_991;
wire n_2275;
wire n_4606;
wire n_3834;
wire n_4303;
wire n_2029;
wire n_1912;
wire n_3923;
wire n_5603;
wire n_938;
wire n_1891;
wire n_5348;
wire n_1000;
wire n_4868;
wire n_4072;
wire n_2792;
wire n_4465;
wire n_2596;
wire n_5217;
wire n_3986;
wire n_5558;
wire n_3725;
wire n_4026;
wire n_4245;
wire n_5520;
wire n_2524;
wire n_3894;
wire n_1702;
wire n_4852;
wire n_3202;
wire n_4290;
wire n_4945;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1082;
wire n_1725;
wire n_5654;
wire n_2318;
wire n_866;
wire n_2819;
wire n_1722;
wire n_2229;
wire n_1644;
wire n_3547;
wire n_4014;
wire n_2551;
wire n_2255;
wire n_5554;
wire n_1252;
wire n_3045;
wire n_773;
wire n_5135;
wire n_4599;
wire n_2706;
wire n_4222;
wire n_718;
wire n_1434;
wire n_1905;
wire n_1569;
wire n_5448;
wire n_2573;
wire n_2336;
wire n_5412;
wire n_1662;
wire n_3249;
wire n_3483;
wire n_4046;
wire n_4701;
wire n_1925;
wire n_782;
wire n_2915;
wire n_4869;
wire n_3213;
wire n_5533;
wire n_4047;
wire n_1244;
wire n_1796;
wire n_2719;
wire n_2876;
wire n_4063;
wire n_5224;
wire n_2778;
wire n_1574;
wire n_3033;
wire n_893;
wire n_1582;
wire n_1981;
wire n_2824;
wire n_5327;
wire n_4417;
wire n_796;
wire n_1374;
wire n_2089;
wire n_4688;
wire n_4939;
wire n_1486;
wire n_3619;
wire n_4013;
wire n_3434;
wire n_4342;
wire n_691;
wire n_4903;
wire n_2131;
wire n_3853;
wire n_4382;
wire n_2509;
wire n_4085;
wire n_5486;
wire n_2135;
wire n_4475;
wire n_5432;
wire n_1463;
wire n_4626;
wire n_4997;
wire n_5065;
wire n_924;
wire n_781;
wire n_2013;
wire n_4638;
wire n_2786;
wire n_4058;
wire n_4090;
wire n_4819;
wire n_2436;
wire n_3517;
wire n_1706;
wire n_2461;
wire n_3719;
wire n_1214;
wire n_3526;
wire n_3888;
wire n_3198;
wire n_1853;
wire n_764;
wire n_1503;
wire n_5295;
wire n_1181;
wire n_1999;
wire n_4841;
wire n_4683;
wire n_5173;
wire n_2873;
wire n_2084;
wire n_3330;
wire n_3514;
wire n_5655;
wire n_3383;
wire n_1835;
wire n_3965;
wire n_1457;
wire n_3905;
wire n_3797;
wire n_1836;
wire n_3416;
wire n_4600;
wire n_1453;
wire n_3943;
wire n_3145;
wire n_2908;
wire n_4106;
wire n_2156;
wire n_1184;
wire n_754;
wire n_2323;
wire n_1073;
wire n_4549;
wire n_1277;
wire n_1746;
wire n_1062;
wire n_4702;
wire n_5102;
wire n_4954;
wire n_740;
wire n_1974;
wire n_4491;
wire n_2906;
wire n_3283;
wire n_4331;
wire n_4159;
wire n_3451;
wire n_4734;
wire n_2832;
wire n_1688;
wire n_2370;
wire n_1944;
wire n_2914;
wire n_5656;
wire n_1988;
wire n_5678;
wire n_1718;
wire n_4515;
wire n_2149;
wire n_2277;
wire n_2539;
wire n_5555;
wire n_2078;
wire n_1145;
wire n_4809;
wire n_787;
wire n_4012;
wire n_1195;
wire n_2049;
wire n_1522;
wire n_5212;
wire n_4760;
wire n_1207;
wire n_3606;
wire n_2232;
wire n_1847;
wire n_4320;
wire n_5084;
wire n_5251;
wire n_1314;
wire n_1512;
wire n_884;
wire n_4980;
wire n_3324;
wire n_2192;
wire n_5407;
wire n_2988;
wire n_4560;
wire n_3230;
wire n_3793;
wire n_859;
wire n_5042;
wire n_4768;
wire n_1889;
wire n_693;
wire n_5368;
wire n_929;
wire n_3207;
wire n_3641;
wire n_3828;
wire n_1850;
wire n_3183;
wire n_3607;
wire n_1637;
wire n_2427;
wire n_3613;
wire n_2885;
wire n_2098;
wire n_2616;
wire n_1751;
wire n_5310;
wire n_2769;
wire n_1548;
wire n_4987;
wire n_3013;
wire n_4572;
wire n_1396;
wire n_2739;
wire n_3962;
wire n_4988;
wire n_2902;
wire n_4360;
wire n_1544;
wire n_4540;
wire n_2094;
wire n_5588;
wire n_3854;
wire n_1354;
wire n_2349;
wire n_3652;
wire n_3449;
wire n_1021;
wire n_3089;
wire n_4854;
wire n_1595;
wire n_1142;
wire n_5477;
wire n_2727;
wire n_942;
wire n_5234;
wire n_1416;
wire n_1599;
wire n_4747;
wire n_3472;
wire n_2527;
wire n_3126;
wire n_2759;
wire n_5007;
wire n_4881;
wire n_2038;
wire n_3958;
wire n_4495;
wire n_4737;
wire n_1838;
wire n_4357;
wire n_2806;
wire n_4502;
wire n_3191;
wire n_1716;
wire n_5334;
wire n_3562;
wire n_2281;
wire n_5253;
wire n_3588;
wire n_1590;
wire n_3280;
wire n_4115;
wire n_5274;
wire n_5418;
wire n_5019;
wire n_1819;
wire n_3095;
wire n_947;
wire n_3698;
wire n_4513;
wire n_1179;
wire n_696;
wire n_1442;
wire n_4775;
wire n_2620;
wire n_1833;
wire n_1691;
wire n_2549;
wire n_2499;
wire n_804;
wire n_1656;
wire n_1382;
wire n_3093;
wire n_2970;
wire n_3885;
wire n_955;
wire n_4264;
wire n_2166;
wire n_3192;
wire n_4709;
wire n_1562;
wire n_3250;
wire n_4223;
wire n_3538;
wire n_3915;
wire n_3839;
wire n_5490;
wire n_5694;
wire n_1972;
wire n_4718;
wire n_3717;
wire n_5489;
wire n_3407;
wire n_3875;
wire n_4029;
wire n_4206;
wire n_2415;
wire n_4099;
wire n_3120;
wire n_2922;
wire n_3193;
wire n_2871;
wire n_5342;
wire n_4794;
wire n_4843;
wire n_5580;
wire n_5215;
wire n_3937;
wire n_4763;
wire n_1418;
wire n_4170;
wire n_5561;
wire n_2462;
wire n_2155;
wire n_2439;
wire n_4838;
wire n_4795;
wire n_3604;
wire n_5430;
wire n_824;
wire n_5659;
wire n_4272;
wire n_5195;
wire n_3176;
wire n_3792;
wire n_4267;
wire n_2083;
wire n_815;
wire n_5598;
wire n_2753;
wire n_1340;
wire n_3021;
wire n_4352;
wire n_2712;
wire n_1433;
wire n_3805;
wire n_3912;
wire n_3950;
wire n_2898;
wire n_1825;
wire n_3567;
wire n_2682;
wire n_5585;
wire n_5112;
wire n_5326;
wire n_1627;
wire n_2903;
wire n_5303;
wire n_3812;
wire n_3127;
wire n_1731;
wire n_799;
wire n_1147;
wire n_2378;
wire n_5530;
wire n_965;
wire n_934;
wire n_2213;
wire n_4056;
wire n_4806;
wire n_1674;
wire n_4015;
wire n_2924;
wire n_4445;
wire n_4462;
wire n_5299;
wire n_4219;
wire n_4484;
wire n_4723;
wire n_2142;
wire n_4517;
wire n_2896;
wire n_1913;
wire n_2069;
wire n_4043;
wire n_1042;
wire n_3170;
wire n_2311;
wire n_1455;
wire n_2287;
wire n_836;
wire n_3415;
wire n_3464;
wire n_3414;
wire n_4234;
wire n_760;
wire n_1483;
wire n_1363;
wire n_1111;
wire n_970;
wire n_3467;
wire n_713;
wire n_3179;
wire n_5522;
wire n_4836;
wire n_3889;
wire n_5262;
wire n_3262;
wire n_5319;
wire n_927;
wire n_3699;
wire n_706;
wire n_2120;
wire n_1419;
wire n_3816;
wire n_3528;
wire n_4207;
wire n_2404;
wire n_2168;
wire n_2757;
wire n_4725;
wire n_2312;
wire n_1826;
wire n_4880;
wire n_2834;
wire n_4051;
wire n_3660;
wire n_4563;
wire n_2996;
wire n_5335;
wire n_1259;
wire n_2801;
wire n_1177;
wire n_4334;
wire n_5284;
wire n_4978;
wire n_3246;
wire n_3299;
wire n_980;
wire n_1618;
wire n_1869;
wire n_3623;
wire n_905;
wire n_2718;
wire n_4707;
wire n_2687;
wire n_4923;
wire n_4911;
wire n_3876;
wire n_5516;
wire n_3615;
wire n_1802;
wire n_2811;
wire n_3019;
wire n_5168;
wire n_3200;
wire n_3642;
wire n_2146;
wire n_4274;
wire n_5583;
wire n_3276;
wire n_5433;
wire n_3682;
wire n_5429;
wire n_5698;
wire n_4007;
wire n_1456;
wire n_1879;
wire n_2129;
wire n_814;
wire n_5120;
wire n_3572;
wire n_2975;
wire n_2399;
wire n_1134;
wire n_3471;
wire n_4075;
wire n_1484;
wire n_2027;
wire n_2932;
wire n_3118;
wire n_5560;
wire n_4441;
wire n_3039;
wire n_3922;
wire n_2195;
wire n_5455;
wire n_1467;
wire n_5209;
wire n_5704;
wire n_4458;
wire n_2159;
wire n_4889;
wire n_3831;
wire n_1744;
wire n_4523;
wire n_3618;
wire n_3705;
wire n_3022;
wire n_1709;
wire n_5099;
wire n_3286;
wire n_5619;
wire n_2023;
wire n_3974;
wire n_3443;
wire n_2599;
wire n_3988;
wire n_5022;
wire n_2075;
wire n_1726;
wire n_2031;
wire n_3761;
wire n_3996;
wire n_5353;
wire n_4771;
wire n_2853;
wire n_3350;
wire n_1098;
wire n_3009;
wire n_777;
wire n_5219;
wire n_920;
wire n_3951;
wire n_5518;
wire n_3035;
wire n_4261;
wire n_1132;
wire n_1823;
wire n_5236;
wire n_4236;
wire n_3942;
wire n_3023;
wire n_2254;
wire n_3290;
wire n_1402;
wire n_3957;
wire n_3418;
wire n_1607;
wire n_5673;
wire n_861;
wire n_1666;
wire n_5103;
wire n_4648;
wire n_2214;
wire n_2256;
wire n_3326;
wire n_2732;
wire n_1883;
wire n_4094;
wire n_2776;
wire n_3224;
wire n_1969;
wire n_5671;
wire n_2949;
wire n_4269;
wire n_1927;
wire n_1222;
wire n_3803;
wire n_5239;
wire n_1919;
wire n_2994;
wire n_1791;
wire n_2124;
wire n_1894;
wire n_1460;
wire n_4913;
wire n_2449;
wire n_4428;
wire n_745;
wire n_1572;
wire n_4463;
wire n_5357;
wire n_3648;
wire n_1975;
wire n_5421;
wire n_1388;
wire n_1266;
wire n_4396;
wire n_1990;
wire n_3491;
wire n_2690;
wire n_3090;
wire n_2474;
wire n_2623;
wire n_1075;
wire n_1890;
wire n_4034;
wire n_4228;
wire n_1227;
wire n_3166;
wire n_3649;
wire n_3065;
wire n_5045;
wire n_5237;
wire n_3924;
wire n_3997;
wire n_3564;
wire n_862;
wire n_2637;
wire n_3795;
wire n_4931;
wire n_2306;
wire n_2071;
wire n_3953;
wire n_4400;
wire n_2414;
wire n_2082;
wire n_2959;
wire n_5434;
wire n_1532;
wire n_1030;
wire n_5181;
wire n_3208;
wire n_1342;
wire n_2737;
wire n_3282;
wire n_852;
wire n_2916;
wire n_1060;
wire n_4424;
wire n_4351;
wire n_4192;
wire n_1748;
wire n_1301;
wire n_3400;
wire n_1466;
wire n_2581;
wire n_1783;
wire n_5146;
wire n_4646;
wire n_4221;
wire n_1037;
wire n_3650;
wire n_1329;
wire n_1993;
wire n_1545;
wire n_4035;
wire n_1480;
wire n_3670;
wire n_2540;
wire n_4190;
wire n_1605;
wire n_3060;
wire n_2984;
wire n_4009;
wire n_2489;
wire n_5013;
wire n_4145;
wire n_5577;
wire n_876;
wire n_5017;
wire n_736;
wire n_2265;
wire n_3524;
wire n_2627;
wire n_1327;
wire n_1475;
wire n_2106;
wire n_4717;
wire n_4739;
wire n_3174;
wire n_3314;
wire n_854;
wire n_2091;
wire n_4312;
wire n_5424;
wire n_3789;
wire n_1658;
wire n_1072;
wire n_1305;
wire n_4750;
wire n_2348;
wire n_1873;
wire n_2667;
wire n_2725;
wire n_3746;
wire n_4537;
wire n_1046;
wire n_3694;
wire n_771;
wire n_5456;
wire n_3893;
wire n_4847;
wire n_2307;
wire n_3702;
wire n_1984;
wire n_3453;
wire n_1556;
wire n_5345;
wire n_2815;
wire n_4427;
wire n_1824;
wire n_1492;
wire n_4065;
wire n_4705;
wire n_819;
wire n_1971;
wire n_2945;
wire n_3543;
wire n_1324;
wire n_1776;
wire n_3448;
wire n_4279;
wire n_2936;
wire n_3609;
wire n_4330;
wire n_4152;
wire n_5537;
wire n_2698;
wire n_5572;
wire n_4783;
wire n_3017;
wire n_2329;
wire n_2570;
wire n_1642;
wire n_2789;
wire n_5409;
wire n_2525;
wire n_2890;
wire n_4539;
wire n_3455;
wire n_807;
wire n_5142;
wire n_3907;
wire n_4603;
wire n_5010;
wire n_4332;
wire n_1987;
wire n_4052;
wire n_3357;
wire n_3388;
wire n_2368;
wire n_802;
wire n_5401;
wire n_4595;
wire n_960;
wire n_2352;
wire n_5201;
wire n_790;
wire n_5551;
wire n_5416;
wire n_4404;
wire n_2377;
wire n_2652;
wire n_5498;
wire n_5543;
wire n_4054;
wire n_1286;
wire n_4617;
wire n_1685;
wire n_2477;
wire n_4611;
wire n_2279;
wire n_3169;
wire n_2222;
wire n_1052;
wire n_4732;
wire n_2203;
wire n_2076;
wire n_1426;
wire n_4969;
wire n_5252;
wire n_4641;
wire n_5063;
wire n_4399;
wire n_4140;
wire n_5171;
wire n_2607;
wire n_3343;
wire n_4712;
wire n_3309;
wire n_2796;
wire n_858;
wire n_5393;
wire n_4817;
wire n_2136;
wire n_3134;
wire n_4909;
wire n_4755;
wire n_2771;
wire n_2403;
wire n_2947;
wire n_5643;
wire n_928;
wire n_3769;
wire n_1565;
wire n_4437;
wire n_3055;
wire n_4070;
wire n_5346;
wire n_748;
wire n_1045;
wire n_1881;
wire n_2635;
wire n_2999;
wire n_988;
wire n_4139;
wire n_4769;
wire n_1958;
wire n_4867;
wire n_3667;
wire n_2713;
wire n_1422;
wire n_1965;
wire n_5167;
wire n_5257;
wire n_4450;
wire n_2934;
wire n_5104;
wire n_2210;
wire n_4368;
wire n_3141;
wire n_2053;
wire n_5272;
wire n_3476;
wire n_1049;
wire n_4430;
wire n_3238;
wire n_2450;
wire n_5338;
wire n_1356;
wire n_1773;
wire n_3175;
wire n_4544;
wire n_2666;
wire n_5578;
wire n_728;
wire n_4191;
wire n_4409;
wire n_2401;
wire n_3255;
wire n_2588;
wire n_935;
wire n_2886;
wire n_4961;
wire n_3827;
wire n_2478;
wire n_911;
wire n_3509;
wire n_1403;
wire n_5395;
wire n_3006;
wire n_4531;
wire n_3770;
wire n_3456;
wire n_4532;
wire n_3790;
wire n_907;
wire n_847;
wire n_747;
wire n_1135;
wire n_2566;
wire n_5095;
wire n_3101;
wire n_3662;
wire n_5199;
wire n_4257;
wire n_4282;
wire n_4341;
wire n_1694;
wire n_1695;
wire n_4027;
wire n_4309;
wire n_4650;
wire n_5480;
wire n_3077;
wire n_4944;
wire n_3478;
wire n_3062;
wire n_1774;
wire n_4994;
wire n_3533;
wire n_5175;
wire n_1994;
wire n_3978;
wire n_3836;
wire n_3409;
wire n_4381;
wire n_3583;
wire n_4316;
wire n_4860;
wire n_4469;
wire n_3540;
wire n_4930;
wire n_5352;
wire n_1157;
wire n_3563;
wire n_1739;
wire n_2642;
wire n_3310;
wire n_4423;
wire n_3689;
wire n_1789;
wire n_763;
wire n_2174;
wire n_5668;
wire n_3442;
wire n_3972;
wire n_2315;
wire n_4209;
wire n_4703;
wire n_1687;
wire n_4934;
wire n_2638;
wire n_2046;
wire n_1756;
wire n_4350;
wire n_1606;
wire n_5600;
wire n_1587;
wire n_2340;
wire n_4804;
wire n_2444;
wire n_4888;
wire n_1014;
wire n_1427;
wire n_2977;
wire n_3991;
wire n_4936;
wire n_2199;
wire n_4669;
wire n_5228;
wire n_1100;
wire n_1617;
wire n_2600;
wire n_3436;
wire n_1962;
wire n_3806;
wire n_4759;
wire n_2114;
wire n_3329;
wire n_2927;
wire n_3833;
wire n_1175;
wire n_4887;
wire n_3751;
wire n_3402;
wire n_1621;
wire n_5186;
wire n_4585;
wire n_1785;
wire n_3406;
wire n_3664;
wire n_4218;
wire n_4687;
wire n_1381;
wire n_3686;
wire n_1183;
wire n_4720;
wire n_2889;
wire n_2141;
wire n_1758;
wire n_1110;
wire n_5604;
wire n_3470;
wire n_5221;
wire n_1407;
wire n_2865;
wire n_973;
wire n_5591;
wire n_4762;
wire n_3844;
wire n_3259;
wire n_2572;
wire n_4490;
wire n_1248;
wire n_1176;
wire n_3677;
wire n_1054;
wire n_5387;
wire n_3292;
wire n_3989;
wire n_4644;
wire n_4752;
wire n_4746;
wire n_1057;
wire n_4131;
wire n_5449;
wire n_4215;
wire n_978;
wire n_2488;
wire n_1509;
wire n_828;
wire n_4158;
wire n_3079;
wire n_5190;
wire n_3269;
wire n_5325;
wire n_4231;
wire n_5047;
wire n_2591;
wire n_5004;
wire n_4926;
wire n_2050;
wire n_2197;
wire n_4872;
wire n_4778;
wire n_5344;
wire n_2550;
wire n_1536;
wire n_3177;
wire n_4667;
wire n_1471;
wire n_3440;
wire n_3658;
wire n_3404;
wire n_2291;
wire n_3346;
wire n_2816;
wire n_1620;
wire n_2542;
wire n_2165;
wire n_4837;
wire n_4210;
wire n_788;
wire n_2169;
wire n_5634;
wire n_5133;
wire n_5305;
wire n_2175;
wire n_1625;
wire n_5689;
wire n_4578;
wire n_5644;
wire n_3644;
wire n_2176;
wire n_1412;
wire n_3059;
wire n_1922;
wire n_940;
wire n_1537;
wire n_4877;
wire n_2065;
wire n_4470;
wire n_4187;
wire n_1904;
wire n_4998;
wire n_5576;
wire n_2395;
wire n_2868;
wire n_1530;
wire n_4057;
wire n_1170;
wire n_2724;
wire n_2258;
wire n_898;
wire n_3328;
wire n_2012;
wire n_3182;
wire n_2967;
wire n_5343;
wire n_1093;
wire n_4021;
wire n_3379;
wire n_4379;
wire n_2268;
wire n_3469;
wire n_1452;
wire n_2835;
wire n_2111;
wire n_3743;
wire n_5542;
wire n_2948;
wire n_5015;
wire n_3099;
wire n_5527;
wire n_2897;
wire n_4812;
wire n_4497;
wire n_2583;
wire n_3155;
wire n_4300;
wire n_2024;
wire n_1770;
wire n_701;
wire n_1003;
wire n_4472;
wire n_2699;
wire n_3901;
wire n_5180;
wire n_1640;
wire n_2973;
wire n_2710;
wire n_2505;
wire n_4519;
wire n_5025;
wire n_2397;
wire n_3878;
wire n_4197;
wire n_2721;
wire n_1892;
wire n_2615;
wire n_4787;
wire n_1212;
wire n_4310;
wire n_4566;
wire n_3933;
wire n_4371;
wire n_1902;
wire n_2784;
wire n_3898;
wire n_694;
wire n_4749;
wire n_1845;
wire n_921;
wire n_5545;
wire n_2104;
wire n_2552;
wire n_1470;
wire n_1533;
wire n_5083;
wire n_3253;
wire n_2088;
wire n_1275;
wire n_4238;
wire n_904;
wire n_2005;
wire n_1696;
wire n_2108;
wire n_3824;
wire n_2246;
wire n_3846;
wire n_5122;
wire n_1497;
wire n_4189;
wire n_2472;
wire n_2705;
wire n_4479;
wire n_3845;
wire n_3203;
wire n_4986;
wire n_1316;
wire n_4668;
wire n_950;
wire n_711;
wire n_4168;
wire n_1369;
wire n_4298;
wire n_4743;
wire n_1781;
wire n_4250;
wire n_3143;
wire n_3690;
wire n_3229;
wire n_2188;
wire n_2430;
wire n_2504;
wire n_5637;
wire n_4211;
wire n_3094;
wire n_741;
wire n_5185;
wire n_2964;
wire n_5032;
wire n_865;
wire n_5034;
wire n_3312;
wire n_1041;
wire n_2451;
wire n_2913;
wire n_993;
wire n_1862;
wire n_3752;
wire n_3672;
wire n_922;
wire n_1004;
wire n_2839;
wire n_3237;
wire n_4128;
wire n_4036;
wire n_5269;
wire n_3655;
wire n_2955;
wire n_1764;
wire n_4807;
wire n_5115;
wire n_902;
wire n_1723;
wire n_3918;
wire n_5324;
wire n_4101;
wire n_4915;
wire n_3866;
wire n_1946;
wire n_4383;
wire n_4830;
wire n_4391;
wire n_4095;
wire n_1310;
wire n_4485;
wire n_3593;
wire n_5163;
wire n_1229;
wire n_2582;
wire n_3327;
wire n_4356;
wire n_1896;
wire n_1516;
wire n_4890;
wire n_2485;
wire n_2563;
wire n_4224;
wire n_1670;
wire n_1799;
wire n_5507;
wire n_4573;
wire n_1328;
wire n_4943;
wire n_2875;
wire n_3519;
wire n_2209;
wire n_4042;
wire n_4244;
wire n_1928;
wire n_5642;
wire n_4708;
wire n_4883;
wire n_4553;
wire n_1634;
wire n_1203;
wire n_1699;
wire n_5226;
wire n_2081;
wire n_937;
wire n_1474;
wire n_1631;
wire n_1794;
wire n_5696;
wire n_1375;
wire n_3053;
wire n_5014;
wire n_3772;
wire n_2891;
wire n_4335;
wire n_3128;
wire n_5677;
wire n_4277;
wire n_4614;
wire n_4629;
wire n_1002;
wire n_4516;
wire n_5235;
wire n_1129;
wire n_1464;
wire n_2798;
wire n_3217;
wire n_1249;
wire n_3821;
wire n_3201;
wire n_3503;
wire n_1870;
wire n_4467;
wire n_5521;
wire n_2654;
wire n_3935;
wire n_1861;
wire n_1228;
wire n_2319;
wire n_2965;
wire n_4955;
wire n_5410;
wire n_1251;
wire n_1989;
wire n_2689;
wire n_1762;
wire n_3798;
wire n_3080;
wire n_5241;
wire n_4248;
wire n_1672;
wire n_2228;
wire n_4645;
wire n_5331;
wire n_3308;
wire n_841;
wire n_3204;
wire n_4134;
wire n_5018;
wire n_3428;
wire n_2851;
wire n_4017;
wire n_2345;
wire n_1730;
wire n_5258;

CKINVDCx5p33_ASAP7_75t_R g691 ( 
.A(n_449),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_616),
.Y(n_692)
);

CKINVDCx5p33_ASAP7_75t_R g693 ( 
.A(n_88),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_329),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_14),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_49),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_309),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_539),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_278),
.Y(n_699)
);

BUFx3_ASAP7_75t_L g700 ( 
.A(n_300),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_411),
.Y(n_701)
);

CKINVDCx20_ASAP7_75t_R g702 ( 
.A(n_292),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_425),
.Y(n_703)
);

CKINVDCx20_ASAP7_75t_R g704 ( 
.A(n_113),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_84),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_275),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_626),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_478),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_638),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_489),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_276),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_123),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_688),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_319),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_566),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_188),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_296),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_627),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_151),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_281),
.Y(n_720)
);

CKINVDCx5p33_ASAP7_75t_R g721 ( 
.A(n_35),
.Y(n_721)
);

CKINVDCx20_ASAP7_75t_R g722 ( 
.A(n_370),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_642),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_35),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_492),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_331),
.Y(n_726)
);

CKINVDCx14_ASAP7_75t_R g727 ( 
.A(n_566),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_139),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_680),
.Y(n_729)
);

INVx2_ASAP7_75t_L g730 ( 
.A(n_321),
.Y(n_730)
);

CKINVDCx5p33_ASAP7_75t_R g731 ( 
.A(n_227),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_209),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_648),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_349),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_308),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_27),
.Y(n_736)
);

CKINVDCx20_ASAP7_75t_R g737 ( 
.A(n_240),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_674),
.Y(n_738)
);

CKINVDCx5p33_ASAP7_75t_R g739 ( 
.A(n_91),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_129),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_123),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_127),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_157),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_449),
.Y(n_744)
);

CKINVDCx20_ASAP7_75t_R g745 ( 
.A(n_626),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_531),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_410),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_621),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_19),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_110),
.Y(n_750)
);

BUFx2_ASAP7_75t_SL g751 ( 
.A(n_641),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_579),
.Y(n_752)
);

CKINVDCx20_ASAP7_75t_R g753 ( 
.A(n_111),
.Y(n_753)
);

CKINVDCx5p33_ASAP7_75t_R g754 ( 
.A(n_90),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_359),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_480),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_668),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_466),
.Y(n_758)
);

CKINVDCx5p33_ASAP7_75t_R g759 ( 
.A(n_38),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_91),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_76),
.Y(n_761)
);

CKINVDCx20_ASAP7_75t_R g762 ( 
.A(n_439),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_564),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_434),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_317),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_511),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_247),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_628),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_75),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_54),
.Y(n_770)
);

CKINVDCx5p33_ASAP7_75t_R g771 ( 
.A(n_343),
.Y(n_771)
);

BUFx2_ASAP7_75t_SL g772 ( 
.A(n_110),
.Y(n_772)
);

CKINVDCx5p33_ASAP7_75t_R g773 ( 
.A(n_673),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_527),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_412),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_265),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_597),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_307),
.Y(n_778)
);

INVx3_ASAP7_75t_L g779 ( 
.A(n_300),
.Y(n_779)
);

CKINVDCx20_ASAP7_75t_R g780 ( 
.A(n_5),
.Y(n_780)
);

CKINVDCx5p33_ASAP7_75t_R g781 ( 
.A(n_271),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_671),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_227),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_23),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_588),
.Y(n_785)
);

CKINVDCx5p33_ASAP7_75t_R g786 ( 
.A(n_572),
.Y(n_786)
);

CKINVDCx20_ASAP7_75t_R g787 ( 
.A(n_569),
.Y(n_787)
);

BUFx3_ASAP7_75t_L g788 ( 
.A(n_544),
.Y(n_788)
);

CKINVDCx5p33_ASAP7_75t_R g789 ( 
.A(n_316),
.Y(n_789)
);

CKINVDCx5p33_ASAP7_75t_R g790 ( 
.A(n_48),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_652),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_331),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_524),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_63),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_29),
.Y(n_795)
);

BUFx6f_ASAP7_75t_L g796 ( 
.A(n_259),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_73),
.Y(n_797)
);

CKINVDCx5p33_ASAP7_75t_R g798 ( 
.A(n_10),
.Y(n_798)
);

CKINVDCx5p33_ASAP7_75t_R g799 ( 
.A(n_167),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_646),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_115),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_47),
.Y(n_802)
);

INVx1_ASAP7_75t_SL g803 ( 
.A(n_624),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_133),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_23),
.Y(n_805)
);

CKINVDCx5p33_ASAP7_75t_R g806 ( 
.A(n_162),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_572),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_480),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_216),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_57),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_217),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_184),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_663),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_653),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_475),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_137),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_143),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_279),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_296),
.Y(n_819)
);

CKINVDCx20_ASAP7_75t_R g820 ( 
.A(n_29),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_683),
.Y(n_821)
);

INVx2_ASAP7_75t_L g822 ( 
.A(n_658),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_619),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_24),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_71),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_471),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_591),
.Y(n_827)
);

INVx2_ASAP7_75t_SL g828 ( 
.A(n_202),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_463),
.Y(n_829)
);

CKINVDCx5p33_ASAP7_75t_R g830 ( 
.A(n_48),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_678),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_102),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_218),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_137),
.Y(n_834)
);

CKINVDCx20_ASAP7_75t_R g835 ( 
.A(n_573),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_676),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_681),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_478),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_84),
.Y(n_839)
);

BUFx6f_ASAP7_75t_L g840 ( 
.A(n_339),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_224),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_320),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_235),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_409),
.Y(n_844)
);

BUFx6f_ASAP7_75t_L g845 ( 
.A(n_134),
.Y(n_845)
);

CKINVDCx5p33_ASAP7_75t_R g846 ( 
.A(n_92),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_370),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_15),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_210),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_577),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_112),
.Y(n_851)
);

CKINVDCx20_ASAP7_75t_R g852 ( 
.A(n_434),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_525),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_621),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_192),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_147),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_423),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_1),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_532),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_348),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_684),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_238),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_504),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_465),
.Y(n_864)
);

CKINVDCx5p33_ASAP7_75t_R g865 ( 
.A(n_486),
.Y(n_865)
);

INVx2_ASAP7_75t_SL g866 ( 
.A(n_549),
.Y(n_866)
);

CKINVDCx16_ASAP7_75t_R g867 ( 
.A(n_535),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_333),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_585),
.Y(n_869)
);

CKINVDCx20_ASAP7_75t_R g870 ( 
.A(n_289),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_502),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_685),
.Y(n_872)
);

INVx1_ASAP7_75t_SL g873 ( 
.A(n_613),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_479),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_237),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_50),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_187),
.Y(n_877)
);

INVx2_ASAP7_75t_SL g878 ( 
.A(n_312),
.Y(n_878)
);

BUFx2_ASAP7_75t_SL g879 ( 
.A(n_398),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_512),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_264),
.Y(n_881)
);

BUFx6f_ASAP7_75t_L g882 ( 
.A(n_155),
.Y(n_882)
);

CKINVDCx5p33_ASAP7_75t_R g883 ( 
.A(n_636),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_148),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_638),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_606),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_219),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_424),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_173),
.Y(n_889)
);

INVx2_ASAP7_75t_SL g890 ( 
.A(n_99),
.Y(n_890)
);

BUFx6f_ASAP7_75t_SL g891 ( 
.A(n_2),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_412),
.Y(n_892)
);

INVx2_ASAP7_75t_SL g893 ( 
.A(n_495),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_106),
.Y(n_894)
);

BUFx8_ASAP7_75t_SL g895 ( 
.A(n_419),
.Y(n_895)
);

CKINVDCx5p33_ASAP7_75t_R g896 ( 
.A(n_349),
.Y(n_896)
);

BUFx3_ASAP7_75t_L g897 ( 
.A(n_316),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_617),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_206),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_666),
.Y(n_900)
);

INVx2_ASAP7_75t_SL g901 ( 
.A(n_226),
.Y(n_901)
);

CKINVDCx20_ASAP7_75t_R g902 ( 
.A(n_557),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_2),
.Y(n_903)
);

CKINVDCx20_ASAP7_75t_R g904 ( 
.A(n_198),
.Y(n_904)
);

CKINVDCx5p33_ASAP7_75t_R g905 ( 
.A(n_342),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_440),
.Y(n_906)
);

BUFx3_ASAP7_75t_L g907 ( 
.A(n_452),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_58),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_342),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_166),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_215),
.Y(n_911)
);

BUFx3_ASAP7_75t_L g912 ( 
.A(n_248),
.Y(n_912)
);

INVx1_ASAP7_75t_SL g913 ( 
.A(n_160),
.Y(n_913)
);

BUFx6f_ASAP7_75t_L g914 ( 
.A(n_288),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_665),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_22),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_433),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_446),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_323),
.Y(n_919)
);

BUFx6f_ASAP7_75t_L g920 ( 
.A(n_259),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_391),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_469),
.Y(n_922)
);

INVxp33_ASAP7_75t_L g923 ( 
.A(n_422),
.Y(n_923)
);

CKINVDCx5p33_ASAP7_75t_R g924 ( 
.A(n_670),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_338),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_662),
.Y(n_926)
);

CKINVDCx20_ASAP7_75t_R g927 ( 
.A(n_233),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_97),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_437),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_250),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_291),
.Y(n_931)
);

CKINVDCx20_ASAP7_75t_R g932 ( 
.A(n_328),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_97),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_580),
.Y(n_934)
);

BUFx2_ASAP7_75t_SL g935 ( 
.A(n_204),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_675),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_345),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_679),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_468),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_190),
.Y(n_940)
);

CKINVDCx5p33_ASAP7_75t_R g941 ( 
.A(n_126),
.Y(n_941)
);

BUFx10_ASAP7_75t_L g942 ( 
.A(n_126),
.Y(n_942)
);

BUFx5_ASAP7_75t_L g943 ( 
.A(n_441),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_590),
.Y(n_944)
);

BUFx10_ASAP7_75t_L g945 ( 
.A(n_19),
.Y(n_945)
);

CKINVDCx20_ASAP7_75t_R g946 ( 
.A(n_99),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_512),
.Y(n_947)
);

CKINVDCx5p33_ASAP7_75t_R g948 ( 
.A(n_690),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_217),
.Y(n_949)
);

BUFx10_ASAP7_75t_L g950 ( 
.A(n_257),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_115),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_76),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_151),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_167),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_461),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_42),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_534),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_600),
.Y(n_958)
);

CKINVDCx5p33_ASAP7_75t_R g959 ( 
.A(n_334),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_34),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_444),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_537),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_396),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_326),
.Y(n_964)
);

CKINVDCx20_ASAP7_75t_R g965 ( 
.A(n_604),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_357),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_586),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_74),
.Y(n_968)
);

INVx1_ASAP7_75t_SL g969 ( 
.A(n_231),
.Y(n_969)
);

BUFx3_ASAP7_75t_L g970 ( 
.A(n_506),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_561),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_420),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_563),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_223),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_362),
.Y(n_975)
);

BUFx2_ASAP7_75t_L g976 ( 
.A(n_361),
.Y(n_976)
);

CKINVDCx5p33_ASAP7_75t_R g977 ( 
.A(n_651),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_350),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_630),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_252),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_492),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_441),
.Y(n_982)
);

INVx3_ASAP7_75t_L g983 ( 
.A(n_304),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_284),
.Y(n_984)
);

CKINVDCx20_ASAP7_75t_R g985 ( 
.A(n_261),
.Y(n_985)
);

CKINVDCx5p33_ASAP7_75t_R g986 ( 
.A(n_436),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_240),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_225),
.Y(n_988)
);

CKINVDCx20_ASAP7_75t_R g989 ( 
.A(n_510),
.Y(n_989)
);

INVx1_ASAP7_75t_SL g990 ( 
.A(n_7),
.Y(n_990)
);

CKINVDCx16_ASAP7_75t_R g991 ( 
.A(n_588),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_507),
.Y(n_992)
);

BUFx8_ASAP7_75t_SL g993 ( 
.A(n_64),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_413),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_192),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_667),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_321),
.Y(n_997)
);

CKINVDCx5p33_ASAP7_75t_R g998 ( 
.A(n_216),
.Y(n_998)
);

BUFx10_ASAP7_75t_L g999 ( 
.A(n_419),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_340),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_540),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_246),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_602),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_241),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_647),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_498),
.Y(n_1006)
);

CKINVDCx5p33_ASAP7_75t_R g1007 ( 
.A(n_686),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_100),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_682),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_283),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_664),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_131),
.Y(n_1012)
);

INVx2_ASAP7_75t_L g1013 ( 
.A(n_233),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_241),
.Y(n_1014)
);

CKINVDCx20_ASAP7_75t_R g1015 ( 
.A(n_491),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_90),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_290),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_579),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_485),
.Y(n_1019)
);

CKINVDCx20_ASAP7_75t_R g1020 ( 
.A(n_485),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_585),
.Y(n_1021)
);

BUFx3_ASAP7_75t_L g1022 ( 
.A(n_557),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_176),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_183),
.Y(n_1024)
);

BUFx2_ASAP7_75t_L g1025 ( 
.A(n_425),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_394),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_426),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_565),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_537),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_380),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_58),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_417),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_636),
.Y(n_1033)
);

CKINVDCx20_ASAP7_75t_R g1034 ( 
.A(n_657),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_515),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_372),
.Y(n_1036)
);

BUFx10_ASAP7_75t_L g1037 ( 
.A(n_501),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_401),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_380),
.Y(n_1039)
);

CKINVDCx16_ASAP7_75t_R g1040 ( 
.A(n_536),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_536),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_421),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_563),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_440),
.Y(n_1044)
);

CKINVDCx16_ASAP7_75t_R g1045 ( 
.A(n_206),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_661),
.Y(n_1046)
);

CKINVDCx20_ASAP7_75t_R g1047 ( 
.A(n_334),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_98),
.Y(n_1048)
);

BUFx2_ASAP7_75t_SL g1049 ( 
.A(n_144),
.Y(n_1049)
);

BUFx10_ASAP7_75t_L g1050 ( 
.A(n_0),
.Y(n_1050)
);

INVx2_ASAP7_75t_L g1051 ( 
.A(n_625),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_203),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_346),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_200),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_468),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_153),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_486),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_543),
.Y(n_1058)
);

CKINVDCx5p33_ASAP7_75t_R g1059 ( 
.A(n_272),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_619),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_135),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_533),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_354),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_643),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_28),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_654),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_71),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_297),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_629),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_507),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_524),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_268),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_338),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_357),
.Y(n_1074)
);

CKINVDCx5p33_ASAP7_75t_R g1075 ( 
.A(n_511),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_335),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_656),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_78),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_257),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_41),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_379),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_385),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_292),
.Y(n_1083)
);

INVx1_ASAP7_75t_SL g1084 ( 
.A(n_436),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_286),
.Y(n_1085)
);

INVx1_ASAP7_75t_SL g1086 ( 
.A(n_389),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_325),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_128),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_247),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_519),
.Y(n_1090)
);

CKINVDCx5p33_ASAP7_75t_R g1091 ( 
.A(n_125),
.Y(n_1091)
);

CKINVDCx20_ASAP7_75t_R g1092 ( 
.A(n_134),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_31),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_42),
.Y(n_1094)
);

BUFx2_ASAP7_75t_L g1095 ( 
.A(n_41),
.Y(n_1095)
);

INVx1_ASAP7_75t_SL g1096 ( 
.A(n_583),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_533),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_531),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_448),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_472),
.Y(n_1100)
);

INVx2_ASAP7_75t_L g1101 ( 
.A(n_145),
.Y(n_1101)
);

INVx1_ASAP7_75t_SL g1102 ( 
.A(n_677),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_60),
.Y(n_1103)
);

INVx1_ASAP7_75t_L g1104 ( 
.A(n_464),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_659),
.Y(n_1105)
);

CKINVDCx5p33_ASAP7_75t_R g1106 ( 
.A(n_650),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_463),
.Y(n_1107)
);

INVxp67_ASAP7_75t_SL g1108 ( 
.A(n_33),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_339),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_385),
.Y(n_1110)
);

BUFx6f_ASAP7_75t_L g1111 ( 
.A(n_594),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_224),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_104),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_469),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_118),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_169),
.Y(n_1116)
);

CKINVDCx5p33_ASAP7_75t_R g1117 ( 
.A(n_107),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_36),
.Y(n_1118)
);

CKINVDCx5p33_ASAP7_75t_R g1119 ( 
.A(n_9),
.Y(n_1119)
);

BUFx10_ASAP7_75t_L g1120 ( 
.A(n_275),
.Y(n_1120)
);

BUFx3_ASAP7_75t_L g1121 ( 
.A(n_152),
.Y(n_1121)
);

BUFx3_ASAP7_75t_L g1122 ( 
.A(n_687),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_89),
.Y(n_1123)
);

INVx2_ASAP7_75t_SL g1124 ( 
.A(n_574),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_230),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_248),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_116),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_313),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_211),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_359),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_278),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_249),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_190),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_477),
.Y(n_1134)
);

CKINVDCx20_ASAP7_75t_R g1135 ( 
.A(n_632),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_142),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_153),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_238),
.Y(n_1138)
);

CKINVDCx16_ASAP7_75t_R g1139 ( 
.A(n_336),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_479),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_637),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_613),
.Y(n_1142)
);

INVx2_ASAP7_75t_L g1143 ( 
.A(n_556),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_644),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_184),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_187),
.Y(n_1146)
);

CKINVDCx5p33_ASAP7_75t_R g1147 ( 
.A(n_222),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_26),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_561),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_604),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_159),
.Y(n_1151)
);

INVx2_ASAP7_75t_L g1152 ( 
.A(n_131),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_615),
.Y(n_1153)
);

INVx1_ASAP7_75t_L g1154 ( 
.A(n_94),
.Y(n_1154)
);

BUFx2_ASAP7_75t_L g1155 ( 
.A(n_36),
.Y(n_1155)
);

CKINVDCx5p33_ASAP7_75t_R g1156 ( 
.A(n_4),
.Y(n_1156)
);

INVxp67_ASAP7_75t_L g1157 ( 
.A(n_299),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_174),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_317),
.Y(n_1159)
);

CKINVDCx5p33_ASAP7_75t_R g1160 ( 
.A(n_502),
.Y(n_1160)
);

CKINVDCx5p33_ASAP7_75t_R g1161 ( 
.A(n_347),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_279),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_303),
.Y(n_1163)
);

CKINVDCx5p33_ASAP7_75t_R g1164 ( 
.A(n_113),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_348),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_408),
.Y(n_1166)
);

BUFx6f_ASAP7_75t_L g1167 ( 
.A(n_164),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_109),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_130),
.Y(n_1169)
);

INVx1_ASAP7_75t_L g1170 ( 
.A(n_249),
.Y(n_1170)
);

CKINVDCx5p33_ASAP7_75t_R g1171 ( 
.A(n_162),
.Y(n_1171)
);

CKINVDCx5p33_ASAP7_75t_R g1172 ( 
.A(n_366),
.Y(n_1172)
);

CKINVDCx5p33_ASAP7_75t_R g1173 ( 
.A(n_148),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_445),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_180),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_672),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_474),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_170),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_201),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_11),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_288),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_669),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_655),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_545),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_293),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_689),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_264),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_429),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_59),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_139),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_522),
.Y(n_1191)
);

BUFx3_ASAP7_75t_L g1192 ( 
.A(n_423),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_414),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_302),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_250),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_138),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_565),
.Y(n_1197)
);

CKINVDCx20_ASAP7_75t_R g1198 ( 
.A(n_442),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_432),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_518),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_660),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_62),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_466),
.Y(n_1203)
);

CKINVDCx16_ASAP7_75t_R g1204 ( 
.A(n_26),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_630),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_366),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_506),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_78),
.Y(n_1208)
);

CKINVDCx5p33_ASAP7_75t_R g1209 ( 
.A(n_411),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_74),
.Y(n_1210)
);

INVxp67_ASAP7_75t_L g1211 ( 
.A(n_155),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_285),
.Y(n_1212)
);

CKINVDCx16_ASAP7_75t_R g1213 ( 
.A(n_467),
.Y(n_1213)
);

BUFx10_ASAP7_75t_L g1214 ( 
.A(n_193),
.Y(n_1214)
);

CKINVDCx5p33_ASAP7_75t_R g1215 ( 
.A(n_194),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_603),
.Y(n_1216)
);

INVx2_ASAP7_75t_L g1217 ( 
.A(n_645),
.Y(n_1217)
);

NOR2xp33_ASAP7_75t_L g1218 ( 
.A(n_923),
.B(n_779),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_727),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_779),
.Y(n_1220)
);

HB1xp67_ASAP7_75t_L g1221 ( 
.A(n_976),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_779),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_943),
.Y(n_1223)
);

INVx2_ASAP7_75t_SL g1224 ( 
.A(n_700),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_779),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_908),
.Y(n_1226)
);

CKINVDCx5p33_ASAP7_75t_R g1227 ( 
.A(n_895),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_908),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_891),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_908),
.Y(n_1230)
);

CKINVDCx20_ASAP7_75t_R g1231 ( 
.A(n_867),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_891),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_908),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_982),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_891),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_982),
.Y(n_1236)
);

BUFx3_ASAP7_75t_L g1237 ( 
.A(n_1122),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_982),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_993),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_891),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_982),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_983),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_943),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_983),
.Y(n_1244)
);

CKINVDCx20_ASAP7_75t_R g1245 ( 
.A(n_867),
.Y(n_1245)
);

BUFx5_ASAP7_75t_L g1246 ( 
.A(n_713),
.Y(n_1246)
);

BUFx2_ASAP7_75t_L g1247 ( 
.A(n_976),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_983),
.Y(n_1248)
);

CKINVDCx16_ASAP7_75t_R g1249 ( 
.A(n_991),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_983),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1025),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_700),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_991),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_943),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_1034),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_702),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_700),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_704),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_1040),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_788),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_788),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_788),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_1040),
.Y(n_1263)
);

CKINVDCx20_ASAP7_75t_R g1264 ( 
.A(n_1045),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_871),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_871),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_1045),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_871),
.Y(n_1268)
);

CKINVDCx20_ASAP7_75t_R g1269 ( 
.A(n_1139),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_897),
.Y(n_1270)
);

BUFx2_ASAP7_75t_SL g1271 ( 
.A(n_1122),
.Y(n_1271)
);

BUFx3_ASAP7_75t_L g1272 ( 
.A(n_1122),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_897),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_897),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_907),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_907),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_907),
.Y(n_1277)
);

CKINVDCx20_ASAP7_75t_R g1278 ( 
.A(n_1139),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_912),
.Y(n_1279)
);

INVx2_ASAP7_75t_L g1280 ( 
.A(n_943),
.Y(n_1280)
);

CKINVDCx5p33_ASAP7_75t_R g1281 ( 
.A(n_1187),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_912),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_912),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_713),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_970),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_970),
.Y(n_1286)
);

INVx2_ASAP7_75t_L g1287 ( 
.A(n_943),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_970),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1022),
.Y(n_1289)
);

INVx1_ASAP7_75t_L g1290 ( 
.A(n_1022),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1022),
.Y(n_1291)
);

INVx1_ASAP7_75t_SL g1292 ( 
.A(n_722),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1039),
.Y(n_1293)
);

BUFx5_ASAP7_75t_L g1294 ( 
.A(n_782),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1039),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1039),
.Y(n_1296)
);

CKINVDCx20_ASAP7_75t_R g1297 ( 
.A(n_1187),
.Y(n_1297)
);

CKINVDCx20_ASAP7_75t_R g1298 ( 
.A(n_1204),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1121),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_943),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1121),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1204),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1121),
.Y(n_1303)
);

INVxp33_ASAP7_75t_L g1304 ( 
.A(n_1132),
.Y(n_1304)
);

INVxp67_ASAP7_75t_L g1305 ( 
.A(n_1025),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1192),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1192),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1192),
.Y(n_1308)
);

INVxp33_ASAP7_75t_L g1309 ( 
.A(n_1073),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1073),
.Y(n_1310)
);

INVxp33_ASAP7_75t_L g1311 ( 
.A(n_1095),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1205),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1205),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1205),
.Y(n_1314)
);

BUFx3_ASAP7_75t_L g1315 ( 
.A(n_782),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1095),
.B(n_0),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_726),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_726),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_726),
.Y(n_1319)
);

INVxp33_ASAP7_75t_L g1320 ( 
.A(n_1155),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_783),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_783),
.Y(n_1322)
);

CKINVDCx20_ASAP7_75t_R g1323 ( 
.A(n_1213),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_783),
.Y(n_1324)
);

BUFx8_ASAP7_75t_SL g1325 ( 
.A(n_1155),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_880),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_1213),
.Y(n_1327)
);

INVx2_ASAP7_75t_L g1328 ( 
.A(n_943),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_691),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_693),
.Y(n_1330)
);

CKINVDCx16_ASAP7_75t_R g1331 ( 
.A(n_942),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_694),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_880),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_696),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_880),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_934),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_737),
.Y(n_1337)
);

INVx1_ASAP7_75t_SL g1338 ( 
.A(n_745),
.Y(n_1338)
);

CKINVDCx16_ASAP7_75t_R g1339 ( 
.A(n_942),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_943),
.Y(n_1340)
);

INVxp67_ASAP7_75t_L g1341 ( 
.A(n_1200),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1200),
.Y(n_1342)
);

INVxp33_ASAP7_75t_L g1343 ( 
.A(n_730),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_934),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_934),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_697),
.Y(n_1346)
);

BUFx3_ASAP7_75t_L g1347 ( 
.A(n_821),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_698),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1109),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_943),
.Y(n_1350)
);

INVxp67_ASAP7_75t_SL g1351 ( 
.A(n_1217),
.Y(n_1351)
);

INVx1_ASAP7_75t_SL g1352 ( 
.A(n_748),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1109),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1109),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1217),
.Y(n_1355)
);

INVxp67_ASAP7_75t_L g1356 ( 
.A(n_751),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1217),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_692),
.Y(n_1358)
);

NOR2xp33_ASAP7_75t_L g1359 ( 
.A(n_821),
.B(n_3),
.Y(n_1359)
);

CKINVDCx5p33_ASAP7_75t_R g1360 ( 
.A(n_701),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_942),
.Y(n_1361)
);

INVxp67_ASAP7_75t_L g1362 ( 
.A(n_751),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_692),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_861),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_695),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_695),
.Y(n_1366)
);

CKINVDCx20_ASAP7_75t_R g1367 ( 
.A(n_753),
.Y(n_1367)
);

INVxp67_ASAP7_75t_SL g1368 ( 
.A(n_796),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_699),
.Y(n_1369)
);

INVxp67_ASAP7_75t_L g1370 ( 
.A(n_772),
.Y(n_1370)
);

CKINVDCx20_ASAP7_75t_R g1371 ( 
.A(n_762),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_699),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_707),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_707),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_796),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_710),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_710),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_703),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_712),
.Y(n_1379)
);

BUFx6f_ASAP7_75t_L g1380 ( 
.A(n_796),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_705),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_712),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_714),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_714),
.Y(n_1384)
);

CKINVDCx14_ASAP7_75t_R g1385 ( 
.A(n_733),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_719),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_719),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_723),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_723),
.Y(n_1389)
);

CKINVDCx16_ASAP7_75t_R g1390 ( 
.A(n_942),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_724),
.Y(n_1391)
);

INVx1_ASAP7_75t_SL g1392 ( 
.A(n_780),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_724),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_734),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_734),
.Y(n_1395)
);

BUFx10_ASAP7_75t_L g1396 ( 
.A(n_796),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_796),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_741),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_741),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_742),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_742),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_749),
.Y(n_1402)
);

INVxp33_ASAP7_75t_SL g1403 ( 
.A(n_706),
.Y(n_1403)
);

INVxp67_ASAP7_75t_SL g1404 ( 
.A(n_796),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_749),
.Y(n_1405)
);

INVxp67_ASAP7_75t_SL g1406 ( 
.A(n_840),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_708),
.Y(n_1407)
);

CKINVDCx5p33_ASAP7_75t_R g1408 ( 
.A(n_709),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_760),
.Y(n_1409)
);

NOR2xp67_ASAP7_75t_L g1410 ( 
.A(n_828),
.B(n_866),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_840),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_760),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_767),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_767),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_768),
.Y(n_1415)
);

INVx2_ASAP7_75t_L g1416 ( 
.A(n_840),
.Y(n_1416)
);

INVxp33_ASAP7_75t_L g1417 ( 
.A(n_730),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_768),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_769),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_711),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_769),
.Y(n_1421)
);

INVxp67_ASAP7_75t_SL g1422 ( 
.A(n_840),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_715),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_793),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_793),
.Y(n_1425)
);

CKINVDCx14_ASAP7_75t_R g1426 ( 
.A(n_738),
.Y(n_1426)
);

CKINVDCx14_ASAP7_75t_R g1427 ( 
.A(n_757),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_795),
.Y(n_1428)
);

INVxp67_ASAP7_75t_L g1429 ( 
.A(n_772),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_716),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_840),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_795),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_802),
.Y(n_1433)
);

INVxp67_ASAP7_75t_SL g1434 ( 
.A(n_840),
.Y(n_1434)
);

INVxp33_ASAP7_75t_SL g1435 ( 
.A(n_717),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_802),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_787),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_845),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_804),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_804),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_805),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_805),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_718),
.Y(n_1443)
);

INVxp33_ASAP7_75t_L g1444 ( 
.A(n_732),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_809),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_809),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_845),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_720),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_721),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_810),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_845),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_810),
.Y(n_1452)
);

CKINVDCx20_ASAP7_75t_R g1453 ( 
.A(n_815),
.Y(n_1453)
);

INVxp67_ASAP7_75t_L g1454 ( 
.A(n_879),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_816),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_845),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_816),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_817),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_817),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_725),
.Y(n_1460)
);

INVxp33_ASAP7_75t_SL g1461 ( 
.A(n_728),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_818),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_818),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_823),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_823),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_845),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_845),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_824),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_882),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_882),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_824),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_731),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_825),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_735),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_825),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_826),
.Y(n_1476)
);

INVxp33_ASAP7_75t_SL g1477 ( 
.A(n_736),
.Y(n_1477)
);

CKINVDCx20_ASAP7_75t_R g1478 ( 
.A(n_820),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_826),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_739),
.Y(n_1480)
);

INVx2_ASAP7_75t_SL g1481 ( 
.A(n_945),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_829),
.Y(n_1482)
);

BUFx3_ASAP7_75t_L g1483 ( 
.A(n_861),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_829),
.Y(n_1484)
);

BUFx2_ASAP7_75t_L g1485 ( 
.A(n_740),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_743),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_882),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_832),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_832),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_834),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_744),
.Y(n_1491)
);

INVx1_ASAP7_75t_SL g1492 ( 
.A(n_835),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_834),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_844),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_746),
.Y(n_1495)
);

CKINVDCx20_ASAP7_75t_R g1496 ( 
.A(n_852),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_844),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_848),
.Y(n_1498)
);

CKINVDCx16_ASAP7_75t_R g1499 ( 
.A(n_945),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_882),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_747),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_848),
.Y(n_1502)
);

CKINVDCx20_ASAP7_75t_R g1503 ( 
.A(n_870),
.Y(n_1503)
);

CKINVDCx20_ASAP7_75t_R g1504 ( 
.A(n_899),
.Y(n_1504)
);

HB1xp67_ASAP7_75t_L g1505 ( 
.A(n_750),
.Y(n_1505)
);

BUFx2_ASAP7_75t_L g1506 ( 
.A(n_752),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_754),
.Y(n_1507)
);

NOR2xp67_ASAP7_75t_L g1508 ( 
.A(n_828),
.B(n_1),
.Y(n_1508)
);

BUFx3_ASAP7_75t_L g1509 ( 
.A(n_872),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_851),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_851),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_854),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_854),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_856),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_856),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_858),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_756),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_858),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_860),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_902),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_860),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_862),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_862),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_758),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_864),
.Y(n_1525)
);

BUFx2_ASAP7_75t_L g1526 ( 
.A(n_759),
.Y(n_1526)
);

NOR2xp67_ASAP7_75t_L g1527 ( 
.A(n_866),
.B(n_3),
.Y(n_1527)
);

NOR2xp33_ASAP7_75t_L g1528 ( 
.A(n_872),
.B(n_5),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_904),
.Y(n_1529)
);

CKINVDCx16_ASAP7_75t_R g1530 ( 
.A(n_945),
.Y(n_1530)
);

CKINVDCx5p33_ASAP7_75t_R g1531 ( 
.A(n_761),
.Y(n_1531)
);

CKINVDCx16_ASAP7_75t_R g1532 ( 
.A(n_945),
.Y(n_1532)
);

NOR2xp67_ASAP7_75t_L g1533 ( 
.A(n_878),
.B(n_4),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_763),
.Y(n_1534)
);

CKINVDCx16_ASAP7_75t_R g1535 ( 
.A(n_950),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_864),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_868),
.Y(n_1537)
);

CKINVDCx5p33_ASAP7_75t_R g1538 ( 
.A(n_764),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_868),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_765),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_874),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_921),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_874),
.Y(n_1543)
);

INVx3_ASAP7_75t_L g1544 ( 
.A(n_882),
.Y(n_1544)
);

INVx2_ASAP7_75t_L g1545 ( 
.A(n_882),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_877),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_877),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_766),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_770),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_885),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_885),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_886),
.Y(n_1552)
);

CKINVDCx20_ASAP7_75t_R g1553 ( 
.A(n_927),
.Y(n_1553)
);

INVxp67_ASAP7_75t_L g1554 ( 
.A(n_879),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_886),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_887),
.Y(n_1556)
);

CKINVDCx16_ASAP7_75t_R g1557 ( 
.A(n_950),
.Y(n_1557)
);

CKINVDCx16_ASAP7_75t_R g1558 ( 
.A(n_950),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_887),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_889),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_889),
.Y(n_1561)
);

CKINVDCx5p33_ASAP7_75t_R g1562 ( 
.A(n_771),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_935),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_894),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_936),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_914),
.Y(n_1566)
);

INVx1_ASAP7_75t_L g1567 ( 
.A(n_894),
.Y(n_1567)
);

CKINVDCx16_ASAP7_75t_R g1568 ( 
.A(n_950),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_910),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_910),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_911),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_L g1572 ( 
.A(n_914),
.Y(n_1572)
);

INVx2_ASAP7_75t_L g1573 ( 
.A(n_914),
.Y(n_1573)
);

CKINVDCx20_ASAP7_75t_R g1574 ( 
.A(n_932),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_774),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_911),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_918),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_918),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_925),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_925),
.Y(n_1580)
);

CKINVDCx5p33_ASAP7_75t_R g1581 ( 
.A(n_775),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_929),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_929),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_936),
.B(n_7),
.Y(n_1584)
);

INVxp33_ASAP7_75t_SL g1585 ( 
.A(n_776),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_930),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_946),
.Y(n_1587)
);

INVxp67_ASAP7_75t_SL g1588 ( 
.A(n_914),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_930),
.Y(n_1589)
);

CKINVDCx5p33_ASAP7_75t_R g1590 ( 
.A(n_777),
.Y(n_1590)
);

INVxp67_ASAP7_75t_L g1591 ( 
.A(n_935),
.Y(n_1591)
);

CKINVDCx5p33_ASAP7_75t_R g1592 ( 
.A(n_778),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_933),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_933),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_937),
.Y(n_1595)
);

BUFx3_ASAP7_75t_L g1596 ( 
.A(n_1011),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_781),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_937),
.Y(n_1598)
);

INVxp67_ASAP7_75t_SL g1599 ( 
.A(n_914),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_939),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_939),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_944),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_944),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_949),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_949),
.Y(n_1605)
);

INVxp67_ASAP7_75t_L g1606 ( 
.A(n_1049),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_914),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_951),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1011),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_920),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_951),
.Y(n_1611)
);

CKINVDCx5p33_ASAP7_75t_R g1612 ( 
.A(n_784),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_955),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_955),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_956),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_956),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_960),
.Y(n_1617)
);

INVxp67_ASAP7_75t_L g1618 ( 
.A(n_1049),
.Y(n_1618)
);

CKINVDCx5p33_ASAP7_75t_R g1619 ( 
.A(n_785),
.Y(n_1619)
);

BUFx3_ASAP7_75t_L g1620 ( 
.A(n_1046),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_960),
.Y(n_1621)
);

CKINVDCx5p33_ASAP7_75t_R g1622 ( 
.A(n_786),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_789),
.Y(n_1623)
);

BUFx6f_ASAP7_75t_L g1624 ( 
.A(n_920),
.Y(n_1624)
);

INVxp33_ASAP7_75t_L g1625 ( 
.A(n_732),
.Y(n_1625)
);

CKINVDCx5p33_ASAP7_75t_R g1626 ( 
.A(n_790),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_961),
.Y(n_1627)
);

INVx3_ASAP7_75t_L g1628 ( 
.A(n_920),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_792),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_961),
.Y(n_1630)
);

BUFx3_ASAP7_75t_L g1631 ( 
.A(n_1046),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_999),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_967),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_967),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_971),
.Y(n_1635)
);

INVx1_ASAP7_75t_SL g1636 ( 
.A(n_965),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_971),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_972),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_794),
.Y(n_1639)
);

CKINVDCx5p33_ASAP7_75t_R g1640 ( 
.A(n_797),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_972),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_978),
.Y(n_1642)
);

CKINVDCx20_ASAP7_75t_R g1643 ( 
.A(n_985),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1220),
.Y(n_1644)
);

CKINVDCx20_ASAP7_75t_R g1645 ( 
.A(n_1367),
.Y(n_1645)
);

CKINVDCx5p33_ASAP7_75t_R g1646 ( 
.A(n_1255),
.Y(n_1646)
);

CKINVDCx5p33_ASAP7_75t_R g1647 ( 
.A(n_1227),
.Y(n_1647)
);

BUFx2_ASAP7_75t_SL g1648 ( 
.A(n_1231),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1222),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1380),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1225),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1226),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1228),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1239),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1230),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1385),
.B(n_1201),
.Y(n_1656)
);

CKINVDCx20_ASAP7_75t_R g1657 ( 
.A(n_1367),
.Y(n_1657)
);

NOR2xp33_ASAP7_75t_L g1658 ( 
.A(n_1385),
.B(n_1201),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1233),
.Y(n_1659)
);

CKINVDCx5p33_ASAP7_75t_R g1660 ( 
.A(n_1256),
.Y(n_1660)
);

CKINVDCx5p33_ASAP7_75t_R g1661 ( 
.A(n_1258),
.Y(n_1661)
);

CKINVDCx20_ASAP7_75t_R g1662 ( 
.A(n_1371),
.Y(n_1662)
);

CKINVDCx5p33_ASAP7_75t_R g1663 ( 
.A(n_1292),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1426),
.B(n_938),
.Y(n_1664)
);

CKINVDCx5p33_ASAP7_75t_R g1665 ( 
.A(n_1337),
.Y(n_1665)
);

BUFx6f_ASAP7_75t_L g1666 ( 
.A(n_1380),
.Y(n_1666)
);

CKINVDCx5p33_ASAP7_75t_R g1667 ( 
.A(n_1338),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1352),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1234),
.Y(n_1669)
);

NOR2xp33_ASAP7_75t_L g1670 ( 
.A(n_1426),
.B(n_1102),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1271),
.B(n_729),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1380),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1343),
.B(n_999),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1236),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1238),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1241),
.Y(n_1676)
);

CKINVDCx20_ASAP7_75t_R g1677 ( 
.A(n_1371),
.Y(n_1677)
);

INVxp67_ASAP7_75t_SL g1678 ( 
.A(n_1237),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1242),
.Y(n_1679)
);

CKINVDCx5p33_ASAP7_75t_R g1680 ( 
.A(n_1392),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1244),
.Y(n_1681)
);

CKINVDCx20_ASAP7_75t_R g1682 ( 
.A(n_1437),
.Y(n_1682)
);

CKINVDCx20_ASAP7_75t_R g1683 ( 
.A(n_1437),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1248),
.Y(n_1684)
);

INVxp67_ASAP7_75t_SL g1685 ( 
.A(n_1237),
.Y(n_1685)
);

CKINVDCx5p33_ASAP7_75t_R g1686 ( 
.A(n_1492),
.Y(n_1686)
);

INVxp67_ASAP7_75t_SL g1687 ( 
.A(n_1272),
.Y(n_1687)
);

INVxp67_ASAP7_75t_SL g1688 ( 
.A(n_1272),
.Y(n_1688)
);

CKINVDCx16_ASAP7_75t_R g1689 ( 
.A(n_1331),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1250),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1380),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1229),
.B(n_729),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1427),
.Y(n_1693)
);

BUFx6f_ASAP7_75t_L g1694 ( 
.A(n_1451),
.Y(n_1694)
);

CKINVDCx5p33_ASAP7_75t_R g1695 ( 
.A(n_1427),
.Y(n_1695)
);

CKINVDCx5p33_ASAP7_75t_R g1696 ( 
.A(n_1360),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1351),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1252),
.Y(n_1698)
);

CKINVDCx5p33_ASAP7_75t_R g1699 ( 
.A(n_1636),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1257),
.Y(n_1700)
);

CKINVDCx5p33_ASAP7_75t_R g1701 ( 
.A(n_1378),
.Y(n_1701)
);

CKINVDCx5p33_ASAP7_75t_R g1702 ( 
.A(n_1381),
.Y(n_1702)
);

CKINVDCx5p33_ASAP7_75t_R g1703 ( 
.A(n_1407),
.Y(n_1703)
);

CKINVDCx20_ASAP7_75t_R g1704 ( 
.A(n_1453),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1260),
.Y(n_1705)
);

NOR2xp33_ASAP7_75t_L g1706 ( 
.A(n_1229),
.B(n_822),
.Y(n_1706)
);

CKINVDCx5p33_ASAP7_75t_R g1707 ( 
.A(n_1581),
.Y(n_1707)
);

BUFx3_ASAP7_75t_L g1708 ( 
.A(n_1396),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1261),
.Y(n_1709)
);

CKINVDCx5p33_ASAP7_75t_R g1710 ( 
.A(n_1590),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1396),
.Y(n_1711)
);

INVxp67_ASAP7_75t_L g1712 ( 
.A(n_1485),
.Y(n_1712)
);

CKINVDCx20_ASAP7_75t_R g1713 ( 
.A(n_1453),
.Y(n_1713)
);

CKINVDCx5p33_ASAP7_75t_R g1714 ( 
.A(n_1592),
.Y(n_1714)
);

CKINVDCx5p33_ASAP7_75t_R g1715 ( 
.A(n_1329),
.Y(n_1715)
);

CKINVDCx20_ASAP7_75t_R g1716 ( 
.A(n_1478),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1262),
.Y(n_1717)
);

INVxp33_ASAP7_75t_SL g1718 ( 
.A(n_1219),
.Y(n_1718)
);

CKINVDCx5p33_ASAP7_75t_R g1719 ( 
.A(n_1329),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1232),
.B(n_822),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1265),
.Y(n_1721)
);

CKINVDCx5p33_ASAP7_75t_R g1722 ( 
.A(n_1330),
.Y(n_1722)
);

INVxp67_ASAP7_75t_SL g1723 ( 
.A(n_1368),
.Y(n_1723)
);

CKINVDCx5p33_ASAP7_75t_R g1724 ( 
.A(n_1330),
.Y(n_1724)
);

INVxp67_ASAP7_75t_SL g1725 ( 
.A(n_1404),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1266),
.Y(n_1726)
);

CKINVDCx5p33_ASAP7_75t_R g1727 ( 
.A(n_1332),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1268),
.Y(n_1728)
);

BUFx2_ASAP7_75t_SL g1729 ( 
.A(n_1231),
.Y(n_1729)
);

HB1xp67_ASAP7_75t_L g1730 ( 
.A(n_1249),
.Y(n_1730)
);

CKINVDCx20_ASAP7_75t_R g1731 ( 
.A(n_1478),
.Y(n_1731)
);

INVxp67_ASAP7_75t_SL g1732 ( 
.A(n_1406),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1451),
.Y(n_1733)
);

CKINVDCx20_ASAP7_75t_R g1734 ( 
.A(n_1496),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1270),
.Y(n_1735)
);

INVxp67_ASAP7_75t_SL g1736 ( 
.A(n_1422),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1273),
.Y(n_1737)
);

CKINVDCx5p33_ASAP7_75t_R g1738 ( 
.A(n_1332),
.Y(n_1738)
);

CKINVDCx5p33_ASAP7_75t_R g1739 ( 
.A(n_1334),
.Y(n_1739)
);

CKINVDCx5p33_ASAP7_75t_R g1740 ( 
.A(n_1232),
.Y(n_1740)
);

BUFx6f_ASAP7_75t_L g1741 ( 
.A(n_1451),
.Y(n_1741)
);

CKINVDCx20_ASAP7_75t_R g1742 ( 
.A(n_1496),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1235),
.B(n_837),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1263),
.Y(n_1744)
);

CKINVDCx16_ASAP7_75t_R g1745 ( 
.A(n_1339),
.Y(n_1745)
);

INVx1_ASAP7_75t_L g1746 ( 
.A(n_1274),
.Y(n_1746)
);

CKINVDCx5p33_ASAP7_75t_R g1747 ( 
.A(n_1334),
.Y(n_1747)
);

INVxp67_ASAP7_75t_SL g1748 ( 
.A(n_1434),
.Y(n_1748)
);

CKINVDCx5p33_ASAP7_75t_R g1749 ( 
.A(n_1346),
.Y(n_1749)
);

CKINVDCx20_ASAP7_75t_R g1750 ( 
.A(n_1503),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1275),
.Y(n_1751)
);

CKINVDCx5p33_ASAP7_75t_R g1752 ( 
.A(n_1346),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1451),
.Y(n_1753)
);

CKINVDCx5p33_ASAP7_75t_R g1754 ( 
.A(n_1348),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1276),
.Y(n_1755)
);

HB1xp67_ASAP7_75t_L g1756 ( 
.A(n_1263),
.Y(n_1756)
);

CKINVDCx20_ASAP7_75t_R g1757 ( 
.A(n_1503),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_L g1758 ( 
.A(n_1235),
.B(n_837),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1277),
.Y(n_1759)
);

INVxp33_ASAP7_75t_L g1760 ( 
.A(n_1218),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1279),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1282),
.Y(n_1762)
);

NOR2xp33_ASAP7_75t_L g1763 ( 
.A(n_1240),
.B(n_1219),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1469),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1283),
.Y(n_1765)
);

NOR2xp67_ASAP7_75t_L g1766 ( 
.A(n_1240),
.B(n_773),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1285),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1286),
.Y(n_1768)
);

CKINVDCx20_ASAP7_75t_R g1769 ( 
.A(n_1504),
.Y(n_1769)
);

CKINVDCx5p33_ASAP7_75t_R g1770 ( 
.A(n_1348),
.Y(n_1770)
);

BUFx2_ASAP7_75t_SL g1771 ( 
.A(n_1245),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1288),
.Y(n_1772)
);

INVx2_ASAP7_75t_L g1773 ( 
.A(n_1469),
.Y(n_1773)
);

CKINVDCx5p33_ASAP7_75t_R g1774 ( 
.A(n_1408),
.Y(n_1774)
);

CKINVDCx20_ASAP7_75t_R g1775 ( 
.A(n_1504),
.Y(n_1775)
);

CKINVDCx20_ASAP7_75t_R g1776 ( 
.A(n_1520),
.Y(n_1776)
);

CKINVDCx5p33_ASAP7_75t_R g1777 ( 
.A(n_1408),
.Y(n_1777)
);

CKINVDCx5p33_ASAP7_75t_R g1778 ( 
.A(n_1420),
.Y(n_1778)
);

CKINVDCx5p33_ASAP7_75t_R g1779 ( 
.A(n_1420),
.Y(n_1779)
);

CKINVDCx5p33_ASAP7_75t_R g1780 ( 
.A(n_1423),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1267),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1289),
.Y(n_1782)
);

CKINVDCx5p33_ASAP7_75t_R g1783 ( 
.A(n_1423),
.Y(n_1783)
);

INVxp33_ASAP7_75t_L g1784 ( 
.A(n_1221),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1290),
.Y(n_1785)
);

INVxp67_ASAP7_75t_L g1786 ( 
.A(n_1506),
.Y(n_1786)
);

CKINVDCx20_ASAP7_75t_R g1787 ( 
.A(n_1520),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1529),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1291),
.Y(n_1789)
);

CKINVDCx20_ASAP7_75t_R g1790 ( 
.A(n_1529),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1293),
.Y(n_1791)
);

CKINVDCx20_ASAP7_75t_R g1792 ( 
.A(n_1542),
.Y(n_1792)
);

CKINVDCx20_ASAP7_75t_R g1793 ( 
.A(n_1542),
.Y(n_1793)
);

XNOR2xp5_ASAP7_75t_L g1794 ( 
.A(n_1553),
.B(n_1574),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1295),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1430),
.Y(n_1796)
);

CKINVDCx20_ASAP7_75t_R g1797 ( 
.A(n_1553),
.Y(n_1797)
);

INVxp33_ASAP7_75t_SL g1798 ( 
.A(n_1259),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1296),
.Y(n_1799)
);

CKINVDCx20_ASAP7_75t_R g1800 ( 
.A(n_1574),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1299),
.Y(n_1801)
);

CKINVDCx5p33_ASAP7_75t_R g1802 ( 
.A(n_1430),
.Y(n_1802)
);

CKINVDCx5p33_ASAP7_75t_R g1803 ( 
.A(n_1443),
.Y(n_1803)
);

CKINVDCx16_ASAP7_75t_R g1804 ( 
.A(n_1361),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1301),
.Y(n_1805)
);

INVx1_ASAP7_75t_SL g1806 ( 
.A(n_1245),
.Y(n_1806)
);

CKINVDCx16_ASAP7_75t_R g1807 ( 
.A(n_1390),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1303),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1306),
.Y(n_1809)
);

INVxp67_ASAP7_75t_SL g1810 ( 
.A(n_1588),
.Y(n_1810)
);

INVxp67_ASAP7_75t_L g1811 ( 
.A(n_1507),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1307),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1308),
.Y(n_1813)
);

CKINVDCx5p33_ASAP7_75t_R g1814 ( 
.A(n_1443),
.Y(n_1814)
);

CKINVDCx5p33_ASAP7_75t_R g1815 ( 
.A(n_1448),
.Y(n_1815)
);

INVx2_ASAP7_75t_L g1816 ( 
.A(n_1469),
.Y(n_1816)
);

NOR2xp33_ASAP7_75t_L g1817 ( 
.A(n_1481),
.B(n_791),
.Y(n_1817)
);

CKINVDCx5p33_ASAP7_75t_R g1818 ( 
.A(n_1448),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1449),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1312),
.Y(n_1820)
);

CKINVDCx5p33_ASAP7_75t_R g1821 ( 
.A(n_1449),
.Y(n_1821)
);

CKINVDCx16_ASAP7_75t_R g1822 ( 
.A(n_1499),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1587),
.Y(n_1823)
);

INVxp67_ASAP7_75t_L g1824 ( 
.A(n_1526),
.Y(n_1824)
);

BUFx6f_ASAP7_75t_SL g1825 ( 
.A(n_1481),
.Y(n_1825)
);

CKINVDCx5p33_ASAP7_75t_R g1826 ( 
.A(n_1460),
.Y(n_1826)
);

CKINVDCx20_ASAP7_75t_R g1827 ( 
.A(n_1587),
.Y(n_1827)
);

CKINVDCx5p33_ASAP7_75t_R g1828 ( 
.A(n_1460),
.Y(n_1828)
);

CKINVDCx20_ASAP7_75t_R g1829 ( 
.A(n_1643),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1469),
.Y(n_1830)
);

INVx2_ASAP7_75t_L g1831 ( 
.A(n_1572),
.Y(n_1831)
);

INVxp67_ASAP7_75t_L g1832 ( 
.A(n_1472),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1313),
.Y(n_1833)
);

HB1xp67_ASAP7_75t_L g1834 ( 
.A(n_1267),
.Y(n_1834)
);

INVxp67_ASAP7_75t_SL g1835 ( 
.A(n_1599),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1474),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1314),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1358),
.Y(n_1838)
);

INVx1_ASAP7_75t_L g1839 ( 
.A(n_1363),
.Y(n_1839)
);

HB1xp67_ASAP7_75t_L g1840 ( 
.A(n_1281),
.Y(n_1840)
);

CKINVDCx20_ASAP7_75t_R g1841 ( 
.A(n_1643),
.Y(n_1841)
);

HB1xp67_ASAP7_75t_L g1842 ( 
.A(n_1281),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1365),
.Y(n_1843)
);

CKINVDCx20_ASAP7_75t_R g1844 ( 
.A(n_1253),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1366),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1369),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1632),
.B(n_813),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1372),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1373),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1374),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1376),
.Y(n_1851)
);

CKINVDCx5p33_ASAP7_75t_R g1852 ( 
.A(n_1474),
.Y(n_1852)
);

INVxp67_ASAP7_75t_L g1853 ( 
.A(n_1491),
.Y(n_1853)
);

CKINVDCx5p33_ASAP7_75t_R g1854 ( 
.A(n_1480),
.Y(n_1854)
);

CKINVDCx20_ASAP7_75t_R g1855 ( 
.A(n_1253),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1302),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1377),
.Y(n_1857)
);

CKINVDCx16_ASAP7_75t_R g1858 ( 
.A(n_1530),
.Y(n_1858)
);

NOR2xp33_ASAP7_75t_L g1859 ( 
.A(n_1632),
.B(n_1403),
.Y(n_1859)
);

CKINVDCx5p33_ASAP7_75t_R g1860 ( 
.A(n_1480),
.Y(n_1860)
);

CKINVDCx5p33_ASAP7_75t_R g1861 ( 
.A(n_1486),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1379),
.Y(n_1862)
);

CKINVDCx5p33_ASAP7_75t_R g1863 ( 
.A(n_1486),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1224),
.B(n_814),
.Y(n_1864)
);

CKINVDCx5p33_ASAP7_75t_R g1865 ( 
.A(n_1495),
.Y(n_1865)
);

CKINVDCx16_ASAP7_75t_R g1866 ( 
.A(n_1532),
.Y(n_1866)
);

CKINVDCx16_ASAP7_75t_R g1867 ( 
.A(n_1535),
.Y(n_1867)
);

CKINVDCx5p33_ASAP7_75t_R g1868 ( 
.A(n_1495),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1382),
.Y(n_1869)
);

CKINVDCx5p33_ASAP7_75t_R g1870 ( 
.A(n_1501),
.Y(n_1870)
);

CKINVDCx20_ASAP7_75t_R g1871 ( 
.A(n_1264),
.Y(n_1871)
);

NOR2xp67_ASAP7_75t_L g1872 ( 
.A(n_1501),
.B(n_1517),
.Y(n_1872)
);

CKINVDCx5p33_ASAP7_75t_R g1873 ( 
.A(n_1517),
.Y(n_1873)
);

CKINVDCx5p33_ASAP7_75t_R g1874 ( 
.A(n_1524),
.Y(n_1874)
);

OAI21x1_ASAP7_75t_L g1875 ( 
.A1(n_1223),
.A2(n_801),
.B(n_755),
.Y(n_1875)
);

CKINVDCx5p33_ASAP7_75t_R g1876 ( 
.A(n_1524),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1383),
.Y(n_1877)
);

BUFx3_ASAP7_75t_L g1878 ( 
.A(n_1396),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1384),
.Y(n_1879)
);

CKINVDCx20_ASAP7_75t_R g1880 ( 
.A(n_1264),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1386),
.Y(n_1881)
);

INVxp67_ASAP7_75t_L g1882 ( 
.A(n_1505),
.Y(n_1882)
);

INVxp33_ASAP7_75t_SL g1883 ( 
.A(n_1531),
.Y(n_1883)
);

INVxp67_ASAP7_75t_SL g1884 ( 
.A(n_1356),
.Y(n_1884)
);

CKINVDCx5p33_ASAP7_75t_R g1885 ( 
.A(n_1531),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1302),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1224),
.B(n_831),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1387),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1572),
.Y(n_1889)
);

CKINVDCx5p33_ASAP7_75t_R g1890 ( 
.A(n_1534),
.Y(n_1890)
);

NOR2xp67_ASAP7_75t_L g1891 ( 
.A(n_1534),
.B(n_836),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1388),
.Y(n_1892)
);

HB1xp67_ASAP7_75t_L g1893 ( 
.A(n_1327),
.Y(n_1893)
);

CKINVDCx16_ASAP7_75t_R g1894 ( 
.A(n_1557),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1389),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1391),
.Y(n_1896)
);

CKINVDCx5p33_ASAP7_75t_R g1897 ( 
.A(n_1325),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1393),
.Y(n_1898)
);

CKINVDCx5p33_ASAP7_75t_R g1899 ( 
.A(n_1538),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1597),
.Y(n_1900)
);

CKINVDCx5p33_ASAP7_75t_R g1901 ( 
.A(n_1538),
.Y(n_1901)
);

CKINVDCx20_ASAP7_75t_R g1902 ( 
.A(n_1269),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1394),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1327),
.Y(n_1904)
);

CKINVDCx20_ASAP7_75t_R g1905 ( 
.A(n_1269),
.Y(n_1905)
);

INVxp67_ASAP7_75t_SL g1906 ( 
.A(n_1362),
.Y(n_1906)
);

CKINVDCx20_ASAP7_75t_R g1907 ( 
.A(n_1278),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1572),
.Y(n_1908)
);

BUFx2_ASAP7_75t_L g1909 ( 
.A(n_1278),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1246),
.B(n_1294),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1395),
.Y(n_1911)
);

NAND2xp5_ASAP7_75t_L g1912 ( 
.A(n_1246),
.B(n_900),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1398),
.Y(n_1913)
);

NOR2xp67_ASAP7_75t_L g1914 ( 
.A(n_1540),
.B(n_915),
.Y(n_1914)
);

INVxp67_ASAP7_75t_L g1915 ( 
.A(n_1325),
.Y(n_1915)
);

CKINVDCx20_ASAP7_75t_R g1916 ( 
.A(n_1297),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1399),
.Y(n_1917)
);

NAND2xp5_ASAP7_75t_L g1918 ( 
.A(n_1246),
.B(n_924),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1572),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1540),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1400),
.Y(n_1921)
);

NOR2xp33_ASAP7_75t_R g1922 ( 
.A(n_1548),
.B(n_926),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1401),
.Y(n_1923)
);

CKINVDCx5p33_ASAP7_75t_R g1924 ( 
.A(n_1548),
.Y(n_1924)
);

INVxp67_ASAP7_75t_L g1925 ( 
.A(n_1247),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1246),
.B(n_948),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1402),
.Y(n_1927)
);

NOR2xp33_ASAP7_75t_L g1928 ( 
.A(n_1403),
.B(n_977),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1405),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1409),
.Y(n_1930)
);

NOR2xp33_ASAP7_75t_R g1931 ( 
.A(n_1549),
.B(n_996),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1435),
.B(n_1007),
.Y(n_1932)
);

CKINVDCx5p33_ASAP7_75t_R g1933 ( 
.A(n_1549),
.Y(n_1933)
);

CKINVDCx5p33_ASAP7_75t_R g1934 ( 
.A(n_1562),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1624),
.Y(n_1935)
);

INVxp67_ASAP7_75t_SL g1936 ( 
.A(n_1370),
.Y(n_1936)
);

INVxp67_ASAP7_75t_L g1937 ( 
.A(n_1342),
.Y(n_1937)
);

INVx1_ASAP7_75t_L g1938 ( 
.A(n_1412),
.Y(n_1938)
);

INVxp67_ASAP7_75t_SL g1939 ( 
.A(n_1429),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1558),
.B(n_999),
.Y(n_1940)
);

CKINVDCx5p33_ASAP7_75t_R g1941 ( 
.A(n_1562),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1624),
.Y(n_1942)
);

CKINVDCx5p33_ASAP7_75t_R g1943 ( 
.A(n_1575),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1413),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1624),
.Y(n_1945)
);

CKINVDCx20_ASAP7_75t_R g1946 ( 
.A(n_1297),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1414),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1415),
.Y(n_1948)
);

CKINVDCx5p33_ASAP7_75t_R g1949 ( 
.A(n_1575),
.Y(n_1949)
);

CKINVDCx5p33_ASAP7_75t_R g1950 ( 
.A(n_1612),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1418),
.Y(n_1951)
);

CKINVDCx5p33_ASAP7_75t_R g1952 ( 
.A(n_1612),
.Y(n_1952)
);

CKINVDCx20_ASAP7_75t_R g1953 ( 
.A(n_1298),
.Y(n_1953)
);

BUFx3_ASAP7_75t_L g1954 ( 
.A(n_1544),
.Y(n_1954)
);

CKINVDCx5p33_ASAP7_75t_R g1955 ( 
.A(n_1619),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1419),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1624),
.Y(n_1957)
);

INVxp67_ASAP7_75t_SL g1958 ( 
.A(n_1454),
.Y(n_1958)
);

INVxp33_ASAP7_75t_L g1959 ( 
.A(n_1309),
.Y(n_1959)
);

CKINVDCx20_ASAP7_75t_R g1960 ( 
.A(n_1298),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1421),
.Y(n_1961)
);

CKINVDCx5p33_ASAP7_75t_R g1962 ( 
.A(n_1619),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1424),
.Y(n_1963)
);

CKINVDCx5p33_ASAP7_75t_R g1964 ( 
.A(n_1622),
.Y(n_1964)
);

OR2x2_ASAP7_75t_L g1965 ( 
.A(n_1251),
.B(n_978),
.Y(n_1965)
);

INVxp67_ASAP7_75t_SL g1966 ( 
.A(n_1554),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1435),
.B(n_1009),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1425),
.Y(n_1968)
);

BUFx2_ASAP7_75t_L g1969 ( 
.A(n_1323),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1544),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1428),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_L g1972 ( 
.A(n_1246),
.B(n_1066),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1432),
.Y(n_1973)
);

CKINVDCx20_ASAP7_75t_R g1974 ( 
.A(n_1323),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1246),
.B(n_1077),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1433),
.Y(n_1976)
);

CKINVDCx5p33_ASAP7_75t_R g1977 ( 
.A(n_1622),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1623),
.Y(n_1978)
);

NOR2xp33_ASAP7_75t_L g1979 ( 
.A(n_1461),
.B(n_1105),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1461),
.B(n_1106),
.Y(n_1980)
);

CKINVDCx5p33_ASAP7_75t_R g1981 ( 
.A(n_1623),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_L g1982 ( 
.A(n_1477),
.B(n_1176),
.Y(n_1982)
);

BUFx2_ASAP7_75t_L g1983 ( 
.A(n_1696),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_L g1984 ( 
.A1(n_1760),
.A2(n_1316),
.B1(n_1591),
.B2(n_1563),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1723),
.Y(n_1985)
);

BUFx6f_ASAP7_75t_L g1986 ( 
.A(n_1954),
.Y(n_1986)
);

BUFx6f_ASAP7_75t_L g1987 ( 
.A(n_1954),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1959),
.B(n_1568),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1725),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1732),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_L g1991 ( 
.A(n_1656),
.B(n_1246),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1736),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1875),
.Y(n_1993)
);

AND2x2_ASAP7_75t_SL g1994 ( 
.A(n_1689),
.B(n_1359),
.Y(n_1994)
);

CKINVDCx5p33_ASAP7_75t_R g1995 ( 
.A(n_1701),
.Y(n_1995)
);

INVx6_ASAP7_75t_L g1996 ( 
.A(n_1708),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1970),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1748),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_L g1999 ( 
.A(n_1693),
.B(n_1294),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1678),
.B(n_1284),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1810),
.Y(n_2001)
);

INVx1_ASAP7_75t_L g2002 ( 
.A(n_1835),
.Y(n_2002)
);

CKINVDCx5p33_ASAP7_75t_R g2003 ( 
.A(n_1702),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1838),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1839),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1970),
.Y(n_2006)
);

CKINVDCx5p33_ASAP7_75t_R g2007 ( 
.A(n_1703),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1843),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1845),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_SL g2010 ( 
.A(n_1740),
.B(n_1294),
.Y(n_2010)
);

INVx2_ASAP7_75t_L g2011 ( 
.A(n_1875),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1959),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1658),
.B(n_1294),
.Y(n_2013)
);

BUFx6f_ASAP7_75t_L g2014 ( 
.A(n_1666),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1650),
.Y(n_2015)
);

INVx3_ASAP7_75t_L g2016 ( 
.A(n_1708),
.Y(n_2016)
);

CKINVDCx5p33_ASAP7_75t_R g2017 ( 
.A(n_1707),
.Y(n_2017)
);

INVx1_ASAP7_75t_L g2018 ( 
.A(n_1846),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1848),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1849),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1850),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_L g2022 ( 
.A(n_1685),
.B(n_1294),
.Y(n_2022)
);

NAND2xp5_ASAP7_75t_L g2023 ( 
.A(n_1687),
.B(n_1294),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1740),
.B(n_1294),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1851),
.Y(n_2025)
);

INVx2_ASAP7_75t_L g2026 ( 
.A(n_1650),
.Y(n_2026)
);

BUFx6f_ASAP7_75t_L g2027 ( 
.A(n_1666),
.Y(n_2027)
);

BUFx2_ASAP7_75t_L g2028 ( 
.A(n_1696),
.Y(n_2028)
);

AND2x6_ASAP7_75t_L g2029 ( 
.A(n_1673),
.B(n_1284),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1857),
.Y(n_2030)
);

NAND2xp33_ASAP7_75t_L g2031 ( 
.A(n_1693),
.B(n_1695),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1862),
.Y(n_2032)
);

XOR2x2_ASAP7_75t_L g2033 ( 
.A(n_1794),
.B(n_1477),
.Y(n_2033)
);

INVx1_ASAP7_75t_L g2034 ( 
.A(n_1869),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1877),
.Y(n_2035)
);

INVx6_ASAP7_75t_L g2036 ( 
.A(n_1878),
.Y(n_2036)
);

CKINVDCx20_ASAP7_75t_R g2037 ( 
.A(n_1645),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1879),
.Y(n_2038)
);

INVx2_ASAP7_75t_L g2039 ( 
.A(n_1672),
.Y(n_2039)
);

CKINVDCx5p33_ASAP7_75t_R g2040 ( 
.A(n_1647),
.Y(n_2040)
);

INVx3_ASAP7_75t_L g2041 ( 
.A(n_1878),
.Y(n_2041)
);

CKINVDCx20_ASAP7_75t_R g2042 ( 
.A(n_1645),
.Y(n_2042)
);

INVx4_ASAP7_75t_L g2043 ( 
.A(n_1695),
.Y(n_2043)
);

INVx1_ASAP7_75t_L g2044 ( 
.A(n_1881),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1672),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1691),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1691),
.Y(n_2047)
);

AND2x2_ASAP7_75t_L g2048 ( 
.A(n_1712),
.B(n_1309),
.Y(n_2048)
);

INVx2_ASAP7_75t_L g2049 ( 
.A(n_1733),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1888),
.Y(n_2050)
);

BUFx6f_ASAP7_75t_L g2051 ( 
.A(n_1666),
.Y(n_2051)
);

INVx1_ASAP7_75t_L g2052 ( 
.A(n_1892),
.Y(n_2052)
);

INVx2_ASAP7_75t_L g2053 ( 
.A(n_1733),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1895),
.Y(n_2054)
);

INVx1_ASAP7_75t_L g2055 ( 
.A(n_1896),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1688),
.B(n_1631),
.Y(n_2056)
);

HB1xp67_ASAP7_75t_L g2057 ( 
.A(n_1925),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1711),
.B(n_1585),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1898),
.Y(n_2059)
);

BUFx6f_ASAP7_75t_L g2060 ( 
.A(n_1666),
.Y(n_2060)
);

CKINVDCx5p33_ASAP7_75t_R g2061 ( 
.A(n_1654),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1903),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1911),
.Y(n_2063)
);

INVx3_ASAP7_75t_L g2064 ( 
.A(n_1644),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_L g2065 ( 
.A(n_1706),
.B(n_1315),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1720),
.B(n_1315),
.Y(n_2066)
);

INVx3_ASAP7_75t_L g2067 ( 
.A(n_1649),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1758),
.B(n_1347),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1913),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1753),
.Y(n_2070)
);

NAND2xp5_ASAP7_75t_L g2071 ( 
.A(n_1664),
.B(n_1347),
.Y(n_2071)
);

BUFx6f_ASAP7_75t_L g2072 ( 
.A(n_1694),
.Y(n_2072)
);

INVx3_ASAP7_75t_L g2073 ( 
.A(n_1651),
.Y(n_2073)
);

BUFx6f_ASAP7_75t_L g2074 ( 
.A(n_1694),
.Y(n_2074)
);

HB1xp67_ASAP7_75t_L g2075 ( 
.A(n_1730),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_1753),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1670),
.B(n_1364),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1711),
.B(n_1585),
.Y(n_2078)
);

AND2x2_ASAP7_75t_L g2079 ( 
.A(n_1786),
.B(n_1311),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1817),
.B(n_1364),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1917),
.Y(n_2081)
);

AND2x6_ASAP7_75t_L g2082 ( 
.A(n_1859),
.B(n_1483),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_1921),
.Y(n_2083)
);

AND2x2_ASAP7_75t_SL g2084 ( 
.A(n_1745),
.B(n_1528),
.Y(n_2084)
);

BUFx6f_ASAP7_75t_L g2085 ( 
.A(n_1694),
.Y(n_2085)
);

INVx1_ASAP7_75t_L g2086 ( 
.A(n_1923),
.Y(n_2086)
);

BUFx2_ASAP7_75t_L g2087 ( 
.A(n_1715),
.Y(n_2087)
);

BUFx6f_ASAP7_75t_L g2088 ( 
.A(n_1694),
.Y(n_2088)
);

BUFx2_ASAP7_75t_L g2089 ( 
.A(n_1719),
.Y(n_2089)
);

AND2x4_ASAP7_75t_L g2090 ( 
.A(n_1697),
.B(n_1631),
.Y(n_2090)
);

INVx2_ASAP7_75t_L g2091 ( 
.A(n_1764),
.Y(n_2091)
);

BUFx6f_ASAP7_75t_L g2092 ( 
.A(n_1741),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1847),
.B(n_1483),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1927),
.Y(n_2094)
);

BUFx6f_ASAP7_75t_L g2095 ( 
.A(n_1741),
.Y(n_2095)
);

INVx1_ASAP7_75t_L g2096 ( 
.A(n_1929),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_1660),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1930),
.Y(n_2098)
);

CKINVDCx5p33_ASAP7_75t_R g2099 ( 
.A(n_1710),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_1938),
.Y(n_2100)
);

HB1xp67_ASAP7_75t_L g2101 ( 
.A(n_1937),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1944),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_1947),
.Y(n_2103)
);

BUFx6f_ASAP7_75t_L g2104 ( 
.A(n_1741),
.Y(n_2104)
);

AND2x4_ASAP7_75t_L g2105 ( 
.A(n_1884),
.B(n_1509),
.Y(n_2105)
);

CKINVDCx5p33_ASAP7_75t_R g2106 ( 
.A(n_1714),
.Y(n_2106)
);

CKINVDCx5p33_ASAP7_75t_R g2107 ( 
.A(n_1661),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1948),
.Y(n_2108)
);

CKINVDCx5p33_ASAP7_75t_R g2109 ( 
.A(n_1663),
.Y(n_2109)
);

INVx1_ASAP7_75t_L g2110 ( 
.A(n_1951),
.Y(n_2110)
);

BUFx12f_ASAP7_75t_L g2111 ( 
.A(n_1897),
.Y(n_2111)
);

INVxp67_ASAP7_75t_L g2112 ( 
.A(n_1665),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_1760),
.B(n_1509),
.Y(n_2113)
);

INVx2_ASAP7_75t_L g2114 ( 
.A(n_1764),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1956),
.Y(n_2115)
);

INVx3_ASAP7_75t_L g2116 ( 
.A(n_1652),
.Y(n_2116)
);

HB1xp67_ASAP7_75t_L g2117 ( 
.A(n_1646),
.Y(n_2117)
);

INVx1_ASAP7_75t_L g2118 ( 
.A(n_1961),
.Y(n_2118)
);

HB1xp67_ASAP7_75t_L g2119 ( 
.A(n_1784),
.Y(n_2119)
);

NAND2xp5_ASAP7_75t_L g2120 ( 
.A(n_1671),
.B(n_1565),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1963),
.Y(n_2121)
);

AND2x2_ASAP7_75t_L g2122 ( 
.A(n_1811),
.B(n_1311),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1968),
.Y(n_2123)
);

CKINVDCx5p33_ASAP7_75t_R g2124 ( 
.A(n_1667),
.Y(n_2124)
);

INVx3_ASAP7_75t_L g2125 ( 
.A(n_1653),
.Y(n_2125)
);

BUFx6f_ASAP7_75t_L g2126 ( 
.A(n_1741),
.Y(n_2126)
);

NAND2xp5_ASAP7_75t_L g2127 ( 
.A(n_1906),
.B(n_1565),
.Y(n_2127)
);

CKINVDCx5p33_ASAP7_75t_R g2128 ( 
.A(n_1897),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_1655),
.Y(n_2129)
);

INVx1_ASAP7_75t_L g2130 ( 
.A(n_1971),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_1773),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_1973),
.Y(n_2132)
);

NAND2xp33_ASAP7_75t_R g2133 ( 
.A(n_1668),
.B(n_1626),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_1773),
.Y(n_2134)
);

OAI22xp5_ASAP7_75t_SL g2135 ( 
.A1(n_1844),
.A2(n_1015),
.B1(n_1020),
.B2(n_989),
.Y(n_2135)
);

AND2x4_ASAP7_75t_L g2136 ( 
.A(n_1936),
.B(n_1596),
.Y(n_2136)
);

BUFx6f_ASAP7_75t_L g2137 ( 
.A(n_1816),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1816),
.Y(n_2138)
);

CKINVDCx16_ASAP7_75t_R g2139 ( 
.A(n_1804),
.Y(n_2139)
);

CKINVDCx20_ASAP7_75t_R g2140 ( 
.A(n_1657),
.Y(n_2140)
);

CKINVDCx16_ASAP7_75t_R g2141 ( 
.A(n_1807),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1976),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1659),
.Y(n_2143)
);

AND2x4_ASAP7_75t_L g2144 ( 
.A(n_1939),
.B(n_1596),
.Y(n_2144)
);

BUFx2_ASAP7_75t_L g2145 ( 
.A(n_1722),
.Y(n_2145)
);

AND2x4_ASAP7_75t_L g2146 ( 
.A(n_1958),
.B(n_1966),
.Y(n_2146)
);

NOR2xp33_ASAP7_75t_SL g2147 ( 
.A(n_1798),
.B(n_1718),
.Y(n_2147)
);

INVxp33_ASAP7_75t_L g2148 ( 
.A(n_1784),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_1669),
.Y(n_2149)
);

OAI21x1_ASAP7_75t_L g2150 ( 
.A1(n_1910),
.A2(n_1243),
.B(n_1223),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_1824),
.B(n_1320),
.Y(n_2151)
);

CKINVDCx16_ASAP7_75t_R g2152 ( 
.A(n_1822),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1692),
.B(n_1609),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1743),
.B(n_1609),
.Y(n_2154)
);

INVx2_ASAP7_75t_L g2155 ( 
.A(n_1830),
.Y(n_2155)
);

CKINVDCx5p33_ASAP7_75t_R g2156 ( 
.A(n_1680),
.Y(n_2156)
);

AND2x4_ASAP7_75t_L g2157 ( 
.A(n_1698),
.B(n_1620),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_1700),
.B(n_1620),
.Y(n_2158)
);

OAI22xp5_ASAP7_75t_L g2159 ( 
.A1(n_1928),
.A2(n_1618),
.B1(n_1606),
.B2(n_1310),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_1674),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_1675),
.Y(n_2161)
);

AND2x2_ASAP7_75t_L g2162 ( 
.A(n_1832),
.B(n_1320),
.Y(n_2162)
);

NAND2xp5_ASAP7_75t_L g2163 ( 
.A(n_1932),
.B(n_1626),
.Y(n_2163)
);

HB1xp67_ASAP7_75t_L g2164 ( 
.A(n_1781),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1967),
.B(n_1629),
.Y(n_2165)
);

INVx3_ASAP7_75t_L g2166 ( 
.A(n_1676),
.Y(n_2166)
);

CKINVDCx20_ASAP7_75t_R g2167 ( 
.A(n_1657),
.Y(n_2167)
);

BUFx6f_ASAP7_75t_L g2168 ( 
.A(n_1830),
.Y(n_2168)
);

INVx2_ASAP7_75t_L g2169 ( 
.A(n_1831),
.Y(n_2169)
);

BUFx6f_ASAP7_75t_L g2170 ( 
.A(n_1831),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_1679),
.Y(n_2171)
);

INVx1_ASAP7_75t_L g2172 ( 
.A(n_1681),
.Y(n_2172)
);

INVx2_ASAP7_75t_L g2173 ( 
.A(n_1889),
.Y(n_2173)
);

INVx3_ASAP7_75t_L g2174 ( 
.A(n_1684),
.Y(n_2174)
);

INVx1_ASAP7_75t_L g2175 ( 
.A(n_1690),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_1979),
.B(n_1629),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_1705),
.Y(n_2177)
);

INVx1_ASAP7_75t_L g2178 ( 
.A(n_1709),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_1889),
.Y(n_2179)
);

CKINVDCx16_ASAP7_75t_R g2180 ( 
.A(n_1858),
.Y(n_2180)
);

INVx1_ASAP7_75t_L g2181 ( 
.A(n_1717),
.Y(n_2181)
);

BUFx3_ASAP7_75t_L g2182 ( 
.A(n_1721),
.Y(n_2182)
);

INVx1_ASAP7_75t_L g2183 ( 
.A(n_1726),
.Y(n_2183)
);

INVx2_ASAP7_75t_L g2184 ( 
.A(n_1908),
.Y(n_2184)
);

INVx1_ASAP7_75t_L g2185 ( 
.A(n_1728),
.Y(n_2185)
);

INVx1_ASAP7_75t_L g2186 ( 
.A(n_1735),
.Y(n_2186)
);

CKINVDCx5p33_ASAP7_75t_R g2187 ( 
.A(n_1686),
.Y(n_2187)
);

OAI22x1_ASAP7_75t_SL g2188 ( 
.A1(n_1662),
.A2(n_1047),
.B1(n_1092),
.B2(n_1032),
.Y(n_2188)
);

OA21x2_ASAP7_75t_L g2189 ( 
.A1(n_1912),
.A2(n_1254),
.B(n_1243),
.Y(n_2189)
);

INVx2_ASAP7_75t_L g2190 ( 
.A(n_1908),
.Y(n_2190)
);

INVx2_ASAP7_75t_L g2191 ( 
.A(n_1919),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_1980),
.B(n_1639),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1737),
.Y(n_2193)
);

AND2x4_ASAP7_75t_L g2194 ( 
.A(n_1746),
.B(n_1410),
.Y(n_2194)
);

OAI21x1_ASAP7_75t_L g2195 ( 
.A1(n_1918),
.A2(n_1280),
.B(n_1254),
.Y(n_2195)
);

NAND2xp5_ASAP7_75t_L g2196 ( 
.A(n_1982),
.B(n_1639),
.Y(n_2196)
);

BUFx6f_ASAP7_75t_SL g2197 ( 
.A(n_1866),
.Y(n_2197)
);

AND2x4_ASAP7_75t_L g2198 ( 
.A(n_1751),
.B(n_1508),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_1965),
.Y(n_2199)
);

AND2x4_ASAP7_75t_L g2200 ( 
.A(n_1755),
.B(n_1527),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_L g2201 ( 
.A(n_1864),
.B(n_1640),
.Y(n_2201)
);

NAND2xp5_ASAP7_75t_SL g2202 ( 
.A(n_1922),
.B(n_1640),
.Y(n_2202)
);

HB1xp67_ASAP7_75t_L g2203 ( 
.A(n_1699),
.Y(n_2203)
);

CKINVDCx20_ASAP7_75t_R g2204 ( 
.A(n_1662),
.Y(n_2204)
);

INVx3_ASAP7_75t_L g2205 ( 
.A(n_1759),
.Y(n_2205)
);

BUFx2_ASAP7_75t_L g2206 ( 
.A(n_1724),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1887),
.B(n_1766),
.Y(n_2207)
);

BUFx2_ASAP7_75t_L g2208 ( 
.A(n_1727),
.Y(n_2208)
);

INVx4_ASAP7_75t_L g2209 ( 
.A(n_1825),
.Y(n_2209)
);

INVx4_ASAP7_75t_L g2210 ( 
.A(n_1825),
.Y(n_2210)
);

AND2x6_ASAP7_75t_L g2211 ( 
.A(n_1763),
.B(n_1584),
.Y(n_2211)
);

BUFx8_ASAP7_75t_L g2212 ( 
.A(n_1909),
.Y(n_2212)
);

INVx3_ASAP7_75t_L g2213 ( 
.A(n_1761),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_1762),
.B(n_1765),
.Y(n_2214)
);

HB1xp67_ASAP7_75t_L g2215 ( 
.A(n_1738),
.Y(n_2215)
);

HB1xp67_ASAP7_75t_L g2216 ( 
.A(n_1739),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1767),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_1768),
.B(n_1533),
.Y(n_2218)
);

CKINVDCx20_ASAP7_75t_R g2219 ( 
.A(n_1677),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1772),
.Y(n_2220)
);

INVx2_ASAP7_75t_L g2221 ( 
.A(n_1919),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1782),
.Y(n_2222)
);

CKINVDCx5p33_ASAP7_75t_R g2223 ( 
.A(n_1747),
.Y(n_2223)
);

INVx3_ASAP7_75t_L g2224 ( 
.A(n_1785),
.Y(n_2224)
);

INVx2_ASAP7_75t_L g2225 ( 
.A(n_1935),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_1789),
.Y(n_2226)
);

CKINVDCx5p33_ASAP7_75t_R g2227 ( 
.A(n_1749),
.Y(n_2227)
);

AND2x4_ASAP7_75t_L g2228 ( 
.A(n_1791),
.B(n_1621),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_1853),
.B(n_1304),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_1795),
.B(n_1343),
.Y(n_2230)
);

AND2x4_ASAP7_75t_L g2231 ( 
.A(n_1799),
.B(n_1627),
.Y(n_2231)
);

NOR2xp33_ASAP7_75t_L g2232 ( 
.A(n_1825),
.B(n_1417),
.Y(n_2232)
);

AND3x1_ASAP7_75t_L g2233 ( 
.A(n_1744),
.B(n_981),
.C(n_980),
.Y(n_2233)
);

INVx3_ASAP7_75t_L g2234 ( 
.A(n_1801),
.Y(n_2234)
);

BUFx3_ASAP7_75t_L g2235 ( 
.A(n_1805),
.Y(n_2235)
);

BUFx6f_ASAP7_75t_L g2236 ( 
.A(n_1935),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1808),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1809),
.Y(n_2238)
);

INVx1_ASAP7_75t_L g2239 ( 
.A(n_1812),
.Y(n_2239)
);

BUFx2_ASAP7_75t_L g2240 ( 
.A(n_1752),
.Y(n_2240)
);

AND2x2_ASAP7_75t_L g2241 ( 
.A(n_1882),
.B(n_1304),
.Y(n_2241)
);

AND2x2_ASAP7_75t_L g2242 ( 
.A(n_1900),
.B(n_1417),
.Y(n_2242)
);

CKINVDCx5p33_ASAP7_75t_R g2243 ( 
.A(n_1754),
.Y(n_2243)
);

BUFx6f_ASAP7_75t_L g2244 ( 
.A(n_1942),
.Y(n_2244)
);

INVx2_ASAP7_75t_L g2245 ( 
.A(n_1942),
.Y(n_2245)
);

INVx2_ASAP7_75t_L g2246 ( 
.A(n_1945),
.Y(n_2246)
);

INVx1_ASAP7_75t_L g2247 ( 
.A(n_1813),
.Y(n_2247)
);

AND2x4_ASAP7_75t_L g2248 ( 
.A(n_1820),
.B(n_1633),
.Y(n_2248)
);

INVx1_ASAP7_75t_L g2249 ( 
.A(n_1833),
.Y(n_2249)
);

BUFx2_ASAP7_75t_L g2250 ( 
.A(n_1770),
.Y(n_2250)
);

INVx2_ASAP7_75t_L g2251 ( 
.A(n_1945),
.Y(n_2251)
);

CKINVDCx5p33_ASAP7_75t_R g2252 ( 
.A(n_1774),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_1837),
.Y(n_2253)
);

INVx2_ASAP7_75t_L g2254 ( 
.A(n_1957),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1957),
.Y(n_2255)
);

INVx1_ASAP7_75t_L g2256 ( 
.A(n_1891),
.Y(n_2256)
);

BUFx6f_ASAP7_75t_L g2257 ( 
.A(n_1926),
.Y(n_2257)
);

INVx2_ASAP7_75t_L g2258 ( 
.A(n_1972),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1914),
.B(n_1444),
.Y(n_2259)
);

BUFx6f_ASAP7_75t_L g2260 ( 
.A(n_1975),
.Y(n_2260)
);

NAND2xp5_ASAP7_75t_L g2261 ( 
.A(n_1931),
.B(n_1872),
.Y(n_2261)
);

INVx1_ASAP7_75t_L g2262 ( 
.A(n_1940),
.Y(n_2262)
);

AND2x4_ASAP7_75t_L g2263 ( 
.A(n_1756),
.B(n_1634),
.Y(n_2263)
);

BUFx6f_ASAP7_75t_L g2264 ( 
.A(n_1777),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_1834),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_1840),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_1842),
.B(n_1444),
.Y(n_2267)
);

NOR2xp33_ASAP7_75t_L g2268 ( 
.A(n_1883),
.B(n_1625),
.Y(n_2268)
);

INVx3_ASAP7_75t_L g2269 ( 
.A(n_1778),
.Y(n_2269)
);

CKINVDCx20_ASAP7_75t_R g2270 ( 
.A(n_1677),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1856),
.Y(n_2271)
);

INVx1_ASAP7_75t_L g2272 ( 
.A(n_1886),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_1981),
.B(n_1625),
.Y(n_2273)
);

AND2x6_ASAP7_75t_L g2274 ( 
.A(n_1806),
.B(n_755),
.Y(n_2274)
);

INVx1_ASAP7_75t_L g2275 ( 
.A(n_1893),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1904),
.Y(n_2276)
);

CKINVDCx5p33_ASAP7_75t_R g2277 ( 
.A(n_1779),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1780),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_1783),
.Y(n_2279)
);

CKINVDCx20_ASAP7_75t_R g2280 ( 
.A(n_1682),
.Y(n_2280)
);

INVx3_ASAP7_75t_L g2281 ( 
.A(n_1796),
.Y(n_2281)
);

CKINVDCx5p33_ASAP7_75t_R g2282 ( 
.A(n_1802),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_1803),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_1814),
.Y(n_2284)
);

AND2x2_ASAP7_75t_L g2285 ( 
.A(n_1815),
.B(n_1305),
.Y(n_2285)
);

OAI21x1_ASAP7_75t_L g2286 ( 
.A1(n_1718),
.A2(n_1287),
.B(n_1280),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_1818),
.Y(n_2287)
);

CKINVDCx5p33_ASAP7_75t_R g2288 ( 
.A(n_1819),
.Y(n_2288)
);

BUFx6f_ASAP7_75t_L g2289 ( 
.A(n_1821),
.Y(n_2289)
);

AND2x6_ASAP7_75t_L g2290 ( 
.A(n_1883),
.B(n_801),
.Y(n_2290)
);

CKINVDCx20_ASAP7_75t_R g2291 ( 
.A(n_1682),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1826),
.Y(n_2292)
);

AND2x6_ASAP7_75t_L g2293 ( 
.A(n_1867),
.B(n_966),
.Y(n_2293)
);

CKINVDCx5p33_ASAP7_75t_R g2294 ( 
.A(n_1828),
.Y(n_2294)
);

INVx3_ASAP7_75t_L g2295 ( 
.A(n_1836),
.Y(n_2295)
);

CKINVDCx5p33_ASAP7_75t_R g2296 ( 
.A(n_1852),
.Y(n_2296)
);

NOR2x1_ASAP7_75t_L g2297 ( 
.A(n_1648),
.B(n_1608),
.Y(n_2297)
);

INVx3_ASAP7_75t_L g2298 ( 
.A(n_1854),
.Y(n_2298)
);

AND2x2_ASAP7_75t_SL g2299 ( 
.A(n_1894),
.B(n_1013),
.Y(n_2299)
);

BUFx6f_ASAP7_75t_L g2300 ( 
.A(n_1860),
.Y(n_2300)
);

NAND2xp5_ASAP7_75t_SL g2301 ( 
.A(n_1861),
.B(n_1863),
.Y(n_2301)
);

INVx3_ASAP7_75t_L g2302 ( 
.A(n_1865),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1868),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1870),
.Y(n_2304)
);

INVx1_ASAP7_75t_L g2305 ( 
.A(n_1873),
.Y(n_2305)
);

BUFx3_ASAP7_75t_L g2306 ( 
.A(n_1874),
.Y(n_2306)
);

INVx1_ASAP7_75t_L g2307 ( 
.A(n_1876),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_1885),
.Y(n_2308)
);

INVx1_ASAP7_75t_L g2309 ( 
.A(n_1890),
.Y(n_2309)
);

INVx1_ASAP7_75t_L g2310 ( 
.A(n_1899),
.Y(n_2310)
);

HB1xp67_ASAP7_75t_L g2311 ( 
.A(n_1901),
.Y(n_2311)
);

BUFx3_ASAP7_75t_L g2312 ( 
.A(n_1920),
.Y(n_2312)
);

BUFx8_ASAP7_75t_L g2313 ( 
.A(n_1969),
.Y(n_2313)
);

OAI22xp5_ASAP7_75t_L g2314 ( 
.A1(n_1924),
.A2(n_1341),
.B1(n_1211),
.B2(n_1157),
.Y(n_2314)
);

INVx2_ASAP7_75t_L g2315 ( 
.A(n_1933),
.Y(n_2315)
);

AOI22xp5_ASAP7_75t_L g2316 ( 
.A1(n_1934),
.A2(n_873),
.B1(n_913),
.B2(n_803),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1941),
.Y(n_2317)
);

AND2x4_ASAP7_75t_L g2318 ( 
.A(n_1943),
.B(n_1617),
.Y(n_2318)
);

BUFx2_ASAP7_75t_L g2319 ( 
.A(n_1949),
.Y(n_2319)
);

CKINVDCx20_ASAP7_75t_R g2320 ( 
.A(n_1683),
.Y(n_2320)
);

INVx1_ASAP7_75t_L g2321 ( 
.A(n_1950),
.Y(n_2321)
);

BUFx2_ASAP7_75t_L g2322 ( 
.A(n_1952),
.Y(n_2322)
);

CKINVDCx20_ASAP7_75t_R g2323 ( 
.A(n_1683),
.Y(n_2323)
);

OAI22xp5_ASAP7_75t_SL g2324 ( 
.A1(n_1844),
.A2(n_1123),
.B1(n_1135),
.B2(n_1070),
.Y(n_2324)
);

INVx4_ASAP7_75t_L g2325 ( 
.A(n_1955),
.Y(n_2325)
);

INVx1_ASAP7_75t_L g2326 ( 
.A(n_1962),
.Y(n_2326)
);

NOR2x1_ASAP7_75t_L g2327 ( 
.A(n_1729),
.B(n_1637),
.Y(n_2327)
);

OAI22xp5_ASAP7_75t_SL g2328 ( 
.A1(n_1855),
.A2(n_1198),
.B1(n_969),
.B2(n_990),
.Y(n_2328)
);

HB1xp67_ASAP7_75t_L g2329 ( 
.A(n_1964),
.Y(n_2329)
);

INVx2_ASAP7_75t_L g2330 ( 
.A(n_1977),
.Y(n_2330)
);

INVx1_ASAP7_75t_L g2331 ( 
.A(n_1978),
.Y(n_2331)
);

INVx1_ASAP7_75t_L g2332 ( 
.A(n_1798),
.Y(n_2332)
);

NAND3xp33_ASAP7_75t_L g2333 ( 
.A(n_1915),
.B(n_799),
.C(n_798),
.Y(n_2333)
);

BUFx2_ASAP7_75t_L g2334 ( 
.A(n_1855),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_1771),
.Y(n_2335)
);

INVx2_ASAP7_75t_L g2336 ( 
.A(n_1871),
.Y(n_2336)
);

BUFx6f_ASAP7_75t_L g2337 ( 
.A(n_1871),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_1880),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1880),
.Y(n_2339)
);

CKINVDCx20_ASAP7_75t_R g2340 ( 
.A(n_1704),
.Y(n_2340)
);

AND2x4_ASAP7_75t_L g2341 ( 
.A(n_1902),
.B(n_1605),
.Y(n_2341)
);

BUFx6f_ASAP7_75t_L g2342 ( 
.A(n_1902),
.Y(n_2342)
);

NAND2xp5_ASAP7_75t_L g2343 ( 
.A(n_1905),
.B(n_1287),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1905),
.Y(n_2344)
);

INVx2_ASAP7_75t_L g2345 ( 
.A(n_1907),
.Y(n_2345)
);

OAI21x1_ASAP7_75t_L g2346 ( 
.A1(n_1907),
.A2(n_1328),
.B(n_1300),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_1916),
.Y(n_2347)
);

AND2x4_ASAP7_75t_L g2348 ( 
.A(n_1916),
.B(n_1611),
.Y(n_2348)
);

CKINVDCx5p33_ASAP7_75t_R g2349 ( 
.A(n_1946),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_1946),
.B(n_1436),
.Y(n_2350)
);

OAI22xp5_ASAP7_75t_SL g2351 ( 
.A1(n_1953),
.A2(n_1084),
.B1(n_1086),
.B2(n_917),
.Y(n_2351)
);

CKINVDCx5p33_ASAP7_75t_R g2352 ( 
.A(n_1704),
.Y(n_2352)
);

NAND2x1_ASAP7_75t_L g2353 ( 
.A(n_1953),
.B(n_1544),
.Y(n_2353)
);

OAI22xp5_ASAP7_75t_L g2354 ( 
.A1(n_1960),
.A2(n_1108),
.B1(n_952),
.B2(n_806),
.Y(n_2354)
);

HB1xp67_ASAP7_75t_L g2355 ( 
.A(n_1960),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_L g2356 ( 
.A(n_1974),
.B(n_1300),
.Y(n_2356)
);

BUFx2_ASAP7_75t_L g2357 ( 
.A(n_1974),
.Y(n_2357)
);

INVx2_ASAP7_75t_L g2358 ( 
.A(n_1713),
.Y(n_2358)
);

BUFx2_ASAP7_75t_L g2359 ( 
.A(n_1713),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_1716),
.B(n_1328),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_1716),
.Y(n_2361)
);

AND2x2_ASAP7_75t_L g2362 ( 
.A(n_1731),
.B(n_1439),
.Y(n_2362)
);

INVx2_ASAP7_75t_L g2363 ( 
.A(n_1731),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_1734),
.Y(n_2364)
);

CKINVDCx5p33_ASAP7_75t_R g2365 ( 
.A(n_1734),
.Y(n_2365)
);

INVx1_ASAP7_75t_L g2366 ( 
.A(n_1742),
.Y(n_2366)
);

CKINVDCx5p33_ASAP7_75t_R g2367 ( 
.A(n_1742),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_1750),
.Y(n_2368)
);

BUFx2_ASAP7_75t_L g2369 ( 
.A(n_1750),
.Y(n_2369)
);

INVx1_ASAP7_75t_L g2370 ( 
.A(n_1757),
.Y(n_2370)
);

INVx1_ASAP7_75t_L g2371 ( 
.A(n_1757),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_L g2372 ( 
.A(n_1769),
.B(n_1340),
.Y(n_2372)
);

AND2x2_ASAP7_75t_L g2373 ( 
.A(n_1769),
.B(n_1440),
.Y(n_2373)
);

BUFx6f_ASAP7_75t_L g2374 ( 
.A(n_1775),
.Y(n_2374)
);

NAND2xp5_ASAP7_75t_L g2375 ( 
.A(n_1775),
.B(n_1340),
.Y(n_2375)
);

AND2x2_ASAP7_75t_L g2376 ( 
.A(n_1776),
.B(n_1441),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_1776),
.B(n_1350),
.Y(n_2377)
);

INVx1_ASAP7_75t_L g2378 ( 
.A(n_2177),
.Y(n_2378)
);

BUFx6f_ASAP7_75t_L g2379 ( 
.A(n_1986),
.Y(n_2379)
);

INVx2_ASAP7_75t_L g2380 ( 
.A(n_2006),
.Y(n_2380)
);

OAI22xp5_ASAP7_75t_L g2381 ( 
.A1(n_2163),
.A2(n_807),
.B1(n_808),
.B2(n_800),
.Y(n_2381)
);

BUFx6f_ASAP7_75t_L g2382 ( 
.A(n_1986),
.Y(n_2382)
);

INVx1_ASAP7_75t_L g2383 ( 
.A(n_2178),
.Y(n_2383)
);

INVx2_ASAP7_75t_L g2384 ( 
.A(n_2006),
.Y(n_2384)
);

BUFx6f_ASAP7_75t_L g2385 ( 
.A(n_1986),
.Y(n_2385)
);

INVx1_ASAP7_75t_L g2386 ( 
.A(n_2181),
.Y(n_2386)
);

INVx1_ASAP7_75t_L g2387 ( 
.A(n_2183),
.Y(n_2387)
);

INVx1_ASAP7_75t_L g2388 ( 
.A(n_2185),
.Y(n_2388)
);

INVx1_ASAP7_75t_L g2389 ( 
.A(n_2186),
.Y(n_2389)
);

INVx2_ASAP7_75t_L g2390 ( 
.A(n_1997),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_2193),
.Y(n_2391)
);

INVx2_ASAP7_75t_L g2392 ( 
.A(n_1997),
.Y(n_2392)
);

INVx1_ASAP7_75t_L g2393 ( 
.A(n_2217),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2220),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2015),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2082),
.B(n_878),
.Y(n_2396)
);

INVx1_ASAP7_75t_L g2397 ( 
.A(n_2222),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2015),
.Y(n_2398)
);

CKINVDCx8_ASAP7_75t_R g2399 ( 
.A(n_2139),
.Y(n_2399)
);

INVx1_ASAP7_75t_L g2400 ( 
.A(n_2226),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2237),
.Y(n_2401)
);

INVx2_ASAP7_75t_L g2402 ( 
.A(n_2026),
.Y(n_2402)
);

INVx2_ASAP7_75t_L g2403 ( 
.A(n_2026),
.Y(n_2403)
);

BUFx8_ASAP7_75t_L g2404 ( 
.A(n_2197),
.Y(n_2404)
);

CKINVDCx8_ASAP7_75t_R g2405 ( 
.A(n_2141),
.Y(n_2405)
);

AND2x2_ASAP7_75t_L g2406 ( 
.A(n_2242),
.B(n_1442),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2267),
.B(n_1445),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2238),
.Y(n_2408)
);

INVx2_ASAP7_75t_L g2409 ( 
.A(n_2039),
.Y(n_2409)
);

BUFx6f_ASAP7_75t_L g2410 ( 
.A(n_1986),
.Y(n_2410)
);

INVx1_ASAP7_75t_L g2411 ( 
.A(n_2239),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2247),
.Y(n_2412)
);

INVx1_ASAP7_75t_L g2413 ( 
.A(n_2249),
.Y(n_2413)
);

NAND2x1p5_ASAP7_75t_L g2414 ( 
.A(n_2209),
.B(n_1317),
.Y(n_2414)
);

OAI22xp5_ASAP7_75t_SL g2415 ( 
.A1(n_2037),
.A2(n_1787),
.B1(n_1790),
.B2(n_1788),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_2253),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_SL g2417 ( 
.A(n_1991),
.B(n_920),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2039),
.Y(n_2418)
);

BUFx2_ASAP7_75t_L g2419 ( 
.A(n_2187),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_2004),
.Y(n_2420)
);

AND2x2_ASAP7_75t_L g2421 ( 
.A(n_2229),
.B(n_1446),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2005),
.Y(n_2422)
);

OA21x2_ASAP7_75t_L g2423 ( 
.A1(n_2011),
.A2(n_1350),
.B(n_1375),
.Y(n_2423)
);

BUFx6f_ASAP7_75t_L g2424 ( 
.A(n_1987),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2045),
.Y(n_2425)
);

INVx1_ASAP7_75t_L g2426 ( 
.A(n_2008),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2082),
.B(n_890),
.Y(n_2427)
);

INVx1_ASAP7_75t_L g2428 ( 
.A(n_2009),
.Y(n_2428)
);

INVx2_ASAP7_75t_L g2429 ( 
.A(n_2045),
.Y(n_2429)
);

INVx1_ASAP7_75t_L g2430 ( 
.A(n_2018),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2019),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2020),
.Y(n_2432)
);

INVx2_ASAP7_75t_L g2433 ( 
.A(n_2046),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_2021),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2025),
.Y(n_2435)
);

AOI22xp5_ASAP7_75t_L g2436 ( 
.A1(n_2290),
.A2(n_1096),
.B1(n_893),
.B2(n_901),
.Y(n_2436)
);

AND2x2_ASAP7_75t_L g2437 ( 
.A(n_2241),
.B(n_1450),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2030),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2046),
.Y(n_2439)
);

INVx1_ASAP7_75t_L g2440 ( 
.A(n_2032),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2082),
.B(n_890),
.Y(n_2441)
);

INVx1_ASAP7_75t_L g2442 ( 
.A(n_2034),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2035),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_2038),
.Y(n_2444)
);

BUFx2_ASAP7_75t_L g2445 ( 
.A(n_2187),
.Y(n_2445)
);

BUFx2_ASAP7_75t_L g2446 ( 
.A(n_2352),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2044),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_2047),
.Y(n_2448)
);

INVx2_ASAP7_75t_L g2449 ( 
.A(n_2047),
.Y(n_2449)
);

INVx1_ASAP7_75t_L g2450 ( 
.A(n_2050),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2082),
.B(n_2113),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2052),
.Y(n_2452)
);

BUFx2_ASAP7_75t_L g2453 ( 
.A(n_2365),
.Y(n_2453)
);

INVx2_ASAP7_75t_L g2454 ( 
.A(n_2049),
.Y(n_2454)
);

INVx1_ASAP7_75t_L g2455 ( 
.A(n_2054),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_L g2456 ( 
.A(n_2082),
.B(n_2071),
.Y(n_2456)
);

INVx3_ASAP7_75t_L g2457 ( 
.A(n_1987),
.Y(n_2457)
);

INVx3_ASAP7_75t_L g2458 ( 
.A(n_1987),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_SL g2459 ( 
.A(n_2013),
.B(n_920),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2077),
.B(n_893),
.Y(n_2460)
);

INVx2_ASAP7_75t_L g2461 ( 
.A(n_2049),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2055),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2059),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_2062),
.Y(n_2464)
);

BUFx6f_ASAP7_75t_L g2465 ( 
.A(n_1987),
.Y(n_2465)
);

BUFx6f_ASAP7_75t_L g2466 ( 
.A(n_1993),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2053),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2000),
.B(n_1452),
.Y(n_2468)
);

INVxp67_ASAP7_75t_L g2469 ( 
.A(n_2203),
.Y(n_2469)
);

HB1xp67_ASAP7_75t_L g2470 ( 
.A(n_2012),
.Y(n_2470)
);

NAND2xp5_ASAP7_75t_L g2471 ( 
.A(n_2065),
.B(n_901),
.Y(n_2471)
);

INVx2_ASAP7_75t_L g2472 ( 
.A(n_2053),
.Y(n_2472)
);

NAND2xp5_ASAP7_75t_SL g2473 ( 
.A(n_2268),
.B(n_920),
.Y(n_2473)
);

INVx2_ASAP7_75t_L g2474 ( 
.A(n_2070),
.Y(n_2474)
);

NAND2xp5_ASAP7_75t_SL g2475 ( 
.A(n_2268),
.B(n_962),
.Y(n_2475)
);

NAND2xp5_ASAP7_75t_L g2476 ( 
.A(n_2066),
.B(n_1044),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2063),
.Y(n_2477)
);

INVx2_ASAP7_75t_L g2478 ( 
.A(n_2070),
.Y(n_2478)
);

INVx3_ASAP7_75t_L g2479 ( 
.A(n_1993),
.Y(n_2479)
);

NAND2xp33_ASAP7_75t_SL g2480 ( 
.A(n_2264),
.B(n_1044),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_SL g2481 ( 
.A(n_2107),
.B(n_2109),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_2069),
.Y(n_2482)
);

INVx2_ASAP7_75t_L g2483 ( 
.A(n_2076),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2081),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2083),
.Y(n_2485)
);

INVxp67_ASAP7_75t_L g2486 ( 
.A(n_2203),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2068),
.B(n_1110),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_2367),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2086),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2094),
.Y(n_2490)
);

INVx2_ASAP7_75t_L g2491 ( 
.A(n_2076),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2096),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2091),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2162),
.B(n_1455),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2098),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_SL g2496 ( 
.A(n_2318),
.B(n_1993),
.Y(n_2496)
);

INVx1_ASAP7_75t_L g2497 ( 
.A(n_2100),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2091),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_L g2499 ( 
.A(n_2080),
.B(n_1110),
.Y(n_2499)
);

INVx3_ASAP7_75t_L g2500 ( 
.A(n_2137),
.Y(n_2500)
);

OAI22xp5_ASAP7_75t_SL g2501 ( 
.A1(n_2037),
.A2(n_1788),
.B1(n_1790),
.B2(n_1787),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_2102),
.Y(n_2502)
);

INVx2_ASAP7_75t_L g2503 ( 
.A(n_2114),
.Y(n_2503)
);

INVxp67_ASAP7_75t_L g2504 ( 
.A(n_2057),
.Y(n_2504)
);

AND2x2_ASAP7_75t_L g2505 ( 
.A(n_2048),
.B(n_1457),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2079),
.B(n_1458),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2103),
.Y(n_2507)
);

INVx2_ASAP7_75t_L g2508 ( 
.A(n_2114),
.Y(n_2508)
);

INVx2_ASAP7_75t_L g2509 ( 
.A(n_2131),
.Y(n_2509)
);

NAND2xp33_ASAP7_75t_SL g2510 ( 
.A(n_2264),
.B(n_1124),
.Y(n_2510)
);

NAND2x1_ASAP7_75t_L g2511 ( 
.A(n_2029),
.B(n_1996),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2137),
.Y(n_2512)
);

INVx1_ASAP7_75t_SL g2513 ( 
.A(n_2124),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2108),
.Y(n_2514)
);

BUFx6f_ASAP7_75t_L g2515 ( 
.A(n_1993),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_2110),
.Y(n_2516)
);

INVx1_ASAP7_75t_SL g2517 ( 
.A(n_2156),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_2318),
.B(n_962),
.Y(n_2518)
);

INVx2_ASAP7_75t_L g2519 ( 
.A(n_2131),
.Y(n_2519)
);

CKINVDCx5p33_ASAP7_75t_R g2520 ( 
.A(n_1995),
.Y(n_2520)
);

AND2x2_ASAP7_75t_L g2521 ( 
.A(n_2122),
.B(n_1459),
.Y(n_2521)
);

BUFx2_ASAP7_75t_L g2522 ( 
.A(n_2075),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_2134),
.Y(n_2523)
);

BUFx6f_ASAP7_75t_L g2524 ( 
.A(n_2014),
.Y(n_2524)
);

INVx8_ASAP7_75t_L g2525 ( 
.A(n_2293),
.Y(n_2525)
);

INVx2_ASAP7_75t_L g2526 ( 
.A(n_2134),
.Y(n_2526)
);

INVx2_ASAP7_75t_L g2527 ( 
.A(n_2138),
.Y(n_2527)
);

INVx1_ASAP7_75t_L g2528 ( 
.A(n_2115),
.Y(n_2528)
);

BUFx2_ASAP7_75t_L g2529 ( 
.A(n_2075),
.Y(n_2529)
);

NAND2xp5_ASAP7_75t_SL g2530 ( 
.A(n_2318),
.B(n_962),
.Y(n_2530)
);

AND2x4_ASAP7_75t_L g2531 ( 
.A(n_2000),
.B(n_2056),
.Y(n_2531)
);

AND2x4_ASAP7_75t_L g2532 ( 
.A(n_2000),
.B(n_1462),
.Y(n_2532)
);

INVx2_ASAP7_75t_L g2533 ( 
.A(n_2138),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2118),
.Y(n_2534)
);

AND2x4_ASAP7_75t_L g2535 ( 
.A(n_2056),
.B(n_1463),
.Y(n_2535)
);

NAND2xp5_ASAP7_75t_L g2536 ( 
.A(n_2093),
.B(n_1124),
.Y(n_2536)
);

AOI22xp5_ASAP7_75t_L g2537 ( 
.A1(n_2290),
.A2(n_2029),
.B1(n_2211),
.B2(n_2146),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_2137),
.Y(n_2538)
);

HB1xp67_ASAP7_75t_L g2539 ( 
.A(n_2012),
.Y(n_2539)
);

NAND2xp5_ASAP7_75t_SL g2540 ( 
.A(n_2209),
.B(n_962),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2121),
.Y(n_2541)
);

NAND2xp5_ASAP7_75t_SL g2542 ( 
.A(n_2210),
.B(n_962),
.Y(n_2542)
);

INVx2_ASAP7_75t_L g2543 ( 
.A(n_2155),
.Y(n_2543)
);

BUFx3_ASAP7_75t_L g2544 ( 
.A(n_2306),
.Y(n_2544)
);

NAND2xp5_ASAP7_75t_L g2545 ( 
.A(n_2146),
.B(n_2105),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2151),
.B(n_1464),
.Y(n_2546)
);

INVx2_ASAP7_75t_L g2547 ( 
.A(n_2155),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2123),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2130),
.Y(n_2549)
);

INVxp67_ASAP7_75t_L g2550 ( 
.A(n_2057),
.Y(n_2550)
);

INVx2_ASAP7_75t_L g2551 ( 
.A(n_2169),
.Y(n_2551)
);

HB1xp67_ASAP7_75t_L g2552 ( 
.A(n_2119),
.Y(n_2552)
);

INVx3_ASAP7_75t_L g2553 ( 
.A(n_2137),
.Y(n_2553)
);

BUFx2_ASAP7_75t_L g2554 ( 
.A(n_2164),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2169),
.Y(n_2555)
);

OAI22xp5_ASAP7_75t_L g2556 ( 
.A1(n_2165),
.A2(n_812),
.B1(n_819),
.B2(n_811),
.Y(n_2556)
);

BUFx6f_ASAP7_75t_L g2557 ( 
.A(n_2014),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2132),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2142),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2210),
.B(n_962),
.Y(n_2560)
);

INVx1_ASAP7_75t_L g2561 ( 
.A(n_2143),
.Y(n_2561)
);

BUFx6f_ASAP7_75t_L g2562 ( 
.A(n_2014),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2149),
.Y(n_2563)
);

INVx3_ASAP7_75t_L g2564 ( 
.A(n_2168),
.Y(n_2564)
);

BUFx2_ASAP7_75t_L g2565 ( 
.A(n_2164),
.Y(n_2565)
);

AOI22xp5_ASAP7_75t_L g2566 ( 
.A1(n_2290),
.A2(n_1183),
.B1(n_1186),
.B2(n_1182),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2146),
.B(n_966),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_SL g2568 ( 
.A(n_2264),
.B(n_973),
.Y(n_2568)
);

INVx2_ASAP7_75t_L g2569 ( 
.A(n_2173),
.Y(n_2569)
);

INVx1_ASAP7_75t_L g2570 ( 
.A(n_2160),
.Y(n_2570)
);

BUFx6f_ASAP7_75t_L g2571 ( 
.A(n_2014),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2173),
.Y(n_2572)
);

INVx2_ASAP7_75t_L g2573 ( 
.A(n_2179),
.Y(n_2573)
);

INVx1_ASAP7_75t_L g2574 ( 
.A(n_2161),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2171),
.Y(n_2575)
);

INVx3_ASAP7_75t_L g2576 ( 
.A(n_2168),
.Y(n_2576)
);

BUFx3_ASAP7_75t_L g2577 ( 
.A(n_2306),
.Y(n_2577)
);

HB1xp67_ASAP7_75t_L g2578 ( 
.A(n_2119),
.Y(n_2578)
);

INVx2_ASAP7_75t_L g2579 ( 
.A(n_2179),
.Y(n_2579)
);

AND2x4_ASAP7_75t_L g2580 ( 
.A(n_2056),
.B(n_1465),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2172),
.Y(n_2581)
);

BUFx6f_ASAP7_75t_L g2582 ( 
.A(n_2027),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2184),
.Y(n_2583)
);

INVxp67_ASAP7_75t_L g2584 ( 
.A(n_2101),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_SL g2585 ( 
.A(n_2264),
.B(n_973),
.Y(n_2585)
);

BUFx6f_ASAP7_75t_L g2586 ( 
.A(n_2027),
.Y(n_2586)
);

OAI22xp33_ASAP7_75t_L g2587 ( 
.A1(n_2147),
.A2(n_1143),
.B1(n_1013),
.B2(n_1051),
.Y(n_2587)
);

INVx2_ASAP7_75t_L g2588 ( 
.A(n_2184),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2175),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2064),
.Y(n_2590)
);

HB1xp67_ASAP7_75t_L g2591 ( 
.A(n_2362),
.Y(n_2591)
);

NAND2xp33_ASAP7_75t_SL g2592 ( 
.A(n_2289),
.B(n_1041),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2190),
.Y(n_2593)
);

INVx1_ASAP7_75t_L g2594 ( 
.A(n_2064),
.Y(n_2594)
);

INVx3_ASAP7_75t_L g2595 ( 
.A(n_2168),
.Y(n_2595)
);

CKINVDCx8_ASAP7_75t_R g2596 ( 
.A(n_2152),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2168),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2067),
.Y(n_2598)
);

INVx1_ASAP7_75t_L g2599 ( 
.A(n_2067),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2073),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2073),
.Y(n_2601)
);

HB1xp67_ASAP7_75t_L g2602 ( 
.A(n_2373),
.Y(n_2602)
);

NAND2xp33_ASAP7_75t_SL g2603 ( 
.A(n_2289),
.B(n_1041),
.Y(n_2603)
);

INVx1_ASAP7_75t_L g2604 ( 
.A(n_2116),
.Y(n_2604)
);

INVx2_ASAP7_75t_L g2605 ( 
.A(n_2190),
.Y(n_2605)
);

HB1xp67_ASAP7_75t_L g2606 ( 
.A(n_2376),
.Y(n_2606)
);

AOI22xp5_ASAP7_75t_L g2607 ( 
.A1(n_2290),
.A2(n_830),
.B1(n_833),
.B2(n_827),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2116),
.Y(n_2608)
);

NOR2xp33_ASAP7_75t_SL g2609 ( 
.A(n_2003),
.B(n_2007),
.Y(n_2609)
);

INVx2_ASAP7_75t_L g2610 ( 
.A(n_2191),
.Y(n_2610)
);

AND2x4_ASAP7_75t_L g2611 ( 
.A(n_2312),
.B(n_1468),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2170),
.Y(n_2612)
);

NAND2xp5_ASAP7_75t_SL g2613 ( 
.A(n_2289),
.B(n_973),
.Y(n_2613)
);

INVx1_ASAP7_75t_L g2614 ( 
.A(n_2125),
.Y(n_2614)
);

INVx1_ASAP7_75t_L g2615 ( 
.A(n_2125),
.Y(n_2615)
);

BUFx6f_ASAP7_75t_SL g2616 ( 
.A(n_2312),
.Y(n_2616)
);

NAND2xp5_ASAP7_75t_SL g2617 ( 
.A(n_2289),
.B(n_2300),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2129),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2129),
.Y(n_2619)
);

INVx3_ASAP7_75t_L g2620 ( 
.A(n_2170),
.Y(n_2620)
);

INVxp67_ASAP7_75t_L g2621 ( 
.A(n_2101),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2191),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2166),
.Y(n_2623)
);

INVx1_ASAP7_75t_L g2624 ( 
.A(n_2166),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2174),
.Y(n_2625)
);

AOI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2290),
.A2(n_839),
.B1(n_841),
.B2(n_838),
.Y(n_2626)
);

AND2x2_ASAP7_75t_L g2627 ( 
.A(n_2285),
.B(n_1471),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2174),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2300),
.B(n_973),
.Y(n_2629)
);

INVx1_ASAP7_75t_L g2630 ( 
.A(n_1985),
.Y(n_2630)
);

NAND2xp5_ASAP7_75t_SL g2631 ( 
.A(n_2300),
.B(n_973),
.Y(n_2631)
);

BUFx6f_ASAP7_75t_L g2632 ( 
.A(n_2027),
.Y(n_2632)
);

NAND2xp5_ASAP7_75t_SL g2633 ( 
.A(n_2300),
.B(n_973),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_1989),
.Y(n_2634)
);

NAND2xp5_ASAP7_75t_L g2635 ( 
.A(n_2105),
.B(n_1051),
.Y(n_2635)
);

NAND2xp33_ASAP7_75t_SL g2636 ( 
.A(n_2325),
.B(n_1056),
.Y(n_2636)
);

NAND2xp5_ASAP7_75t_SL g2637 ( 
.A(n_2010),
.B(n_974),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_1990),
.Y(n_2638)
);

NAND2xp33_ASAP7_75t_SL g2639 ( 
.A(n_2325),
.B(n_1056),
.Y(n_2639)
);

NOR2xp33_ASAP7_75t_L g2640 ( 
.A(n_2176),
.B(n_842),
.Y(n_2640)
);

OAI22xp5_ASAP7_75t_SL g2641 ( 
.A1(n_2042),
.A2(n_1793),
.B1(n_1797),
.B2(n_1792),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2221),
.Y(n_2642)
);

NOR2xp33_ASAP7_75t_L g2643 ( 
.A(n_2192),
.B(n_843),
.Y(n_2643)
);

INVxp67_ASAP7_75t_L g2644 ( 
.A(n_2133),
.Y(n_2644)
);

AND2x2_ASAP7_75t_L g2645 ( 
.A(n_2199),
.B(n_1473),
.Y(n_2645)
);

BUFx6f_ASAP7_75t_L g2646 ( 
.A(n_2027),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2221),
.Y(n_2647)
);

HB1xp67_ASAP7_75t_L g2648 ( 
.A(n_2350),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_SL g2649 ( 
.A(n_2010),
.B(n_974),
.Y(n_2649)
);

INVx2_ASAP7_75t_L g2650 ( 
.A(n_2225),
.Y(n_2650)
);

HB1xp67_ASAP7_75t_L g2651 ( 
.A(n_2341),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2105),
.B(n_1101),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_1992),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_1998),
.Y(n_2654)
);

NOR2xp33_ASAP7_75t_L g2655 ( 
.A(n_2196),
.B(n_846),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2001),
.Y(n_2656)
);

AND2x4_ASAP7_75t_L g2657 ( 
.A(n_2136),
.B(n_1475),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_SL g2658 ( 
.A(n_2024),
.B(n_974),
.Y(n_2658)
);

INVx2_ASAP7_75t_L g2659 ( 
.A(n_2225),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2245),
.Y(n_2660)
);

AND2x2_ASAP7_75t_L g2661 ( 
.A(n_2199),
.B(n_2097),
.Y(n_2661)
);

INVx1_ASAP7_75t_L g2662 ( 
.A(n_2002),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2136),
.B(n_1101),
.Y(n_2663)
);

INVx1_ASAP7_75t_L g2664 ( 
.A(n_2205),
.Y(n_2664)
);

INVx2_ASAP7_75t_L g2665 ( 
.A(n_2245),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2205),
.Y(n_2666)
);

AND2x4_ASAP7_75t_L g2667 ( 
.A(n_2136),
.B(n_1476),
.Y(n_2667)
);

AND2x2_ASAP7_75t_L g2668 ( 
.A(n_2112),
.B(n_1479),
.Y(n_2668)
);

INVx3_ASAP7_75t_L g2669 ( 
.A(n_2170),
.Y(n_2669)
);

BUFx6f_ASAP7_75t_L g2670 ( 
.A(n_2051),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_SL g2671 ( 
.A1(n_2042),
.A2(n_1793),
.B1(n_1797),
.B2(n_1792),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2213),
.Y(n_2672)
);

HB1xp67_ASAP7_75t_L g2673 ( 
.A(n_2341),
.Y(n_2673)
);

AOI22xp5_ASAP7_75t_L g2674 ( 
.A1(n_2029),
.A2(n_849),
.B1(n_850),
.B2(n_847),
.Y(n_2674)
);

AND2x2_ASAP7_75t_L g2675 ( 
.A(n_1988),
.B(n_1482),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2213),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2224),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2170),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2246),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2246),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2224),
.Y(n_2681)
);

INVx2_ASAP7_75t_L g2682 ( 
.A(n_2251),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2234),
.Y(n_2683)
);

AOI22xp5_ASAP7_75t_L g2684 ( 
.A1(n_2029),
.A2(n_855),
.B1(n_857),
.B2(n_853),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2234),
.Y(n_2685)
);

INVx1_ASAP7_75t_L g2686 ( 
.A(n_2214),
.Y(n_2686)
);

AND2x6_ASAP7_75t_L g2687 ( 
.A(n_2011),
.B(n_1128),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2182),
.Y(n_2688)
);

INVx1_ASAP7_75t_L g2689 ( 
.A(n_2182),
.Y(n_2689)
);

INVx1_ASAP7_75t_L g2690 ( 
.A(n_2235),
.Y(n_2690)
);

INVx3_ASAP7_75t_L g2691 ( 
.A(n_2236),
.Y(n_2691)
);

NOR2xp33_ASAP7_75t_L g2692 ( 
.A(n_2058),
.B(n_859),
.Y(n_2692)
);

AND2x6_ASAP7_75t_L g2693 ( 
.A(n_2258),
.B(n_1128),
.Y(n_2693)
);

NAND2xp5_ASAP7_75t_L g2694 ( 
.A(n_2144),
.B(n_1143),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2235),
.Y(n_2695)
);

INVx1_ASAP7_75t_SL g2696 ( 
.A(n_2359),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2228),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2228),
.Y(n_2698)
);

INVx1_ASAP7_75t_L g2699 ( 
.A(n_2228),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2231),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2341),
.Y(n_2701)
);

INVx2_ASAP7_75t_L g2702 ( 
.A(n_2251),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2231),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2231),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2144),
.B(n_1150),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2248),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2248),
.Y(n_2707)
);

INVx1_ASAP7_75t_SL g2708 ( 
.A(n_2369),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2254),
.Y(n_2709)
);

BUFx6f_ASAP7_75t_L g2710 ( 
.A(n_2051),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2248),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2157),
.Y(n_2712)
);

NAND2xp5_ASAP7_75t_L g2713 ( 
.A(n_2144),
.B(n_1150),
.Y(n_2713)
);

INVx1_ASAP7_75t_L g2714 ( 
.A(n_2157),
.Y(n_2714)
);

HB1xp67_ASAP7_75t_L g2715 ( 
.A(n_2348),
.Y(n_2715)
);

INVx2_ASAP7_75t_L g2716 ( 
.A(n_2254),
.Y(n_2716)
);

BUFx6f_ASAP7_75t_L g2717 ( 
.A(n_2051),
.Y(n_2717)
);

AND2x2_ASAP7_75t_L g2718 ( 
.A(n_2148),
.B(n_1484),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2211),
.B(n_1152),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_SL g2720 ( 
.A(n_2024),
.B(n_974),
.Y(n_2720)
);

INVx1_ASAP7_75t_L g2721 ( 
.A(n_2157),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2255),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2348),
.Y(n_2723)
);

AOI22xp5_ASAP7_75t_L g2724 ( 
.A1(n_2029),
.A2(n_865),
.B1(n_869),
.B2(n_863),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2158),
.Y(n_2725)
);

INVx2_ASAP7_75t_L g2726 ( 
.A(n_2286),
.Y(n_2726)
);

HB1xp67_ASAP7_75t_L g2727 ( 
.A(n_2348),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2211),
.B(n_1152),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2236),
.Y(n_2729)
);

INVx1_ASAP7_75t_L g2730 ( 
.A(n_2158),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2158),
.Y(n_2731)
);

INVx2_ASAP7_75t_L g2732 ( 
.A(n_2236),
.Y(n_2732)
);

HB1xp67_ASAP7_75t_L g2733 ( 
.A(n_2263),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2236),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2090),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2293),
.B(n_1488),
.Y(n_2736)
);

NAND2x1_ASAP7_75t_L g2737 ( 
.A(n_1996),
.B(n_1628),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2090),
.Y(n_2738)
);

INVx1_ASAP7_75t_L g2739 ( 
.A(n_2090),
.Y(n_2739)
);

INVx6_ASAP7_75t_L g2740 ( 
.A(n_2043),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2244),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_SL g2742 ( 
.A(n_2016),
.B(n_974),
.Y(n_2742)
);

INVx1_ASAP7_75t_L g2743 ( 
.A(n_2230),
.Y(n_2743)
);

INVx2_ASAP7_75t_L g2744 ( 
.A(n_2244),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2127),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2120),
.Y(n_2746)
);

AND2x2_ASAP7_75t_L g2747 ( 
.A(n_2148),
.B(n_1489),
.Y(n_2747)
);

INVx3_ASAP7_75t_L g2748 ( 
.A(n_2244),
.Y(n_2748)
);

NAND2xp5_ASAP7_75t_SL g2749 ( 
.A(n_2016),
.B(n_2041),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_SL g2750 ( 
.A(n_2041),
.B(n_974),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2211),
.B(n_1174),
.Y(n_2751)
);

INVx1_ASAP7_75t_L g2752 ( 
.A(n_2194),
.Y(n_2752)
);

INVx1_ASAP7_75t_L g2753 ( 
.A(n_2194),
.Y(n_2753)
);

AND2x2_ASAP7_75t_L g2754 ( 
.A(n_2263),
.B(n_1490),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2194),
.Y(n_2755)
);

AND2x2_ASAP7_75t_L g2756 ( 
.A(n_2263),
.B(n_1493),
.Y(n_2756)
);

BUFx6f_ASAP7_75t_L g2757 ( 
.A(n_2051),
.Y(n_2757)
);

BUFx2_ASAP7_75t_L g2758 ( 
.A(n_2140),
.Y(n_2758)
);

INVx2_ASAP7_75t_L g2759 ( 
.A(n_2244),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2022),
.Y(n_2760)
);

INVx2_ASAP7_75t_L g2761 ( 
.A(n_2150),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2023),
.Y(n_2762)
);

INVx2_ASAP7_75t_L g2763 ( 
.A(n_2195),
.Y(n_2763)
);

AND2x6_ASAP7_75t_L g2764 ( 
.A(n_2258),
.B(n_1174),
.Y(n_2764)
);

CKINVDCx5p33_ASAP7_75t_R g2765 ( 
.A(n_2017),
.Y(n_2765)
);

NAND2xp5_ASAP7_75t_SL g2766 ( 
.A(n_2257),
.B(n_2260),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2346),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2153),
.Y(n_2768)
);

HB1xp67_ASAP7_75t_L g2769 ( 
.A(n_2374),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2154),
.Y(n_2770)
);

INVx2_ASAP7_75t_L g2771 ( 
.A(n_2189),
.Y(n_2771)
);

BUFx6f_ASAP7_75t_L g2772 ( 
.A(n_2060),
.Y(n_2772)
);

INVx1_ASAP7_75t_SL g2773 ( 
.A(n_2140),
.Y(n_2773)
);

INVx1_ASAP7_75t_L g2774 ( 
.A(n_2360),
.Y(n_2774)
);

INVx1_ASAP7_75t_L g2775 ( 
.A(n_2372),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2060),
.Y(n_2776)
);

BUFx4f_ASAP7_75t_L g2777 ( 
.A(n_2740),
.Y(n_2777)
);

INVx3_ASAP7_75t_L g2778 ( 
.A(n_2525),
.Y(n_2778)
);

BUFx6f_ASAP7_75t_L g2779 ( 
.A(n_2379),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2686),
.B(n_2211),
.Y(n_2780)
);

HB1xp67_ASAP7_75t_L g2781 ( 
.A(n_2733),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_L g2782 ( 
.A(n_2743),
.B(n_2232),
.Y(n_2782)
);

AND2x4_ASAP7_75t_L g2783 ( 
.A(n_2531),
.B(n_2293),
.Y(n_2783)
);

NAND2xp5_ASAP7_75t_SL g2784 ( 
.A(n_2531),
.B(n_2269),
.Y(n_2784)
);

OR2x2_ASAP7_75t_L g2785 ( 
.A(n_2773),
.B(n_2180),
.Y(n_2785)
);

BUFx3_ASAP7_75t_L g2786 ( 
.A(n_2404),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_SL g2787 ( 
.A(n_2531),
.B(n_2269),
.Y(n_2787)
);

OR2x2_ASAP7_75t_L g2788 ( 
.A(n_2554),
.B(n_2358),
.Y(n_2788)
);

CKINVDCx5p33_ASAP7_75t_R g2789 ( 
.A(n_2520),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2544),
.Y(n_2790)
);

AND2x6_ASAP7_75t_L g2791 ( 
.A(n_2537),
.B(n_2335),
.Y(n_2791)
);

INVx2_ASAP7_75t_L g2792 ( 
.A(n_2380),
.Y(n_2792)
);

BUFx6f_ASAP7_75t_L g2793 ( 
.A(n_2379),
.Y(n_2793)
);

BUFx3_ASAP7_75t_L g2794 ( 
.A(n_2404),
.Y(n_2794)
);

INVx2_ASAP7_75t_L g2795 ( 
.A(n_2380),
.Y(n_2795)
);

INVx3_ASAP7_75t_L g2796 ( 
.A(n_2525),
.Y(n_2796)
);

NAND2xp5_ASAP7_75t_L g2797 ( 
.A(n_2768),
.B(n_2232),
.Y(n_2797)
);

INVx2_ASAP7_75t_L g2798 ( 
.A(n_2384),
.Y(n_2798)
);

BUFx3_ASAP7_75t_L g2799 ( 
.A(n_2404),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2545),
.Y(n_2800)
);

BUFx3_ASAP7_75t_L g2801 ( 
.A(n_2520),
.Y(n_2801)
);

NAND2xp5_ASAP7_75t_L g2802 ( 
.A(n_2770),
.B(n_2273),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2384),
.Y(n_2803)
);

AND2x6_ASAP7_75t_L g2804 ( 
.A(n_2736),
.B(n_2281),
.Y(n_2804)
);

INVx4_ASAP7_75t_L g2805 ( 
.A(n_2525),
.Y(n_2805)
);

INVx2_ASAP7_75t_SL g2806 ( 
.A(n_2544),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2378),
.Y(n_2807)
);

INVx1_ASAP7_75t_L g2808 ( 
.A(n_2383),
.Y(n_2808)
);

BUFx6f_ASAP7_75t_L g2809 ( 
.A(n_2379),
.Y(n_2809)
);

INVx2_ASAP7_75t_L g2810 ( 
.A(n_2395),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2386),
.Y(n_2811)
);

NAND2xp5_ASAP7_75t_L g2812 ( 
.A(n_2774),
.B(n_2201),
.Y(n_2812)
);

INVx2_ASAP7_75t_L g2813 ( 
.A(n_2395),
.Y(n_2813)
);

INVx4_ASAP7_75t_L g2814 ( 
.A(n_2765),
.Y(n_2814)
);

NAND2xp5_ASAP7_75t_L g2815 ( 
.A(n_2775),
.B(n_2375),
.Y(n_2815)
);

INVx5_ASAP7_75t_L g2816 ( 
.A(n_2466),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2387),
.Y(n_2817)
);

NOR2xp33_ASAP7_75t_L g2818 ( 
.A(n_2644),
.B(n_2377),
.Y(n_2818)
);

AND2x2_ASAP7_75t_L g2819 ( 
.A(n_2627),
.B(n_1983),
.Y(n_2819)
);

NOR2xp33_ASAP7_75t_L g2820 ( 
.A(n_2733),
.B(n_2343),
.Y(n_2820)
);

AND2x2_ASAP7_75t_L g2821 ( 
.A(n_2591),
.B(n_2028),
.Y(n_2821)
);

INVx2_ASAP7_75t_L g2822 ( 
.A(n_2398),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_SL g2823 ( 
.A(n_2481),
.B(n_2281),
.Y(n_2823)
);

NAND2xp5_ASAP7_75t_L g2824 ( 
.A(n_2745),
.B(n_2356),
.Y(n_2824)
);

INVx1_ASAP7_75t_L g2825 ( 
.A(n_2388),
.Y(n_2825)
);

INVx3_ASAP7_75t_L g2826 ( 
.A(n_2379),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2389),
.Y(n_2827)
);

NAND2xp5_ASAP7_75t_SL g2828 ( 
.A(n_2609),
.B(n_2295),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_SL g2829 ( 
.A(n_2577),
.B(n_2295),
.Y(n_2829)
);

OR2x6_ASAP7_75t_L g2830 ( 
.A(n_2577),
.B(n_2111),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2746),
.B(n_2257),
.Y(n_2831)
);

NOR2xp33_ASAP7_75t_L g2832 ( 
.A(n_2640),
.B(n_2058),
.Y(n_2832)
);

AO22x2_ASAP7_75t_L g2833 ( 
.A1(n_2771),
.A2(n_2363),
.B1(n_2368),
.B2(n_2358),
.Y(n_2833)
);

BUFx6f_ASAP7_75t_L g2834 ( 
.A(n_2382),
.Y(n_2834)
);

NAND3x1_ASAP7_75t_L g2835 ( 
.A(n_2661),
.B(n_2344),
.C(n_2339),
.Y(n_2835)
);

BUFx6f_ASAP7_75t_L g2836 ( 
.A(n_2382),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2760),
.B(n_2257),
.Y(n_2837)
);

INVx2_ASAP7_75t_L g2838 ( 
.A(n_2398),
.Y(n_2838)
);

INVxp67_ASAP7_75t_L g2839 ( 
.A(n_2522),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2391),
.Y(n_2840)
);

AND2x6_ASAP7_75t_L g2841 ( 
.A(n_2736),
.B(n_2298),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2591),
.B(n_2087),
.Y(n_2842)
);

INVx1_ASAP7_75t_L g2843 ( 
.A(n_2393),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2640),
.B(n_2078),
.Y(n_2844)
);

INVx2_ASAP7_75t_L g2845 ( 
.A(n_2402),
.Y(n_2845)
);

NAND2xp5_ASAP7_75t_SL g2846 ( 
.A(n_2513),
.B(n_2298),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2394),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2397),
.Y(n_2848)
);

INVx2_ASAP7_75t_L g2849 ( 
.A(n_2402),
.Y(n_2849)
);

AND2x2_ASAP7_75t_L g2850 ( 
.A(n_2602),
.B(n_2089),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2400),
.Y(n_2851)
);

AND2x6_ASAP7_75t_L g2852 ( 
.A(n_2736),
.B(n_2302),
.Y(n_2852)
);

BUFx3_ASAP7_75t_L g2853 ( 
.A(n_2765),
.Y(n_2853)
);

NAND2xp5_ASAP7_75t_L g2854 ( 
.A(n_2762),
.B(n_2257),
.Y(n_2854)
);

CKINVDCx5p33_ASAP7_75t_R g2855 ( 
.A(n_2616),
.Y(n_2855)
);

BUFx6f_ASAP7_75t_L g2856 ( 
.A(n_2382),
.Y(n_2856)
);

AOI22xp33_ASAP7_75t_L g2857 ( 
.A1(n_2697),
.A2(n_2328),
.B1(n_2351),
.B2(n_2324),
.Y(n_2857)
);

HB1xp67_ASAP7_75t_L g2858 ( 
.A(n_2529),
.Y(n_2858)
);

INVx2_ASAP7_75t_L g2859 ( 
.A(n_2403),
.Y(n_2859)
);

OR2x2_ASAP7_75t_L g2860 ( 
.A(n_2565),
.B(n_2363),
.Y(n_2860)
);

INVx1_ASAP7_75t_SL g2861 ( 
.A(n_2696),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2401),
.Y(n_2862)
);

AOI22xp5_ASAP7_75t_L g2863 ( 
.A1(n_2643),
.A2(n_2099),
.B1(n_2106),
.B2(n_2223),
.Y(n_2863)
);

A2O1A1Ixp33_ASAP7_75t_L g2864 ( 
.A1(n_2643),
.A2(n_2283),
.B(n_2303),
.C(n_2279),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2408),
.Y(n_2865)
);

INVx2_ASAP7_75t_L g2866 ( 
.A(n_2403),
.Y(n_2866)
);

OR2x2_ASAP7_75t_L g2867 ( 
.A(n_2602),
.B(n_2368),
.Y(n_2867)
);

INVx1_ASAP7_75t_L g2868 ( 
.A(n_2411),
.Y(n_2868)
);

AND2x6_ASAP7_75t_L g2869 ( 
.A(n_2698),
.B(n_2302),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2606),
.B(n_2145),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2412),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2382),
.Y(n_2872)
);

NAND2xp33_ASAP7_75t_SL g2873 ( 
.A(n_2616),
.B(n_2040),
.Y(n_2873)
);

INVx2_ASAP7_75t_L g2874 ( 
.A(n_2409),
.Y(n_2874)
);

NAND2xp5_ASAP7_75t_L g2875 ( 
.A(n_2630),
.B(n_2260),
.Y(n_2875)
);

AND2x4_ASAP7_75t_L g2876 ( 
.A(n_2657),
.B(n_2667),
.Y(n_2876)
);

INVx2_ASAP7_75t_L g2877 ( 
.A(n_2409),
.Y(n_2877)
);

INVx2_ASAP7_75t_SL g2878 ( 
.A(n_2446),
.Y(n_2878)
);

NAND2xp5_ASAP7_75t_L g2879 ( 
.A(n_2634),
.B(n_2260),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2638),
.B(n_2260),
.Y(n_2880)
);

OR2x2_ASAP7_75t_L g2881 ( 
.A(n_2606),
.B(n_2336),
.Y(n_2881)
);

INVxp33_ASAP7_75t_L g2882 ( 
.A(n_2415),
.Y(n_2882)
);

INVx2_ASAP7_75t_L g2883 ( 
.A(n_2418),
.Y(n_2883)
);

OR2x2_ASAP7_75t_L g2884 ( 
.A(n_2648),
.B(n_2336),
.Y(n_2884)
);

AOI22xp33_ASAP7_75t_L g2885 ( 
.A1(n_2699),
.A2(n_2135),
.B1(n_1994),
.B2(n_2084),
.Y(n_2885)
);

INVx1_ASAP7_75t_SL g2886 ( 
.A(n_2708),
.Y(n_2886)
);

INVx4_ASAP7_75t_L g2887 ( 
.A(n_2740),
.Y(n_2887)
);

INVx2_ASAP7_75t_L g2888 ( 
.A(n_2418),
.Y(n_2888)
);

BUFx3_ASAP7_75t_L g2889 ( 
.A(n_2399),
.Y(n_2889)
);

INVxp67_ASAP7_75t_SL g2890 ( 
.A(n_2466),
.Y(n_2890)
);

INVx1_ASAP7_75t_L g2891 ( 
.A(n_2413),
.Y(n_2891)
);

INVx5_ASAP7_75t_L g2892 ( 
.A(n_2466),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2416),
.Y(n_2893)
);

INVx1_ASAP7_75t_L g2894 ( 
.A(n_2420),
.Y(n_2894)
);

AND2x2_ASAP7_75t_L g2895 ( 
.A(n_2648),
.B(n_2206),
.Y(n_2895)
);

OR2x2_ASAP7_75t_L g2896 ( 
.A(n_2552),
.B(n_2338),
.Y(n_2896)
);

AND2x4_ASAP7_75t_L g2897 ( 
.A(n_2657),
.B(n_2293),
.Y(n_2897)
);

INVx3_ASAP7_75t_L g2898 ( 
.A(n_2385),
.Y(n_2898)
);

AND2x2_ASAP7_75t_L g2899 ( 
.A(n_2754),
.B(n_2208),
.Y(n_2899)
);

BUFx6f_ASAP7_75t_L g2900 ( 
.A(n_2385),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2425),
.Y(n_2901)
);

HB1xp67_ASAP7_75t_L g2902 ( 
.A(n_2552),
.Y(n_2902)
);

NAND2xp5_ASAP7_75t_L g2903 ( 
.A(n_2653),
.B(n_2274),
.Y(n_2903)
);

CKINVDCx5p33_ASAP7_75t_R g2904 ( 
.A(n_2399),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2422),
.Y(n_2905)
);

INVx1_ASAP7_75t_L g2906 ( 
.A(n_2426),
.Y(n_2906)
);

NOR2xp33_ASAP7_75t_L g2907 ( 
.A(n_2655),
.B(n_2078),
.Y(n_2907)
);

NAND2xp5_ASAP7_75t_L g2908 ( 
.A(n_2654),
.B(n_2274),
.Y(n_2908)
);

INVx2_ASAP7_75t_L g2909 ( 
.A(n_2425),
.Y(n_2909)
);

BUFx2_ASAP7_75t_L g2910 ( 
.A(n_2758),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_L g2911 ( 
.A(n_2655),
.B(n_2259),
.Y(n_2911)
);

CKINVDCx5p33_ASAP7_75t_R g2912 ( 
.A(n_2405),
.Y(n_2912)
);

INVx3_ASAP7_75t_L g2913 ( 
.A(n_2385),
.Y(n_2913)
);

INVx2_ASAP7_75t_SL g2914 ( 
.A(n_2453),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_SL g2915 ( 
.A(n_2517),
.B(n_2279),
.Y(n_2915)
);

AND2x4_ASAP7_75t_L g2916 ( 
.A(n_2657),
.B(n_2293),
.Y(n_2916)
);

AOI22xp33_ASAP7_75t_L g2917 ( 
.A1(n_2700),
.A2(n_1994),
.B1(n_2084),
.B2(n_2299),
.Y(n_2917)
);

NOR2xp33_ASAP7_75t_SL g2918 ( 
.A(n_2587),
.B(n_2040),
.Y(n_2918)
);

INVx1_ASAP7_75t_L g2919 ( 
.A(n_2428),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2430),
.Y(n_2920)
);

INVxp67_ASAP7_75t_L g2921 ( 
.A(n_2578),
.Y(n_2921)
);

BUFx6f_ASAP7_75t_L g2922 ( 
.A(n_2385),
.Y(n_2922)
);

INVx1_ASAP7_75t_L g2923 ( 
.A(n_2431),
.Y(n_2923)
);

NAND2xp5_ASAP7_75t_L g2924 ( 
.A(n_2656),
.B(n_2274),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2432),
.Y(n_2925)
);

AND2x4_ASAP7_75t_L g2926 ( 
.A(n_2667),
.B(n_2043),
.Y(n_2926)
);

INVx1_ASAP7_75t_L g2927 ( 
.A(n_2434),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_SL g2928 ( 
.A(n_2611),
.B(n_2283),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2435),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2438),
.Y(n_2930)
);

NOR2xp33_ASAP7_75t_SL g2931 ( 
.A(n_2587),
.B(n_2061),
.Y(n_2931)
);

NAND2xp5_ASAP7_75t_SL g2932 ( 
.A(n_2611),
.B(n_2303),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2429),
.Y(n_2933)
);

AOI22xp5_ASAP7_75t_L g2934 ( 
.A1(n_2692),
.A2(n_2227),
.B1(n_2252),
.B2(n_2243),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2410),
.Y(n_2935)
);

INVx2_ASAP7_75t_L g2936 ( 
.A(n_2429),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_SL g2937 ( 
.A(n_2611),
.B(n_2308),
.Y(n_2937)
);

INVx2_ASAP7_75t_L g2938 ( 
.A(n_2433),
.Y(n_2938)
);

BUFx6f_ASAP7_75t_L g2939 ( 
.A(n_2410),
.Y(n_2939)
);

AO22x2_ASAP7_75t_L g2940 ( 
.A1(n_2771),
.A2(n_2338),
.B1(n_2347),
.B2(n_2345),
.Y(n_2940)
);

OR2x2_ASAP7_75t_L g2941 ( 
.A(n_2578),
.B(n_2345),
.Y(n_2941)
);

OR2x2_ASAP7_75t_L g2942 ( 
.A(n_2584),
.B(n_2347),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2488),
.Y(n_2943)
);

INVx1_ASAP7_75t_L g2944 ( 
.A(n_2440),
.Y(n_2944)
);

NAND2xp5_ASAP7_75t_L g2945 ( 
.A(n_2662),
.B(n_2468),
.Y(n_2945)
);

NOR2xp33_ASAP7_75t_L g2946 ( 
.A(n_2470),
.B(n_2308),
.Y(n_2946)
);

CKINVDCx16_ASAP7_75t_R g2947 ( 
.A(n_2501),
.Y(n_2947)
);

INVx1_ASAP7_75t_L g2948 ( 
.A(n_2442),
.Y(n_2948)
);

INVxp67_ASAP7_75t_L g2949 ( 
.A(n_2470),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2539),
.B(n_2496),
.Y(n_2950)
);

NAND2xp5_ASAP7_75t_L g2951 ( 
.A(n_2468),
.B(n_2274),
.Y(n_2951)
);

AND2x6_ASAP7_75t_L g2952 ( 
.A(n_2703),
.B(n_2315),
.Y(n_2952)
);

AOI22xp33_ASAP7_75t_L g2953 ( 
.A1(n_2704),
.A2(n_2299),
.B1(n_2274),
.B2(n_2354),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2756),
.B(n_2421),
.Y(n_2954)
);

INVx1_ASAP7_75t_L g2955 ( 
.A(n_2443),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2539),
.B(n_2315),
.Y(n_2956)
);

INVx2_ASAP7_75t_L g2957 ( 
.A(n_2433),
.Y(n_2957)
);

NAND2x1p5_ASAP7_75t_L g2958 ( 
.A(n_2511),
.B(n_2240),
.Y(n_2958)
);

INVx1_ASAP7_75t_L g2959 ( 
.A(n_2444),
.Y(n_2959)
);

BUFx3_ASAP7_75t_L g2960 ( 
.A(n_2405),
.Y(n_2960)
);

NAND2xp5_ASAP7_75t_SL g2961 ( 
.A(n_2469),
.B(n_2330),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2447),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2419),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2468),
.B(n_1984),
.Y(n_2964)
);

INVx1_ASAP7_75t_L g2965 ( 
.A(n_2450),
.Y(n_2965)
);

INVx1_ASAP7_75t_L g2966 ( 
.A(n_2452),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2439),
.Y(n_2967)
);

INVx3_ASAP7_75t_L g2968 ( 
.A(n_2410),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2439),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2455),
.Y(n_2970)
);

AND2x4_ASAP7_75t_L g2971 ( 
.A(n_2667),
.B(n_2297),
.Y(n_2971)
);

NAND3xp33_ASAP7_75t_L g2972 ( 
.A(n_2719),
.B(n_1999),
.C(n_2330),
.Y(n_2972)
);

BUFx2_ASAP7_75t_L g2973 ( 
.A(n_2445),
.Y(n_2973)
);

BUFx2_ASAP7_75t_L g2974 ( 
.A(n_2486),
.Y(n_2974)
);

INVx1_ASAP7_75t_L g2975 ( 
.A(n_2462),
.Y(n_2975)
);

NAND2xp5_ASAP7_75t_SL g2976 ( 
.A(n_2621),
.B(n_2277),
.Y(n_2976)
);

AND2x6_ASAP7_75t_L g2977 ( 
.A(n_2706),
.B(n_2327),
.Y(n_2977)
);

INVx4_ASAP7_75t_L g2978 ( 
.A(n_2740),
.Y(n_2978)
);

OR2x2_ASAP7_75t_L g2979 ( 
.A(n_2504),
.B(n_2334),
.Y(n_2979)
);

AND2x2_ASAP7_75t_L g2980 ( 
.A(n_2437),
.B(n_2250),
.Y(n_2980)
);

INVx4_ASAP7_75t_SL g2981 ( 
.A(n_2687),
.Y(n_2981)
);

NAND2xp5_ASAP7_75t_SL g2982 ( 
.A(n_2550),
.B(n_2282),
.Y(n_2982)
);

INVx1_ASAP7_75t_L g2983 ( 
.A(n_2463),
.Y(n_2983)
);

AND2x6_ASAP7_75t_L g2984 ( 
.A(n_2707),
.B(n_2262),
.Y(n_2984)
);

OA22x2_ASAP7_75t_L g2985 ( 
.A1(n_2651),
.A2(n_2316),
.B1(n_2364),
.B2(n_2361),
.Y(n_2985)
);

INVx2_ASAP7_75t_L g2986 ( 
.A(n_2448),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2645),
.B(n_2319),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2464),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_SL g2989 ( 
.A(n_2636),
.B(n_2288),
.Y(n_2989)
);

NAND2xp5_ASAP7_75t_L g2990 ( 
.A(n_2532),
.B(n_2207),
.Y(n_2990)
);

NOR2xp33_ASAP7_75t_L g2991 ( 
.A(n_2496),
.B(n_2301),
.Y(n_2991)
);

CKINVDCx5p33_ASAP7_75t_R g2992 ( 
.A(n_2596),
.Y(n_2992)
);

NAND2xp5_ASAP7_75t_SL g2993 ( 
.A(n_2636),
.B(n_2294),
.Y(n_2993)
);

INVx1_ASAP7_75t_L g2994 ( 
.A(n_2477),
.Y(n_2994)
);

INVxp67_ASAP7_75t_L g2995 ( 
.A(n_2668),
.Y(n_2995)
);

BUFx6f_ASAP7_75t_L g2996 ( 
.A(n_2410),
.Y(n_2996)
);

INVx1_ASAP7_75t_L g2997 ( 
.A(n_2482),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2484),
.Y(n_2998)
);

NAND2xp5_ASAP7_75t_SL g2999 ( 
.A(n_2639),
.B(n_2296),
.Y(n_2999)
);

BUFx3_ASAP7_75t_L g3000 ( 
.A(n_2596),
.Y(n_3000)
);

BUFx6f_ASAP7_75t_L g3001 ( 
.A(n_2424),
.Y(n_3001)
);

INVx2_ASAP7_75t_L g3002 ( 
.A(n_2448),
.Y(n_3002)
);

INVx3_ASAP7_75t_L g3003 ( 
.A(n_2424),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2485),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2489),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2424),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2490),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2449),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2532),
.B(n_1999),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2492),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2495),
.Y(n_3011)
);

AO22x2_ASAP7_75t_L g3012 ( 
.A1(n_2752),
.A2(n_2370),
.B1(n_2371),
.B2(n_2366),
.Y(n_3012)
);

INVx2_ASAP7_75t_L g3013 ( 
.A(n_2449),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_L g3014 ( 
.A(n_2532),
.B(n_2256),
.Y(n_3014)
);

NOR2xp33_ASAP7_75t_SL g3015 ( 
.A(n_2451),
.B(n_2061),
.Y(n_3015)
);

INVx2_ASAP7_75t_L g3016 ( 
.A(n_2454),
.Y(n_3016)
);

INVx2_ASAP7_75t_L g3017 ( 
.A(n_2454),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2535),
.B(n_2332),
.Y(n_3018)
);

INVx2_ASAP7_75t_L g3019 ( 
.A(n_2461),
.Y(n_3019)
);

AOI22xp5_ASAP7_75t_L g3020 ( 
.A1(n_2692),
.A2(n_2133),
.B1(n_2301),
.B2(n_2287),
.Y(n_3020)
);

INVx2_ASAP7_75t_SL g3021 ( 
.A(n_2718),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2769),
.Y(n_3022)
);

AOI22xp33_ASAP7_75t_L g3023 ( 
.A1(n_2711),
.A2(n_2033),
.B1(n_2200),
.B2(n_2198),
.Y(n_3023)
);

OR2x6_ASAP7_75t_L g3024 ( 
.A(n_2641),
.B(n_2111),
.Y(n_3024)
);

NAND2xp5_ASAP7_75t_L g3025 ( 
.A(n_2535),
.B(n_2159),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2497),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2461),
.Y(n_3027)
);

INVx6_ASAP7_75t_L g3028 ( 
.A(n_2535),
.Y(n_3028)
);

NAND2xp5_ASAP7_75t_SL g3029 ( 
.A(n_2639),
.B(n_2278),
.Y(n_3029)
);

BUFx2_ASAP7_75t_L g3030 ( 
.A(n_2671),
.Y(n_3030)
);

AND2x4_ASAP7_75t_L g3031 ( 
.A(n_2580),
.B(n_2322),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_SL g3032 ( 
.A(n_2674),
.B(n_2292),
.Y(n_3032)
);

AND2x6_ASAP7_75t_L g3033 ( 
.A(n_2479),
.B(n_2304),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2651),
.B(n_2357),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2673),
.B(n_2349),
.Y(n_3035)
);

INVx1_ASAP7_75t_L g3036 ( 
.A(n_2502),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2580),
.B(n_2305),
.Y(n_3037)
);

INVx2_ASAP7_75t_L g3038 ( 
.A(n_2467),
.Y(n_3038)
);

INVx4_ASAP7_75t_L g3039 ( 
.A(n_2424),
.Y(n_3039)
);

INVx1_ASAP7_75t_L g3040 ( 
.A(n_2507),
.Y(n_3040)
);

NOR2xp33_ASAP7_75t_R g3041 ( 
.A(n_2480),
.B(n_2128),
.Y(n_3041)
);

INVx3_ASAP7_75t_L g3042 ( 
.A(n_2465),
.Y(n_3042)
);

BUFx3_ASAP7_75t_L g3043 ( 
.A(n_2769),
.Y(n_3043)
);

BUFx4f_ASAP7_75t_L g3044 ( 
.A(n_2414),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2514),
.Y(n_3045)
);

AND2x4_ASAP7_75t_L g3046 ( 
.A(n_2580),
.B(n_2117),
.Y(n_3046)
);

INVx2_ASAP7_75t_L g3047 ( 
.A(n_2467),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2516),
.Y(n_3048)
);

BUFx2_ASAP7_75t_L g3049 ( 
.A(n_2673),
.Y(n_3049)
);

BUFx6f_ASAP7_75t_L g3050 ( 
.A(n_2465),
.Y(n_3050)
);

NAND2xp5_ASAP7_75t_L g3051 ( 
.A(n_2407),
.B(n_2307),
.Y(n_3051)
);

INVx1_ASAP7_75t_L g3052 ( 
.A(n_2528),
.Y(n_3052)
);

NAND2xp5_ASAP7_75t_SL g3053 ( 
.A(n_2684),
.B(n_2309),
.Y(n_3053)
);

BUFx3_ASAP7_75t_L g3054 ( 
.A(n_2747),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2472),
.Y(n_3055)
);

INVx1_ASAP7_75t_SL g3056 ( 
.A(n_2505),
.Y(n_3056)
);

INVx2_ASAP7_75t_L g3057 ( 
.A(n_2472),
.Y(n_3057)
);

INVx5_ASAP7_75t_L g3058 ( 
.A(n_2466),
.Y(n_3058)
);

CKINVDCx5p33_ASAP7_75t_R g3059 ( 
.A(n_2701),
.Y(n_3059)
);

BUFx3_ASAP7_75t_L g3060 ( 
.A(n_2506),
.Y(n_3060)
);

INVxp67_ASAP7_75t_L g3061 ( 
.A(n_2494),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2724),
.B(n_2310),
.Y(n_3062)
);

INVx4_ASAP7_75t_L g3063 ( 
.A(n_2465),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2521),
.B(n_2215),
.Y(n_3064)
);

NAND2xp5_ASAP7_75t_SL g3065 ( 
.A(n_2436),
.B(n_2317),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2534),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2590),
.B(n_2321),
.Y(n_3067)
);

BUFx2_ASAP7_75t_L g3068 ( 
.A(n_2701),
.Y(n_3068)
);

INVx1_ASAP7_75t_SL g3069 ( 
.A(n_2546),
.Y(n_3069)
);

OR2x2_ASAP7_75t_L g3070 ( 
.A(n_2715),
.B(n_2349),
.Y(n_3070)
);

INVx1_ASAP7_75t_L g3071 ( 
.A(n_2541),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_2465),
.Y(n_3072)
);

NAND2xp5_ASAP7_75t_L g3073 ( 
.A(n_2594),
.B(n_2326),
.Y(n_3073)
);

OR2x6_ASAP7_75t_L g3074 ( 
.A(n_2715),
.B(n_2374),
.Y(n_3074)
);

INVx3_ASAP7_75t_L g3075 ( 
.A(n_2524),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2675),
.B(n_2215),
.Y(n_3076)
);

BUFx2_ASAP7_75t_L g3077 ( 
.A(n_2723),
.Y(n_3077)
);

INVx1_ASAP7_75t_L g3078 ( 
.A(n_2548),
.Y(n_3078)
);

NAND2xp5_ASAP7_75t_L g3079 ( 
.A(n_2598),
.B(n_2331),
.Y(n_3079)
);

INVx1_ASAP7_75t_L g3080 ( 
.A(n_2549),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2558),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2559),
.Y(n_3082)
);

NOR2xp33_ASAP7_75t_L g3083 ( 
.A(n_2723),
.B(n_2202),
.Y(n_3083)
);

NOR2xp33_ASAP7_75t_L g3084 ( 
.A(n_2727),
.B(n_2202),
.Y(n_3084)
);

INVxp33_ASAP7_75t_L g3085 ( 
.A(n_2727),
.Y(n_3085)
);

INVxp67_ASAP7_75t_SL g3086 ( 
.A(n_2515),
.Y(n_3086)
);

INVx1_ASAP7_75t_L g3087 ( 
.A(n_2561),
.Y(n_3087)
);

AND2x6_ASAP7_75t_L g3088 ( 
.A(n_2479),
.B(n_2265),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2563),
.Y(n_3089)
);

INVx4_ASAP7_75t_L g3090 ( 
.A(n_2524),
.Y(n_3090)
);

NAND2xp5_ASAP7_75t_L g3091 ( 
.A(n_2599),
.B(n_2216),
.Y(n_3091)
);

OR2x6_ASAP7_75t_L g3092 ( 
.A(n_2617),
.B(n_2374),
.Y(n_3092)
);

NAND2xp5_ASAP7_75t_L g3093 ( 
.A(n_2600),
.B(n_2216),
.Y(n_3093)
);

INVx3_ASAP7_75t_L g3094 ( 
.A(n_2524),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2406),
.B(n_2284),
.Y(n_3095)
);

INVx3_ASAP7_75t_L g3096 ( 
.A(n_2524),
.Y(n_3096)
);

INVx5_ASAP7_75t_L g3097 ( 
.A(n_2515),
.Y(n_3097)
);

NAND2xp5_ASAP7_75t_L g3098 ( 
.A(n_2601),
.B(n_2284),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_2570),
.Y(n_3099)
);

BUFx2_ASAP7_75t_L g3100 ( 
.A(n_2480),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2557),
.Y(n_3101)
);

NOR2x1p5_ASAP7_75t_L g3102 ( 
.A(n_2753),
.B(n_2128),
.Y(n_3102)
);

INVx2_ASAP7_75t_L g3103 ( 
.A(n_2474),
.Y(n_3103)
);

AND2x6_ASAP7_75t_L g3104 ( 
.A(n_2479),
.B(n_2266),
.Y(n_3104)
);

BUFx3_ASAP7_75t_L g3105 ( 
.A(n_2737),
.Y(n_3105)
);

BUFx4f_ASAP7_75t_L g3106 ( 
.A(n_2414),
.Y(n_3106)
);

AOI22xp5_ASAP7_75t_L g3107 ( 
.A1(n_2518),
.A2(n_2530),
.B1(n_2556),
.B2(n_2381),
.Y(n_3107)
);

INVxp67_ASAP7_75t_L g3108 ( 
.A(n_2518),
.Y(n_3108)
);

BUFx3_ASAP7_75t_L g3109 ( 
.A(n_2574),
.Y(n_3109)
);

INVx1_ASAP7_75t_SL g3110 ( 
.A(n_2728),
.Y(n_3110)
);

BUFx6f_ASAP7_75t_L g3111 ( 
.A(n_2557),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2575),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2474),
.Y(n_3113)
);

INVx1_ASAP7_75t_SL g3114 ( 
.A(n_2751),
.Y(n_3114)
);

NOR2xp33_ASAP7_75t_L g3115 ( 
.A(n_2688),
.B(n_2261),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2557),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_SL g3117 ( 
.A(n_2607),
.B(n_2311),
.Y(n_3117)
);

INVx2_ASAP7_75t_L g3118 ( 
.A(n_2478),
.Y(n_3118)
);

NAND2x1p5_ASAP7_75t_L g3119 ( 
.A(n_2457),
.B(n_2458),
.Y(n_3119)
);

BUFx4f_ASAP7_75t_L g3120 ( 
.A(n_2735),
.Y(n_3120)
);

NAND3xp33_ASAP7_75t_L g3121 ( 
.A(n_2499),
.B(n_2233),
.C(n_2311),
.Y(n_3121)
);

BUFx6f_ASAP7_75t_L g3122 ( 
.A(n_2557),
.Y(n_3122)
);

BUFx6f_ASAP7_75t_L g3123 ( 
.A(n_2562),
.Y(n_3123)
);

NOR2xp33_ASAP7_75t_L g3124 ( 
.A(n_2689),
.B(n_2690),
.Y(n_3124)
);

INVx2_ASAP7_75t_L g3125 ( 
.A(n_2478),
.Y(n_3125)
);

CKINVDCx20_ASAP7_75t_R g3126 ( 
.A(n_2510),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2483),
.Y(n_3127)
);

NAND2x1p5_ASAP7_75t_L g3128 ( 
.A(n_2457),
.B(n_2458),
.Y(n_3128)
);

AND2x4_ASAP7_75t_L g3129 ( 
.A(n_2755),
.B(n_2117),
.Y(n_3129)
);

INVx5_ASAP7_75t_L g3130 ( 
.A(n_2515),
.Y(n_3130)
);

AND3x2_ASAP7_75t_L g3131 ( 
.A(n_2738),
.B(n_2355),
.C(n_2329),
.Y(n_3131)
);

INVx4_ASAP7_75t_L g3132 ( 
.A(n_2562),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2581),
.Y(n_3133)
);

BUFx3_ASAP7_75t_L g3134 ( 
.A(n_2589),
.Y(n_3134)
);

INVx2_ASAP7_75t_L g3135 ( 
.A(n_2483),
.Y(n_3135)
);

BUFx10_ASAP7_75t_L g3136 ( 
.A(n_2693),
.Y(n_3136)
);

INVx2_ASAP7_75t_L g3137 ( 
.A(n_2491),
.Y(n_3137)
);

BUFx6f_ASAP7_75t_L g3138 ( 
.A(n_2562),
.Y(n_3138)
);

AND2x4_ASAP7_75t_L g3139 ( 
.A(n_2712),
.B(n_2198),
.Y(n_3139)
);

NAND2xp5_ASAP7_75t_SL g3140 ( 
.A(n_2626),
.B(n_2329),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2604),
.B(n_2198),
.Y(n_3141)
);

NAND2xp5_ASAP7_75t_L g3142 ( 
.A(n_2608),
.B(n_2200),
.Y(n_3142)
);

OR2x2_ASAP7_75t_L g3143 ( 
.A(n_2567),
.B(n_2355),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2739),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2722),
.Y(n_3145)
);

BUFx10_ASAP7_75t_L g3146 ( 
.A(n_2693),
.Y(n_3146)
);

INVx2_ASAP7_75t_L g3147 ( 
.A(n_2491),
.Y(n_3147)
);

AND2x4_ASAP7_75t_L g3148 ( 
.A(n_2714),
.B(n_2200),
.Y(n_3148)
);

INVx1_ASAP7_75t_L g3149 ( 
.A(n_2722),
.Y(n_3149)
);

OR2x2_ASAP7_75t_L g3150 ( 
.A(n_2635),
.B(n_2374),
.Y(n_3150)
);

NOR3xp33_ASAP7_75t_L g3151 ( 
.A(n_2617),
.B(n_2314),
.C(n_2031),
.Y(n_3151)
);

NOR2xp33_ASAP7_75t_L g3152 ( 
.A(n_2695),
.B(n_2271),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2390),
.Y(n_3153)
);

INVx4_ASAP7_75t_L g3154 ( 
.A(n_2562),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2390),
.Y(n_3155)
);

AND3x4_ASAP7_75t_L g3156 ( 
.A(n_2510),
.B(n_2204),
.C(n_2167),
.Y(n_3156)
);

NOR2xp33_ASAP7_75t_L g3157 ( 
.A(n_2614),
.B(n_2272),
.Y(n_3157)
);

NOR2xp33_ASAP7_75t_L g3158 ( 
.A(n_2615),
.B(n_2618),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2493),
.Y(n_3159)
);

NAND2x1p5_ASAP7_75t_L g3160 ( 
.A(n_2576),
.B(n_2353),
.Y(n_3160)
);

INVx1_ASAP7_75t_L g3161 ( 
.A(n_2392),
.Y(n_3161)
);

INVx3_ASAP7_75t_L g3162 ( 
.A(n_2571),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_SL g3163 ( 
.A(n_2566),
.B(n_2275),
.Y(n_3163)
);

INVx4_ASAP7_75t_L g3164 ( 
.A(n_2571),
.Y(n_3164)
);

NAND2xp5_ASAP7_75t_L g3165 ( 
.A(n_2619),
.B(n_2218),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2392),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2721),
.Y(n_3167)
);

AND2x2_ASAP7_75t_L g3168 ( 
.A(n_2725),
.B(n_2276),
.Y(n_3168)
);

NOR2xp33_ASAP7_75t_SL g3169 ( 
.A(n_2456),
.B(n_2197),
.Y(n_3169)
);

INVx1_ASAP7_75t_L g3170 ( 
.A(n_2730),
.Y(n_3170)
);

NAND2xp5_ASAP7_75t_L g3171 ( 
.A(n_2623),
.B(n_2218),
.Y(n_3171)
);

INVx3_ASAP7_75t_L g3172 ( 
.A(n_2571),
.Y(n_3172)
);

INVx6_ASAP7_75t_L g3173 ( 
.A(n_2571),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2624),
.B(n_2218),
.Y(n_3174)
);

INVx2_ASAP7_75t_L g3175 ( 
.A(n_2493),
.Y(n_3175)
);

INVx1_ASAP7_75t_SL g3176 ( 
.A(n_2652),
.Y(n_3176)
);

INVx4_ASAP7_75t_L g3177 ( 
.A(n_2582),
.Y(n_3177)
);

HB1xp67_ASAP7_75t_L g3178 ( 
.A(n_2731),
.Y(n_3178)
);

BUFx2_ASAP7_75t_L g3179 ( 
.A(n_2693),
.Y(n_3179)
);

INVx1_ASAP7_75t_L g3180 ( 
.A(n_2625),
.Y(n_3180)
);

NOR2xp33_ASAP7_75t_L g3181 ( 
.A(n_2628),
.B(n_2664),
.Y(n_3181)
);

INVx4_ASAP7_75t_SL g3182 ( 
.A(n_2687),
.Y(n_3182)
);

BUFx3_ASAP7_75t_L g3183 ( 
.A(n_2663),
.Y(n_3183)
);

INVxp67_ASAP7_75t_SL g3184 ( 
.A(n_2515),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_2666),
.B(n_2189),
.Y(n_3185)
);

AND2x6_ASAP7_75t_L g3186 ( 
.A(n_2767),
.B(n_2337),
.Y(n_3186)
);

NOR2xp33_ASAP7_75t_L g3187 ( 
.A(n_2672),
.B(n_1996),
.Y(n_3187)
);

AND2x4_ASAP7_75t_L g3188 ( 
.A(n_2530),
.B(n_2337),
.Y(n_3188)
);

INVx4_ASAP7_75t_L g3189 ( 
.A(n_2582),
.Y(n_3189)
);

INVx2_ASAP7_75t_L g3190 ( 
.A(n_2498),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2676),
.Y(n_3191)
);

BUFx6f_ASAP7_75t_L g3192 ( 
.A(n_2582),
.Y(n_3192)
);

OR2x2_ASAP7_75t_L g3193 ( 
.A(n_2694),
.B(n_2337),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2677),
.Y(n_3194)
);

INVx2_ASAP7_75t_SL g3195 ( 
.A(n_2705),
.Y(n_3195)
);

INVx2_ASAP7_75t_L g3196 ( 
.A(n_2498),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_L g3197 ( 
.A(n_2911),
.B(n_2713),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_SL g3198 ( 
.A(n_2918),
.B(n_2337),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_2911),
.B(n_2460),
.Y(n_3199)
);

OAI22xp5_ASAP7_75t_L g3200 ( 
.A1(n_2832),
.A2(n_2907),
.B1(n_2844),
.B2(n_2995),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_2832),
.B(n_2471),
.Y(n_3201)
);

AOI22xp5_ASAP7_75t_L g3202 ( 
.A1(n_2918),
.A2(n_2031),
.B1(n_2204),
.B2(n_2167),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2807),
.Y(n_3203)
);

INVx4_ASAP7_75t_L g3204 ( 
.A(n_2777),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_SL g3205 ( 
.A(n_2931),
.B(n_2342),
.Y(n_3205)
);

BUFx3_ASAP7_75t_L g3206 ( 
.A(n_2801),
.Y(n_3206)
);

OAI22xp33_ASAP7_75t_L g3207 ( 
.A1(n_2931),
.A2(n_2683),
.B1(n_2685),
.B2(n_2681),
.Y(n_3207)
);

INVx4_ASAP7_75t_L g3208 ( 
.A(n_2777),
.Y(n_3208)
);

INVx2_ASAP7_75t_L g3209 ( 
.A(n_2792),
.Y(n_3209)
);

INVx2_ASAP7_75t_SL g3210 ( 
.A(n_3031),
.Y(n_3210)
);

NAND2xp5_ASAP7_75t_SL g3211 ( 
.A(n_3031),
.B(n_2342),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_2844),
.B(n_2476),
.Y(n_3212)
);

AND2x2_ASAP7_75t_L g3213 ( 
.A(n_2819),
.B(n_2342),
.Y(n_3213)
);

OR2x2_ASAP7_75t_L g3214 ( 
.A(n_3056),
.B(n_2342),
.Y(n_3214)
);

INVx2_ASAP7_75t_L g3215 ( 
.A(n_2795),
.Y(n_3215)
);

NAND2xp5_ASAP7_75t_L g3216 ( 
.A(n_2907),
.B(n_2487),
.Y(n_3216)
);

AOI22xp33_ASAP7_75t_L g3217 ( 
.A1(n_2885),
.A2(n_2693),
.B1(n_2764),
.B2(n_2475),
.Y(n_3217)
);

NAND2xp5_ASAP7_75t_SL g3218 ( 
.A(n_3046),
.B(n_2592),
.Y(n_3218)
);

OAI22xp5_ASAP7_75t_L g3219 ( 
.A1(n_2995),
.A2(n_2749),
.B1(n_2536),
.B2(n_2036),
.Y(n_3219)
);

AOI22xp33_ASAP7_75t_L g3220 ( 
.A1(n_2885),
.A2(n_2693),
.B1(n_2764),
.B2(n_2475),
.Y(n_3220)
);

NAND2xp5_ASAP7_75t_L g3221 ( 
.A(n_2954),
.B(n_2764),
.Y(n_3221)
);

NAND2xp5_ASAP7_75t_L g3222 ( 
.A(n_2820),
.B(n_2764),
.Y(n_3222)
);

NAND2xp5_ASAP7_75t_L g3223 ( 
.A(n_2820),
.B(n_2764),
.Y(n_3223)
);

NAND2xp5_ASAP7_75t_L g3224 ( 
.A(n_3056),
.B(n_2749),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_L g3225 ( 
.A(n_3069),
.B(n_2036),
.Y(n_3225)
);

AOI21xp5_ASAP7_75t_L g3226 ( 
.A1(n_2780),
.A2(n_2761),
.B(n_2763),
.Y(n_3226)
);

NOR2xp33_ASAP7_75t_L g3227 ( 
.A(n_2899),
.B(n_2766),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_2808),
.Y(n_3228)
);

INVx1_ASAP7_75t_L g3229 ( 
.A(n_2811),
.Y(n_3229)
);

NAND2xp5_ASAP7_75t_L g3230 ( 
.A(n_3069),
.B(n_2036),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_2798),
.Y(n_3231)
);

INVx4_ASAP7_75t_L g3232 ( 
.A(n_2887),
.Y(n_3232)
);

AND2x2_ASAP7_75t_L g3233 ( 
.A(n_3076),
.B(n_2987),
.Y(n_3233)
);

INVx1_ASAP7_75t_L g3234 ( 
.A(n_2817),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3061),
.B(n_2473),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3061),
.B(n_2473),
.Y(n_3236)
);

NAND2xp5_ASAP7_75t_L g3237 ( 
.A(n_2818),
.B(n_2592),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_2818),
.B(n_2603),
.Y(n_3238)
);

NAND2xp5_ASAP7_75t_L g3239 ( 
.A(n_2815),
.B(n_2603),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_2825),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_2827),
.Y(n_3241)
);

AOI22xp5_ASAP7_75t_L g3242 ( 
.A1(n_2980),
.A2(n_2270),
.B1(n_2280),
.B2(n_2219),
.Y(n_3242)
);

AND2x4_ASAP7_75t_L g3243 ( 
.A(n_2783),
.B(n_2876),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_2815),
.B(n_2766),
.Y(n_3244)
);

NOR2xp33_ASAP7_75t_L g3245 ( 
.A(n_2812),
.B(n_2396),
.Y(n_3245)
);

NOR3xp33_ASAP7_75t_L g3246 ( 
.A(n_3121),
.B(n_2333),
.C(n_981),
.Y(n_3246)
);

NOR2xp33_ASAP7_75t_L g3247 ( 
.A(n_2812),
.B(n_2427),
.Y(n_3247)
);

INVx8_ASAP7_75t_L g3248 ( 
.A(n_2830),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_2780),
.A2(n_2761),
.B(n_2763),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_2824),
.B(n_2441),
.Y(n_3250)
);

NOR2x1_ASAP7_75t_R g3251 ( 
.A(n_2789),
.B(n_2219),
.Y(n_3251)
);

AOI22xp33_ASAP7_75t_L g3252 ( 
.A1(n_2985),
.A2(n_1037),
.B1(n_1120),
.B2(n_1050),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2824),
.B(n_2503),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2840),
.Y(n_3254)
);

AND2x2_ASAP7_75t_L g3255 ( 
.A(n_3064),
.B(n_1800),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_L g3256 ( 
.A(n_3095),
.B(n_2802),
.Y(n_3256)
);

AND2x6_ASAP7_75t_SL g3257 ( 
.A(n_3024),
.B(n_2270),
.Y(n_3257)
);

NOR2xp33_ASAP7_75t_L g3258 ( 
.A(n_2863),
.B(n_2280),
.Y(n_3258)
);

INVx1_ASAP7_75t_L g3259 ( 
.A(n_2843),
.Y(n_3259)
);

INVx1_ASAP7_75t_L g3260 ( 
.A(n_2847),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_SL g3261 ( 
.A(n_3046),
.B(n_2757),
.Y(n_3261)
);

INVx4_ASAP7_75t_L g3262 ( 
.A(n_2887),
.Y(n_3262)
);

INVx2_ASAP7_75t_SL g3263 ( 
.A(n_2889),
.Y(n_3263)
);

INVx2_ASAP7_75t_L g3264 ( 
.A(n_2803),
.Y(n_3264)
);

NOR3x1_ASAP7_75t_L g3265 ( 
.A(n_2973),
.B(n_984),
.C(n_980),
.Y(n_3265)
);

BUFx6f_ASAP7_75t_L g3266 ( 
.A(n_3111),
.Y(n_3266)
);

INVxp67_ASAP7_75t_L g3267 ( 
.A(n_2858),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_2802),
.B(n_2503),
.Y(n_3268)
);

NAND2xp5_ASAP7_75t_L g3269 ( 
.A(n_3051),
.B(n_2508),
.Y(n_3269)
);

BUFx6f_ASAP7_75t_L g3270 ( 
.A(n_3111),
.Y(n_3270)
);

AOI22xp33_ASAP7_75t_SL g3271 ( 
.A1(n_3030),
.A2(n_2320),
.B1(n_2323),
.B2(n_2291),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_2848),
.Y(n_3272)
);

OAI22xp5_ASAP7_75t_L g3273 ( 
.A1(n_3020),
.A2(n_2776),
.B1(n_2649),
.B2(n_2658),
.Y(n_3273)
);

INVxp33_ASAP7_75t_L g3274 ( 
.A(n_2858),
.Y(n_3274)
);

INVx3_ASAP7_75t_L g3275 ( 
.A(n_2805),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3051),
.B(n_2508),
.Y(n_3276)
);

AOI22xp5_ASAP7_75t_L g3277 ( 
.A1(n_2934),
.A2(n_2320),
.B1(n_2323),
.B2(n_2291),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_2946),
.B(n_2509),
.Y(n_3278)
);

INVx2_ASAP7_75t_SL g3279 ( 
.A(n_2960),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_2946),
.B(n_2509),
.Y(n_3280)
);

INVx2_ASAP7_75t_SL g3281 ( 
.A(n_3000),
.Y(n_3281)
);

XOR2xp5_ASAP7_75t_L g3282 ( 
.A(n_2904),
.B(n_1800),
.Y(n_3282)
);

NAND2xp5_ASAP7_75t_L g3283 ( 
.A(n_2956),
.B(n_2519),
.Y(n_3283)
);

INVx2_ASAP7_75t_SL g3284 ( 
.A(n_2853),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_2956),
.B(n_2519),
.Y(n_3285)
);

HB1xp67_ASAP7_75t_L g3286 ( 
.A(n_2781),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2851),
.Y(n_3287)
);

OR2x6_ASAP7_75t_L g3288 ( 
.A(n_2830),
.B(n_2729),
.Y(n_3288)
);

NAND2xp33_ASAP7_75t_L g3289 ( 
.A(n_3033),
.B(n_2582),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_2810),
.Y(n_3290)
);

INVx2_ASAP7_75t_L g3291 ( 
.A(n_2813),
.Y(n_3291)
);

AOI22xp33_ASAP7_75t_L g3292 ( 
.A1(n_2985),
.A2(n_1037),
.B1(n_1120),
.B2(n_999),
.Y(n_3292)
);

NOR2xp33_ASAP7_75t_L g3293 ( 
.A(n_2839),
.B(n_2340),
.Y(n_3293)
);

AND2x2_ASAP7_75t_L g3294 ( 
.A(n_2821),
.B(n_1823),
.Y(n_3294)
);

NAND2xp5_ASAP7_75t_L g3295 ( 
.A(n_3176),
.B(n_2523),
.Y(n_3295)
);

NOR2xp33_ASAP7_75t_L g3296 ( 
.A(n_2839),
.B(n_2340),
.Y(n_3296)
);

NAND2xp5_ASAP7_75t_L g3297 ( 
.A(n_3176),
.B(n_2523),
.Y(n_3297)
);

INVx5_ASAP7_75t_L g3298 ( 
.A(n_2804),
.Y(n_3298)
);

INVx8_ASAP7_75t_L g3299 ( 
.A(n_2830),
.Y(n_3299)
);

NOR2xp33_ASAP7_75t_L g3300 ( 
.A(n_2861),
.B(n_1823),
.Y(n_3300)
);

NAND2xp5_ASAP7_75t_SL g3301 ( 
.A(n_2926),
.B(n_2757),
.Y(n_3301)
);

NAND2xp5_ASAP7_75t_L g3302 ( 
.A(n_2964),
.B(n_2526),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_2862),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_2842),
.B(n_1827),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_2822),
.Y(n_3305)
);

INVx1_ASAP7_75t_L g3306 ( 
.A(n_2865),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_2868),
.Y(n_3307)
);

OAI21xp5_ASAP7_75t_L g3308 ( 
.A1(n_2972),
.A2(n_2649),
.B(n_2637),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_SL g3309 ( 
.A(n_2926),
.B(n_2757),
.Y(n_3309)
);

NAND2xp5_ASAP7_75t_L g3310 ( 
.A(n_2964),
.B(n_2526),
.Y(n_3310)
);

BUFx6f_ASAP7_75t_L g3311 ( 
.A(n_3111),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2800),
.B(n_2527),
.Y(n_3312)
);

NAND2xp5_ASAP7_75t_SL g3313 ( 
.A(n_2861),
.B(n_2757),
.Y(n_3313)
);

AOI21xp5_ASAP7_75t_L g3314 ( 
.A1(n_2890),
.A2(n_2459),
.B(n_2417),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_3021),
.B(n_2527),
.Y(n_3315)
);

NOR2xp33_ASAP7_75t_L g3316 ( 
.A(n_2782),
.B(n_2637),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_2850),
.B(n_1827),
.Y(n_3317)
);

BUFx6f_ASAP7_75t_L g3318 ( 
.A(n_3116),
.Y(n_3318)
);

INVx2_ASAP7_75t_L g3319 ( 
.A(n_2838),
.Y(n_3319)
);

BUFx6f_ASAP7_75t_L g3320 ( 
.A(n_3116),
.Y(n_3320)
);

INVx2_ASAP7_75t_SL g3321 ( 
.A(n_2786),
.Y(n_3321)
);

INVxp33_ASAP7_75t_L g3322 ( 
.A(n_2785),
.Y(n_3322)
);

INVx1_ASAP7_75t_L g3323 ( 
.A(n_2871),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2891),
.Y(n_3324)
);

NAND2xp5_ASAP7_75t_L g3325 ( 
.A(n_2782),
.B(n_2533),
.Y(n_3325)
);

NAND2xp5_ASAP7_75t_L g3326 ( 
.A(n_3025),
.B(n_2533),
.Y(n_3326)
);

NAND2xp5_ASAP7_75t_SL g3327 ( 
.A(n_2886),
.B(n_2772),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_2845),
.Y(n_3328)
);

AOI22xp33_ASAP7_75t_L g3329 ( 
.A1(n_2953),
.A2(n_1050),
.B1(n_1120),
.B2(n_1037),
.Y(n_3329)
);

O2A1O1Ixp33_ASAP7_75t_L g3330 ( 
.A1(n_2864),
.A2(n_2750),
.B(n_2742),
.C(n_2720),
.Y(n_3330)
);

INVx1_ASAP7_75t_L g3331 ( 
.A(n_2893),
.Y(n_3331)
);

NAND2xp5_ASAP7_75t_L g3332 ( 
.A(n_3025),
.B(n_2543),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_3083),
.B(n_2543),
.Y(n_3333)
);

OAI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3009),
.A2(n_2776),
.B1(n_2720),
.B2(n_2658),
.Y(n_3334)
);

NOR2xp33_ASAP7_75t_L g3335 ( 
.A(n_2797),
.B(n_2576),
.Y(n_3335)
);

AOI22xp33_ASAP7_75t_L g3336 ( 
.A1(n_2953),
.A2(n_1050),
.B1(n_1120),
.B2(n_1037),
.Y(n_3336)
);

NAND2xp5_ASAP7_75t_SL g3337 ( 
.A(n_2886),
.B(n_2717),
.Y(n_3337)
);

NOR2xp33_ASAP7_75t_L g3338 ( 
.A(n_2797),
.B(n_2576),
.Y(n_3338)
);

AOI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_2870),
.A2(n_1841),
.B1(n_1829),
.B2(n_2212),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3083),
.B(n_2547),
.Y(n_3340)
);

AOI22xp33_ASAP7_75t_L g3341 ( 
.A1(n_2857),
.A2(n_2917),
.B1(n_3156),
.B2(n_2882),
.Y(n_3341)
);

NOR2xp33_ASAP7_75t_L g3342 ( 
.A(n_3018),
.B(n_2595),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_L g3343 ( 
.A(n_3084),
.B(n_2547),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3084),
.B(n_2551),
.Y(n_3344)
);

NAND2xp5_ASAP7_75t_SL g3345 ( 
.A(n_2974),
.B(n_2772),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_SL g3346 ( 
.A(n_3129),
.B(n_2814),
.Y(n_3346)
);

NAND2xp5_ASAP7_75t_L g3347 ( 
.A(n_2945),
.B(n_2551),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_2894),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_2945),
.B(n_2555),
.Y(n_3349)
);

INVx1_ASAP7_75t_L g3350 ( 
.A(n_2905),
.Y(n_3350)
);

NAND2xp5_ASAP7_75t_L g3351 ( 
.A(n_2950),
.B(n_2555),
.Y(n_3351)
);

INVx2_ASAP7_75t_L g3352 ( 
.A(n_2849),
.Y(n_3352)
);

NAND2xp5_ASAP7_75t_L g3353 ( 
.A(n_2950),
.B(n_2569),
.Y(n_3353)
);

INVx1_ASAP7_75t_L g3354 ( 
.A(n_2906),
.Y(n_3354)
);

INVx2_ASAP7_75t_L g3355 ( 
.A(n_2859),
.Y(n_3355)
);

INVx2_ASAP7_75t_L g3356 ( 
.A(n_2866),
.Y(n_3356)
);

INVx1_ASAP7_75t_SL g3357 ( 
.A(n_2943),
.Y(n_3357)
);

AOI22xp5_ASAP7_75t_L g3358 ( 
.A1(n_2895),
.A2(n_1841),
.B1(n_1829),
.B2(n_2212),
.Y(n_3358)
);

OAI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3107),
.A2(n_1196),
.B1(n_1188),
.B2(n_1082),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3060),
.B(n_2569),
.Y(n_3360)
);

NAND2xp5_ASAP7_75t_L g3361 ( 
.A(n_2781),
.B(n_2572),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_SL g3362 ( 
.A(n_3129),
.B(n_2772),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3054),
.B(n_2572),
.Y(n_3363)
);

INVx2_ASAP7_75t_SL g3364 ( 
.A(n_2794),
.Y(n_3364)
);

INVx2_ASAP7_75t_SL g3365 ( 
.A(n_2799),
.Y(n_3365)
);

OAI22xp5_ASAP7_75t_SL g3366 ( 
.A1(n_2857),
.A2(n_2188),
.B1(n_876),
.B2(n_881),
.Y(n_3366)
);

O2A1O1Ixp5_ASAP7_75t_L g3367 ( 
.A1(n_2991),
.A2(n_2585),
.B(n_2613),
.C(n_2568),
.Y(n_3367)
);

NAND2xp5_ASAP7_75t_L g3368 ( 
.A(n_2902),
.B(n_2573),
.Y(n_3368)
);

AND2x2_ASAP7_75t_L g3369 ( 
.A(n_2876),
.B(n_1494),
.Y(n_3369)
);

AOI22xp5_ASAP7_75t_SL g3370 ( 
.A1(n_2947),
.A2(n_2313),
.B1(n_883),
.B2(n_884),
.Y(n_3370)
);

NAND2xp5_ASAP7_75t_L g3371 ( 
.A(n_2902),
.B(n_2573),
.Y(n_3371)
);

A2O1A1Ixp33_ASAP7_75t_L g3372 ( 
.A1(n_2991),
.A2(n_2585),
.B(n_2613),
.C(n_2568),
.Y(n_3372)
);

NOR2xp33_ASAP7_75t_L g3373 ( 
.A(n_3028),
.B(n_2313),
.Y(n_3373)
);

INVx2_ASAP7_75t_L g3374 ( 
.A(n_2874),
.Y(n_3374)
);

INVx2_ASAP7_75t_L g3375 ( 
.A(n_2877),
.Y(n_3375)
);

INVx1_ASAP7_75t_L g3376 ( 
.A(n_2919),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_2921),
.B(n_2579),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_2921),
.B(n_2949),
.Y(n_3378)
);

INVx2_ASAP7_75t_L g3379 ( 
.A(n_2883),
.Y(n_3379)
);

AOI22xp33_ASAP7_75t_L g3380 ( 
.A1(n_2917),
.A2(n_1050),
.B1(n_1214),
.B2(n_2579),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_2888),
.Y(n_3381)
);

INVx2_ASAP7_75t_SL g3382 ( 
.A(n_2912),
.Y(n_3382)
);

NAND2xp5_ASAP7_75t_L g3383 ( 
.A(n_2949),
.B(n_2583),
.Y(n_3383)
);

NAND2xp5_ASAP7_75t_L g3384 ( 
.A(n_2990),
.B(n_2583),
.Y(n_3384)
);

BUFx5_ASAP7_75t_L g3385 ( 
.A(n_3033),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_3023),
.A2(n_1214),
.B1(n_2593),
.B2(n_2588),
.Y(n_3386)
);

NAND2x1_ASAP7_75t_L g3387 ( 
.A(n_3173),
.B(n_2595),
.Y(n_3387)
);

NOR2x1p5_ASAP7_75t_L g3388 ( 
.A(n_2814),
.B(n_2776),
.Y(n_3388)
);

INVx1_ASAP7_75t_L g3389 ( 
.A(n_2920),
.Y(n_3389)
);

AOI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3059),
.A2(n_2631),
.B1(n_2633),
.B2(n_2629),
.Y(n_3390)
);

NAND2xp5_ASAP7_75t_L g3391 ( 
.A(n_2990),
.B(n_2588),
.Y(n_3391)
);

INVx2_ASAP7_75t_L g3392 ( 
.A(n_2901),
.Y(n_3392)
);

NAND2xp5_ASAP7_75t_L g3393 ( 
.A(n_3018),
.B(n_2593),
.Y(n_3393)
);

OAI22xp5_ASAP7_75t_L g3394 ( 
.A1(n_3009),
.A2(n_2595),
.B1(n_2512),
.B2(n_2538),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_2923),
.Y(n_3395)
);

NAND2xp5_ASAP7_75t_L g3396 ( 
.A(n_3037),
.B(n_2605),
.Y(n_3396)
);

NAND2xp5_ASAP7_75t_L g3397 ( 
.A(n_3037),
.B(n_2605),
.Y(n_3397)
);

INVx1_ASAP7_75t_L g3398 ( 
.A(n_2925),
.Y(n_3398)
);

NOR2x1p5_ASAP7_75t_L g3399 ( 
.A(n_2992),
.B(n_2500),
.Y(n_3399)
);

NAND2xp5_ASAP7_75t_SL g3400 ( 
.A(n_3015),
.B(n_2772),
.Y(n_3400)
);

AOI22xp5_ASAP7_75t_L g3401 ( 
.A1(n_2943),
.A2(n_2631),
.B1(n_2633),
.B2(n_2629),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3151),
.B(n_2610),
.Y(n_3402)
);

NAND2xp5_ASAP7_75t_L g3403 ( 
.A(n_3151),
.B(n_2610),
.Y(n_3403)
);

INVx3_ASAP7_75t_L g3404 ( 
.A(n_2805),
.Y(n_3404)
);

INVx3_ASAP7_75t_L g3405 ( 
.A(n_2778),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3109),
.B(n_3134),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_2927),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3115),
.B(n_2622),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_SL g3409 ( 
.A(n_3015),
.B(n_2710),
.Y(n_3409)
);

NAND2xp5_ASAP7_75t_L g3410 ( 
.A(n_3115),
.B(n_2622),
.Y(n_3410)
);

INVx3_ASAP7_75t_L g3411 ( 
.A(n_2778),
.Y(n_3411)
);

NAND2xp5_ASAP7_75t_SL g3412 ( 
.A(n_2963),
.B(n_3044),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_2929),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2909),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3035),
.B(n_2729),
.Y(n_3415)
);

NOR2xp33_ASAP7_75t_L g3416 ( 
.A(n_3070),
.B(n_2732),
.Y(n_3416)
);

NAND2xp5_ASAP7_75t_SL g3417 ( 
.A(n_3044),
.B(n_2717),
.Y(n_3417)
);

INVx1_ASAP7_75t_L g3418 ( 
.A(n_2930),
.Y(n_3418)
);

INVx1_ASAP7_75t_L g3419 ( 
.A(n_2944),
.Y(n_3419)
);

NAND2xp5_ASAP7_75t_L g3420 ( 
.A(n_3195),
.B(n_2642),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_2948),
.Y(n_3421)
);

NAND2xp5_ASAP7_75t_SL g3422 ( 
.A(n_3106),
.B(n_2717),
.Y(n_3422)
);

AOI22xp33_ASAP7_75t_L g3423 ( 
.A1(n_3023),
.A2(n_1214),
.B1(n_2647),
.B2(n_2642),
.Y(n_3423)
);

INVx1_ASAP7_75t_L g3424 ( 
.A(n_2955),
.Y(n_3424)
);

OAI22xp5_ASAP7_75t_L g3425 ( 
.A1(n_3067),
.A2(n_2512),
.B1(n_2538),
.B2(n_2500),
.Y(n_3425)
);

INVx2_ASAP7_75t_L g3426 ( 
.A(n_2933),
.Y(n_3426)
);

NAND2xp5_ASAP7_75t_L g3427 ( 
.A(n_3152),
.B(n_2647),
.Y(n_3427)
);

INVx1_ASAP7_75t_L g3428 ( 
.A(n_2959),
.Y(n_3428)
);

NAND2xp5_ASAP7_75t_L g3429 ( 
.A(n_3152),
.B(n_2650),
.Y(n_3429)
);

INVx2_ASAP7_75t_L g3430 ( 
.A(n_2936),
.Y(n_3430)
);

CKINVDCx5p33_ASAP7_75t_R g3431 ( 
.A(n_2855),
.Y(n_3431)
);

NAND2xp5_ASAP7_75t_SL g3432 ( 
.A(n_3106),
.B(n_2586),
.Y(n_3432)
);

NAND2xp5_ASAP7_75t_L g3433 ( 
.A(n_2962),
.B(n_2965),
.Y(n_3433)
);

NAND2xp5_ASAP7_75t_L g3434 ( 
.A(n_2966),
.B(n_2650),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_2970),
.Y(n_3435)
);

INVx2_ASAP7_75t_L g3436 ( 
.A(n_2938),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_SL g3437 ( 
.A(n_3041),
.B(n_2586),
.Y(n_3437)
);

NAND2xp5_ASAP7_75t_L g3438 ( 
.A(n_2975),
.B(n_2659),
.Y(n_3438)
);

AOI22xp33_ASAP7_75t_L g3439 ( 
.A1(n_2971),
.A2(n_1214),
.B1(n_2660),
.B2(n_2659),
.Y(n_3439)
);

A2O1A1Ixp33_ASAP7_75t_L g3440 ( 
.A1(n_2972),
.A2(n_2542),
.B(n_2560),
.C(n_2540),
.Y(n_3440)
);

INVx2_ASAP7_75t_L g3441 ( 
.A(n_2957),
.Y(n_3441)
);

INVxp67_ASAP7_75t_L g3442 ( 
.A(n_2788),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_2983),
.Y(n_3443)
);

NAND2xp5_ASAP7_75t_L g3444 ( 
.A(n_2988),
.B(n_2660),
.Y(n_3444)
);

NAND2xp5_ASAP7_75t_L g3445 ( 
.A(n_2994),
.B(n_2665),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_2997),
.Y(n_3446)
);

NOR2xp33_ASAP7_75t_L g3447 ( 
.A(n_3028),
.B(n_2732),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_2967),
.Y(n_3448)
);

NAND2xp5_ASAP7_75t_L g3449 ( 
.A(n_2998),
.B(n_2665),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3041),
.B(n_2586),
.Y(n_3450)
);

NOR2xp33_ASAP7_75t_L g3451 ( 
.A(n_3028),
.B(n_2734),
.Y(n_3451)
);

BUFx3_ASAP7_75t_L g3452 ( 
.A(n_2910),
.Y(n_3452)
);

AOI22xp33_ASAP7_75t_L g3453 ( 
.A1(n_2971),
.A2(n_2680),
.B1(n_2682),
.B2(n_2679),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3004),
.B(n_2679),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3005),
.Y(n_3455)
);

NAND3xp33_ASAP7_75t_L g3456 ( 
.A(n_3121),
.B(n_3053),
.C(n_3032),
.Y(n_3456)
);

NAND2xp5_ASAP7_75t_L g3457 ( 
.A(n_3007),
.B(n_2680),
.Y(n_3457)
);

NOR2xp33_ASAP7_75t_L g3458 ( 
.A(n_3085),
.B(n_2734),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3010),
.Y(n_3459)
);

OR2x6_ASAP7_75t_L g3460 ( 
.A(n_2783),
.B(n_2741),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_2969),
.Y(n_3461)
);

INVx2_ASAP7_75t_L g3462 ( 
.A(n_2986),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3034),
.B(n_2741),
.Y(n_3463)
);

O2A1O1Ixp5_ASAP7_75t_L g3464 ( 
.A1(n_3062),
.A2(n_2459),
.B(n_2417),
.C(n_2726),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3011),
.Y(n_3465)
);

OAI22x1_ASAP7_75t_L g3466 ( 
.A1(n_3100),
.A2(n_2542),
.B1(n_2560),
.B2(n_2540),
.Y(n_3466)
);

NOR2xp33_ASAP7_75t_L g3467 ( 
.A(n_3150),
.B(n_2744),
.Y(n_3467)
);

INVx1_ASAP7_75t_L g3468 ( 
.A(n_3026),
.Y(n_3468)
);

NAND2xp5_ASAP7_75t_L g3469 ( 
.A(n_3036),
.B(n_2682),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_2878),
.B(n_2586),
.Y(n_3470)
);

NAND2xp5_ASAP7_75t_L g3471 ( 
.A(n_3040),
.B(n_2702),
.Y(n_3471)
);

NAND2xp5_ASAP7_75t_L g3472 ( 
.A(n_3045),
.B(n_2702),
.Y(n_3472)
);

NAND2xp5_ASAP7_75t_L g3473 ( 
.A(n_3048),
.B(n_2709),
.Y(n_3473)
);

NOR2xp33_ASAP7_75t_R g3474 ( 
.A(n_2873),
.B(n_2632),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3052),
.Y(n_3475)
);

OAI22xp5_ASAP7_75t_L g3476 ( 
.A1(n_3067),
.A2(n_2564),
.B1(n_2597),
.B2(n_2553),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3066),
.B(n_2709),
.Y(n_3477)
);

NOR2xp33_ASAP7_75t_L g3478 ( 
.A(n_2979),
.B(n_2744),
.Y(n_3478)
);

AOI21xp5_ASAP7_75t_L g3479 ( 
.A1(n_2890),
.A2(n_2726),
.B(n_2742),
.Y(n_3479)
);

AOI22xp33_ASAP7_75t_L g3480 ( 
.A1(n_3145),
.A2(n_2716),
.B1(n_988),
.B2(n_992),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3071),
.Y(n_3481)
);

NAND2xp33_ASAP7_75t_L g3482 ( 
.A(n_3033),
.B(n_2632),
.Y(n_3482)
);

NAND2xp5_ASAP7_75t_SL g3483 ( 
.A(n_2914),
.B(n_2632),
.Y(n_3483)
);

INVx1_ASAP7_75t_L g3484 ( 
.A(n_3078),
.Y(n_3484)
);

INVxp67_ASAP7_75t_L g3485 ( 
.A(n_2860),
.Y(n_3485)
);

NAND2xp5_ASAP7_75t_L g3486 ( 
.A(n_3080),
.B(n_2716),
.Y(n_3486)
);

NOR2xp33_ASAP7_75t_L g3487 ( 
.A(n_3117),
.B(n_2759),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3081),
.B(n_2553),
.Y(n_3488)
);

NOR3xp33_ASAP7_75t_L g3489 ( 
.A(n_3140),
.B(n_988),
.C(n_984),
.Y(n_3489)
);

HB1xp67_ASAP7_75t_L g3490 ( 
.A(n_3049),
.Y(n_3490)
);

NOR2xp33_ASAP7_75t_L g3491 ( 
.A(n_3193),
.B(n_3068),
.Y(n_3491)
);

INVx3_ASAP7_75t_L g3492 ( 
.A(n_2796),
.Y(n_3492)
);

INVx2_ASAP7_75t_L g3493 ( 
.A(n_3002),
.Y(n_3493)
);

INVx2_ASAP7_75t_L g3494 ( 
.A(n_3008),
.Y(n_3494)
);

NAND2xp5_ASAP7_75t_SL g3495 ( 
.A(n_2978),
.B(n_2632),
.Y(n_3495)
);

NAND2xp5_ASAP7_75t_SL g3496 ( 
.A(n_2978),
.B(n_2646),
.Y(n_3496)
);

NOR2xp33_ASAP7_75t_L g3497 ( 
.A(n_3077),
.B(n_2759),
.Y(n_3497)
);

XOR2xp5_ASAP7_75t_L g3498 ( 
.A(n_3126),
.B(n_2750),
.Y(n_3498)
);

INVx1_ASAP7_75t_SL g3499 ( 
.A(n_2896),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3082),
.B(n_2564),
.Y(n_3500)
);

NAND2xp33_ASAP7_75t_L g3501 ( 
.A(n_3033),
.B(n_2646),
.Y(n_3501)
);

INVx2_ASAP7_75t_L g3502 ( 
.A(n_3013),
.Y(n_3502)
);

OAI221xp5_ASAP7_75t_L g3503 ( 
.A1(n_3091),
.A2(n_997),
.B1(n_1000),
.B2(n_995),
.C(n_992),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3087),
.Y(n_3504)
);

INVx1_ASAP7_75t_SL g3505 ( 
.A(n_2941),
.Y(n_3505)
);

O2A1O1Ixp33_ASAP7_75t_L g3506 ( 
.A1(n_2823),
.A2(n_2828),
.B(n_2961),
.C(n_3065),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3089),
.Y(n_3507)
);

INVx5_ASAP7_75t_L g3508 ( 
.A(n_2804),
.Y(n_3508)
);

INVx2_ASAP7_75t_L g3509 ( 
.A(n_3016),
.Y(n_3509)
);

AND2x2_ASAP7_75t_L g3510 ( 
.A(n_3168),
.B(n_1497),
.Y(n_3510)
);

INVx2_ASAP7_75t_SL g3511 ( 
.A(n_3102),
.Y(n_3511)
);

NAND2xp5_ASAP7_75t_L g3512 ( 
.A(n_3099),
.B(n_2597),
.Y(n_3512)
);

INVx2_ASAP7_75t_L g3513 ( 
.A(n_3017),
.Y(n_3513)
);

AOI22xp33_ASAP7_75t_L g3514 ( 
.A1(n_3149),
.A2(n_997),
.B1(n_1000),
.B2(n_995),
.Y(n_3514)
);

NAND2xp5_ASAP7_75t_L g3515 ( 
.A(n_3112),
.B(n_2612),
.Y(n_3515)
);

AOI22xp5_ASAP7_75t_L g3516 ( 
.A1(n_2976),
.A2(n_2687),
.B1(n_2620),
.B2(n_2669),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3133),
.B(n_2612),
.Y(n_3517)
);

A2O1A1Ixp33_ASAP7_75t_L g3518 ( 
.A1(n_2831),
.A2(n_2669),
.B(n_2678),
.C(n_2620),
.Y(n_3518)
);

AOI22xp33_ASAP7_75t_L g3519 ( 
.A1(n_3012),
.A2(n_1004),
.B1(n_1008),
.B2(n_1002),
.Y(n_3519)
);

AND2x4_ASAP7_75t_SL g3520 ( 
.A(n_2897),
.B(n_2646),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3178),
.B(n_3157),
.Y(n_3521)
);

NAND2xp5_ASAP7_75t_SL g3522 ( 
.A(n_2897),
.B(n_2646),
.Y(n_3522)
);

NOR2xp33_ASAP7_75t_L g3523 ( 
.A(n_2982),
.B(n_2678),
.Y(n_3523)
);

INVx4_ASAP7_75t_L g3524 ( 
.A(n_2804),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3178),
.B(n_2691),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3019),
.Y(n_3526)
);

NOR2xp67_ASAP7_75t_SL g3527 ( 
.A(n_2816),
.B(n_2670),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_SL g3528 ( 
.A(n_2916),
.B(n_2670),
.Y(n_3528)
);

INVx1_ASAP7_75t_L g3529 ( 
.A(n_3144),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_2867),
.B(n_1498),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3167),
.Y(n_3531)
);

NAND2xp5_ASAP7_75t_L g3532 ( 
.A(n_3157),
.B(n_2691),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3027),
.Y(n_3533)
);

AOI22xp33_ASAP7_75t_L g3534 ( 
.A1(n_3012),
.A2(n_1004),
.B1(n_1008),
.B2(n_1002),
.Y(n_3534)
);

BUFx3_ASAP7_75t_L g3535 ( 
.A(n_3024),
.Y(n_3535)
);

NAND3xp33_ASAP7_75t_L g3536 ( 
.A(n_3029),
.B(n_892),
.C(n_875),
.Y(n_3536)
);

NOR2xp33_ASAP7_75t_L g3537 ( 
.A(n_3143),
.B(n_2748),
.Y(n_3537)
);

AOI22xp5_ASAP7_75t_L g3538 ( 
.A1(n_2804),
.A2(n_2687),
.B1(n_2748),
.B2(n_896),
.Y(n_3538)
);

NAND2xp5_ASAP7_75t_L g3539 ( 
.A(n_3183),
.B(n_2687),
.Y(n_3539)
);

BUFx6f_ASAP7_75t_SL g3540 ( 
.A(n_3024),
.Y(n_3540)
);

NOR2xp33_ASAP7_75t_L g3541 ( 
.A(n_2928),
.B(n_2670),
.Y(n_3541)
);

NAND2xp5_ASAP7_75t_SL g3542 ( 
.A(n_2916),
.B(n_2670),
.Y(n_3542)
);

NOR2xp67_ASAP7_75t_L g3543 ( 
.A(n_2790),
.B(n_2710),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3170),
.Y(n_3544)
);

NAND2xp5_ASAP7_75t_L g3545 ( 
.A(n_3139),
.B(n_2710),
.Y(n_3545)
);

INVx3_ASAP7_75t_L g3546 ( 
.A(n_2796),
.Y(n_3546)
);

NOR2xp33_ASAP7_75t_L g3547 ( 
.A(n_3091),
.B(n_2710),
.Y(n_3547)
);

INVx2_ASAP7_75t_SL g3548 ( 
.A(n_2881),
.Y(n_3548)
);

AND2x2_ASAP7_75t_L g3549 ( 
.A(n_2884),
.B(n_2942),
.Y(n_3549)
);

AOI22xp33_ASAP7_75t_L g3550 ( 
.A1(n_3012),
.A2(n_1016),
.B1(n_1017),
.B2(n_1014),
.Y(n_3550)
);

INVx1_ASAP7_75t_L g3551 ( 
.A(n_3180),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_L g3552 ( 
.A(n_3139),
.B(n_2717),
.Y(n_3552)
);

INVx1_ASAP7_75t_L g3553 ( 
.A(n_3191),
.Y(n_3553)
);

INVx1_ASAP7_75t_L g3554 ( 
.A(n_3194),
.Y(n_3554)
);

CKINVDCx5p33_ASAP7_75t_R g3555 ( 
.A(n_3074),
.Y(n_3555)
);

NAND2xp5_ASAP7_75t_L g3556 ( 
.A(n_3148),
.B(n_1502),
.Y(n_3556)
);

INVx2_ASAP7_75t_L g3557 ( 
.A(n_3038),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3148),
.B(n_1510),
.Y(n_3558)
);

HB1xp67_ASAP7_75t_L g3559 ( 
.A(n_3074),
.Y(n_3559)
);

INVx1_ASAP7_75t_L g3560 ( 
.A(n_3124),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3047),
.Y(n_3561)
);

INVx2_ASAP7_75t_L g3562 ( 
.A(n_3055),
.Y(n_3562)
);

NOR2xp33_ASAP7_75t_L g3563 ( 
.A(n_2932),
.B(n_888),
.Y(n_3563)
);

INVx4_ASAP7_75t_L g3564 ( 
.A(n_2841),
.Y(n_3564)
);

NAND2xp5_ASAP7_75t_L g3565 ( 
.A(n_3093),
.B(n_1511),
.Y(n_3565)
);

NOR2xp33_ASAP7_75t_L g3566 ( 
.A(n_2937),
.B(n_898),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3074),
.B(n_1512),
.Y(n_3567)
);

NAND2xp5_ASAP7_75t_L g3568 ( 
.A(n_3093),
.B(n_1513),
.Y(n_3568)
);

NAND2xp5_ASAP7_75t_L g3569 ( 
.A(n_3098),
.B(n_1514),
.Y(n_3569)
);

NAND2xp5_ASAP7_75t_L g3570 ( 
.A(n_3098),
.B(n_1515),
.Y(n_3570)
);

NAND2xp5_ASAP7_75t_L g3571 ( 
.A(n_3188),
.B(n_1516),
.Y(n_3571)
);

AOI21xp5_ASAP7_75t_L g3572 ( 
.A1(n_3086),
.A2(n_2189),
.B(n_2423),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3124),
.Y(n_3573)
);

AOI22xp5_ASAP7_75t_L g3574 ( 
.A1(n_2841),
.A2(n_905),
.B1(n_906),
.B2(n_903),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3200),
.B(n_2791),
.Y(n_3575)
);

CKINVDCx5p33_ASAP7_75t_R g3576 ( 
.A(n_3431),
.Y(n_3576)
);

INVx1_ASAP7_75t_L g3577 ( 
.A(n_3203),
.Y(n_3577)
);

NAND2xp5_ASAP7_75t_L g3578 ( 
.A(n_3256),
.B(n_3022),
.Y(n_3578)
);

INVx5_ASAP7_75t_L g3579 ( 
.A(n_3204),
.Y(n_3579)
);

NAND2xp5_ASAP7_75t_SL g3580 ( 
.A(n_3202),
.B(n_3120),
.Y(n_3580)
);

NAND2xp5_ASAP7_75t_L g3581 ( 
.A(n_3549),
.B(n_3043),
.Y(n_3581)
);

BUFx12f_ASAP7_75t_SL g3582 ( 
.A(n_3204),
.Y(n_3582)
);

INVx1_ASAP7_75t_L g3583 ( 
.A(n_3228),
.Y(n_3583)
);

INVx1_ASAP7_75t_L g3584 ( 
.A(n_3229),
.Y(n_3584)
);

AND2x4_ASAP7_75t_L g3585 ( 
.A(n_3243),
.B(n_2806),
.Y(n_3585)
);

NOR2x1p5_ASAP7_75t_L g3586 ( 
.A(n_3208),
.B(n_3014),
.Y(n_3586)
);

INVx1_ASAP7_75t_L g3587 ( 
.A(n_3234),
.Y(n_3587)
);

INVx1_ASAP7_75t_L g3588 ( 
.A(n_3240),
.Y(n_3588)
);

AOI22xp33_ASAP7_75t_L g3589 ( 
.A1(n_3341),
.A2(n_3188),
.B1(n_2951),
.B2(n_2984),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3241),
.Y(n_3590)
);

INVx2_ASAP7_75t_L g3591 ( 
.A(n_3209),
.Y(n_3591)
);

NOR2x2_ASAP7_75t_L g3592 ( 
.A(n_3251),
.B(n_3288),
.Y(n_3592)
);

INVxp67_ASAP7_75t_L g3593 ( 
.A(n_3300),
.Y(n_3593)
);

BUFx6f_ASAP7_75t_L g3594 ( 
.A(n_3208),
.Y(n_3594)
);

INVx2_ASAP7_75t_L g3595 ( 
.A(n_3215),
.Y(n_3595)
);

BUFx6f_ASAP7_75t_L g3596 ( 
.A(n_3243),
.Y(n_3596)
);

AOI22xp33_ASAP7_75t_L g3597 ( 
.A1(n_3341),
.A2(n_2951),
.B1(n_2984),
.B2(n_2952),
.Y(n_3597)
);

AOI22xp5_ASAP7_75t_L g3598 ( 
.A1(n_3489),
.A2(n_2791),
.B1(n_2852),
.B2(n_2841),
.Y(n_3598)
);

BUFx6f_ASAP7_75t_L g3599 ( 
.A(n_3266),
.Y(n_3599)
);

NAND2xp5_ASAP7_75t_L g3600 ( 
.A(n_3245),
.B(n_3247),
.Y(n_3600)
);

NAND2xp5_ASAP7_75t_L g3601 ( 
.A(n_3245),
.B(n_2791),
.Y(n_3601)
);

INVx3_ASAP7_75t_L g3602 ( 
.A(n_3524),
.Y(n_3602)
);

AND3x1_ASAP7_75t_L g3603 ( 
.A(n_3258),
.B(n_3169),
.C(n_1196),
.Y(n_3603)
);

INVx1_ASAP7_75t_L g3604 ( 
.A(n_3254),
.Y(n_3604)
);

INVx5_ASAP7_75t_L g3605 ( 
.A(n_3298),
.Y(n_3605)
);

INVxp67_ASAP7_75t_L g3606 ( 
.A(n_3233),
.Y(n_3606)
);

BUFx3_ASAP7_75t_L g3607 ( 
.A(n_3206),
.Y(n_3607)
);

INVx2_ASAP7_75t_SL g3608 ( 
.A(n_3248),
.Y(n_3608)
);

NAND2xp5_ASAP7_75t_SL g3609 ( 
.A(n_3298),
.B(n_3120),
.Y(n_3609)
);

AND2x2_ASAP7_75t_L g3610 ( 
.A(n_3255),
.B(n_3131),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3499),
.B(n_3014),
.Y(n_3611)
);

INVx2_ASAP7_75t_L g3612 ( 
.A(n_3231),
.Y(n_3612)
);

NOR3xp33_ASAP7_75t_SL g3613 ( 
.A(n_3346),
.B(n_2846),
.C(n_2989),
.Y(n_3613)
);

NAND2xp5_ASAP7_75t_L g3614 ( 
.A(n_3505),
.B(n_3131),
.Y(n_3614)
);

NAND2xp5_ASAP7_75t_L g3615 ( 
.A(n_3199),
.B(n_2984),
.Y(n_3615)
);

AOI22xp33_ASAP7_75t_L g3616 ( 
.A1(n_3366),
.A2(n_2984),
.B1(n_2952),
.B2(n_2833),
.Y(n_3616)
);

HB1xp67_ASAP7_75t_L g3617 ( 
.A(n_3490),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3442),
.B(n_2915),
.Y(n_3618)
);

NAND2xp33_ASAP7_75t_R g3619 ( 
.A(n_3474),
.B(n_3092),
.Y(n_3619)
);

NAND2xp5_ASAP7_75t_L g3620 ( 
.A(n_3442),
.B(n_3163),
.Y(n_3620)
);

AND2x2_ASAP7_75t_L g3621 ( 
.A(n_3369),
.B(n_3092),
.Y(n_3621)
);

AND2x4_ASAP7_75t_L g3622 ( 
.A(n_3399),
.B(n_3092),
.Y(n_3622)
);

NAND2x1p5_ASAP7_75t_L g3623 ( 
.A(n_3298),
.B(n_2816),
.Y(n_3623)
);

AND2x4_ASAP7_75t_SL g3624 ( 
.A(n_3524),
.B(n_2779),
.Y(n_3624)
);

OAI21xp5_ASAP7_75t_L g3625 ( 
.A1(n_3316),
.A2(n_2854),
.B(n_2837),
.Y(n_3625)
);

AO21x1_ASAP7_75t_L g3626 ( 
.A1(n_3359),
.A2(n_2854),
.B(n_2837),
.Y(n_3626)
);

NAND2xp5_ASAP7_75t_SL g3627 ( 
.A(n_3298),
.B(n_3508),
.Y(n_3627)
);

INVx1_ASAP7_75t_L g3628 ( 
.A(n_3259),
.Y(n_3628)
);

BUFx3_ASAP7_75t_L g3629 ( 
.A(n_3452),
.Y(n_3629)
);

INVx2_ASAP7_75t_L g3630 ( 
.A(n_3264),
.Y(n_3630)
);

INVx1_ASAP7_75t_L g3631 ( 
.A(n_3260),
.Y(n_3631)
);

BUFx2_ASAP7_75t_L g3632 ( 
.A(n_3210),
.Y(n_3632)
);

AND2x2_ASAP7_75t_L g3633 ( 
.A(n_3294),
.B(n_3073),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_SL g3634 ( 
.A(n_3508),
.B(n_3169),
.Y(n_3634)
);

AND2x4_ASAP7_75t_L g3635 ( 
.A(n_3520),
.B(n_2841),
.Y(n_3635)
);

INVx1_ASAP7_75t_L g3636 ( 
.A(n_3272),
.Y(n_3636)
);

INVx6_ASAP7_75t_L g3637 ( 
.A(n_3248),
.Y(n_3637)
);

AOI22xp33_ASAP7_75t_L g3638 ( 
.A1(n_3329),
.A2(n_3336),
.B1(n_3317),
.B2(n_3304),
.Y(n_3638)
);

NOR2xp33_ASAP7_75t_L g3639 ( 
.A(n_3293),
.B(n_2993),
.Y(n_3639)
);

INVx1_ASAP7_75t_L g3640 ( 
.A(n_3287),
.Y(n_3640)
);

BUFx3_ASAP7_75t_L g3641 ( 
.A(n_3284),
.Y(n_3641)
);

INVx1_ASAP7_75t_L g3642 ( 
.A(n_3303),
.Y(n_3642)
);

NAND2xp5_ASAP7_75t_L g3643 ( 
.A(n_3485),
.B(n_3073),
.Y(n_3643)
);

INVx2_ASAP7_75t_L g3644 ( 
.A(n_3290),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3288),
.B(n_2852),
.Y(n_3645)
);

NAND2xp5_ASAP7_75t_L g3646 ( 
.A(n_3485),
.B(n_3079),
.Y(n_3646)
);

INVx2_ASAP7_75t_L g3647 ( 
.A(n_3291),
.Y(n_3647)
);

INVx2_ASAP7_75t_SL g3648 ( 
.A(n_3248),
.Y(n_3648)
);

NAND3xp33_ASAP7_75t_SL g3649 ( 
.A(n_3277),
.B(n_2999),
.C(n_916),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3306),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3307),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3323),
.Y(n_3652)
);

AND3x1_ASAP7_75t_L g3653 ( 
.A(n_3296),
.B(n_1188),
.C(n_1016),
.Y(n_3653)
);

NAND2xp5_ASAP7_75t_SL g3654 ( 
.A(n_3508),
.B(n_2816),
.Y(n_3654)
);

AND2x4_ASAP7_75t_L g3655 ( 
.A(n_3288),
.B(n_2852),
.Y(n_3655)
);

BUFx4f_ASAP7_75t_L g3656 ( 
.A(n_3299),
.Y(n_3656)
);

CKINVDCx5p33_ASAP7_75t_R g3657 ( 
.A(n_3257),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3201),
.B(n_3079),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3324),
.Y(n_3659)
);

AOI22xp5_ASAP7_75t_L g3660 ( 
.A1(n_3489),
.A2(n_2791),
.B1(n_2852),
.B2(n_2952),
.Y(n_3660)
);

INVx2_ASAP7_75t_SL g3661 ( 
.A(n_3299),
.Y(n_3661)
);

INVx1_ASAP7_75t_L g3662 ( 
.A(n_3331),
.Y(n_3662)
);

BUFx3_ASAP7_75t_L g3663 ( 
.A(n_3263),
.Y(n_3663)
);

AND2x2_ASAP7_75t_L g3664 ( 
.A(n_3213),
.B(n_1518),
.Y(n_3664)
);

NAND2xp5_ASAP7_75t_L g3665 ( 
.A(n_3212),
.B(n_3216),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3348),
.Y(n_3666)
);

NAND2xp5_ASAP7_75t_L g3667 ( 
.A(n_3521),
.B(n_2784),
.Y(n_3667)
);

INVx1_ASAP7_75t_L g3668 ( 
.A(n_3350),
.Y(n_3668)
);

INVx2_ASAP7_75t_L g3669 ( 
.A(n_3305),
.Y(n_3669)
);

BUFx2_ASAP7_75t_L g3670 ( 
.A(n_3357),
.Y(n_3670)
);

OAI22xp5_ASAP7_75t_L g3671 ( 
.A1(n_3560),
.A2(n_3142),
.B1(n_3165),
.B2(n_3141),
.Y(n_3671)
);

NAND2xp5_ASAP7_75t_L g3672 ( 
.A(n_3548),
.B(n_3197),
.Y(n_3672)
);

INVx1_ASAP7_75t_L g3673 ( 
.A(n_3354),
.Y(n_3673)
);

AND2x4_ASAP7_75t_L g3674 ( 
.A(n_3564),
.B(n_3388),
.Y(n_3674)
);

INVx1_ASAP7_75t_L g3675 ( 
.A(n_3376),
.Y(n_3675)
);

BUFx6f_ASAP7_75t_L g3676 ( 
.A(n_3266),
.Y(n_3676)
);

OAI22xp5_ASAP7_75t_L g3677 ( 
.A1(n_3573),
.A2(n_3142),
.B1(n_3165),
.B2(n_3141),
.Y(n_3677)
);

INVx1_ASAP7_75t_L g3678 ( 
.A(n_3389),
.Y(n_3678)
);

NAND2xp5_ASAP7_75t_SL g3679 ( 
.A(n_3508),
.B(n_3097),
.Y(n_3679)
);

INVx1_ASAP7_75t_L g3680 ( 
.A(n_3395),
.Y(n_3680)
);

AND2x4_ASAP7_75t_L g3681 ( 
.A(n_3564),
.B(n_3460),
.Y(n_3681)
);

AOI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3359),
.A2(n_2952),
.B1(n_2869),
.B2(n_2835),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3398),
.Y(n_3683)
);

NOR3xp33_ASAP7_75t_SL g3684 ( 
.A(n_3378),
.B(n_2829),
.C(n_919),
.Y(n_3684)
);

NAND2xp5_ASAP7_75t_L g3685 ( 
.A(n_3530),
.B(n_2787),
.Y(n_3685)
);

AND2x2_ASAP7_75t_L g3686 ( 
.A(n_3286),
.B(n_1519),
.Y(n_3686)
);

O2A1O1Ixp33_ASAP7_75t_L g3687 ( 
.A1(n_3503),
.A2(n_3174),
.B(n_3171),
.C(n_3158),
.Y(n_3687)
);

BUFx3_ASAP7_75t_L g3688 ( 
.A(n_3279),
.Y(n_3688)
);

INVx2_ASAP7_75t_L g3689 ( 
.A(n_3319),
.Y(n_3689)
);

INVx3_ASAP7_75t_L g3690 ( 
.A(n_3266),
.Y(n_3690)
);

NAND2xp5_ASAP7_75t_SL g3691 ( 
.A(n_3207),
.B(n_2816),
.Y(n_3691)
);

NAND2xp5_ASAP7_75t_L g3692 ( 
.A(n_3510),
.B(n_2831),
.Y(n_3692)
);

BUFx3_ASAP7_75t_L g3693 ( 
.A(n_3281),
.Y(n_3693)
);

INVx2_ASAP7_75t_L g3694 ( 
.A(n_3328),
.Y(n_3694)
);

INVx4_ASAP7_75t_L g3695 ( 
.A(n_3299),
.Y(n_3695)
);

NAND2xp5_ASAP7_75t_L g3696 ( 
.A(n_3286),
.B(n_3491),
.Y(n_3696)
);

INVx1_ASAP7_75t_L g3697 ( 
.A(n_3407),
.Y(n_3697)
);

AND2x2_ASAP7_75t_L g3698 ( 
.A(n_3490),
.B(n_1521),
.Y(n_3698)
);

INVx1_ASAP7_75t_L g3699 ( 
.A(n_3413),
.Y(n_3699)
);

CKINVDCx5p33_ASAP7_75t_R g3700 ( 
.A(n_3540),
.Y(n_3700)
);

INVx1_ASAP7_75t_L g3701 ( 
.A(n_3418),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3419),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3421),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3491),
.B(n_2869),
.Y(n_3704)
);

OR2x2_ASAP7_75t_L g3705 ( 
.A(n_3242),
.B(n_3171),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3424),
.Y(n_3706)
);

INVx5_ASAP7_75t_L g3707 ( 
.A(n_3460),
.Y(n_3707)
);

AND2x4_ASAP7_75t_L g3708 ( 
.A(n_3460),
.B(n_2981),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3352),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3428),
.Y(n_3710)
);

AOI22xp33_ASAP7_75t_SL g3711 ( 
.A1(n_3370),
.A2(n_2940),
.B1(n_2833),
.B2(n_2977),
.Y(n_3711)
);

NAND2xp5_ASAP7_75t_SL g3712 ( 
.A(n_3207),
.B(n_3130),
.Y(n_3712)
);

NOR2xp33_ASAP7_75t_L g3713 ( 
.A(n_3274),
.B(n_3174),
.Y(n_3713)
);

AND2x2_ASAP7_75t_L g3714 ( 
.A(n_3267),
.B(n_3567),
.Y(n_3714)
);

AOI21xp33_ASAP7_75t_L g3715 ( 
.A1(n_3329),
.A2(n_2940),
.B(n_2833),
.Y(n_3715)
);

BUFx4f_ASAP7_75t_SL g3716 ( 
.A(n_3382),
.Y(n_3716)
);

NAND2xp5_ASAP7_75t_SL g3717 ( 
.A(n_3247),
.B(n_2892),
.Y(n_3717)
);

NAND2xp5_ASAP7_75t_L g3718 ( 
.A(n_3267),
.B(n_2869),
.Y(n_3718)
);

INVx1_ASAP7_75t_L g3719 ( 
.A(n_3435),
.Y(n_3719)
);

OAI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3339),
.A2(n_2879),
.B1(n_2880),
.B2(n_2875),
.Y(n_3720)
);

NAND2xp5_ASAP7_75t_L g3721 ( 
.A(n_3227),
.B(n_3463),
.Y(n_3721)
);

NAND2xp5_ASAP7_75t_SL g3722 ( 
.A(n_3406),
.B(n_2892),
.Y(n_3722)
);

INVx3_ASAP7_75t_L g3723 ( 
.A(n_3270),
.Y(n_3723)
);

NAND2x1p5_ASAP7_75t_L g3724 ( 
.A(n_3527),
.B(n_2892),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3443),
.Y(n_3725)
);

BUFx6f_ASAP7_75t_L g3726 ( 
.A(n_3270),
.Y(n_3726)
);

NAND2x1p5_ASAP7_75t_L g3727 ( 
.A(n_3232),
.B(n_2892),
.Y(n_3727)
);

INVx3_ASAP7_75t_L g3728 ( 
.A(n_3270),
.Y(n_3728)
);

INVx1_ASAP7_75t_L g3729 ( 
.A(n_3446),
.Y(n_3729)
);

NAND2xp5_ASAP7_75t_L g3730 ( 
.A(n_3227),
.B(n_2869),
.Y(n_3730)
);

INVx2_ASAP7_75t_SL g3731 ( 
.A(n_3214),
.Y(n_3731)
);

BUFx3_ASAP7_75t_L g3732 ( 
.A(n_3321),
.Y(n_3732)
);

NAND2xp5_ASAP7_75t_SL g3733 ( 
.A(n_3237),
.B(n_3058),
.Y(n_3733)
);

AND2x4_ASAP7_75t_L g3734 ( 
.A(n_3511),
.B(n_2981),
.Y(n_3734)
);

INVx3_ASAP7_75t_L g3735 ( 
.A(n_3311),
.Y(n_3735)
);

NAND2xp5_ASAP7_75t_L g3736 ( 
.A(n_3463),
.B(n_2875),
.Y(n_3736)
);

AND2x2_ASAP7_75t_L g3737 ( 
.A(n_3271),
.B(n_1522),
.Y(n_3737)
);

NAND2xp5_ASAP7_75t_SL g3738 ( 
.A(n_3238),
.B(n_3058),
.Y(n_3738)
);

OR2x2_ASAP7_75t_L g3739 ( 
.A(n_3322),
.B(n_2879),
.Y(n_3739)
);

NAND2xp5_ASAP7_75t_SL g3740 ( 
.A(n_3271),
.B(n_3058),
.Y(n_3740)
);

NAND2xp5_ASAP7_75t_L g3741 ( 
.A(n_3253),
.B(n_2880),
.Y(n_3741)
);

INVx1_ASAP7_75t_L g3742 ( 
.A(n_3455),
.Y(n_3742)
);

INVx2_ASAP7_75t_L g3743 ( 
.A(n_3355),
.Y(n_3743)
);

NAND2xp33_ASAP7_75t_L g3744 ( 
.A(n_3385),
.B(n_3088),
.Y(n_3744)
);

AND2x4_ASAP7_75t_L g3745 ( 
.A(n_3261),
.B(n_2981),
.Y(n_3745)
);

AND2x4_ASAP7_75t_L g3746 ( 
.A(n_3535),
.B(n_3182),
.Y(n_3746)
);

NAND2xp5_ASAP7_75t_SL g3747 ( 
.A(n_3342),
.B(n_3130),
.Y(n_3747)
);

INVx4_ASAP7_75t_L g3748 ( 
.A(n_3232),
.Y(n_3748)
);

INVx1_ASAP7_75t_L g3749 ( 
.A(n_3459),
.Y(n_3749)
);

NAND2xp5_ASAP7_75t_L g3750 ( 
.A(n_3268),
.B(n_3110),
.Y(n_3750)
);

INVx2_ASAP7_75t_SL g3751 ( 
.A(n_3364),
.Y(n_3751)
);

NAND2xp5_ASAP7_75t_L g3752 ( 
.A(n_3335),
.B(n_3110),
.Y(n_3752)
);

INVx2_ASAP7_75t_L g3753 ( 
.A(n_3356),
.Y(n_3753)
);

AOI22xp5_ASAP7_75t_L g3754 ( 
.A1(n_3336),
.A2(n_2977),
.B1(n_3108),
.B2(n_2908),
.Y(n_3754)
);

INVx2_ASAP7_75t_L g3755 ( 
.A(n_3374),
.Y(n_3755)
);

BUFx2_ASAP7_75t_L g3756 ( 
.A(n_3282),
.Y(n_3756)
);

AND2x4_ASAP7_75t_L g3757 ( 
.A(n_3218),
.B(n_3182),
.Y(n_3757)
);

NAND2xp5_ASAP7_75t_L g3758 ( 
.A(n_3335),
.B(n_3338),
.Y(n_3758)
);

NAND2xp5_ASAP7_75t_L g3759 ( 
.A(n_3338),
.B(n_3114),
.Y(n_3759)
);

NOR2xp33_ASAP7_75t_R g3760 ( 
.A(n_3540),
.B(n_3116),
.Y(n_3760)
);

BUFx6f_ASAP7_75t_L g3761 ( 
.A(n_3311),
.Y(n_3761)
);

INVx1_ASAP7_75t_L g3762 ( 
.A(n_3465),
.Y(n_3762)
);

INVx1_ASAP7_75t_L g3763 ( 
.A(n_3468),
.Y(n_3763)
);

NAND2xp5_ASAP7_75t_SL g3764 ( 
.A(n_3342),
.B(n_3547),
.Y(n_3764)
);

NOR2xp33_ASAP7_75t_L g3765 ( 
.A(n_3358),
.B(n_2958),
.Y(n_3765)
);

BUFx3_ASAP7_75t_L g3766 ( 
.A(n_3365),
.Y(n_3766)
);

OR2x2_ASAP7_75t_L g3767 ( 
.A(n_3556),
.B(n_3153),
.Y(n_3767)
);

NAND2xp5_ASAP7_75t_SL g3768 ( 
.A(n_3547),
.B(n_3058),
.Y(n_3768)
);

NAND2xp5_ASAP7_75t_L g3769 ( 
.A(n_3478),
.B(n_2977),
.Y(n_3769)
);

NAND2xp5_ASAP7_75t_L g3770 ( 
.A(n_3565),
.B(n_2977),
.Y(n_3770)
);

INVx1_ASAP7_75t_L g3771 ( 
.A(n_3475),
.Y(n_3771)
);

BUFx12f_ASAP7_75t_L g3772 ( 
.A(n_3555),
.Y(n_3772)
);

AND2x6_ASAP7_75t_L g3773 ( 
.A(n_3538),
.B(n_3075),
.Y(n_3773)
);

INVx1_ASAP7_75t_L g3774 ( 
.A(n_3481),
.Y(n_3774)
);

AOI22xp33_ASAP7_75t_L g3775 ( 
.A1(n_3519),
.A2(n_2940),
.B1(n_2908),
.B2(n_2924),
.Y(n_3775)
);

NAND2xp5_ASAP7_75t_L g3776 ( 
.A(n_3568),
.B(n_3158),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3484),
.Y(n_3777)
);

INVx2_ASAP7_75t_L g3778 ( 
.A(n_3375),
.Y(n_3778)
);

NOR2x1p5_ASAP7_75t_L g3779 ( 
.A(n_3558),
.B(n_2903),
.Y(n_3779)
);

AND2x4_ASAP7_75t_L g3780 ( 
.A(n_3559),
.B(n_3182),
.Y(n_3780)
);

AND2x4_ASAP7_75t_L g3781 ( 
.A(n_3559),
.B(n_3090),
.Y(n_3781)
);

NOR2xp33_ASAP7_75t_L g3782 ( 
.A(n_3211),
.B(n_2958),
.Y(n_3782)
);

INVx1_ASAP7_75t_L g3783 ( 
.A(n_3504),
.Y(n_3783)
);

INVx3_ASAP7_75t_L g3784 ( 
.A(n_3311),
.Y(n_3784)
);

INVx1_ASAP7_75t_L g3785 ( 
.A(n_3507),
.Y(n_3785)
);

INVx2_ASAP7_75t_L g3786 ( 
.A(n_3379),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3381),
.Y(n_3787)
);

NOR2x1p5_ASAP7_75t_L g3788 ( 
.A(n_3225),
.B(n_2903),
.Y(n_3788)
);

BUFx2_ASAP7_75t_L g3789 ( 
.A(n_3318),
.Y(n_3789)
);

BUFx6f_ASAP7_75t_L g3790 ( 
.A(n_3318),
.Y(n_3790)
);

AND2x2_ASAP7_75t_L g3791 ( 
.A(n_3498),
.B(n_1523),
.Y(n_3791)
);

NAND2xp5_ASAP7_75t_L g3792 ( 
.A(n_3569),
.B(n_3181),
.Y(n_3792)
);

INVx2_ASAP7_75t_L g3793 ( 
.A(n_3392),
.Y(n_3793)
);

NAND2xp5_ASAP7_75t_SL g3794 ( 
.A(n_3316),
.B(n_3097),
.Y(n_3794)
);

OAI21xp5_ASAP7_75t_L g3795 ( 
.A1(n_3402),
.A2(n_3185),
.B(n_3181),
.Y(n_3795)
);

HB1xp67_ASAP7_75t_L g3796 ( 
.A(n_3497),
.Y(n_3796)
);

NAND2xp5_ASAP7_75t_L g3797 ( 
.A(n_3570),
.B(n_3088),
.Y(n_3797)
);

NOR2xp33_ASAP7_75t_SL g3798 ( 
.A(n_3385),
.B(n_3136),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3433),
.Y(n_3799)
);

AOI22xp5_ASAP7_75t_L g3800 ( 
.A1(n_3456),
.A2(n_3108),
.B1(n_2924),
.B2(n_3104),
.Y(n_3800)
);

INVx2_ASAP7_75t_SL g3801 ( 
.A(n_3412),
.Y(n_3801)
);

NAND2xp5_ASAP7_75t_L g3802 ( 
.A(n_3537),
.B(n_3088),
.Y(n_3802)
);

INVxp67_ASAP7_75t_L g3803 ( 
.A(n_3415),
.Y(n_3803)
);

NAND2xp5_ASAP7_75t_L g3804 ( 
.A(n_3537),
.B(n_3088),
.Y(n_3804)
);

AND2x4_ASAP7_75t_L g3805 ( 
.A(n_3362),
.B(n_3090),
.Y(n_3805)
);

AND2x2_ASAP7_75t_SL g3806 ( 
.A(n_3519),
.B(n_3534),
.Y(n_3806)
);

NAND2xp5_ASAP7_75t_SL g3807 ( 
.A(n_3250),
.B(n_3097),
.Y(n_3807)
);

NAND2xp5_ASAP7_75t_L g3808 ( 
.A(n_3415),
.B(n_3104),
.Y(n_3808)
);

INVx3_ASAP7_75t_L g3809 ( 
.A(n_3318),
.Y(n_3809)
);

NAND2xp5_ASAP7_75t_L g3810 ( 
.A(n_3416),
.B(n_3104),
.Y(n_3810)
);

NAND2xp5_ASAP7_75t_L g3811 ( 
.A(n_3416),
.B(n_3497),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3551),
.Y(n_3812)
);

AOI22xp33_ASAP7_75t_L g3813 ( 
.A1(n_3534),
.A2(n_3114),
.B1(n_3186),
.B2(n_3103),
.Y(n_3813)
);

NAND2x1p5_ASAP7_75t_L g3814 ( 
.A(n_3262),
.B(n_3097),
.Y(n_3814)
);

INVx2_ASAP7_75t_L g3815 ( 
.A(n_3414),
.Y(n_3815)
);

NAND2xp5_ASAP7_75t_L g3816 ( 
.A(n_3269),
.B(n_3104),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3553),
.Y(n_3817)
);

BUFx6f_ASAP7_75t_L g3818 ( 
.A(n_3320),
.Y(n_3818)
);

NAND2xp5_ASAP7_75t_L g3819 ( 
.A(n_3326),
.B(n_3155),
.Y(n_3819)
);

NAND2xp5_ASAP7_75t_L g3820 ( 
.A(n_3276),
.B(n_3161),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3426),
.Y(n_3821)
);

INVx2_ASAP7_75t_SL g3822 ( 
.A(n_3373),
.Y(n_3822)
);

AOI22xp5_ASAP7_75t_L g3823 ( 
.A1(n_3380),
.A2(n_3187),
.B1(n_3186),
.B2(n_3179),
.Y(n_3823)
);

INVx3_ASAP7_75t_L g3824 ( 
.A(n_3320),
.Y(n_3824)
);

BUFx3_ASAP7_75t_L g3825 ( 
.A(n_3320),
.Y(n_3825)
);

INVxp67_ASAP7_75t_L g3826 ( 
.A(n_3458),
.Y(n_3826)
);

AOI22xp33_ASAP7_75t_L g3827 ( 
.A1(n_3550),
.A2(n_3186),
.B1(n_3113),
.B2(n_3118),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3554),
.Y(n_3828)
);

BUFx3_ASAP7_75t_L g3829 ( 
.A(n_3360),
.Y(n_3829)
);

INVx5_ASAP7_75t_L g3830 ( 
.A(n_3262),
.Y(n_3830)
);

AND2x2_ASAP7_75t_L g3831 ( 
.A(n_3265),
.B(n_1525),
.Y(n_3831)
);

INVx3_ASAP7_75t_SL g3832 ( 
.A(n_3437),
.Y(n_3832)
);

NOR2xp33_ASAP7_75t_L g3833 ( 
.A(n_3230),
.B(n_3187),
.Y(n_3833)
);

NAND2xp5_ASAP7_75t_SL g3834 ( 
.A(n_3506),
.B(n_3130),
.Y(n_3834)
);

OR2x6_ASAP7_75t_L g3835 ( 
.A(n_3545),
.B(n_3160),
.Y(n_3835)
);

BUFx12f_ASAP7_75t_L g3836 ( 
.A(n_3523),
.Y(n_3836)
);

NAND2xp5_ASAP7_75t_SL g3837 ( 
.A(n_3506),
.B(n_3130),
.Y(n_3837)
);

NAND2xp5_ASAP7_75t_L g3838 ( 
.A(n_3368),
.B(n_3166),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3529),
.Y(n_3839)
);

CKINVDCx5p33_ASAP7_75t_R g3840 ( 
.A(n_3458),
.Y(n_3840)
);

AOI21xp5_ASAP7_75t_L g3841 ( 
.A1(n_3289),
.A2(n_3184),
.B(n_3086),
.Y(n_3841)
);

NAND2xp5_ASAP7_75t_SL g3842 ( 
.A(n_3552),
.B(n_3122),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3531),
.Y(n_3843)
);

AO22x1_ASAP7_75t_L g3844 ( 
.A1(n_3246),
.A2(n_3186),
.B1(n_3105),
.B2(n_922),
.Y(n_3844)
);

AOI22xp5_ASAP7_75t_L g3845 ( 
.A1(n_3380),
.A2(n_928),
.B1(n_987),
.B2(n_958),
.Y(n_3845)
);

NAND2xp5_ASAP7_75t_SL g3846 ( 
.A(n_3239),
.B(n_3122),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3544),
.Y(n_3847)
);

NAND2xp5_ASAP7_75t_L g3848 ( 
.A(n_3371),
.B(n_3057),
.Y(n_3848)
);

AND2x2_ASAP7_75t_L g3849 ( 
.A(n_3252),
.B(n_1536),
.Y(n_3849)
);

INVx2_ASAP7_75t_SL g3850 ( 
.A(n_3450),
.Y(n_3850)
);

NAND2xp5_ASAP7_75t_L g3851 ( 
.A(n_3325),
.B(n_3125),
.Y(n_3851)
);

AND2x4_ASAP7_75t_L g3852 ( 
.A(n_3522),
.B(n_3132),
.Y(n_3852)
);

NAND2xp5_ASAP7_75t_SL g3853 ( 
.A(n_3278),
.B(n_3122),
.Y(n_3853)
);

OAI21xp33_ASAP7_75t_SL g3854 ( 
.A1(n_3532),
.A2(n_3184),
.B(n_3185),
.Y(n_3854)
);

CKINVDCx5p33_ASAP7_75t_R g3855 ( 
.A(n_3563),
.Y(n_3855)
);

NAND2xp5_ASAP7_75t_L g3856 ( 
.A(n_3244),
.B(n_3127),
.Y(n_3856)
);

NAND2xp5_ASAP7_75t_L g3857 ( 
.A(n_3377),
.B(n_3135),
.Y(n_3857)
);

NAND2xp33_ASAP7_75t_SL g3858 ( 
.A(n_3275),
.B(n_3123),
.Y(n_3858)
);

AOI22xp33_ASAP7_75t_L g3859 ( 
.A1(n_3550),
.A2(n_3137),
.B1(n_3159),
.B2(n_3147),
.Y(n_3859)
);

NAND2xp5_ASAP7_75t_L g3860 ( 
.A(n_3383),
.B(n_3175),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3332),
.B(n_3190),
.Y(n_3861)
);

INVx4_ASAP7_75t_L g3862 ( 
.A(n_3275),
.Y(n_3862)
);

NAND2xp5_ASAP7_75t_L g3863 ( 
.A(n_3302),
.B(n_3196),
.Y(n_3863)
);

BUFx3_ASAP7_75t_L g3864 ( 
.A(n_3363),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3361),
.Y(n_3865)
);

NOR2xp33_ASAP7_75t_L g3866 ( 
.A(n_3224),
.B(n_2968),
.Y(n_3866)
);

NAND2xp5_ASAP7_75t_L g3867 ( 
.A(n_3280),
.B(n_2968),
.Y(n_3867)
);

INVx3_ASAP7_75t_L g3868 ( 
.A(n_3404),
.Y(n_3868)
);

AND2x2_ASAP7_75t_L g3869 ( 
.A(n_3252),
.B(n_3292),
.Y(n_3869)
);

AND2x6_ASAP7_75t_L g3870 ( 
.A(n_3310),
.B(n_3162),
.Y(n_3870)
);

AOI22xp33_ASAP7_75t_L g3871 ( 
.A1(n_3386),
.A2(n_3160),
.B1(n_3146),
.B2(n_3136),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3430),
.Y(n_3872)
);

AOI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3386),
.A2(n_3423),
.B1(n_3292),
.B2(n_3198),
.Y(n_3873)
);

AOI22xp33_ASAP7_75t_L g3874 ( 
.A1(n_3423),
.A2(n_3146),
.B1(n_1017),
.B2(n_1019),
.Y(n_3874)
);

NAND2xp5_ASAP7_75t_L g3875 ( 
.A(n_3283),
.B(n_2872),
.Y(n_3875)
);

INVx2_ASAP7_75t_L g3876 ( 
.A(n_3436),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3441),
.Y(n_3877)
);

NAND2xp5_ASAP7_75t_SL g3878 ( 
.A(n_3600),
.B(n_3403),
.Y(n_3878)
);

NAND2xp5_ASAP7_75t_L g3879 ( 
.A(n_3600),
.B(n_3285),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3665),
.B(n_3205),
.Y(n_3880)
);

OR2x2_ASAP7_75t_L g3881 ( 
.A(n_3696),
.B(n_3617),
.Y(n_3881)
);

NAND2xp5_ASAP7_75t_SL g3882 ( 
.A(n_3758),
.B(n_3222),
.Y(n_3882)
);

NAND2xp5_ASAP7_75t_SL g3883 ( 
.A(n_3758),
.B(n_3223),
.Y(n_3883)
);

NAND2xp5_ASAP7_75t_SL g3884 ( 
.A(n_3601),
.B(n_3385),
.Y(n_3884)
);

NAND2xp5_ASAP7_75t_SL g3885 ( 
.A(n_3840),
.B(n_3427),
.Y(n_3885)
);

NAND2xp5_ASAP7_75t_SL g3886 ( 
.A(n_3721),
.B(n_3429),
.Y(n_3886)
);

AND2x2_ASAP7_75t_L g3887 ( 
.A(n_3633),
.B(n_3246),
.Y(n_3887)
);

NAND2xp5_ASAP7_75t_SL g3888 ( 
.A(n_3811),
.B(n_3333),
.Y(n_3888)
);

NAND2xp5_ASAP7_75t_SL g3889 ( 
.A(n_3776),
.B(n_3340),
.Y(n_3889)
);

NAND2xp5_ASAP7_75t_SL g3890 ( 
.A(n_3792),
.B(n_3343),
.Y(n_3890)
);

NAND2xp5_ASAP7_75t_SL g3891 ( 
.A(n_3601),
.B(n_3344),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_SL g3892 ( 
.A(n_3720),
.B(n_3487),
.Y(n_3892)
);

NAND2xp5_ASAP7_75t_SL g3893 ( 
.A(n_3803),
.B(n_3408),
.Y(n_3893)
);

NAND2xp5_ASAP7_75t_SL g3894 ( 
.A(n_3682),
.B(n_3410),
.Y(n_3894)
);

NAND2xp33_ASAP7_75t_SL g3895 ( 
.A(n_3748),
.B(n_3404),
.Y(n_3895)
);

NAND2xp5_ASAP7_75t_SL g3896 ( 
.A(n_3682),
.B(n_3385),
.Y(n_3896)
);

NAND2xp5_ASAP7_75t_SL g3897 ( 
.A(n_3603),
.B(n_3385),
.Y(n_3897)
);

NAND2xp5_ASAP7_75t_SL g3898 ( 
.A(n_3603),
.B(n_3385),
.Y(n_3898)
);

NAND2xp5_ASAP7_75t_SL g3899 ( 
.A(n_3598),
.B(n_3351),
.Y(n_3899)
);

NAND2xp33_ASAP7_75t_SL g3900 ( 
.A(n_3748),
.B(n_3613),
.Y(n_3900)
);

NAND2xp5_ASAP7_75t_L g3901 ( 
.A(n_3658),
.B(n_3514),
.Y(n_3901)
);

NAND2xp5_ASAP7_75t_SL g3902 ( 
.A(n_3598),
.B(n_3353),
.Y(n_3902)
);

NAND2xp5_ASAP7_75t_SL g3903 ( 
.A(n_3752),
.B(n_3390),
.Y(n_3903)
);

NAND2xp5_ASAP7_75t_SL g3904 ( 
.A(n_3752),
.B(n_3516),
.Y(n_3904)
);

NAND2xp5_ASAP7_75t_SL g3905 ( 
.A(n_3759),
.B(n_3539),
.Y(n_3905)
);

NAND2xp5_ASAP7_75t_L g3906 ( 
.A(n_3672),
.B(n_3514),
.Y(n_3906)
);

NAND2xp33_ASAP7_75t_SL g3907 ( 
.A(n_3576),
.B(n_3387),
.Y(n_3907)
);

NAND2xp33_ASAP7_75t_SL g3908 ( 
.A(n_3862),
.B(n_3525),
.Y(n_3908)
);

NAND2xp33_ASAP7_75t_SL g3909 ( 
.A(n_3862),
.B(n_3405),
.Y(n_3909)
);

NAND2xp5_ASAP7_75t_SL g3910 ( 
.A(n_3759),
.B(n_3615),
.Y(n_3910)
);

NAND2xp5_ASAP7_75t_SL g3911 ( 
.A(n_3660),
.B(n_3400),
.Y(n_3911)
);

NAND2xp5_ASAP7_75t_SL g3912 ( 
.A(n_3660),
.B(n_3409),
.Y(n_3912)
);

NAND2xp5_ASAP7_75t_SL g3913 ( 
.A(n_3855),
.B(n_3217),
.Y(n_3913)
);

NAND2xp33_ASAP7_75t_SL g3914 ( 
.A(n_3760),
.B(n_3405),
.Y(n_3914)
);

NAND2xp5_ASAP7_75t_SL g3915 ( 
.A(n_3797),
.B(n_3653),
.Y(n_3915)
);

NAND2xp5_ASAP7_75t_SL g3916 ( 
.A(n_3653),
.B(n_3217),
.Y(n_3916)
);

NAND2xp5_ASAP7_75t_L g3917 ( 
.A(n_3643),
.B(n_3396),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3646),
.B(n_3397),
.Y(n_3918)
);

NAND2xp5_ASAP7_75t_SL g3919 ( 
.A(n_3692),
.B(n_3220),
.Y(n_3919)
);

NAND2xp5_ASAP7_75t_SL g3920 ( 
.A(n_3736),
.B(n_3220),
.Y(n_3920)
);

NAND2xp5_ASAP7_75t_L g3921 ( 
.A(n_3796),
.B(n_3295),
.Y(n_3921)
);

NAND2xp5_ASAP7_75t_SL g3922 ( 
.A(n_3770),
.B(n_3543),
.Y(n_3922)
);

NAND2xp5_ASAP7_75t_SL g3923 ( 
.A(n_3808),
.B(n_3401),
.Y(n_3923)
);

NAND2xp5_ASAP7_75t_SL g3924 ( 
.A(n_3810),
.B(n_3467),
.Y(n_3924)
);

NAND2xp5_ASAP7_75t_SL g3925 ( 
.A(n_3832),
.B(n_3467),
.Y(n_3925)
);

NAND2xp5_ASAP7_75t_SL g3926 ( 
.A(n_3833),
.B(n_3221),
.Y(n_3926)
);

NAND2xp5_ASAP7_75t_SL g3927 ( 
.A(n_3822),
.B(n_3541),
.Y(n_3927)
);

NAND2xp33_ASAP7_75t_SL g3928 ( 
.A(n_3674),
.B(n_3411),
.Y(n_3928)
);

NAND2xp33_ASAP7_75t_SL g3929 ( 
.A(n_3674),
.B(n_3411),
.Y(n_3929)
);

NAND2xp33_ASAP7_75t_SL g3930 ( 
.A(n_3684),
.B(n_3492),
.Y(n_3930)
);

NAND2xp5_ASAP7_75t_SL g3931 ( 
.A(n_3769),
.B(n_3447),
.Y(n_3931)
);

NAND2xp5_ASAP7_75t_SL g3932 ( 
.A(n_3605),
.B(n_3447),
.Y(n_3932)
);

NAND2xp5_ASAP7_75t_SL g3933 ( 
.A(n_3605),
.B(n_3802),
.Y(n_3933)
);

NAND2xp5_ASAP7_75t_SL g3934 ( 
.A(n_3605),
.B(n_3451),
.Y(n_3934)
);

NAND2xp33_ASAP7_75t_SL g3935 ( 
.A(n_3594),
.B(n_3492),
.Y(n_3935)
);

NAND2xp5_ASAP7_75t_SL g3936 ( 
.A(n_3804),
.B(n_3451),
.Y(n_3936)
);

AND2x2_ASAP7_75t_L g3937 ( 
.A(n_3714),
.B(n_3566),
.Y(n_3937)
);

NAND2xp5_ASAP7_75t_L g3938 ( 
.A(n_3799),
.B(n_3297),
.Y(n_3938)
);

NAND2xp5_ASAP7_75t_SL g3939 ( 
.A(n_3850),
.B(n_3730),
.Y(n_3939)
);

AND2x4_ASAP7_75t_L g3940 ( 
.A(n_3681),
.B(n_3528),
.Y(n_3940)
);

NAND2xp5_ASAP7_75t_SL g3941 ( 
.A(n_3765),
.B(n_3235),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_SL g3942 ( 
.A(n_3625),
.B(n_3826),
.Y(n_3942)
);

NAND2xp5_ASAP7_75t_SL g3943 ( 
.A(n_3625),
.B(n_3704),
.Y(n_3943)
);

NAND2xp33_ASAP7_75t_SL g3944 ( 
.A(n_3594),
.B(n_3546),
.Y(n_3944)
);

NAND2xp5_ASAP7_75t_SL g3945 ( 
.A(n_3602),
.B(n_3236),
.Y(n_3945)
);

NAND2xp33_ASAP7_75t_SL g3946 ( 
.A(n_3594),
.B(n_3546),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3865),
.B(n_3393),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_SL g3948 ( 
.A(n_3602),
.B(n_2779),
.Y(n_3948)
);

NAND2xp5_ASAP7_75t_SL g3949 ( 
.A(n_3671),
.B(n_2779),
.Y(n_3949)
);

NAND2xp5_ASAP7_75t_SL g3950 ( 
.A(n_3671),
.B(n_2793),
.Y(n_3950)
);

NAND2xp5_ASAP7_75t_SL g3951 ( 
.A(n_3677),
.B(n_2793),
.Y(n_3951)
);

NAND2xp33_ASAP7_75t_SL g3952 ( 
.A(n_3586),
.B(n_3219),
.Y(n_3952)
);

XOR2xp5_ASAP7_75t_L g3953 ( 
.A(n_3700),
.B(n_3574),
.Y(n_3953)
);

NAND2xp5_ASAP7_75t_L g3954 ( 
.A(n_3578),
.B(n_3571),
.Y(n_3954)
);

NAND2xp33_ASAP7_75t_SL g3955 ( 
.A(n_3575),
.B(n_3301),
.Y(n_3955)
);

NAND2xp5_ASAP7_75t_SL g3956 ( 
.A(n_3677),
.B(n_2793),
.Y(n_3956)
);

NAND2xp5_ASAP7_75t_SL g3957 ( 
.A(n_3764),
.B(n_2809),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_SL g3958 ( 
.A(n_3836),
.B(n_3639),
.Y(n_3958)
);

NAND2xp5_ASAP7_75t_SL g3959 ( 
.A(n_3575),
.B(n_2809),
.Y(n_3959)
);

NAND2xp5_ASAP7_75t_SL g3960 ( 
.A(n_3620),
.B(n_2809),
.Y(n_3960)
);

NAND2xp5_ASAP7_75t_L g3961 ( 
.A(n_3686),
.B(n_3420),
.Y(n_3961)
);

NAND2xp33_ASAP7_75t_SL g3962 ( 
.A(n_3868),
.B(n_3309),
.Y(n_3962)
);

NAND2xp33_ASAP7_75t_SL g3963 ( 
.A(n_3868),
.B(n_3488),
.Y(n_3963)
);

NAND2xp33_ASAP7_75t_SL g3964 ( 
.A(n_3718),
.B(n_3667),
.Y(n_3964)
);

NAND2xp5_ASAP7_75t_SL g3965 ( 
.A(n_3622),
.B(n_2834),
.Y(n_3965)
);

NAND2xp5_ASAP7_75t_SL g3966 ( 
.A(n_3622),
.B(n_2834),
.Y(n_3966)
);

NAND2xp5_ASAP7_75t_L g3967 ( 
.A(n_3606),
.B(n_3698),
.Y(n_3967)
);

NAND2xp5_ASAP7_75t_SL g3968 ( 
.A(n_3816),
.B(n_2834),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_SL g3969 ( 
.A(n_3580),
.B(n_3830),
.Y(n_3969)
);

NAND2xp5_ASAP7_75t_SL g3970 ( 
.A(n_3830),
.B(n_2836),
.Y(n_3970)
);

NAND2xp33_ASAP7_75t_SL g3971 ( 
.A(n_3695),
.B(n_3500),
.Y(n_3971)
);

NAND2xp5_ASAP7_75t_SL g3972 ( 
.A(n_3830),
.B(n_2836),
.Y(n_3972)
);

AND2x2_ASAP7_75t_L g3973 ( 
.A(n_3664),
.B(n_1014),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_SL g3974 ( 
.A(n_3705),
.B(n_2836),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_SL g3975 ( 
.A(n_3757),
.B(n_2856),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_SL g3976 ( 
.A(n_3757),
.B(n_2856),
.Y(n_3976)
);

NAND2xp5_ASAP7_75t_SL g3977 ( 
.A(n_3806),
.B(n_2856),
.Y(n_3977)
);

NAND2xp5_ASAP7_75t_SL g3978 ( 
.A(n_3781),
.B(n_2900),
.Y(n_3978)
);

NAND2xp5_ASAP7_75t_L g3979 ( 
.A(n_3611),
.B(n_3315),
.Y(n_3979)
);

NAND2xp5_ASAP7_75t_SL g3980 ( 
.A(n_3781),
.B(n_2900),
.Y(n_3980)
);

OR2x2_ASAP7_75t_L g3981 ( 
.A(n_3581),
.B(n_3345),
.Y(n_3981)
);

NAND2xp5_ASAP7_75t_SL g3982 ( 
.A(n_3579),
.B(n_2900),
.Y(n_3982)
);

NAND2xp5_ASAP7_75t_L g3983 ( 
.A(n_3670),
.B(n_3347),
.Y(n_3983)
);

NAND2xp5_ASAP7_75t_SL g3984 ( 
.A(n_3579),
.B(n_2922),
.Y(n_3984)
);

NAND2xp33_ASAP7_75t_SL g3985 ( 
.A(n_3695),
.B(n_3512),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3791),
.B(n_1019),
.Y(n_3986)
);

NAND2xp5_ASAP7_75t_SL g3987 ( 
.A(n_3579),
.B(n_2922),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3681),
.B(n_3542),
.Y(n_3988)
);

NAND2xp5_ASAP7_75t_SL g3989 ( 
.A(n_3599),
.B(n_2922),
.Y(n_3989)
);

NAND2xp33_ASAP7_75t_SL g3990 ( 
.A(n_3619),
.B(n_3515),
.Y(n_3990)
);

NAND2xp5_ASAP7_75t_SL g3991 ( 
.A(n_3599),
.B(n_2935),
.Y(n_3991)
);

NAND2xp5_ASAP7_75t_SL g3992 ( 
.A(n_3599),
.B(n_2935),
.Y(n_3992)
);

NAND2xp5_ASAP7_75t_SL g3993 ( 
.A(n_3676),
.B(n_2935),
.Y(n_3993)
);

NAND2xp5_ASAP7_75t_SL g3994 ( 
.A(n_3676),
.B(n_2939),
.Y(n_3994)
);

NAND2xp33_ASAP7_75t_SL g3995 ( 
.A(n_3657),
.B(n_3517),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_SL g3996 ( 
.A(n_3676),
.B(n_2939),
.Y(n_3996)
);

AND2x4_ASAP7_75t_L g3997 ( 
.A(n_3645),
.B(n_3313),
.Y(n_3997)
);

NAND2xp5_ASAP7_75t_SL g3998 ( 
.A(n_3726),
.B(n_2939),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_SL g3999 ( 
.A(n_3726),
.B(n_2996),
.Y(n_3999)
);

NAND2xp5_ASAP7_75t_SL g4000 ( 
.A(n_3726),
.B(n_2996),
.Y(n_4000)
);

NAND2xp5_ASAP7_75t_SL g4001 ( 
.A(n_3761),
.B(n_2996),
.Y(n_4001)
);

NAND2xp5_ASAP7_75t_SL g4002 ( 
.A(n_3761),
.B(n_3001),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3761),
.B(n_3001),
.Y(n_4003)
);

NAND2xp33_ASAP7_75t_SL g4004 ( 
.A(n_3801),
.B(n_3417),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_SL g4005 ( 
.A(n_3790),
.B(n_3001),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_SL g4006 ( 
.A(n_3790),
.B(n_3818),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_SL g4007 ( 
.A(n_3790),
.B(n_3006),
.Y(n_4007)
);

NAND2xp5_ASAP7_75t_SL g4008 ( 
.A(n_3818),
.B(n_3006),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_SL g4009 ( 
.A(n_3818),
.B(n_3006),
.Y(n_4009)
);

NAND2xp33_ASAP7_75t_SL g4010 ( 
.A(n_3645),
.B(n_3422),
.Y(n_4010)
);

NAND2xp5_ASAP7_75t_SL g4011 ( 
.A(n_3823),
.B(n_3717),
.Y(n_4011)
);

NAND2xp5_ASAP7_75t_L g4012 ( 
.A(n_3739),
.B(n_3349),
.Y(n_4012)
);

NAND2xp5_ASAP7_75t_SL g4013 ( 
.A(n_3823),
.B(n_3050),
.Y(n_4013)
);

NAND2xp5_ASAP7_75t_SL g4014 ( 
.A(n_3782),
.B(n_3795),
.Y(n_4014)
);

NAND2xp5_ASAP7_75t_SL g4015 ( 
.A(n_3795),
.B(n_3050),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_SL g4016 ( 
.A(n_3805),
.B(n_3050),
.Y(n_4016)
);

NAND2xp5_ASAP7_75t_SL g4017 ( 
.A(n_3805),
.B(n_3072),
.Y(n_4017)
);

NAND2xp5_ASAP7_75t_SL g4018 ( 
.A(n_3687),
.B(n_3072),
.Y(n_4018)
);

NAND2xp33_ASAP7_75t_L g4019 ( 
.A(n_3724),
.B(n_3123),
.Y(n_4019)
);

NAND2xp33_ASAP7_75t_SL g4020 ( 
.A(n_3655),
.B(n_3432),
.Y(n_4020)
);

NAND2xp33_ASAP7_75t_SL g4021 ( 
.A(n_3655),
.B(n_3138),
.Y(n_4021)
);

NAND2xp5_ASAP7_75t_SL g4022 ( 
.A(n_3597),
.B(n_3072),
.Y(n_4022)
);

NAND2xp5_ASAP7_75t_SL g4023 ( 
.A(n_3593),
.B(n_3123),
.Y(n_4023)
);

NAND2xp5_ASAP7_75t_SL g4024 ( 
.A(n_3616),
.B(n_3138),
.Y(n_4024)
);

NAND2xp5_ASAP7_75t_SL g4025 ( 
.A(n_3866),
.B(n_3138),
.Y(n_4025)
);

NAND2xp5_ASAP7_75t_SL g4026 ( 
.A(n_3852),
.B(n_3192),
.Y(n_4026)
);

NAND2xp5_ASAP7_75t_SL g4027 ( 
.A(n_3852),
.B(n_3192),
.Y(n_4027)
);

NAND2xp33_ASAP7_75t_SL g4028 ( 
.A(n_3608),
.B(n_3192),
.Y(n_4028)
);

NAND2xp5_ASAP7_75t_SL g4029 ( 
.A(n_3858),
.B(n_3425),
.Y(n_4029)
);

NAND2xp5_ASAP7_75t_SL g4030 ( 
.A(n_3800),
.B(n_3476),
.Y(n_4030)
);

NAND2xp5_ASAP7_75t_SL g4031 ( 
.A(n_3800),
.B(n_3439),
.Y(n_4031)
);

NAND2xp33_ASAP7_75t_SL g4032 ( 
.A(n_3648),
.B(n_3132),
.Y(n_4032)
);

NAND2xp33_ASAP7_75t_SL g4033 ( 
.A(n_3661),
.B(n_3154),
.Y(n_4033)
);

NAND2xp5_ASAP7_75t_L g4034 ( 
.A(n_3713),
.B(n_3434),
.Y(n_4034)
);

NAND2xp33_ASAP7_75t_SL g4035 ( 
.A(n_3609),
.B(n_3154),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_SL g4036 ( 
.A(n_3754),
.B(n_3439),
.Y(n_4036)
);

NAND2xp5_ASAP7_75t_SL g4037 ( 
.A(n_3754),
.B(n_3273),
.Y(n_4037)
);

AND2x4_ASAP7_75t_L g4038 ( 
.A(n_3708),
.B(n_3327),
.Y(n_4038)
);

NAND2xp5_ASAP7_75t_SL g4039 ( 
.A(n_3626),
.B(n_3337),
.Y(n_4039)
);

NAND2xp5_ASAP7_75t_SL g4040 ( 
.A(n_3747),
.B(n_3039),
.Y(n_4040)
);

NAND2xp5_ASAP7_75t_SL g4041 ( 
.A(n_3741),
.B(n_3039),
.Y(n_4041)
);

NAND2xp33_ASAP7_75t_SL g4042 ( 
.A(n_3691),
.B(n_3712),
.Y(n_4042)
);

NAND2xp5_ASAP7_75t_L g4043 ( 
.A(n_3737),
.B(n_3438),
.Y(n_4043)
);

NAND2xp5_ASAP7_75t_SL g4044 ( 
.A(n_3741),
.B(n_3063),
.Y(n_4044)
);

NAND2xp5_ASAP7_75t_SL g4045 ( 
.A(n_3768),
.B(n_3063),
.Y(n_4045)
);

NAND2xp33_ASAP7_75t_SL g4046 ( 
.A(n_3685),
.B(n_3164),
.Y(n_4046)
);

NAND2xp5_ASAP7_75t_SL g4047 ( 
.A(n_3829),
.B(n_3164),
.Y(n_4047)
);

NAND2xp33_ASAP7_75t_SL g4048 ( 
.A(n_3751),
.B(n_3177),
.Y(n_4048)
);

NAND2xp5_ASAP7_75t_SL g4049 ( 
.A(n_3864),
.B(n_3177),
.Y(n_4049)
);

NAND2xp5_ASAP7_75t_SL g4050 ( 
.A(n_3794),
.B(n_3189),
.Y(n_4050)
);

NAND2xp5_ASAP7_75t_L g4051 ( 
.A(n_3869),
.B(n_3444),
.Y(n_4051)
);

NAND2xp33_ASAP7_75t_SL g4052 ( 
.A(n_3635),
.B(n_3189),
.Y(n_4052)
);

NAND2xp5_ASAP7_75t_SL g4053 ( 
.A(n_3873),
.B(n_3470),
.Y(n_4053)
);

NAND2xp5_ASAP7_75t_SL g4054 ( 
.A(n_3610),
.B(n_3483),
.Y(n_4054)
);

NAND2xp33_ASAP7_75t_SL g4055 ( 
.A(n_3635),
.B(n_3075),
.Y(n_4055)
);

NAND2xp5_ASAP7_75t_SL g4056 ( 
.A(n_3690),
.B(n_2826),
.Y(n_4056)
);

NAND2xp5_ASAP7_75t_L g4057 ( 
.A(n_3731),
.B(n_3445),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_SL g4058 ( 
.A(n_3690),
.B(n_2826),
.Y(n_4058)
);

NAND2xp5_ASAP7_75t_SL g4059 ( 
.A(n_3723),
.B(n_2872),
.Y(n_4059)
);

AND2x4_ASAP7_75t_L g4060 ( 
.A(n_3708),
.B(n_2898),
.Y(n_4060)
);

NAND2xp5_ASAP7_75t_L g4061 ( 
.A(n_3750),
.B(n_3449),
.Y(n_4061)
);

NAND2xp5_ASAP7_75t_SL g4062 ( 
.A(n_3723),
.B(n_2898),
.Y(n_4062)
);

AND2x4_ASAP7_75t_L g4063 ( 
.A(n_3780),
.B(n_2913),
.Y(n_4063)
);

NAND2xp5_ASAP7_75t_SL g4064 ( 
.A(n_3728),
.B(n_2913),
.Y(n_4064)
);

NAND2xp5_ASAP7_75t_SL g4065 ( 
.A(n_3728),
.B(n_3735),
.Y(n_4065)
);

NAND2xp33_ASAP7_75t_SL g4066 ( 
.A(n_3596),
.B(n_3094),
.Y(n_4066)
);

NAND2xp33_ASAP7_75t_SL g4067 ( 
.A(n_3596),
.B(n_3094),
.Y(n_4067)
);

NAND2xp5_ASAP7_75t_SL g4068 ( 
.A(n_3735),
.B(n_3003),
.Y(n_4068)
);

NAND2xp5_ASAP7_75t_SL g4069 ( 
.A(n_3784),
.B(n_3003),
.Y(n_4069)
);

NAND2xp5_ASAP7_75t_L g4070 ( 
.A(n_3750),
.B(n_3454),
.Y(n_4070)
);

NAND2xp5_ASAP7_75t_SL g4071 ( 
.A(n_3784),
.B(n_3042),
.Y(n_4071)
);

NAND2xp5_ASAP7_75t_SL g4072 ( 
.A(n_3809),
.B(n_3042),
.Y(n_4072)
);

NAND2xp5_ASAP7_75t_SL g4073 ( 
.A(n_3809),
.B(n_3394),
.Y(n_4073)
);

NAND2xp5_ASAP7_75t_L g4074 ( 
.A(n_3638),
.B(n_3457),
.Y(n_4074)
);

NAND2xp5_ASAP7_75t_L g4075 ( 
.A(n_3849),
.B(n_3469),
.Y(n_4075)
);

NAND2xp5_ASAP7_75t_SL g4076 ( 
.A(n_3824),
.B(n_3384),
.Y(n_4076)
);

NAND2xp5_ASAP7_75t_SL g4077 ( 
.A(n_3824),
.B(n_3391),
.Y(n_4077)
);

NAND2xp5_ASAP7_75t_SL g4078 ( 
.A(n_3745),
.B(n_3096),
.Y(n_4078)
);

NAND2xp33_ASAP7_75t_SL g4079 ( 
.A(n_3596),
.B(n_3096),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_SL g4080 ( 
.A(n_3745),
.B(n_3101),
.Y(n_4080)
);

NAND2xp5_ASAP7_75t_SL g4081 ( 
.A(n_3656),
.B(n_3101),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_SL g4082 ( 
.A(n_3656),
.B(n_3621),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_SL g4083 ( 
.A(n_3707),
.B(n_3162),
.Y(n_4083)
);

NAND2xp5_ASAP7_75t_SL g4084 ( 
.A(n_3707),
.B(n_3854),
.Y(n_4084)
);

AND2x4_ASAP7_75t_L g4085 ( 
.A(n_3780),
.B(n_3172),
.Y(n_4085)
);

NAND2xp5_ASAP7_75t_L g4086 ( 
.A(n_3632),
.B(n_3577),
.Y(n_4086)
);

NAND2xp5_ASAP7_75t_SL g4087 ( 
.A(n_3707),
.B(n_3172),
.Y(n_4087)
);

NAND2xp5_ASAP7_75t_SL g4088 ( 
.A(n_3854),
.B(n_3480),
.Y(n_4088)
);

NAND2xp33_ASAP7_75t_SL g4089 ( 
.A(n_3627),
.B(n_3734),
.Y(n_4089)
);

NAND2xp5_ASAP7_75t_SL g4090 ( 
.A(n_3589),
.B(n_3480),
.Y(n_4090)
);

NAND2xp33_ASAP7_75t_SL g4091 ( 
.A(n_3734),
.B(n_3495),
.Y(n_4091)
);

NAND2xp5_ASAP7_75t_SL g4092 ( 
.A(n_3834),
.B(n_3471),
.Y(n_4092)
);

NAND2xp33_ASAP7_75t_SL g4093 ( 
.A(n_3654),
.B(n_3496),
.Y(n_4093)
);

NAND2xp5_ASAP7_75t_SL g4094 ( 
.A(n_3837),
.B(n_3472),
.Y(n_4094)
);

NAND2xp5_ASAP7_75t_L g4095 ( 
.A(n_3583),
.B(n_3473),
.Y(n_4095)
);

AND2x4_ASAP7_75t_L g4096 ( 
.A(n_3746),
.B(n_3448),
.Y(n_4096)
);

AND2x2_ASAP7_75t_L g4097 ( 
.A(n_3831),
.B(n_1021),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_SL g4098 ( 
.A(n_3789),
.B(n_3477),
.Y(n_4098)
);

NAND2xp5_ASAP7_75t_L g4099 ( 
.A(n_3584),
.B(n_3587),
.Y(n_4099)
);

AND2x2_ASAP7_75t_SL g4100 ( 
.A(n_3744),
.B(n_3482),
.Y(n_4100)
);

NAND2xp5_ASAP7_75t_SL g4101 ( 
.A(n_3807),
.B(n_3486),
.Y(n_4101)
);

NAND2xp5_ASAP7_75t_L g4102 ( 
.A(n_3588),
.B(n_3590),
.Y(n_4102)
);

NAND2xp5_ASAP7_75t_SL g4103 ( 
.A(n_3711),
.B(n_3466),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3604),
.B(n_3461),
.Y(n_4104)
);

NAND2xp5_ASAP7_75t_SL g4105 ( 
.A(n_3663),
.B(n_3334),
.Y(n_4105)
);

NAND2xp5_ASAP7_75t_SL g4106 ( 
.A(n_3688),
.B(n_3312),
.Y(n_4106)
);

NAND2xp5_ASAP7_75t_L g4107 ( 
.A(n_3628),
.B(n_3462),
.Y(n_4107)
);

NAND2xp5_ASAP7_75t_SL g4108 ( 
.A(n_3693),
.B(n_3372),
.Y(n_4108)
);

NAND2xp33_ASAP7_75t_SL g4109 ( 
.A(n_3679),
.B(n_3779),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_SL g4110 ( 
.A(n_3813),
.B(n_3119),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_SL g4111 ( 
.A(n_3767),
.B(n_3119),
.Y(n_4111)
);

NAND2xp5_ASAP7_75t_SL g4112 ( 
.A(n_3618),
.B(n_3128),
.Y(n_4112)
);

AND2x4_ASAP7_75t_L g4113 ( 
.A(n_3746),
.B(n_3493),
.Y(n_4113)
);

NAND2xp5_ASAP7_75t_SL g4114 ( 
.A(n_3740),
.B(n_3128),
.Y(n_4114)
);

NAND2xp33_ASAP7_75t_SL g4115 ( 
.A(n_3634),
.B(n_909),
.Y(n_4115)
);

NAND2xp5_ASAP7_75t_SL g4116 ( 
.A(n_3841),
.B(n_3518),
.Y(n_4116)
);

NAND2xp5_ASAP7_75t_SL g4117 ( 
.A(n_3838),
.B(n_3453),
.Y(n_4117)
);

NAND2xp5_ASAP7_75t_SL g4118 ( 
.A(n_3629),
.B(n_3453),
.Y(n_4118)
);

NAND2xp33_ASAP7_75t_SL g4119 ( 
.A(n_3788),
.B(n_931),
.Y(n_4119)
);

NAND2xp5_ASAP7_75t_SL g4120 ( 
.A(n_3825),
.B(n_3367),
.Y(n_4120)
);

NAND2xp5_ASAP7_75t_SL g4121 ( 
.A(n_3641),
.B(n_3367),
.Y(n_4121)
);

NAND2xp5_ASAP7_75t_L g4122 ( 
.A(n_3631),
.B(n_3494),
.Y(n_4122)
);

NAND2xp5_ASAP7_75t_L g4123 ( 
.A(n_3636),
.B(n_3502),
.Y(n_4123)
);

NAND2xp5_ASAP7_75t_L g4124 ( 
.A(n_3640),
.B(n_3509),
.Y(n_4124)
);

NAND2xp5_ASAP7_75t_SL g4125 ( 
.A(n_3867),
.B(n_3875),
.Y(n_4125)
);

NAND2xp5_ASAP7_75t_L g4126 ( 
.A(n_3642),
.B(n_3513),
.Y(n_4126)
);

NAND2xp5_ASAP7_75t_SL g4127 ( 
.A(n_3585),
.B(n_3536),
.Y(n_4127)
);

NAND2xp5_ASAP7_75t_SL g4128 ( 
.A(n_3585),
.B(n_3308),
.Y(n_4128)
);

NAND2xp33_ASAP7_75t_SL g4129 ( 
.A(n_3733),
.B(n_940),
.Y(n_4129)
);

NAND2xp5_ASAP7_75t_SL g4130 ( 
.A(n_3820),
.B(n_3330),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_SL g4131 ( 
.A(n_3738),
.B(n_3330),
.Y(n_4131)
);

NAND2xp33_ASAP7_75t_SL g4132 ( 
.A(n_3756),
.B(n_3716),
.Y(n_4132)
);

NAND2xp33_ASAP7_75t_SL g4133 ( 
.A(n_3650),
.B(n_941),
.Y(n_4133)
);

NAND2xp5_ASAP7_75t_L g4134 ( 
.A(n_3651),
.B(n_3526),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_SL g4135 ( 
.A(n_3827),
.B(n_3440),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_SL g4136 ( 
.A(n_3798),
.B(n_3846),
.Y(n_4136)
);

NAND2xp5_ASAP7_75t_L g4137 ( 
.A(n_3652),
.B(n_3533),
.Y(n_4137)
);

NAND2xp5_ASAP7_75t_SL g4138 ( 
.A(n_3798),
.B(n_3819),
.Y(n_4138)
);

NAND2xp5_ASAP7_75t_L g4139 ( 
.A(n_3659),
.B(n_3557),
.Y(n_4139)
);

NAND2xp5_ASAP7_75t_L g4140 ( 
.A(n_3662),
.B(n_3561),
.Y(n_4140)
);

NAND2xp5_ASAP7_75t_SL g4141 ( 
.A(n_3819),
.B(n_3464),
.Y(n_4141)
);

NAND2xp5_ASAP7_75t_L g4142 ( 
.A(n_3881),
.B(n_3666),
.Y(n_4142)
);

O2A1O1Ixp33_ASAP7_75t_L g4143 ( 
.A1(n_3892),
.A2(n_3649),
.B(n_1023),
.C(n_1027),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4099),
.Y(n_4144)
);

INVx1_ASAP7_75t_L g4145 ( 
.A(n_4141),
.Y(n_4145)
);

O2A1O1Ixp33_ASAP7_75t_L g4146 ( 
.A1(n_4108),
.A2(n_1023),
.B(n_1027),
.C(n_1021),
.Y(n_4146)
);

INVx2_ASAP7_75t_L g4147 ( 
.A(n_4102),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4104),
.Y(n_4148)
);

BUFx2_ASAP7_75t_L g4149 ( 
.A(n_4086),
.Y(n_4149)
);

CKINVDCx20_ASAP7_75t_R g4150 ( 
.A(n_4132),
.Y(n_4150)
);

INVx2_ASAP7_75t_SL g4151 ( 
.A(n_3967),
.Y(n_4151)
);

INVx1_ASAP7_75t_SL g4152 ( 
.A(n_3958),
.Y(n_4152)
);

INVx1_ASAP7_75t_L g4153 ( 
.A(n_4107),
.Y(n_4153)
);

INVx3_ASAP7_75t_L g4154 ( 
.A(n_3997),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_3937),
.B(n_3668),
.Y(n_4155)
);

INVx3_ASAP7_75t_L g4156 ( 
.A(n_3997),
.Y(n_4156)
);

O2A1O1Ixp5_ASAP7_75t_SL g4157 ( 
.A1(n_4121),
.A2(n_3675),
.B(n_3678),
.C(n_3673),
.Y(n_4157)
);

INVx1_ASAP7_75t_L g4158 ( 
.A(n_4122),
.Y(n_4158)
);

BUFx6f_ASAP7_75t_L g4159 ( 
.A(n_4063),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4123),
.Y(n_4160)
);

O2A1O1Ixp33_ASAP7_75t_SL g4161 ( 
.A1(n_3878),
.A2(n_1030),
.B(n_1033),
.C(n_1029),
.Y(n_4161)
);

NAND2xp5_ASAP7_75t_L g4162 ( 
.A(n_3878),
.B(n_3680),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_3887),
.B(n_3683),
.Y(n_4163)
);

AOI21xp5_ASAP7_75t_L g4164 ( 
.A1(n_4037),
.A2(n_3501),
.B(n_3844),
.Y(n_4164)
);

BUFx2_ASAP7_75t_L g4165 ( 
.A(n_3907),
.Y(n_4165)
);

HB1xp67_ASAP7_75t_L g4166 ( 
.A(n_3910),
.Y(n_4166)
);

AOI21x1_ASAP7_75t_L g4167 ( 
.A1(n_4039),
.A2(n_3853),
.B(n_3572),
.Y(n_4167)
);

OAI21xp5_ASAP7_75t_L g4168 ( 
.A1(n_4018),
.A2(n_3845),
.B(n_3464),
.Y(n_4168)
);

BUFx2_ASAP7_75t_L g4169 ( 
.A(n_3981),
.Y(n_4169)
);

NAND2xp5_ASAP7_75t_L g4170 ( 
.A(n_3983),
.B(n_3697),
.Y(n_4170)
);

AOI21xp33_ASAP7_75t_L g4171 ( 
.A1(n_4036),
.A2(n_3614),
.B(n_3845),
.Y(n_4171)
);

OR2x6_ASAP7_75t_L g4172 ( 
.A(n_4082),
.B(n_3637),
.Y(n_4172)
);

CKINVDCx8_ASAP7_75t_R g4173 ( 
.A(n_4096),
.Y(n_4173)
);

INVx2_ASAP7_75t_L g4174 ( 
.A(n_4124),
.Y(n_4174)
);

AND2x2_ASAP7_75t_L g4175 ( 
.A(n_3973),
.B(n_3699),
.Y(n_4175)
);

AOI21x1_ASAP7_75t_L g4176 ( 
.A1(n_3915),
.A2(n_4120),
.B(n_4105),
.Y(n_4176)
);

INVx4_ASAP7_75t_L g4177 ( 
.A(n_4063),
.Y(n_4177)
);

AND2x4_ASAP7_75t_L g4178 ( 
.A(n_3997),
.B(n_3701),
.Y(n_4178)
);

INVx2_ASAP7_75t_SL g4179 ( 
.A(n_4063),
.Y(n_4179)
);

INVx1_ASAP7_75t_L g4180 ( 
.A(n_4126),
.Y(n_4180)
);

OAI22x1_ASAP7_75t_L g4181 ( 
.A1(n_3913),
.A2(n_3702),
.B1(n_3706),
.B2(n_3703),
.Y(n_4181)
);

NOR2xp33_ASAP7_75t_L g4182 ( 
.A(n_3885),
.B(n_3607),
.Y(n_4182)
);

OAI21xp5_ASAP7_75t_L g4183 ( 
.A1(n_3916),
.A2(n_3870),
.B(n_3314),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4134),
.Y(n_4184)
);

HB1xp67_ASAP7_75t_L g4185 ( 
.A(n_4125),
.Y(n_4185)
);

AOI21xp5_ASAP7_75t_L g4186 ( 
.A1(n_3963),
.A2(n_3479),
.B(n_3249),
.Y(n_4186)
);

NOR2xp33_ASAP7_75t_L g4187 ( 
.A(n_3953),
.B(n_3732),
.Y(n_4187)
);

A2O1A1Ixp33_ASAP7_75t_L g4188 ( 
.A1(n_4133),
.A2(n_3715),
.B(n_3874),
.C(n_3719),
.Y(n_4188)
);

INVxp67_ASAP7_75t_L g4189 ( 
.A(n_3961),
.Y(n_4189)
);

OAI22xp33_ASAP7_75t_L g4190 ( 
.A1(n_4031),
.A2(n_3835),
.B1(n_3715),
.B2(n_3766),
.Y(n_4190)
);

INVx2_ASAP7_75t_L g4191 ( 
.A(n_4137),
.Y(n_4191)
);

AOI22xp33_ASAP7_75t_L g4192 ( 
.A1(n_4090),
.A2(n_3877),
.B1(n_3562),
.B2(n_3595),
.Y(n_4192)
);

INVx1_ASAP7_75t_SL g4193 ( 
.A(n_3995),
.Y(n_4193)
);

NAND2xp5_ASAP7_75t_SL g4194 ( 
.A(n_4100),
.B(n_3722),
.Y(n_4194)
);

NOR2xp33_ASAP7_75t_L g4195 ( 
.A(n_3942),
.B(n_3582),
.Y(n_4195)
);

NOR2xp67_ASAP7_75t_SL g4196 ( 
.A(n_3969),
.B(n_3772),
.Y(n_4196)
);

AOI21x1_ASAP7_75t_L g4197 ( 
.A1(n_4116),
.A2(n_4130),
.B(n_4073),
.Y(n_4197)
);

INVx2_ASAP7_75t_L g4198 ( 
.A(n_4139),
.Y(n_4198)
);

INVx5_ASAP7_75t_L g4199 ( 
.A(n_4085),
.Y(n_4199)
);

INVx1_ASAP7_75t_L g4200 ( 
.A(n_4140),
.Y(n_4200)
);

NOR2xp33_ASAP7_75t_L g4201 ( 
.A(n_3879),
.B(n_947),
.Y(n_4201)
);

AOI22xp5_ASAP7_75t_L g4202 ( 
.A1(n_4119),
.A2(n_4042),
.B1(n_3977),
.B2(n_3941),
.Y(n_4202)
);

NAND2xp5_ASAP7_75t_L g4203 ( 
.A(n_3921),
.B(n_3710),
.Y(n_4203)
);

INVx2_ASAP7_75t_SL g4204 ( 
.A(n_4085),
.Y(n_4204)
);

CKINVDCx5p33_ASAP7_75t_R g4205 ( 
.A(n_3986),
.Y(n_4205)
);

BUFx12f_ASAP7_75t_L g4206 ( 
.A(n_4097),
.Y(n_4206)
);

INVx2_ASAP7_75t_L g4207 ( 
.A(n_4095),
.Y(n_4207)
);

NOR2xp67_ASAP7_75t_SL g4208 ( 
.A(n_3901),
.B(n_3637),
.Y(n_4208)
);

AND2x4_ASAP7_75t_L g4209 ( 
.A(n_4038),
.B(n_3725),
.Y(n_4209)
);

INVx1_ASAP7_75t_L g4210 ( 
.A(n_4057),
.Y(n_4210)
);

OAI22xp5_ASAP7_75t_L g4211 ( 
.A1(n_4030),
.A2(n_3871),
.B1(n_3775),
.B2(n_3835),
.Y(n_4211)
);

NOR2xp33_ASAP7_75t_L g4212 ( 
.A(n_3893),
.B(n_3926),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4051),
.Y(n_4213)
);

INVx1_ASAP7_75t_L g4214 ( 
.A(n_3891),
.Y(n_4214)
);

INVx2_ASAP7_75t_L g4215 ( 
.A(n_3938),
.Y(n_4215)
);

INVx1_ASAP7_75t_L g4216 ( 
.A(n_3959),
.Y(n_4216)
);

NAND2xp5_ASAP7_75t_L g4217 ( 
.A(n_3917),
.B(n_3729),
.Y(n_4217)
);

AOI21xp5_ASAP7_75t_L g4218 ( 
.A1(n_4100),
.A2(n_3479),
.B(n_3249),
.Y(n_4218)
);

INVx1_ASAP7_75t_L g4219 ( 
.A(n_3947),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_3918),
.B(n_3742),
.Y(n_4220)
);

INVx1_ASAP7_75t_L g4221 ( 
.A(n_3974),
.Y(n_4221)
);

INVx4_ASAP7_75t_L g4222 ( 
.A(n_4085),
.Y(n_4222)
);

INVx1_ASAP7_75t_L g4223 ( 
.A(n_3943),
.Y(n_4223)
);

O2A1O1Ixp33_ASAP7_75t_L g4224 ( 
.A1(n_4127),
.A2(n_1030),
.B(n_1042),
.C(n_1029),
.Y(n_4224)
);

NAND2xp5_ASAP7_75t_SL g4225 ( 
.A(n_3900),
.B(n_3848),
.Y(n_4225)
);

A2O1A1Ixp33_ASAP7_75t_L g4226 ( 
.A1(n_4088),
.A2(n_3847),
.B(n_3762),
.C(n_3763),
.Y(n_4226)
);

AND2x4_ASAP7_75t_L g4227 ( 
.A(n_4038),
.B(n_3749),
.Y(n_4227)
);

INVx2_ASAP7_75t_SL g4228 ( 
.A(n_4060),
.Y(n_4228)
);

HB1xp67_ASAP7_75t_L g4229 ( 
.A(n_4015),
.Y(n_4229)
);

INVx1_ASAP7_75t_L g4230 ( 
.A(n_3880),
.Y(n_4230)
);

NOR2xp33_ASAP7_75t_L g4231 ( 
.A(n_3927),
.B(n_953),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_SL g4232 ( 
.A(n_4109),
.B(n_3771),
.Y(n_4232)
);

NAND2xp5_ASAP7_75t_SL g4233 ( 
.A(n_3928),
.B(n_3774),
.Y(n_4233)
);

INVx4_ASAP7_75t_L g4234 ( 
.A(n_4060),
.Y(n_4234)
);

INVx2_ASAP7_75t_L g4235 ( 
.A(n_4096),
.Y(n_4235)
);

OAI22xp5_ASAP7_75t_L g4236 ( 
.A1(n_4135),
.A2(n_3835),
.B1(n_3777),
.B2(n_3785),
.Y(n_4236)
);

INVx2_ASAP7_75t_SL g4237 ( 
.A(n_4060),
.Y(n_4237)
);

INVx2_ASAP7_75t_L g4238 ( 
.A(n_4096),
.Y(n_4238)
);

AND2x2_ASAP7_75t_L g4239 ( 
.A(n_4014),
.B(n_3783),
.Y(n_4239)
);

INVx3_ASAP7_75t_L g4240 ( 
.A(n_4038),
.Y(n_4240)
);

INVx2_ASAP7_75t_L g4241 ( 
.A(n_4113),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4034),
.B(n_3812),
.Y(n_4242)
);

INVx2_ASAP7_75t_L g4243 ( 
.A(n_4113),
.Y(n_4243)
);

BUFx6f_ASAP7_75t_L g4244 ( 
.A(n_4113),
.Y(n_4244)
);

INVx3_ASAP7_75t_L g4245 ( 
.A(n_3940),
.Y(n_4245)
);

INVx2_ASAP7_75t_L g4246 ( 
.A(n_4061),
.Y(n_4246)
);

NAND2xp5_ASAP7_75t_L g4247 ( 
.A(n_4070),
.B(n_3954),
.Y(n_4247)
);

AOI21x1_ASAP7_75t_L g4248 ( 
.A1(n_4053),
.A2(n_3572),
.B(n_3856),
.Y(n_4248)
);

NOR2xp33_ASAP7_75t_L g4249 ( 
.A(n_4106),
.B(n_954),
.Y(n_4249)
);

BUFx12f_ASAP7_75t_L g4250 ( 
.A(n_3940),
.Y(n_4250)
);

INVx1_ASAP7_75t_L g4251 ( 
.A(n_3939),
.Y(n_4251)
);

OAI22xp5_ASAP7_75t_L g4252 ( 
.A1(n_4135),
.A2(n_3828),
.B1(n_3839),
.B2(n_3817),
.Y(n_4252)
);

AOI22xp33_ASAP7_75t_SL g4253 ( 
.A1(n_4074),
.A2(n_4043),
.B1(n_3906),
.B2(n_4075),
.Y(n_4253)
);

INVx2_ASAP7_75t_L g4254 ( 
.A(n_4012),
.Y(n_4254)
);

INVx3_ASAP7_75t_L g4255 ( 
.A(n_3940),
.Y(n_4255)
);

AOI22xp5_ASAP7_75t_L g4256 ( 
.A1(n_4103),
.A2(n_3773),
.B1(n_3870),
.B2(n_3843),
.Y(n_4256)
);

INVx1_ASAP7_75t_SL g4257 ( 
.A(n_3914),
.Y(n_4257)
);

INVx1_ASAP7_75t_L g4258 ( 
.A(n_3882),
.Y(n_4258)
);

CKINVDCx5p33_ASAP7_75t_R g4259 ( 
.A(n_3930),
.Y(n_4259)
);

INVx2_ASAP7_75t_L g4260 ( 
.A(n_3905),
.Y(n_4260)
);

AO22x1_ASAP7_75t_L g4261 ( 
.A1(n_3988),
.A2(n_3870),
.B1(n_3773),
.B2(n_3592),
.Y(n_4261)
);

AOI21xp5_ASAP7_75t_L g4262 ( 
.A1(n_3908),
.A2(n_3226),
.B(n_3314),
.Y(n_4262)
);

BUFx6f_ASAP7_75t_L g4263 ( 
.A(n_3988),
.Y(n_4263)
);

CKINVDCx11_ASAP7_75t_R g4264 ( 
.A(n_3988),
.Y(n_4264)
);

INVx2_ASAP7_75t_L g4265 ( 
.A(n_3960),
.Y(n_4265)
);

INVxp67_ASAP7_75t_L g4266 ( 
.A(n_3925),
.Y(n_4266)
);

INVx1_ASAP7_75t_L g4267 ( 
.A(n_3882),
.Y(n_4267)
);

NOR2xp33_ASAP7_75t_L g4268 ( 
.A(n_4023),
.B(n_957),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_3883),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_3883),
.Y(n_4270)
);

INVx2_ASAP7_75t_L g4271 ( 
.A(n_4076),
.Y(n_4271)
);

OAI21xp5_ASAP7_75t_L g4272 ( 
.A1(n_4131),
.A2(n_3870),
.B(n_3773),
.Y(n_4272)
);

INVx2_ASAP7_75t_L g4273 ( 
.A(n_4077),
.Y(n_4273)
);

INVx1_ASAP7_75t_SL g4274 ( 
.A(n_3935),
.Y(n_4274)
);

OAI22xp5_ASAP7_75t_L g4275 ( 
.A1(n_3894),
.A2(n_3814),
.B1(n_3727),
.B2(n_1042),
.Y(n_4275)
);

INVx4_ASAP7_75t_L g4276 ( 
.A(n_3944),
.Y(n_4276)
);

NAND2xp5_ASAP7_75t_SL g4277 ( 
.A(n_3929),
.B(n_3857),
.Y(n_4277)
);

AOI21xp5_ASAP7_75t_L g4278 ( 
.A1(n_3971),
.A2(n_3226),
.B(n_3861),
.Y(n_4278)
);

AOI22xp5_ASAP7_75t_L g4279 ( 
.A1(n_4115),
.A2(n_3773),
.B1(n_963),
.B2(n_964),
.Y(n_4279)
);

AOI21xp5_ASAP7_75t_L g4280 ( 
.A1(n_3985),
.A2(n_3863),
.B(n_3861),
.Y(n_4280)
);

AOI21xp5_ASAP7_75t_L g4281 ( 
.A1(n_4029),
.A2(n_3863),
.B(n_3851),
.Y(n_4281)
);

A2O1A1Ixp33_ASAP7_75t_L g4282 ( 
.A1(n_3952),
.A2(n_1043),
.B(n_1048),
.C(n_1033),
.Y(n_4282)
);

INVxp67_ASAP7_75t_L g4283 ( 
.A(n_3979),
.Y(n_4283)
);

BUFx6f_ASAP7_75t_L g4284 ( 
.A(n_3965),
.Y(n_4284)
);

CKINVDCx6p67_ASAP7_75t_R g4285 ( 
.A(n_4006),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4011),
.B(n_1043),
.Y(n_4286)
);

INVx1_ASAP7_75t_SL g4287 ( 
.A(n_3946),
.Y(n_4287)
);

BUFx4f_ASAP7_75t_SL g4288 ( 
.A(n_3966),
.Y(n_4288)
);

BUFx10_ASAP7_75t_L g4289 ( 
.A(n_4129),
.Y(n_4289)
);

OR2x6_ASAP7_75t_L g4290 ( 
.A(n_4118),
.B(n_3623),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_3949),
.Y(n_4291)
);

A2O1A1Ixp33_ASAP7_75t_L g4292 ( 
.A1(n_3920),
.A2(n_1053),
.B(n_1055),
.C(n_1048),
.Y(n_4292)
);

NOR2x1_ASAP7_75t_SL g4293 ( 
.A(n_4084),
.B(n_3842),
.Y(n_4293)
);

NAND2xp5_ASAP7_75t_L g4294 ( 
.A(n_3903),
.B(n_3860),
.Y(n_4294)
);

CKINVDCx5p33_ASAP7_75t_R g4295 ( 
.A(n_3990),
.Y(n_4295)
);

AOI22xp33_ASAP7_75t_L g4296 ( 
.A1(n_3919),
.A2(n_3612),
.B1(n_3630),
.B2(n_3591),
.Y(n_4296)
);

INVx2_ASAP7_75t_SL g4297 ( 
.A(n_4065),
.Y(n_4297)
);

INVx1_ASAP7_75t_L g4298 ( 
.A(n_3950),
.Y(n_4298)
);

INVx1_ASAP7_75t_L g4299 ( 
.A(n_3884),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4111),
.Y(n_4300)
);

OR2x6_ASAP7_75t_L g4301 ( 
.A(n_4054),
.B(n_3644),
.Y(n_4301)
);

OAI22xp5_ASAP7_75t_L g4302 ( 
.A1(n_3951),
.A2(n_1055),
.B1(n_1061),
.B2(n_1053),
.Y(n_4302)
);

BUFx6f_ASAP7_75t_L g4303 ( 
.A(n_3978),
.Y(n_4303)
);

O2A1O1Ixp33_ASAP7_75t_L g4304 ( 
.A1(n_3889),
.A2(n_3890),
.B(n_3886),
.C(n_3888),
.Y(n_4304)
);

OAI22xp5_ASAP7_75t_L g4305 ( 
.A1(n_3956),
.A2(n_1063),
.B1(n_1080),
.B2(n_1061),
.Y(n_4305)
);

INVx2_ASAP7_75t_L g4306 ( 
.A(n_4098),
.Y(n_4306)
);

INVx5_ASAP7_75t_L g4307 ( 
.A(n_4021),
.Y(n_4307)
);

INVx2_ASAP7_75t_L g4308 ( 
.A(n_3968),
.Y(n_4308)
);

NAND2xp5_ASAP7_75t_L g4309 ( 
.A(n_3924),
.B(n_3647),
.Y(n_4309)
);

AOI21xp5_ASAP7_75t_L g4310 ( 
.A1(n_4138),
.A2(n_3624),
.B(n_3859),
.Y(n_4310)
);

INVx3_ASAP7_75t_L g4311 ( 
.A(n_3964),
.Y(n_4311)
);

BUFx12f_ASAP7_75t_L g4312 ( 
.A(n_4028),
.Y(n_4312)
);

INVx1_ASAP7_75t_L g4313 ( 
.A(n_3884),
.Y(n_4313)
);

AND2x4_ASAP7_75t_L g4314 ( 
.A(n_3933),
.B(n_3669),
.Y(n_4314)
);

AOI21xp5_ASAP7_75t_L g4315 ( 
.A1(n_4138),
.A2(n_2423),
.B(n_3689),
.Y(n_4315)
);

CKINVDCx20_ASAP7_75t_R g4316 ( 
.A(n_4089),
.Y(n_4316)
);

AOI21xp5_ASAP7_75t_L g4317 ( 
.A1(n_3909),
.A2(n_2423),
.B(n_3694),
.Y(n_4317)
);

NAND2xp5_ASAP7_75t_L g4318 ( 
.A(n_3899),
.B(n_3902),
.Y(n_4318)
);

NAND2x1p5_ASAP7_75t_L g4319 ( 
.A(n_4081),
.B(n_3793),
.Y(n_4319)
);

OAI22xp5_ASAP7_75t_L g4320 ( 
.A1(n_4128),
.A2(n_1080),
.B1(n_1082),
.B2(n_1063),
.Y(n_4320)
);

AOI22xp5_ASAP7_75t_L g4321 ( 
.A1(n_4010),
.A2(n_4020),
.B1(n_3911),
.B2(n_3912),
.Y(n_4321)
);

INVx2_ASAP7_75t_L g4322 ( 
.A(n_3923),
.Y(n_4322)
);

NAND2xp5_ASAP7_75t_L g4323 ( 
.A(n_3904),
.B(n_3709),
.Y(n_4323)
);

O2A1O1Ixp33_ASAP7_75t_L g4324 ( 
.A1(n_3957),
.A2(n_1097),
.B(n_1103),
.C(n_1098),
.Y(n_4324)
);

NOR2xp33_ASAP7_75t_L g4325 ( 
.A(n_3931),
.B(n_959),
.Y(n_4325)
);

NAND2xp5_ASAP7_75t_L g4326 ( 
.A(n_3936),
.B(n_3743),
.Y(n_4326)
);

AOI22xp5_ASAP7_75t_L g4327 ( 
.A1(n_4024),
.A2(n_975),
.B1(n_979),
.B2(n_968),
.Y(n_4327)
);

AND2x4_ASAP7_75t_L g4328 ( 
.A(n_3980),
.B(n_3753),
.Y(n_4328)
);

BUFx2_ASAP7_75t_L g4329 ( 
.A(n_3955),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4013),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4025),
.B(n_3755),
.Y(n_4331)
);

NOR2xp33_ASAP7_75t_L g4332 ( 
.A(n_4112),
.B(n_986),
.Y(n_4332)
);

NOR2xp33_ASAP7_75t_L g4333 ( 
.A(n_4041),
.B(n_994),
.Y(n_4333)
);

NAND2xp5_ASAP7_75t_L g4334 ( 
.A(n_4117),
.B(n_3778),
.Y(n_4334)
);

OAI22xp5_ASAP7_75t_SL g4335 ( 
.A1(n_3895),
.A2(n_1097),
.B1(n_1098),
.B2(n_1083),
.Y(n_4335)
);

INVx2_ASAP7_75t_L g4336 ( 
.A(n_3922),
.Y(n_4336)
);

NAND2xp5_ASAP7_75t_SL g4337 ( 
.A(n_4048),
.B(n_4046),
.Y(n_4337)
);

NOR2xp67_ASAP7_75t_L g4338 ( 
.A(n_4136),
.B(n_1318),
.Y(n_4338)
);

NAND2xp5_ASAP7_75t_SL g4339 ( 
.A(n_4055),
.B(n_3786),
.Y(n_4339)
);

CKINVDCx20_ASAP7_75t_R g4340 ( 
.A(n_4066),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_3945),
.Y(n_4341)
);

INVx2_ASAP7_75t_SL g4342 ( 
.A(n_4047),
.Y(n_4342)
);

BUFx6f_ASAP7_75t_L g4343 ( 
.A(n_3975),
.Y(n_4343)
);

NOR2xp33_ASAP7_75t_L g4344 ( 
.A(n_4044),
.B(n_998),
.Y(n_4344)
);

AND2x2_ASAP7_75t_L g4345 ( 
.A(n_4016),
.B(n_4017),
.Y(n_4345)
);

NOR3xp33_ASAP7_75t_L g4346 ( 
.A(n_4004),
.B(n_1103),
.C(n_1083),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4101),
.Y(n_4347)
);

AND2x4_ASAP7_75t_L g4348 ( 
.A(n_3932),
.B(n_3787),
.Y(n_4348)
);

INVx1_ASAP7_75t_L g4349 ( 
.A(n_4092),
.Y(n_4349)
);

CKINVDCx5p33_ASAP7_75t_R g4350 ( 
.A(n_4091),
.Y(n_4350)
);

INVx2_ASAP7_75t_L g4351 ( 
.A(n_4094),
.Y(n_4351)
);

NAND2x1_ASAP7_75t_SL g4352 ( 
.A(n_4052),
.B(n_1319),
.Y(n_4352)
);

CKINVDCx6p67_ASAP7_75t_R g4353 ( 
.A(n_3970),
.Y(n_4353)
);

INVx1_ASAP7_75t_L g4354 ( 
.A(n_4136),
.Y(n_4354)
);

AOI21xp5_ASAP7_75t_L g4355 ( 
.A1(n_3896),
.A2(n_3821),
.B(n_3815),
.Y(n_4355)
);

AND2x4_ASAP7_75t_L g4356 ( 
.A(n_3934),
.B(n_3872),
.Y(n_4356)
);

INVx2_ASAP7_75t_SL g4357 ( 
.A(n_4049),
.Y(n_4357)
);

AOI22xp33_ASAP7_75t_L g4358 ( 
.A1(n_4110),
.A2(n_3876),
.B1(n_1107),
.B2(n_1112),
.Y(n_4358)
);

NOR2xp33_ASAP7_75t_SL g4359 ( 
.A(n_4067),
.B(n_3173),
.Y(n_4359)
);

OAI22xp5_ASAP7_75t_L g4360 ( 
.A1(n_4022),
.A2(n_1107),
.B1(n_1112),
.B2(n_1104),
.Y(n_4360)
);

OR2x2_ASAP7_75t_L g4361 ( 
.A(n_4026),
.B(n_1321),
.Y(n_4361)
);

BUFx6f_ASAP7_75t_L g4362 ( 
.A(n_3976),
.Y(n_4362)
);

INVx1_ASAP7_75t_L g4363 ( 
.A(n_4114),
.Y(n_4363)
);

AOI21xp5_ASAP7_75t_L g4364 ( 
.A1(n_4019),
.A2(n_1114),
.B(n_1104),
.Y(n_4364)
);

INVx2_ASAP7_75t_L g4365 ( 
.A(n_4027),
.Y(n_4365)
);

BUFx3_ASAP7_75t_L g4366 ( 
.A(n_4079),
.Y(n_4366)
);

BUFx8_ASAP7_75t_L g4367 ( 
.A(n_4032),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4078),
.Y(n_4368)
);

INVx2_ASAP7_75t_L g4369 ( 
.A(n_4080),
.Y(n_4369)
);

INVx3_ASAP7_75t_SL g4370 ( 
.A(n_3989),
.Y(n_4370)
);

AOI21xp5_ASAP7_75t_L g4371 ( 
.A1(n_3962),
.A2(n_4093),
.B(n_3898),
.Y(n_4371)
);

HB1xp67_ASAP7_75t_L g4372 ( 
.A(n_4050),
.Y(n_4372)
);

INVx3_ASAP7_75t_L g4373 ( 
.A(n_4033),
.Y(n_4373)
);

O2A1O1Ixp33_ASAP7_75t_L g4374 ( 
.A1(n_4040),
.A2(n_1126),
.B(n_1127),
.C(n_1114),
.Y(n_4374)
);

INVx2_ASAP7_75t_L g4375 ( 
.A(n_4056),
.Y(n_4375)
);

BUFx3_ASAP7_75t_L g4376 ( 
.A(n_3991),
.Y(n_4376)
);

A2O1A1Ixp33_ASAP7_75t_L g4377 ( 
.A1(n_3897),
.A2(n_1127),
.B(n_1129),
.C(n_1126),
.Y(n_4377)
);

INVx3_ASAP7_75t_L g4378 ( 
.A(n_4035),
.Y(n_4378)
);

INVx2_ASAP7_75t_L g4379 ( 
.A(n_4058),
.Y(n_4379)
);

BUFx6f_ASAP7_75t_L g4380 ( 
.A(n_3972),
.Y(n_4380)
);

BUFx3_ASAP7_75t_L g4381 ( 
.A(n_3992),
.Y(n_4381)
);

A2O1A1Ixp33_ASAP7_75t_L g4382 ( 
.A1(n_4045),
.A2(n_1130),
.B(n_1131),
.C(n_1129),
.Y(n_4382)
);

BUFx6f_ASAP7_75t_L g4383 ( 
.A(n_3982),
.Y(n_4383)
);

OAI22xp5_ASAP7_75t_L g4384 ( 
.A1(n_3948),
.A2(n_1131),
.B1(n_1144),
.B2(n_1130),
.Y(n_4384)
);

BUFx3_ASAP7_75t_L g4385 ( 
.A(n_3993),
.Y(n_4385)
);

OR2x6_ASAP7_75t_L g4386 ( 
.A(n_4083),
.B(n_3173),
.Y(n_4386)
);

NAND2xp5_ASAP7_75t_L g4387 ( 
.A(n_3994),
.B(n_1144),
.Y(n_4387)
);

INVx4_ASAP7_75t_L g4388 ( 
.A(n_3996),
.Y(n_4388)
);

OR2x6_ASAP7_75t_L g4389 ( 
.A(n_4087),
.B(n_1322),
.Y(n_4389)
);

INVx4_ASAP7_75t_L g4390 ( 
.A(n_4259),
.Y(n_4390)
);

A2O1A1Ixp33_ASAP7_75t_L g4391 ( 
.A1(n_4279),
.A2(n_1154),
.B(n_1158),
.C(n_1151),
.Y(n_4391)
);

AOI22xp33_ASAP7_75t_L g4392 ( 
.A1(n_4171),
.A2(n_1151),
.B1(n_1158),
.B2(n_1154),
.Y(n_4392)
);

BUFx2_ASAP7_75t_L g4393 ( 
.A(n_4149),
.Y(n_4393)
);

AOI22xp5_ASAP7_75t_L g4394 ( 
.A1(n_4321),
.A2(n_4062),
.B1(n_4064),
.B2(n_4059),
.Y(n_4394)
);

INVx1_ASAP7_75t_L g4395 ( 
.A(n_4258),
.Y(n_4395)
);

INVx2_ASAP7_75t_L g4396 ( 
.A(n_4144),
.Y(n_4396)
);

AND2x2_ASAP7_75t_L g4397 ( 
.A(n_4163),
.B(n_3998),
.Y(n_4397)
);

A2O1A1Ixp33_ASAP7_75t_L g4398 ( 
.A1(n_4164),
.A2(n_4143),
.B(n_4201),
.C(n_4256),
.Y(n_4398)
);

INVx5_ASAP7_75t_L g4399 ( 
.A(n_4307),
.Y(n_4399)
);

AOI21xp5_ASAP7_75t_L g4400 ( 
.A1(n_4337),
.A2(n_3987),
.B(n_3984),
.Y(n_4400)
);

AOI21xp5_ASAP7_75t_L g4401 ( 
.A1(n_4311),
.A2(n_4000),
.B(n_3999),
.Y(n_4401)
);

O2A1O1Ixp33_ASAP7_75t_SL g4402 ( 
.A1(n_4150),
.A2(n_1169),
.B(n_1170),
.C(n_1168),
.Y(n_4402)
);

AOI21x1_ASAP7_75t_L g4403 ( 
.A1(n_4197),
.A2(n_4002),
.B(n_4001),
.Y(n_4403)
);

INVx1_ASAP7_75t_SL g4404 ( 
.A(n_4205),
.Y(n_4404)
);

AOI221xp5_ASAP7_75t_L g4405 ( 
.A1(n_4146),
.A2(n_1170),
.B1(n_1177),
.B2(n_1169),
.C(n_1168),
.Y(n_4405)
);

BUFx2_ASAP7_75t_L g4406 ( 
.A(n_4165),
.Y(n_4406)
);

INVx3_ASAP7_75t_L g4407 ( 
.A(n_4159),
.Y(n_4407)
);

INVx1_ASAP7_75t_SL g4408 ( 
.A(n_4206),
.Y(n_4408)
);

A2O1A1Ixp33_ASAP7_75t_L g4409 ( 
.A1(n_4202),
.A2(n_1178),
.B(n_1179),
.C(n_1177),
.Y(n_4409)
);

O2A1O1Ixp33_ASAP7_75t_L g4410 ( 
.A1(n_4282),
.A2(n_1179),
.B(n_1185),
.C(n_1178),
.Y(n_4410)
);

INVxp67_ASAP7_75t_L g4411 ( 
.A(n_4169),
.Y(n_4411)
);

AOI21xp5_ASAP7_75t_L g4412 ( 
.A1(n_4311),
.A2(n_4005),
.B(n_4003),
.Y(n_4412)
);

NOR2xp33_ASAP7_75t_L g4413 ( 
.A(n_4187),
.B(n_6),
.Y(n_4413)
);

INVx1_ASAP7_75t_L g4414 ( 
.A(n_4267),
.Y(n_4414)
);

O2A1O1Ixp5_ASAP7_75t_L g4415 ( 
.A1(n_4176),
.A2(n_4008),
.B(n_4009),
.C(n_4007),
.Y(n_4415)
);

NOR2xp33_ASAP7_75t_L g4416 ( 
.A(n_4193),
.B(n_6),
.Y(n_4416)
);

OAI21x1_ASAP7_75t_L g4417 ( 
.A1(n_4262),
.A2(n_4069),
.B(n_4068),
.Y(n_4417)
);

O2A1O1Ixp33_ASAP7_75t_SL g4418 ( 
.A1(n_4257),
.A2(n_1193),
.B(n_1202),
.C(n_1185),
.Y(n_4418)
);

OA21x2_ASAP7_75t_L g4419 ( 
.A1(n_4183),
.A2(n_4072),
.B(n_4071),
.Y(n_4419)
);

INVx5_ASAP7_75t_L g4420 ( 
.A(n_4307),
.Y(n_4420)
);

AOI21xp5_ASAP7_75t_L g4421 ( 
.A1(n_4371),
.A2(n_1202),
.B(n_1193),
.Y(n_4421)
);

INVx1_ASAP7_75t_L g4422 ( 
.A(n_4269),
.Y(n_4422)
);

O2A1O1Ixp33_ASAP7_75t_SL g4423 ( 
.A1(n_4232),
.A2(n_1212),
.B(n_1203),
.C(n_1537),
.Y(n_4423)
);

AOI21xp5_ASAP7_75t_L g4424 ( 
.A1(n_4233),
.A2(n_1212),
.B(n_1203),
.Y(n_4424)
);

NAND2xp5_ASAP7_75t_L g4425 ( 
.A(n_4239),
.B(n_1111),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4329),
.A2(n_1541),
.B(n_1539),
.Y(n_4426)
);

INVx3_ASAP7_75t_L g4427 ( 
.A(n_4159),
.Y(n_4427)
);

INVx1_ASAP7_75t_L g4428 ( 
.A(n_4270),
.Y(n_4428)
);

OAI22xp5_ASAP7_75t_L g4429 ( 
.A1(n_4316),
.A2(n_1167),
.B1(n_1111),
.B2(n_1003),
.Y(n_4429)
);

INVx2_ASAP7_75t_SL g4430 ( 
.A(n_4155),
.Y(n_4430)
);

OAI21x1_ASAP7_75t_L g4431 ( 
.A1(n_4186),
.A2(n_1326),
.B(n_1324),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4147),
.Y(n_4432)
);

AND2x4_ASAP7_75t_L g4433 ( 
.A(n_4240),
.B(n_1333),
.Y(n_4433)
);

INVxp67_ASAP7_75t_L g4434 ( 
.A(n_4182),
.Y(n_4434)
);

AND2x6_ASAP7_75t_SL g4435 ( 
.A(n_4195),
.B(n_1543),
.Y(n_4435)
);

BUFx3_ASAP7_75t_L g4436 ( 
.A(n_4151),
.Y(n_4436)
);

INVx1_ASAP7_75t_L g4437 ( 
.A(n_4162),
.Y(n_4437)
);

AO21x2_ASAP7_75t_L g4438 ( 
.A1(n_4315),
.A2(n_1336),
.B(n_1335),
.Y(n_4438)
);

INVx2_ASAP7_75t_L g4439 ( 
.A(n_4174),
.Y(n_4439)
);

AO31x2_ASAP7_75t_L g4440 ( 
.A1(n_4293),
.A2(n_1345),
.A3(n_1349),
.B(n_1344),
.Y(n_4440)
);

AOI21xp5_ASAP7_75t_L g4441 ( 
.A1(n_4272),
.A2(n_1547),
.B(n_1546),
.Y(n_4441)
);

AOI21xp5_ASAP7_75t_L g4442 ( 
.A1(n_4278),
.A2(n_1551),
.B(n_1550),
.Y(n_4442)
);

BUFx2_ASAP7_75t_L g4443 ( 
.A(n_4367),
.Y(n_4443)
);

A2O1A1Ixp33_ASAP7_75t_L g4444 ( 
.A1(n_4325),
.A2(n_1354),
.B(n_1355),
.C(n_1353),
.Y(n_4444)
);

NAND2xp5_ASAP7_75t_L g4445 ( 
.A(n_4230),
.B(n_1111),
.Y(n_4445)
);

AOI21xp5_ASAP7_75t_L g4446 ( 
.A1(n_4277),
.A2(n_1555),
.B(n_1552),
.Y(n_4446)
);

AOI21xp5_ASAP7_75t_L g4447 ( 
.A1(n_4225),
.A2(n_1559),
.B(n_1556),
.Y(n_4447)
);

OAI21x1_ASAP7_75t_L g4448 ( 
.A1(n_4317),
.A2(n_1357),
.B(n_1375),
.Y(n_4448)
);

OAI21x1_ASAP7_75t_L g4449 ( 
.A1(n_4248),
.A2(n_4157),
.B(n_4167),
.Y(n_4449)
);

INVx2_ASAP7_75t_L g4450 ( 
.A(n_4191),
.Y(n_4450)
);

AOI21xp5_ASAP7_75t_L g4451 ( 
.A1(n_4280),
.A2(n_4194),
.B(n_4261),
.Y(n_4451)
);

NAND3x1_ASAP7_75t_L g4452 ( 
.A(n_4212),
.B(n_1561),
.C(n_1560),
.Y(n_4452)
);

INVx3_ASAP7_75t_L g4453 ( 
.A(n_4159),
.Y(n_4453)
);

INVx2_ASAP7_75t_L g4454 ( 
.A(n_4198),
.Y(n_4454)
);

AO31x2_ASAP7_75t_L g4455 ( 
.A1(n_4293),
.A2(n_1411),
.A3(n_1416),
.B(n_1397),
.Y(n_4455)
);

OAI22x1_ASAP7_75t_L g4456 ( 
.A1(n_4152),
.A2(n_1005),
.B1(n_1010),
.B2(n_1001),
.Y(n_4456)
);

AOI21xp5_ASAP7_75t_L g4457 ( 
.A1(n_4261),
.A2(n_4218),
.B(n_4318),
.Y(n_4457)
);

AO32x2_ASAP7_75t_L g4458 ( 
.A1(n_4252),
.A2(n_1569),
.A3(n_1570),
.B1(n_1567),
.B2(n_1564),
.Y(n_4458)
);

OAI21xp5_ASAP7_75t_L g4459 ( 
.A1(n_4346),
.A2(n_1642),
.B(n_1576),
.Y(n_4459)
);

AOI21xp5_ASAP7_75t_L g4460 ( 
.A1(n_4378),
.A2(n_1577),
.B(n_1571),
.Y(n_4460)
);

OAI22xp5_ASAP7_75t_L g4461 ( 
.A1(n_4335),
.A2(n_1167),
.B1(n_1111),
.B2(n_1012),
.Y(n_4461)
);

AOI22xp5_ASAP7_75t_L g4462 ( 
.A1(n_4211),
.A2(n_1579),
.B1(n_1580),
.B2(n_1578),
.Y(n_4462)
);

O2A1O1Ixp33_ASAP7_75t_L g4463 ( 
.A1(n_4292),
.A2(n_4320),
.B(n_4286),
.C(n_4304),
.Y(n_4463)
);

AOI21xp5_ASAP7_75t_L g4464 ( 
.A1(n_4378),
.A2(n_1583),
.B(n_1582),
.Y(n_4464)
);

BUFx12f_ASAP7_75t_L g4465 ( 
.A(n_4289),
.Y(n_4465)
);

AOI21xp5_ASAP7_75t_L g4466 ( 
.A1(n_4168),
.A2(n_1589),
.B(n_1586),
.Y(n_4466)
);

INVx2_ASAP7_75t_L g4467 ( 
.A(n_4148),
.Y(n_4467)
);

INVx2_ASAP7_75t_L g4468 ( 
.A(n_4153),
.Y(n_4468)
);

AOI21xp5_ASAP7_75t_L g4469 ( 
.A1(n_4276),
.A2(n_1594),
.B(n_1593),
.Y(n_4469)
);

OA21x2_ASAP7_75t_L g4470 ( 
.A1(n_4226),
.A2(n_4145),
.B(n_4354),
.Y(n_4470)
);

AO31x2_ASAP7_75t_L g4471 ( 
.A1(n_4181),
.A2(n_1411),
.A3(n_1416),
.B(n_1397),
.Y(n_4471)
);

O2A1O1Ixp33_ASAP7_75t_SL g4472 ( 
.A1(n_4274),
.A2(n_1598),
.B(n_1600),
.C(n_1595),
.Y(n_4472)
);

INVx1_ASAP7_75t_L g4473 ( 
.A(n_4142),
.Y(n_4473)
);

AOI21xp5_ASAP7_75t_L g4474 ( 
.A1(n_4276),
.A2(n_1602),
.B(n_1601),
.Y(n_4474)
);

AOI21xp5_ASAP7_75t_L g4475 ( 
.A1(n_4287),
.A2(n_1604),
.B(n_1603),
.Y(n_4475)
);

BUFx12f_ASAP7_75t_L g4476 ( 
.A(n_4289),
.Y(n_4476)
);

OAI21xp5_ASAP7_75t_SL g4477 ( 
.A1(n_4373),
.A2(n_4231),
.B(n_4268),
.Y(n_4477)
);

CKINVDCx5p33_ASAP7_75t_R g4478 ( 
.A(n_4283),
.Y(n_4478)
);

AOI21xp5_ASAP7_75t_L g4479 ( 
.A1(n_4307),
.A2(n_1614),
.B(n_1613),
.Y(n_4479)
);

INVx1_ASAP7_75t_L g4480 ( 
.A(n_4158),
.Y(n_4480)
);

AOI21xp5_ASAP7_75t_L g4481 ( 
.A1(n_4281),
.A2(n_1616),
.B(n_1615),
.Y(n_4481)
);

AOI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_4373),
.A2(n_1635),
.B(n_1630),
.Y(n_4482)
);

NAND2xp5_ASAP7_75t_L g4483 ( 
.A(n_4247),
.B(n_1111),
.Y(n_4483)
);

INVx1_ASAP7_75t_L g4484 ( 
.A(n_4160),
.Y(n_4484)
);

INVx2_ASAP7_75t_L g4485 ( 
.A(n_4180),
.Y(n_4485)
);

O2A1O1Ixp5_ASAP7_75t_L g4486 ( 
.A1(n_4145),
.A2(n_1438),
.B(n_1447),
.C(n_1431),
.Y(n_4486)
);

AO32x2_ASAP7_75t_L g4487 ( 
.A1(n_4236),
.A2(n_1641),
.A3(n_1638),
.B1(n_1447),
.B2(n_1456),
.Y(n_4487)
);

INVx2_ASAP7_75t_SL g4488 ( 
.A(n_4175),
.Y(n_4488)
);

BUFx3_ASAP7_75t_L g4489 ( 
.A(n_4264),
.Y(n_4489)
);

AOI21xp5_ASAP7_75t_L g4490 ( 
.A1(n_4350),
.A2(n_4339),
.B(n_4366),
.Y(n_4490)
);

OAI22x1_ASAP7_75t_L g4491 ( 
.A1(n_4189),
.A2(n_1018),
.B1(n_1026),
.B2(n_1006),
.Y(n_4491)
);

OAI21xp5_ASAP7_75t_L g4492 ( 
.A1(n_4249),
.A2(n_1028),
.B(n_1024),
.Y(n_4492)
);

NAND2xp5_ASAP7_75t_L g4493 ( 
.A(n_4166),
.B(n_1111),
.Y(n_4493)
);

AOI21xp5_ASAP7_75t_L g4494 ( 
.A1(n_4310),
.A2(n_1167),
.B(n_1035),
.Y(n_4494)
);

BUFx8_ASAP7_75t_L g4495 ( 
.A(n_4312),
.Y(n_4495)
);

HB1xp67_ASAP7_75t_L g4496 ( 
.A(n_4185),
.Y(n_4496)
);

AO21x2_ASAP7_75t_L g4497 ( 
.A1(n_4338),
.A2(n_4323),
.B(n_4334),
.Y(n_4497)
);

NAND2xp5_ASAP7_75t_L g4498 ( 
.A(n_4223),
.B(n_1167),
.Y(n_4498)
);

AO31x2_ASAP7_75t_L g4499 ( 
.A1(n_4300),
.A2(n_1431),
.A3(n_1456),
.B(n_1438),
.Y(n_4499)
);

INVx3_ASAP7_75t_SL g4500 ( 
.A(n_4295),
.Y(n_4500)
);

AO31x2_ASAP7_75t_L g4501 ( 
.A1(n_4265),
.A2(n_1466),
.A3(n_1470),
.B(n_1467),
.Y(n_4501)
);

NOR2xp33_ASAP7_75t_L g4502 ( 
.A(n_4266),
.B(n_8),
.Y(n_4502)
);

NAND2xp5_ASAP7_75t_L g4503 ( 
.A(n_4246),
.B(n_1167),
.Y(n_4503)
);

NOR2xp33_ASAP7_75t_L g4504 ( 
.A(n_4177),
.B(n_8),
.Y(n_4504)
);

INVxp67_ASAP7_75t_SL g4505 ( 
.A(n_4299),
.Y(n_4505)
);

A2O1A1Ixp33_ASAP7_75t_L g4506 ( 
.A1(n_4327),
.A2(n_1036),
.B(n_1038),
.C(n_1031),
.Y(n_4506)
);

AO31x2_ASAP7_75t_L g4507 ( 
.A1(n_4355),
.A2(n_1466),
.A3(n_1470),
.B(n_1467),
.Y(n_4507)
);

AOI21xp5_ASAP7_75t_L g4508 ( 
.A1(n_4302),
.A2(n_1167),
.B(n_1054),
.Y(n_4508)
);

BUFx6f_ASAP7_75t_L g4509 ( 
.A(n_4244),
.Y(n_4509)
);

O2A1O1Ixp5_ASAP7_75t_L g4510 ( 
.A1(n_4208),
.A2(n_1500),
.B(n_1545),
.C(n_1487),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_L g4511 ( 
.A(n_4214),
.B(n_9),
.Y(n_4511)
);

AOI21xp5_ASAP7_75t_L g4512 ( 
.A1(n_4305),
.A2(n_1057),
.B(n_1052),
.Y(n_4512)
);

O2A1O1Ixp33_ASAP7_75t_L g4513 ( 
.A1(n_4161),
.A2(n_1500),
.B(n_1545),
.C(n_1487),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4219),
.B(n_10),
.Y(n_4514)
);

A2O1A1Ixp33_ASAP7_75t_L g4515 ( 
.A1(n_4188),
.A2(n_1059),
.B(n_1060),
.C(n_1058),
.Y(n_4515)
);

OR2x6_ASAP7_75t_L g4516 ( 
.A(n_4172),
.B(n_1566),
.Y(n_4516)
);

INVx1_ASAP7_75t_L g4517 ( 
.A(n_4184),
.Y(n_4517)
);

NOR2xp33_ASAP7_75t_L g4518 ( 
.A(n_4177),
.B(n_11),
.Y(n_4518)
);

OAI22xp5_ASAP7_75t_L g4519 ( 
.A1(n_4340),
.A2(n_1064),
.B1(n_1065),
.B2(n_1062),
.Y(n_4519)
);

OAI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4288),
.A2(n_4253),
.B1(n_4353),
.B2(n_4285),
.Y(n_4520)
);

INVxp67_ASAP7_75t_SL g4521 ( 
.A(n_4299),
.Y(n_4521)
);

NOR2xp67_ASAP7_75t_L g4522 ( 
.A(n_4242),
.B(n_1566),
.Y(n_4522)
);

AOI21xp5_ASAP7_75t_L g4523 ( 
.A1(n_4359),
.A2(n_1068),
.B(n_1067),
.Y(n_4523)
);

INVx1_ASAP7_75t_L g4524 ( 
.A(n_4200),
.Y(n_4524)
);

NAND2xp33_ASAP7_75t_L g4525 ( 
.A(n_4380),
.B(n_1069),
.Y(n_4525)
);

BUFx3_ASAP7_75t_L g4526 ( 
.A(n_4367),
.Y(n_4526)
);

AOI21xp5_ASAP7_75t_L g4527 ( 
.A1(n_4349),
.A2(n_1072),
.B(n_1071),
.Y(n_4527)
);

NAND2xp5_ASAP7_75t_L g4528 ( 
.A(n_4260),
.B(n_12),
.Y(n_4528)
);

INVx1_ASAP7_75t_L g4529 ( 
.A(n_4207),
.Y(n_4529)
);

NAND2xp5_ASAP7_75t_L g4530 ( 
.A(n_4217),
.B(n_12),
.Y(n_4530)
);

NAND2xp5_ASAP7_75t_SL g4531 ( 
.A(n_4322),
.B(n_1573),
.Y(n_4531)
);

OAI21x1_ASAP7_75t_L g4532 ( 
.A1(n_4352),
.A2(n_1607),
.B(n_1573),
.Y(n_4532)
);

NAND2xp5_ASAP7_75t_L g4533 ( 
.A(n_4220),
.B(n_13),
.Y(n_4533)
);

O2A1O1Ixp33_ASAP7_75t_L g4534 ( 
.A1(n_4224),
.A2(n_1610),
.B(n_1607),
.C(n_1628),
.Y(n_4534)
);

OAI21x1_ASAP7_75t_L g4535 ( 
.A1(n_4351),
.A2(n_1610),
.B(n_1628),
.Y(n_4535)
);

NAND2xp5_ASAP7_75t_L g4536 ( 
.A(n_4170),
.B(n_13),
.Y(n_4536)
);

INVx1_ASAP7_75t_L g4537 ( 
.A(n_4203),
.Y(n_4537)
);

AOI221x1_ASAP7_75t_L g4538 ( 
.A1(n_4251),
.A2(n_2074),
.B1(n_2085),
.B2(n_2072),
.C(n_2060),
.Y(n_4538)
);

INVx1_ASAP7_75t_L g4539 ( 
.A(n_4341),
.Y(n_4539)
);

AOI21xp5_ASAP7_75t_L g4540 ( 
.A1(n_4294),
.A2(n_1076),
.B(n_1075),
.Y(n_4540)
);

AO31x2_ASAP7_75t_L g4541 ( 
.A1(n_4291),
.A2(n_2072),
.A3(n_2074),
.B(n_2060),
.Y(n_4541)
);

A2O1A1Ixp33_ASAP7_75t_L g4542 ( 
.A1(n_4332),
.A2(n_1078),
.B(n_1081),
.C(n_1079),
.Y(n_4542)
);

NOR2xp33_ASAP7_75t_L g4543 ( 
.A(n_4222),
.B(n_14),
.Y(n_4543)
);

OAI21x1_ASAP7_75t_L g4544 ( 
.A1(n_4347),
.A2(n_2074),
.B(n_2072),
.Y(n_4544)
);

AOI21xp5_ASAP7_75t_L g4545 ( 
.A1(n_4298),
.A2(n_1087),
.B(n_1074),
.Y(n_4545)
);

NAND2xp5_ASAP7_75t_L g4546 ( 
.A(n_4210),
.B(n_15),
.Y(n_4546)
);

NAND2x1p5_ASAP7_75t_L g4547 ( 
.A(n_4196),
.B(n_4199),
.Y(n_4547)
);

INVxp67_ASAP7_75t_SL g4548 ( 
.A(n_4313),
.Y(n_4548)
);

AOI21x1_ASAP7_75t_L g4549 ( 
.A1(n_4387),
.A2(n_1088),
.B(n_1085),
.Y(n_4549)
);

OAI21x1_ASAP7_75t_L g4550 ( 
.A1(n_4308),
.A2(n_4309),
.B(n_4326),
.Y(n_4550)
);

OAI21x1_ASAP7_75t_L g4551 ( 
.A1(n_4216),
.A2(n_2074),
.B(n_2072),
.Y(n_4551)
);

INVx1_ASAP7_75t_L g4552 ( 
.A(n_4229),
.Y(n_4552)
);

AO31x2_ASAP7_75t_L g4553 ( 
.A1(n_4336),
.A2(n_1090),
.A3(n_1091),
.B(n_1089),
.Y(n_4553)
);

INVx3_ASAP7_75t_L g4554 ( 
.A(n_4222),
.Y(n_4554)
);

O2A1O1Ixp33_ASAP7_75t_SL g4555 ( 
.A1(n_4372),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_4555)
);

AOI21x1_ASAP7_75t_L g4556 ( 
.A1(n_4364),
.A2(n_1094),
.B(n_1093),
.Y(n_4556)
);

AO31x2_ASAP7_75t_L g4557 ( 
.A1(n_4363),
.A2(n_1100),
.A3(n_1113),
.B(n_1099),
.Y(n_4557)
);

CKINVDCx5p33_ASAP7_75t_R g4558 ( 
.A(n_4254),
.Y(n_4558)
);

INVx2_ASAP7_75t_L g4559 ( 
.A(n_4306),
.Y(n_4559)
);

INVx2_ASAP7_75t_L g4560 ( 
.A(n_4331),
.Y(n_4560)
);

A2O1A1Ixp33_ASAP7_75t_L g4561 ( 
.A1(n_4333),
.A2(n_1116),
.B(n_1118),
.C(n_1115),
.Y(n_4561)
);

O2A1O1Ixp33_ASAP7_75t_L g4562 ( 
.A1(n_4377),
.A2(n_1119),
.B(n_1125),
.C(n_1117),
.Y(n_4562)
);

O2A1O1Ixp33_ASAP7_75t_SL g4563 ( 
.A1(n_4297),
.A2(n_18),
.B(n_16),
.C(n_17),
.Y(n_4563)
);

O2A1O1Ixp33_ASAP7_75t_L g4564 ( 
.A1(n_4382),
.A2(n_1207),
.B(n_1208),
.C(n_1206),
.Y(n_4564)
);

OR2x6_ASAP7_75t_L g4565 ( 
.A(n_4172),
.B(n_2085),
.Y(n_4565)
);

OAI21xp5_ASAP7_75t_L g4566 ( 
.A1(n_4344),
.A2(n_1134),
.B(n_1133),
.Y(n_4566)
);

BUFx6f_ASAP7_75t_L g4567 ( 
.A(n_4244),
.Y(n_4567)
);

AOI21xp5_ASAP7_75t_L g4568 ( 
.A1(n_4275),
.A2(n_1137),
.B(n_1136),
.Y(n_4568)
);

AOI22xp33_ASAP7_75t_L g4569 ( 
.A1(n_4190),
.A2(n_1140),
.B1(n_1141),
.B2(n_1138),
.Y(n_4569)
);

AOI21xp5_ASAP7_75t_L g4570 ( 
.A1(n_4199),
.A2(n_1145),
.B(n_1142),
.Y(n_4570)
);

INVx1_ASAP7_75t_L g4571 ( 
.A(n_4330),
.Y(n_4571)
);

AOI21xp5_ASAP7_75t_L g4572 ( 
.A1(n_4199),
.A2(n_1147),
.B(n_1146),
.Y(n_4572)
);

AND2x2_ASAP7_75t_L g4573 ( 
.A(n_4240),
.B(n_20),
.Y(n_4573)
);

INVx1_ASAP7_75t_L g4574 ( 
.A(n_4221),
.Y(n_4574)
);

INVx1_ASAP7_75t_SL g4575 ( 
.A(n_4370),
.Y(n_4575)
);

HB1xp67_ASAP7_75t_L g4576 ( 
.A(n_4271),
.Y(n_4576)
);

O2A1O1Ixp5_ASAP7_75t_SL g4577 ( 
.A1(n_4245),
.A2(n_1149),
.B(n_1153),
.C(n_1148),
.Y(n_4577)
);

AO31x2_ASAP7_75t_L g4578 ( 
.A1(n_4273),
.A2(n_2088),
.A3(n_2092),
.B(n_2085),
.Y(n_4578)
);

NAND2xp5_ASAP7_75t_L g4579 ( 
.A(n_4213),
.B(n_20),
.Y(n_4579)
);

AOI221xp5_ASAP7_75t_L g4580 ( 
.A1(n_4324),
.A2(n_1160),
.B1(n_1161),
.B2(n_1159),
.C(n_1156),
.Y(n_4580)
);

AO31x2_ASAP7_75t_L g4581 ( 
.A1(n_4215),
.A2(n_4235),
.A3(n_4241),
.B(n_4238),
.Y(n_4581)
);

OA21x2_ASAP7_75t_L g4582 ( 
.A1(n_4365),
.A2(n_1163),
.B(n_1162),
.Y(n_4582)
);

AOI22xp33_ASAP7_75t_L g4583 ( 
.A1(n_4192),
.A2(n_1165),
.B1(n_1166),
.B2(n_1164),
.Y(n_4583)
);

A2O1A1Ixp33_ASAP7_75t_L g4584 ( 
.A1(n_4374),
.A2(n_1172),
.B(n_1173),
.C(n_1171),
.Y(n_4584)
);

OA21x2_ASAP7_75t_L g4585 ( 
.A1(n_4296),
.A2(n_1180),
.B(n_1175),
.Y(n_4585)
);

BUFx3_ASAP7_75t_L g4586 ( 
.A(n_4250),
.Y(n_4586)
);

OAI22xp5_ASAP7_75t_L g4587 ( 
.A1(n_4358),
.A2(n_1184),
.B1(n_1189),
.B2(n_1181),
.Y(n_4587)
);

AOI21xp5_ASAP7_75t_L g4588 ( 
.A1(n_4290),
.A2(n_1191),
.B(n_1190),
.Y(n_4588)
);

INVx2_ASAP7_75t_L g4589 ( 
.A(n_4209),
.Y(n_4589)
);

AOI21xp5_ASAP7_75t_L g4590 ( 
.A1(n_4290),
.A2(n_1195),
.B(n_1194),
.Y(n_4590)
);

NOR2x1_ASAP7_75t_SL g4591 ( 
.A(n_4234),
.B(n_2085),
.Y(n_4591)
);

INVx1_ASAP7_75t_L g4592 ( 
.A(n_4209),
.Y(n_4592)
);

OAI21xp5_ASAP7_75t_L g4593 ( 
.A1(n_4384),
.A2(n_1199),
.B(n_1197),
.Y(n_4593)
);

OAI21x1_ASAP7_75t_L g4594 ( 
.A1(n_4375),
.A2(n_2092),
.B(n_2088),
.Y(n_4594)
);

AO22x2_ASAP7_75t_L g4595 ( 
.A1(n_4243),
.A2(n_24),
.B1(n_21),
.B2(n_22),
.Y(n_4595)
);

A2O1A1Ixp33_ASAP7_75t_L g4596 ( 
.A1(n_4360),
.A2(n_1210),
.B(n_1216),
.C(n_1215),
.Y(n_4596)
);

NAND2x1p5_ASAP7_75t_L g4597 ( 
.A(n_4234),
.B(n_2088),
.Y(n_4597)
);

AOI21xp33_ASAP7_75t_L g4598 ( 
.A1(n_4361),
.A2(n_1209),
.B(n_21),
.Y(n_4598)
);

OAI21x1_ASAP7_75t_L g4599 ( 
.A1(n_4379),
.A2(n_2092),
.B(n_2088),
.Y(n_4599)
);

A2O1A1Ixp33_ASAP7_75t_L g4600 ( 
.A1(n_4178),
.A2(n_28),
.B(n_25),
.C(n_27),
.Y(n_4600)
);

INVx2_ASAP7_75t_L g4601 ( 
.A(n_4227),
.Y(n_4601)
);

NOR2xp67_ASAP7_75t_L g4602 ( 
.A(n_4388),
.B(n_25),
.Y(n_4602)
);

HB1xp67_ASAP7_75t_L g4603 ( 
.A(n_4227),
.Y(n_4603)
);

INVx2_ASAP7_75t_L g4604 ( 
.A(n_4178),
.Y(n_4604)
);

NAND2xp5_ASAP7_75t_L g4605 ( 
.A(n_4342),
.B(n_30),
.Y(n_4605)
);

BUFx3_ASAP7_75t_L g4606 ( 
.A(n_4244),
.Y(n_4606)
);

AOI21xp5_ASAP7_75t_L g4607 ( 
.A1(n_4357),
.A2(n_2095),
.B(n_2092),
.Y(n_4607)
);

AOI211x1_ASAP7_75t_L g4608 ( 
.A1(n_4345),
.A2(n_32),
.B(n_30),
.C(n_31),
.Y(n_4608)
);

AOI21xp5_ASAP7_75t_L g4609 ( 
.A1(n_4388),
.A2(n_2104),
.B(n_2095),
.Y(n_4609)
);

A2O1A1Ixp33_ASAP7_75t_L g4610 ( 
.A1(n_4368),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_4610)
);

INVx2_ASAP7_75t_SL g4611 ( 
.A(n_4376),
.Y(n_4611)
);

NAND2xp5_ASAP7_75t_L g4612 ( 
.A(n_4369),
.B(n_37),
.Y(n_4612)
);

INVx1_ASAP7_75t_L g4613 ( 
.A(n_4245),
.Y(n_4613)
);

AND2x4_ASAP7_75t_L g4614 ( 
.A(n_4154),
.B(n_37),
.Y(n_4614)
);

OA21x2_ASAP7_75t_L g4615 ( 
.A1(n_4314),
.A2(n_38),
.B(n_39),
.Y(n_4615)
);

INVx1_ASAP7_75t_L g4616 ( 
.A(n_4255),
.Y(n_4616)
);

OAI21x1_ASAP7_75t_L g4617 ( 
.A1(n_4319),
.A2(n_2104),
.B(n_2095),
.Y(n_4617)
);

INVxp67_ASAP7_75t_SL g4618 ( 
.A(n_4154),
.Y(n_4618)
);

AND2x2_ASAP7_75t_L g4619 ( 
.A(n_4156),
.B(n_39),
.Y(n_4619)
);

INVx2_ASAP7_75t_SL g4620 ( 
.A(n_4381),
.Y(n_4620)
);

NAND3xp33_ASAP7_75t_L g4621 ( 
.A(n_4303),
.B(n_2104),
.C(n_2095),
.Y(n_4621)
);

BUFx3_ASAP7_75t_L g4622 ( 
.A(n_4263),
.Y(n_4622)
);

AND3x2_ASAP7_75t_L g4623 ( 
.A(n_4314),
.B(n_40),
.C(n_43),
.Y(n_4623)
);

OAI21xp33_ASAP7_75t_L g4624 ( 
.A1(n_4385),
.A2(n_40),
.B(n_43),
.Y(n_4624)
);

INVxp67_ASAP7_75t_L g4625 ( 
.A(n_4343),
.Y(n_4625)
);

AO31x2_ASAP7_75t_L g4626 ( 
.A1(n_4301),
.A2(n_46),
.A3(n_44),
.B(n_45),
.Y(n_4626)
);

NOR2xp33_ASAP7_75t_SL g4627 ( 
.A(n_4173),
.B(n_2104),
.Y(n_4627)
);

AO31x2_ASAP7_75t_L g4628 ( 
.A1(n_4301),
.A2(n_46),
.A3(n_44),
.B(n_45),
.Y(n_4628)
);

AOI21xp5_ASAP7_75t_L g4629 ( 
.A1(n_4389),
.A2(n_2126),
.B(n_47),
.Y(n_4629)
);

OAI21x1_ASAP7_75t_L g4630 ( 
.A1(n_4255),
.A2(n_2126),
.B(n_649),
.Y(n_4630)
);

INVx1_ASAP7_75t_L g4631 ( 
.A(n_4156),
.Y(n_4631)
);

NOR2xp33_ASAP7_75t_L g4632 ( 
.A(n_4179),
.B(n_49),
.Y(n_4632)
);

AND2x2_ASAP7_75t_L g4633 ( 
.A(n_4204),
.B(n_4228),
.Y(n_4633)
);

AO31x2_ASAP7_75t_L g4634 ( 
.A1(n_4348),
.A2(n_2126),
.A3(n_52),
.B(n_50),
.Y(n_4634)
);

NOR2xp67_ASAP7_75t_L g4635 ( 
.A(n_4399),
.B(n_4237),
.Y(n_4635)
);

AO21x2_ASAP7_75t_L g4636 ( 
.A1(n_4503),
.A2(n_4356),
.B(n_4348),
.Y(n_4636)
);

OAI21x1_ASAP7_75t_SL g4637 ( 
.A1(n_4490),
.A2(n_4383),
.B(n_4380),
.Y(n_4637)
);

CKINVDCx16_ASAP7_75t_R g4638 ( 
.A(n_4489),
.Y(n_4638)
);

CKINVDCx5p33_ASAP7_75t_R g4639 ( 
.A(n_4465),
.Y(n_4639)
);

AOI22xp33_ASAP7_75t_L g4640 ( 
.A1(n_4585),
.A2(n_4356),
.B1(n_4328),
.B2(n_4263),
.Y(n_4640)
);

CKINVDCx5p33_ASAP7_75t_R g4641 ( 
.A(n_4476),
.Y(n_4641)
);

INVx1_ASAP7_75t_L g4642 ( 
.A(n_4395),
.Y(n_4642)
);

INVx2_ASAP7_75t_SL g4643 ( 
.A(n_4436),
.Y(n_4643)
);

OA21x2_ASAP7_75t_L g4644 ( 
.A1(n_4449),
.A2(n_4328),
.B(n_4263),
.Y(n_4644)
);

OAI22xp5_ASAP7_75t_L g4645 ( 
.A1(n_4569),
.A2(n_4389),
.B1(n_4383),
.B2(n_4380),
.Y(n_4645)
);

INVx1_ASAP7_75t_L g4646 ( 
.A(n_4414),
.Y(n_4646)
);

OAI21x1_ASAP7_75t_L g4647 ( 
.A1(n_4451),
.A2(n_4383),
.B(n_4362),
.Y(n_4647)
);

AOI21xp5_ASAP7_75t_L g4648 ( 
.A1(n_4457),
.A2(n_4386),
.B(n_4303),
.Y(n_4648)
);

INVx6_ASAP7_75t_L g4649 ( 
.A(n_4495),
.Y(n_4649)
);

HB1xp67_ASAP7_75t_L g4650 ( 
.A(n_4496),
.Y(n_4650)
);

INVx2_ASAP7_75t_L g4651 ( 
.A(n_4571),
.Y(n_4651)
);

HB1xp67_ASAP7_75t_L g4652 ( 
.A(n_4393),
.Y(n_4652)
);

NAND2xp5_ASAP7_75t_L g4653 ( 
.A(n_4437),
.B(n_4303),
.Y(n_4653)
);

INVx1_ASAP7_75t_L g4654 ( 
.A(n_4422),
.Y(n_4654)
);

INVx1_ASAP7_75t_L g4655 ( 
.A(n_4428),
.Y(n_4655)
);

INVx1_ASAP7_75t_L g4656 ( 
.A(n_4480),
.Y(n_4656)
);

INVx1_ASAP7_75t_L g4657 ( 
.A(n_4484),
.Y(n_4657)
);

AOI22xp33_ASAP7_75t_SL g4658 ( 
.A1(n_4585),
.A2(n_4284),
.B1(n_4362),
.B2(n_4343),
.Y(n_4658)
);

BUFx6f_ASAP7_75t_L g4659 ( 
.A(n_4399),
.Y(n_4659)
);

AO21x2_ASAP7_75t_L g4660 ( 
.A1(n_4445),
.A2(n_4362),
.B(n_4343),
.Y(n_4660)
);

AND2x4_ASAP7_75t_L g4661 ( 
.A(n_4603),
.B(n_4618),
.Y(n_4661)
);

OAI21x1_ASAP7_75t_L g4662 ( 
.A1(n_4551),
.A2(n_4284),
.B(n_4386),
.Y(n_4662)
);

OAI21x1_ASAP7_75t_L g4663 ( 
.A1(n_4544),
.A2(n_4599),
.B(n_4594),
.Y(n_4663)
);

INVx4_ASAP7_75t_L g4664 ( 
.A(n_4526),
.Y(n_4664)
);

CKINVDCx5p33_ASAP7_75t_R g4665 ( 
.A(n_4478),
.Y(n_4665)
);

OAI21x1_ASAP7_75t_L g4666 ( 
.A1(n_4417),
.A2(n_4284),
.B(n_51),
.Y(n_4666)
);

AOI221xp5_ASAP7_75t_L g4667 ( 
.A1(n_4595),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.C(n_54),
.Y(n_4667)
);

CKINVDCx5p33_ASAP7_75t_R g4668 ( 
.A(n_4558),
.Y(n_4668)
);

BUFx3_ASAP7_75t_L g4669 ( 
.A(n_4443),
.Y(n_4669)
);

OAI21xp5_ASAP7_75t_L g4670 ( 
.A1(n_4515),
.A2(n_53),
.B(n_55),
.Y(n_4670)
);

INVx1_ASAP7_75t_L g4671 ( 
.A(n_4517),
.Y(n_4671)
);

AO21x2_ASAP7_75t_L g4672 ( 
.A1(n_4498),
.A2(n_55),
.B(n_56),
.Y(n_4672)
);

INVxp67_ASAP7_75t_L g4673 ( 
.A(n_4406),
.Y(n_4673)
);

AOI221xp5_ASAP7_75t_L g4674 ( 
.A1(n_4595),
.A2(n_59),
.B1(n_56),
.B2(n_57),
.C(n_60),
.Y(n_4674)
);

INVx1_ASAP7_75t_L g4675 ( 
.A(n_4524),
.Y(n_4675)
);

INVx1_ASAP7_75t_L g4676 ( 
.A(n_4539),
.Y(n_4676)
);

INVx2_ASAP7_75t_L g4677 ( 
.A(n_4550),
.Y(n_4677)
);

INVx3_ASAP7_75t_L g4678 ( 
.A(n_4399),
.Y(n_4678)
);

OR2x6_ASAP7_75t_L g4679 ( 
.A(n_4547),
.B(n_2126),
.Y(n_4679)
);

INVx1_ASAP7_75t_L g4680 ( 
.A(n_4574),
.Y(n_4680)
);

INVx2_ASAP7_75t_L g4681 ( 
.A(n_4559),
.Y(n_4681)
);

INVx1_ASAP7_75t_L g4682 ( 
.A(n_4505),
.Y(n_4682)
);

AND2x4_ASAP7_75t_L g4683 ( 
.A(n_4552),
.B(n_61),
.Y(n_4683)
);

BUFx10_ASAP7_75t_L g4684 ( 
.A(n_4416),
.Y(n_4684)
);

INVx2_ASAP7_75t_L g4685 ( 
.A(n_4467),
.Y(n_4685)
);

OAI21x1_ASAP7_75t_L g4686 ( 
.A1(n_4609),
.A2(n_61),
.B(n_62),
.Y(n_4686)
);

AOI21xp5_ASAP7_75t_L g4687 ( 
.A1(n_4398),
.A2(n_63),
.B(n_64),
.Y(n_4687)
);

OAI21xp5_ASAP7_75t_L g4688 ( 
.A1(n_4421),
.A2(n_65),
.B(n_66),
.Y(n_4688)
);

BUFx12f_ASAP7_75t_L g4689 ( 
.A(n_4435),
.Y(n_4689)
);

NAND2xp5_ASAP7_75t_L g4690 ( 
.A(n_4411),
.B(n_65),
.Y(n_4690)
);

CKINVDCx12_ASAP7_75t_R g4691 ( 
.A(n_4516),
.Y(n_4691)
);

OA21x2_ASAP7_75t_L g4692 ( 
.A1(n_4521),
.A2(n_66),
.B(n_67),
.Y(n_4692)
);

OR2x2_ASAP7_75t_L g4693 ( 
.A(n_4488),
.B(n_67),
.Y(n_4693)
);

AOI22xp33_ASAP7_75t_L g4694 ( 
.A1(n_4582),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_4694)
);

NAND2xp5_ASAP7_75t_L g4695 ( 
.A(n_4473),
.B(n_68),
.Y(n_4695)
);

NAND2xp5_ASAP7_75t_L g4696 ( 
.A(n_4430),
.B(n_69),
.Y(n_4696)
);

OAI21x1_ASAP7_75t_SL g4697 ( 
.A1(n_4520),
.A2(n_70),
.B(n_72),
.Y(n_4697)
);

AND2x2_ASAP7_75t_L g4698 ( 
.A(n_4575),
.B(n_72),
.Y(n_4698)
);

INVx2_ASAP7_75t_L g4699 ( 
.A(n_4468),
.Y(n_4699)
);

INVx2_ASAP7_75t_L g4700 ( 
.A(n_4485),
.Y(n_4700)
);

OAI21x1_ASAP7_75t_L g4701 ( 
.A1(n_4448),
.A2(n_73),
.B(n_75),
.Y(n_4701)
);

OAI21x1_ASAP7_75t_L g4702 ( 
.A1(n_4403),
.A2(n_77),
.B(n_79),
.Y(n_4702)
);

OAI21x1_ASAP7_75t_L g4703 ( 
.A1(n_4431),
.A2(n_77),
.B(n_79),
.Y(n_4703)
);

OA21x2_ASAP7_75t_L g4704 ( 
.A1(n_4548),
.A2(n_80),
.B(n_81),
.Y(n_4704)
);

AND2x2_ASAP7_75t_L g4705 ( 
.A(n_4611),
.B(n_80),
.Y(n_4705)
);

AOI22xp5_ASAP7_75t_L g4706 ( 
.A1(n_4624),
.A2(n_83),
.B1(n_81),
.B2(n_82),
.Y(n_4706)
);

OAI21x1_ASAP7_75t_L g4707 ( 
.A1(n_4401),
.A2(n_82),
.B(n_83),
.Y(n_4707)
);

BUFx3_ASAP7_75t_L g4708 ( 
.A(n_4404),
.Y(n_4708)
);

NAND2xp5_ASAP7_75t_L g4709 ( 
.A(n_4537),
.B(n_85),
.Y(n_4709)
);

OAI21x1_ASAP7_75t_L g4710 ( 
.A1(n_4412),
.A2(n_85),
.B(n_86),
.Y(n_4710)
);

NOR2xp33_ASAP7_75t_L g4711 ( 
.A(n_4500),
.B(n_4390),
.Y(n_4711)
);

OAI22xp5_ASAP7_75t_L g4712 ( 
.A1(n_4477),
.A2(n_88),
.B1(n_86),
.B2(n_87),
.Y(n_4712)
);

INVx2_ASAP7_75t_L g4713 ( 
.A(n_4560),
.Y(n_4713)
);

INVx2_ASAP7_75t_L g4714 ( 
.A(n_4396),
.Y(n_4714)
);

CKINVDCx6p67_ASAP7_75t_R g4715 ( 
.A(n_4408),
.Y(n_4715)
);

OAI22xp5_ASAP7_75t_L g4716 ( 
.A1(n_4600),
.A2(n_92),
.B1(n_87),
.B2(n_89),
.Y(n_4716)
);

OAI21x1_ASAP7_75t_L g4717 ( 
.A1(n_4535),
.A2(n_93),
.B(n_94),
.Y(n_4717)
);

OAI21x1_ASAP7_75t_L g4718 ( 
.A1(n_4607),
.A2(n_93),
.B(n_95),
.Y(n_4718)
);

BUFx3_ASAP7_75t_L g4719 ( 
.A(n_4620),
.Y(n_4719)
);

AOI21xp5_ASAP7_75t_L g4720 ( 
.A1(n_4400),
.A2(n_4472),
.B(n_4423),
.Y(n_4720)
);

NOR2xp33_ASAP7_75t_L g4721 ( 
.A(n_4413),
.B(n_95),
.Y(n_4721)
);

OAI21xp5_ASAP7_75t_L g4722 ( 
.A1(n_4452),
.A2(n_96),
.B(n_98),
.Y(n_4722)
);

OAI21x1_ASAP7_75t_L g4723 ( 
.A1(n_4493),
.A2(n_96),
.B(n_100),
.Y(n_4723)
);

INVx1_ASAP7_75t_L g4724 ( 
.A(n_4576),
.Y(n_4724)
);

INVx2_ASAP7_75t_L g4725 ( 
.A(n_4439),
.Y(n_4725)
);

NAND2xp5_ASAP7_75t_L g4726 ( 
.A(n_4397),
.B(n_101),
.Y(n_4726)
);

NAND2xp5_ASAP7_75t_L g4727 ( 
.A(n_4425),
.B(n_101),
.Y(n_4727)
);

BUFx5_ASAP7_75t_L g4728 ( 
.A(n_4433),
.Y(n_4728)
);

AND2x2_ASAP7_75t_L g4729 ( 
.A(n_4613),
.B(n_102),
.Y(n_4729)
);

OAI21x1_ASAP7_75t_L g4730 ( 
.A1(n_4617),
.A2(n_103),
.B(n_104),
.Y(n_4730)
);

OA21x2_ASAP7_75t_L g4731 ( 
.A1(n_4483),
.A2(n_103),
.B(n_105),
.Y(n_4731)
);

INVx1_ASAP7_75t_L g4732 ( 
.A(n_4470),
.Y(n_4732)
);

INVx1_ASAP7_75t_SL g4733 ( 
.A(n_4633),
.Y(n_4733)
);

OAI21x1_ASAP7_75t_L g4734 ( 
.A1(n_4415),
.A2(n_105),
.B(n_106),
.Y(n_4734)
);

OAI21x1_ASAP7_75t_L g4735 ( 
.A1(n_4630),
.A2(n_107),
.B(n_108),
.Y(n_4735)
);

INVx2_ASAP7_75t_L g4736 ( 
.A(n_4450),
.Y(n_4736)
);

INVx2_ASAP7_75t_L g4737 ( 
.A(n_4454),
.Y(n_4737)
);

AO31x2_ASAP7_75t_L g4738 ( 
.A1(n_4538),
.A2(n_111),
.A3(n_108),
.B(n_109),
.Y(n_4738)
);

OAI21x1_ASAP7_75t_SL g4739 ( 
.A1(n_4591),
.A2(n_112),
.B(n_114),
.Y(n_4739)
);

OAI21x1_ASAP7_75t_SL g4740 ( 
.A1(n_4612),
.A2(n_114),
.B(n_116),
.Y(n_4740)
);

INVx1_ASAP7_75t_L g4741 ( 
.A(n_4470),
.Y(n_4741)
);

BUFx2_ASAP7_75t_L g4742 ( 
.A(n_4616),
.Y(n_4742)
);

NOR2x1_ASAP7_75t_SL g4743 ( 
.A(n_4420),
.B(n_117),
.Y(n_4743)
);

AOI221xp5_ASAP7_75t_L g4744 ( 
.A1(n_4608),
.A2(n_4555),
.B1(n_4409),
.B2(n_4598),
.C(n_4563),
.Y(n_4744)
);

OAI21x1_ASAP7_75t_L g4745 ( 
.A1(n_4486),
.A2(n_117),
.B(n_118),
.Y(n_4745)
);

OAI21x1_ASAP7_75t_L g4746 ( 
.A1(n_4494),
.A2(n_4442),
.B(n_4615),
.Y(n_4746)
);

INVx1_ASAP7_75t_L g4747 ( 
.A(n_4432),
.Y(n_4747)
);

AND2x4_ASAP7_75t_L g4748 ( 
.A(n_4631),
.B(n_119),
.Y(n_4748)
);

AOI22xp33_ASAP7_75t_L g4749 ( 
.A1(n_4582),
.A2(n_121),
.B1(n_119),
.B2(n_120),
.Y(n_4749)
);

AOI21xp33_ASAP7_75t_L g4750 ( 
.A1(n_4615),
.A2(n_120),
.B(n_121),
.Y(n_4750)
);

INVx2_ASAP7_75t_L g4751 ( 
.A(n_4581),
.Y(n_4751)
);

AND2x4_ASAP7_75t_L g4752 ( 
.A(n_4592),
.B(n_122),
.Y(n_4752)
);

INVx2_ASAP7_75t_L g4753 ( 
.A(n_4581),
.Y(n_4753)
);

NAND2x1p5_ASAP7_75t_L g4754 ( 
.A(n_4420),
.B(n_122),
.Y(n_4754)
);

INVx1_ASAP7_75t_L g4755 ( 
.A(n_4529),
.Y(n_4755)
);

A2O1A1Ixp33_ASAP7_75t_L g4756 ( 
.A1(n_4588),
.A2(n_127),
.B(n_124),
.C(n_125),
.Y(n_4756)
);

BUFx16f_ASAP7_75t_R g4757 ( 
.A(n_4614),
.Y(n_4757)
);

INVx2_ASAP7_75t_L g4758 ( 
.A(n_4581),
.Y(n_4758)
);

INVx2_ASAP7_75t_SL g4759 ( 
.A(n_4586),
.Y(n_4759)
);

OAI21x1_ASAP7_75t_L g4760 ( 
.A1(n_4419),
.A2(n_124),
.B(n_128),
.Y(n_4760)
);

OA21x2_ASAP7_75t_L g4761 ( 
.A1(n_4625),
.A2(n_129),
.B(n_130),
.Y(n_4761)
);

NAND2xp5_ASAP7_75t_L g4762 ( 
.A(n_4536),
.B(n_132),
.Y(n_4762)
);

OAI21x1_ASAP7_75t_L g4763 ( 
.A1(n_4419),
.A2(n_132),
.B(n_133),
.Y(n_4763)
);

OAI21x1_ASAP7_75t_L g4764 ( 
.A1(n_4466),
.A2(n_135),
.B(n_136),
.Y(n_4764)
);

INVxp67_ASAP7_75t_SL g4765 ( 
.A(n_4522),
.Y(n_4765)
);

OAI21x1_ASAP7_75t_L g4766 ( 
.A1(n_4532),
.A2(n_136),
.B(n_138),
.Y(n_4766)
);

INVx2_ASAP7_75t_L g4767 ( 
.A(n_4497),
.Y(n_4767)
);

OAI21x1_ASAP7_75t_L g4768 ( 
.A1(n_4510),
.A2(n_140),
.B(n_141),
.Y(n_4768)
);

OAI22xp5_ASAP7_75t_L g4769 ( 
.A1(n_4610),
.A2(n_142),
.B1(n_140),
.B2(n_141),
.Y(n_4769)
);

AOI21xp33_ASAP7_75t_L g4770 ( 
.A1(n_4511),
.A2(n_143),
.B(n_144),
.Y(n_4770)
);

AO32x2_ASAP7_75t_L g4771 ( 
.A1(n_4429),
.A2(n_4519),
.A3(n_4461),
.B1(n_4601),
.B2(n_4589),
.Y(n_4771)
);

OAI22xp5_ASAP7_75t_L g4772 ( 
.A1(n_4462),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_4772)
);

AND2x4_ASAP7_75t_L g4773 ( 
.A(n_4604),
.B(n_146),
.Y(n_4773)
);

AOI22xp33_ASAP7_75t_L g4774 ( 
.A1(n_4456),
.A2(n_4392),
.B1(n_4623),
.B2(n_4545),
.Y(n_4774)
);

OAI21x1_ASAP7_75t_L g4775 ( 
.A1(n_4629),
.A2(n_4597),
.B(n_4531),
.Y(n_4775)
);

INVx2_ASAP7_75t_SL g4776 ( 
.A(n_4622),
.Y(n_4776)
);

OAI21x1_ASAP7_75t_L g4777 ( 
.A1(n_4528),
.A2(n_4427),
.B(n_4407),
.Y(n_4777)
);

NAND2xp5_ASAP7_75t_L g4778 ( 
.A(n_4530),
.B(n_149),
.Y(n_4778)
);

AOI21x1_ASAP7_75t_L g4779 ( 
.A1(n_4602),
.A2(n_149),
.B(n_150),
.Y(n_4779)
);

NAND2x1p5_ASAP7_75t_L g4780 ( 
.A(n_4420),
.B(n_4614),
.Y(n_4780)
);

CKINVDCx20_ASAP7_75t_R g4781 ( 
.A(n_4606),
.Y(n_4781)
);

NAND2xp5_ASAP7_75t_SL g4782 ( 
.A(n_4434),
.B(n_150),
.Y(n_4782)
);

AND2x4_ASAP7_75t_L g4783 ( 
.A(n_4554),
.B(n_152),
.Y(n_4783)
);

INVx1_ASAP7_75t_L g4784 ( 
.A(n_4541),
.Y(n_4784)
);

A2O1A1Ixp33_ASAP7_75t_L g4785 ( 
.A1(n_4590),
.A2(n_157),
.B(n_154),
.C(n_156),
.Y(n_4785)
);

OAI21x1_ASAP7_75t_L g4786 ( 
.A1(n_4453),
.A2(n_154),
.B(n_156),
.Y(n_4786)
);

INVx3_ASAP7_75t_L g4787 ( 
.A(n_4433),
.Y(n_4787)
);

OAI21x1_ASAP7_75t_L g4788 ( 
.A1(n_4481),
.A2(n_158),
.B(n_159),
.Y(n_4788)
);

INVx8_ASAP7_75t_L g4789 ( 
.A(n_4565),
.Y(n_4789)
);

OAI21x1_ASAP7_75t_L g4790 ( 
.A1(n_4424),
.A2(n_158),
.B(n_160),
.Y(n_4790)
);

OAI21x1_ASAP7_75t_SL g4791 ( 
.A1(n_4533),
.A2(n_161),
.B(n_163),
.Y(n_4791)
);

INVx1_ASAP7_75t_L g4792 ( 
.A(n_4541),
.Y(n_4792)
);

AOI21xp5_ASAP7_75t_L g4793 ( 
.A1(n_4463),
.A2(n_161),
.B(n_163),
.Y(n_4793)
);

AOI221xp5_ASAP7_75t_L g4794 ( 
.A1(n_4391),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.C(n_168),
.Y(n_4794)
);

INVx3_ASAP7_75t_L g4795 ( 
.A(n_4509),
.Y(n_4795)
);

INVx1_ASAP7_75t_L g4796 ( 
.A(n_4541),
.Y(n_4796)
);

OAI21x1_ASAP7_75t_L g4797 ( 
.A1(n_4546),
.A2(n_165),
.B(n_168),
.Y(n_4797)
);

AND2x2_ASAP7_75t_SL g4798 ( 
.A(n_4627),
.B(n_169),
.Y(n_4798)
);

CKINVDCx16_ASAP7_75t_R g4799 ( 
.A(n_4573),
.Y(n_4799)
);

INVxp67_ASAP7_75t_SL g4800 ( 
.A(n_4509),
.Y(n_4800)
);

OA21x2_ASAP7_75t_L g4801 ( 
.A1(n_4514),
.A2(n_170),
.B(n_171),
.Y(n_4801)
);

OAI21x1_ASAP7_75t_L g4802 ( 
.A1(n_4479),
.A2(n_171),
.B(n_172),
.Y(n_4802)
);

INVx2_ASAP7_75t_L g4803 ( 
.A(n_4501),
.Y(n_4803)
);

INVx2_ASAP7_75t_L g4804 ( 
.A(n_4501),
.Y(n_4804)
);

NAND2xp5_ASAP7_75t_L g4805 ( 
.A(n_4579),
.B(n_172),
.Y(n_4805)
);

AOI22xp33_ASAP7_75t_L g4806 ( 
.A1(n_4508),
.A2(n_4583),
.B1(n_4405),
.B2(n_4540),
.Y(n_4806)
);

INVx2_ASAP7_75t_SL g4807 ( 
.A(n_4567),
.Y(n_4807)
);

A2O1A1Ixp33_ASAP7_75t_SL g4808 ( 
.A1(n_4504),
.A2(n_175),
.B(n_173),
.C(n_174),
.Y(n_4808)
);

OAI21x1_ASAP7_75t_L g4809 ( 
.A1(n_4426),
.A2(n_175),
.B(n_176),
.Y(n_4809)
);

INVx3_ASAP7_75t_L g4810 ( 
.A(n_4567),
.Y(n_4810)
);

OAI21x1_ASAP7_75t_L g4811 ( 
.A1(n_4441),
.A2(n_177),
.B(n_178),
.Y(n_4811)
);

NAND2xp5_ASAP7_75t_L g4812 ( 
.A(n_4502),
.B(n_177),
.Y(n_4812)
);

NOR3xp33_ASAP7_75t_SL g4813 ( 
.A(n_4518),
.B(n_178),
.C(n_179),
.Y(n_4813)
);

OAI21x1_ASAP7_75t_L g4814 ( 
.A1(n_4482),
.A2(n_4464),
.B(n_4460),
.Y(n_4814)
);

OAI21x1_ASAP7_75t_L g4815 ( 
.A1(n_4605),
.A2(n_179),
.B(n_180),
.Y(n_4815)
);

NAND2xp5_ASAP7_75t_L g4816 ( 
.A(n_4619),
.B(n_181),
.Y(n_4816)
);

INVx2_ASAP7_75t_L g4817 ( 
.A(n_4501),
.Y(n_4817)
);

AO21x2_ASAP7_75t_L g4818 ( 
.A1(n_4438),
.A2(n_181),
.B(n_182),
.Y(n_4818)
);

OAI21x1_ASAP7_75t_L g4819 ( 
.A1(n_4469),
.A2(n_182),
.B(n_183),
.Y(n_4819)
);

INVx1_ASAP7_75t_L g4820 ( 
.A(n_4634),
.Y(n_4820)
);

OAI21x1_ASAP7_75t_L g4821 ( 
.A1(n_4474),
.A2(n_185),
.B(n_186),
.Y(n_4821)
);

BUFx2_ASAP7_75t_L g4822 ( 
.A(n_4565),
.Y(n_4822)
);

AO32x2_ASAP7_75t_L g4823 ( 
.A1(n_4487),
.A2(n_188),
.A3(n_185),
.B1(n_186),
.B2(n_189),
.Y(n_4823)
);

OAI21x1_ASAP7_75t_L g4824 ( 
.A1(n_4577),
.A2(n_189),
.B(n_191),
.Y(n_4824)
);

OAI21x1_ASAP7_75t_L g4825 ( 
.A1(n_4621),
.A2(n_4475),
.B(n_4446),
.Y(n_4825)
);

INVx1_ASAP7_75t_L g4826 ( 
.A(n_4634),
.Y(n_4826)
);

OAI21xp5_ASAP7_75t_L g4827 ( 
.A1(n_4492),
.A2(n_191),
.B(n_193),
.Y(n_4827)
);

AOI21x1_ASAP7_75t_L g4828 ( 
.A1(n_4549),
.A2(n_194),
.B(n_195),
.Y(n_4828)
);

OA21x2_ASAP7_75t_L g4829 ( 
.A1(n_4543),
.A2(n_195),
.B(n_196),
.Y(n_4829)
);

O2A1O1Ixp33_ASAP7_75t_SL g4830 ( 
.A1(n_4782),
.A2(n_4561),
.B(n_4542),
.C(n_4506),
.Y(n_4830)
);

INVx1_ASAP7_75t_L g4831 ( 
.A(n_4642),
.Y(n_4831)
);

OAI22xp5_ASAP7_75t_L g4832 ( 
.A1(n_4706),
.A2(n_4394),
.B1(n_4632),
.B2(n_4516),
.Y(n_4832)
);

INVx1_ASAP7_75t_L g4833 ( 
.A(n_4642),
.Y(n_4833)
);

CKINVDCx6p67_ASAP7_75t_R g4834 ( 
.A(n_4715),
.Y(n_4834)
);

OAI22xp33_ASAP7_75t_L g4835 ( 
.A1(n_4706),
.A2(n_4458),
.B1(n_4566),
.B2(n_4634),
.Y(n_4835)
);

OAI22xp5_ASAP7_75t_L g4836 ( 
.A1(n_4687),
.A2(n_4527),
.B1(n_4584),
.B2(n_4596),
.Y(n_4836)
);

NOR2x1_ASAP7_75t_R g4837 ( 
.A(n_4649),
.B(n_4402),
.Y(n_4837)
);

AOI22xp33_ASAP7_75t_L g4838 ( 
.A1(n_4829),
.A2(n_4525),
.B1(n_4491),
.B2(n_4570),
.Y(n_4838)
);

INVx4_ASAP7_75t_L g4839 ( 
.A(n_4649),
.Y(n_4839)
);

AOI22xp33_ASAP7_75t_L g4840 ( 
.A1(n_4829),
.A2(n_4572),
.B1(n_4593),
.B2(n_4580),
.Y(n_4840)
);

AND2x4_ASAP7_75t_L g4841 ( 
.A(n_4661),
.B(n_4440),
.Y(n_4841)
);

NAND3xp33_ASAP7_75t_L g4842 ( 
.A(n_4793),
.B(n_4418),
.C(n_4410),
.Y(n_4842)
);

AND2x2_ASAP7_75t_L g4843 ( 
.A(n_4733),
.B(n_4557),
.Y(n_4843)
);

AOI22xp33_ASAP7_75t_L g4844 ( 
.A1(n_4658),
.A2(n_4674),
.B1(n_4667),
.B2(n_4670),
.Y(n_4844)
);

INVx1_ASAP7_75t_L g4845 ( 
.A(n_4646),
.Y(n_4845)
);

AND2x4_ASAP7_75t_L g4846 ( 
.A(n_4661),
.B(n_4440),
.Y(n_4846)
);

O2A1O1Ixp5_ASAP7_75t_L g4847 ( 
.A1(n_4721),
.A2(n_4812),
.B(n_4712),
.C(n_4724),
.Y(n_4847)
);

INVx6_ASAP7_75t_L g4848 ( 
.A(n_4638),
.Y(n_4848)
);

NAND2xp5_ASAP7_75t_L g4849 ( 
.A(n_4650),
.B(n_4557),
.Y(n_4849)
);

BUFx6f_ASAP7_75t_L g4850 ( 
.A(n_4659),
.Y(n_4850)
);

OAI221xp5_ASAP7_75t_L g4851 ( 
.A1(n_4774),
.A2(n_4444),
.B1(n_4523),
.B2(n_4568),
.C(n_4564),
.Y(n_4851)
);

NAND2xp5_ASAP7_75t_L g4852 ( 
.A(n_4724),
.B(n_4440),
.Y(n_4852)
);

INVx1_ASAP7_75t_L g4853 ( 
.A(n_4646),
.Y(n_4853)
);

OAI21x1_ASAP7_75t_L g4854 ( 
.A1(n_4732),
.A2(n_4741),
.B(n_4767),
.Y(n_4854)
);

INVx1_ASAP7_75t_L g4855 ( 
.A(n_4654),
.Y(n_4855)
);

AOI21xp5_ASAP7_75t_L g4856 ( 
.A1(n_4648),
.A2(n_4447),
.B(n_4534),
.Y(n_4856)
);

AOI221xp5_ASAP7_75t_L g4857 ( 
.A1(n_4750),
.A2(n_4587),
.B1(n_4512),
.B2(n_4562),
.C(n_4459),
.Y(n_4857)
);

OAI22xp33_ASAP7_75t_L g4858 ( 
.A1(n_4799),
.A2(n_4458),
.B1(n_4556),
.B2(n_4626),
.Y(n_4858)
);

BUFx6f_ASAP7_75t_L g4859 ( 
.A(n_4659),
.Y(n_4859)
);

INVx1_ASAP7_75t_L g4860 ( 
.A(n_4654),
.Y(n_4860)
);

BUFx3_ASAP7_75t_L g4861 ( 
.A(n_4668),
.Y(n_4861)
);

INVx4_ASAP7_75t_L g4862 ( 
.A(n_4665),
.Y(n_4862)
);

AOI221xp5_ASAP7_75t_L g4863 ( 
.A1(n_4770),
.A2(n_4513),
.B1(n_4628),
.B2(n_4626),
.C(n_4553),
.Y(n_4863)
);

INVx1_ASAP7_75t_L g4864 ( 
.A(n_4655),
.Y(n_4864)
);

A2O1A1Ixp33_ASAP7_75t_L g4865 ( 
.A1(n_4722),
.A2(n_4458),
.B(n_4628),
.C(n_4553),
.Y(n_4865)
);

INVx1_ASAP7_75t_L g4866 ( 
.A(n_4655),
.Y(n_4866)
);

INVx3_ASAP7_75t_L g4867 ( 
.A(n_4638),
.Y(n_4867)
);

AOI22xp33_ASAP7_75t_L g4868 ( 
.A1(n_4744),
.A2(n_4487),
.B1(n_4471),
.B2(n_4455),
.Y(n_4868)
);

BUFx2_ASAP7_75t_L g4869 ( 
.A(n_4781),
.Y(n_4869)
);

AOI221xp5_ASAP7_75t_L g4870 ( 
.A1(n_4769),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.C(n_199),
.Y(n_4870)
);

AND2x4_ASAP7_75t_L g4871 ( 
.A(n_4822),
.B(n_4455),
.Y(n_4871)
);

INVx1_ASAP7_75t_L g4872 ( 
.A(n_4676),
.Y(n_4872)
);

AOI21xp5_ASAP7_75t_L g4873 ( 
.A1(n_4720),
.A2(n_4487),
.B(n_4455),
.Y(n_4873)
);

INVx3_ASAP7_75t_L g4874 ( 
.A(n_4669),
.Y(n_4874)
);

NAND2xp5_ASAP7_75t_L g4875 ( 
.A(n_4652),
.B(n_4471),
.Y(n_4875)
);

BUFx2_ASAP7_75t_L g4876 ( 
.A(n_4673),
.Y(n_4876)
);

INVx1_ASAP7_75t_L g4877 ( 
.A(n_4676),
.Y(n_4877)
);

INVx2_ASAP7_75t_L g4878 ( 
.A(n_4751),
.Y(n_4878)
);

OAI22xp5_ASAP7_75t_L g4879 ( 
.A1(n_4813),
.A2(n_200),
.B1(n_197),
.B2(n_199),
.Y(n_4879)
);

OAI22xp5_ASAP7_75t_L g4880 ( 
.A1(n_4799),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_4880)
);

INVx4_ASAP7_75t_L g4881 ( 
.A(n_4639),
.Y(n_4881)
);

A2O1A1Ixp33_ASAP7_75t_L g4882 ( 
.A1(n_4827),
.A2(n_207),
.B(n_204),
.C(n_205),
.Y(n_4882)
);

CKINVDCx16_ASAP7_75t_R g4883 ( 
.A(n_4689),
.Y(n_4883)
);

OR2x6_ASAP7_75t_SL g4884 ( 
.A(n_4641),
.B(n_4507),
.Y(n_4884)
);

AOI22xp33_ASAP7_75t_L g4885 ( 
.A1(n_4640),
.A2(n_4507),
.B1(n_4499),
.B2(n_4578),
.Y(n_4885)
);

OAI22xp33_ASAP7_75t_L g4886 ( 
.A1(n_4704),
.A2(n_4578),
.B1(n_4507),
.B2(n_4499),
.Y(n_4886)
);

OA21x2_ASAP7_75t_L g4887 ( 
.A1(n_4732),
.A2(n_4499),
.B(n_4578),
.Y(n_4887)
);

BUFx2_ASAP7_75t_L g4888 ( 
.A(n_4719),
.Y(n_4888)
);

AND2x2_ASAP7_75t_L g4889 ( 
.A(n_4733),
.B(n_4643),
.Y(n_4889)
);

OR2x6_ASAP7_75t_L g4890 ( 
.A(n_4789),
.B(n_205),
.Y(n_4890)
);

BUFx2_ASAP7_75t_L g4891 ( 
.A(n_4742),
.Y(n_4891)
);

AOI22xp33_ASAP7_75t_L g4892 ( 
.A1(n_4741),
.A2(n_209),
.B1(n_207),
.B2(n_208),
.Y(n_4892)
);

INVxp67_ASAP7_75t_SL g4893 ( 
.A(n_4682),
.Y(n_4893)
);

NOR2x1_ASAP7_75t_SL g4894 ( 
.A(n_4757),
.B(n_4679),
.Y(n_4894)
);

OAI21xp5_ASAP7_75t_L g4895 ( 
.A1(n_4704),
.A2(n_208),
.B(n_210),
.Y(n_4895)
);

BUFx8_ASAP7_75t_L g4896 ( 
.A(n_4698),
.Y(n_4896)
);

AND2x4_ASAP7_75t_L g4897 ( 
.A(n_4787),
.B(n_211),
.Y(n_4897)
);

INVx1_ASAP7_75t_L g4898 ( 
.A(n_4680),
.Y(n_4898)
);

INVx2_ASAP7_75t_L g4899 ( 
.A(n_4753),
.Y(n_4899)
);

INVx2_ASAP7_75t_L g4900 ( 
.A(n_4758),
.Y(n_4900)
);

AO31x2_ASAP7_75t_L g4901 ( 
.A1(n_4820),
.A2(n_4826),
.A3(n_4677),
.B(n_4792),
.Y(n_4901)
);

INVx4_ASAP7_75t_SL g4902 ( 
.A(n_4783),
.Y(n_4902)
);

AOI22xp33_ASAP7_75t_SL g4903 ( 
.A1(n_4692),
.A2(n_214),
.B1(n_212),
.B2(n_213),
.Y(n_4903)
);

AND2x4_ASAP7_75t_L g4904 ( 
.A(n_4787),
.B(n_212),
.Y(n_4904)
);

AND2x4_ASAP7_75t_L g4905 ( 
.A(n_4635),
.B(n_213),
.Y(n_4905)
);

OR2x6_ASAP7_75t_L g4906 ( 
.A(n_4789),
.B(n_214),
.Y(n_4906)
);

INVx3_ASAP7_75t_L g4907 ( 
.A(n_4664),
.Y(n_4907)
);

AOI22xp33_ASAP7_75t_SL g4908 ( 
.A1(n_4692),
.A2(n_219),
.B1(n_215),
.B2(n_218),
.Y(n_4908)
);

OAI22xp5_ASAP7_75t_L g4909 ( 
.A1(n_4798),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_4909)
);

AOI22xp33_ASAP7_75t_L g4910 ( 
.A1(n_4820),
.A2(n_223),
.B1(n_220),
.B2(n_221),
.Y(n_4910)
);

INVx2_ASAP7_75t_L g4911 ( 
.A(n_4651),
.Y(n_4911)
);

OAI22xp33_ASAP7_75t_L g4912 ( 
.A1(n_4761),
.A2(n_228),
.B1(n_225),
.B2(n_226),
.Y(n_4912)
);

NOR2xp33_ASAP7_75t_L g4913 ( 
.A(n_4664),
.B(n_228),
.Y(n_4913)
);

OAI21x1_ASAP7_75t_L g4914 ( 
.A1(n_4647),
.A2(n_229),
.B(n_230),
.Y(n_4914)
);

OAI22xp33_ASAP7_75t_L g4915 ( 
.A1(n_4761),
.A2(n_232),
.B1(n_229),
.B2(n_231),
.Y(n_4915)
);

OAI22xp5_ASAP7_75t_L g4916 ( 
.A1(n_4780),
.A2(n_235),
.B1(n_232),
.B2(n_234),
.Y(n_4916)
);

CKINVDCx5p33_ASAP7_75t_R g4917 ( 
.A(n_4708),
.Y(n_4917)
);

INVx2_ASAP7_75t_L g4918 ( 
.A(n_4680),
.Y(n_4918)
);

INVx1_ASAP7_75t_L g4919 ( 
.A(n_4656),
.Y(n_4919)
);

A2O1A1Ixp33_ASAP7_75t_L g4920 ( 
.A1(n_4694),
.A2(n_237),
.B(n_234),
.C(n_236),
.Y(n_4920)
);

OR2x6_ASAP7_75t_L g4921 ( 
.A(n_4789),
.B(n_236),
.Y(n_4921)
);

OR2x2_ASAP7_75t_L g4922 ( 
.A(n_4682),
.B(n_239),
.Y(n_4922)
);

INVx1_ASAP7_75t_L g4923 ( 
.A(n_4656),
.Y(n_4923)
);

INVx2_ASAP7_75t_L g4924 ( 
.A(n_4681),
.Y(n_4924)
);

AOI22xp33_ASAP7_75t_L g4925 ( 
.A1(n_4826),
.A2(n_4801),
.B1(n_4716),
.B2(n_4749),
.Y(n_4925)
);

INVx1_ASAP7_75t_L g4926 ( 
.A(n_4657),
.Y(n_4926)
);

OAI22xp5_ASAP7_75t_L g4927 ( 
.A1(n_4754),
.A2(n_4757),
.B1(n_4693),
.B2(n_4783),
.Y(n_4927)
);

NOR2x1_ASAP7_75t_SL g4928 ( 
.A(n_4679),
.B(n_239),
.Y(n_4928)
);

INVx3_ASAP7_75t_L g4929 ( 
.A(n_4776),
.Y(n_4929)
);

AND2x2_ASAP7_75t_L g4930 ( 
.A(n_4657),
.B(n_242),
.Y(n_4930)
);

INVx3_ASAP7_75t_L g4931 ( 
.A(n_4759),
.Y(n_4931)
);

CKINVDCx11_ASAP7_75t_R g4932 ( 
.A(n_4684),
.Y(n_4932)
);

AOI22xp33_ASAP7_75t_L g4933 ( 
.A1(n_4801),
.A2(n_244),
.B1(n_242),
.B2(n_243),
.Y(n_4933)
);

HB1xp67_ASAP7_75t_L g4934 ( 
.A(n_4671),
.Y(n_4934)
);

AOI21xp33_ASAP7_75t_L g4935 ( 
.A1(n_4808),
.A2(n_243),
.B(n_244),
.Y(n_4935)
);

OAI22xp5_ASAP7_75t_L g4936 ( 
.A1(n_4679),
.A2(n_4748),
.B1(n_4726),
.B2(n_4806),
.Y(n_4936)
);

AND2x4_ASAP7_75t_L g4937 ( 
.A(n_4635),
.B(n_245),
.Y(n_4937)
);

CKINVDCx5p33_ASAP7_75t_R g4938 ( 
.A(n_4711),
.Y(n_4938)
);

AND2x2_ASAP7_75t_L g4939 ( 
.A(n_4671),
.B(n_245),
.Y(n_4939)
);

BUFx2_ASAP7_75t_R g4940 ( 
.A(n_4690),
.Y(n_4940)
);

NOR2xp33_ASAP7_75t_L g4941 ( 
.A(n_4684),
.B(n_246),
.Y(n_4941)
);

AND2x2_ASAP7_75t_L g4942 ( 
.A(n_4675),
.B(n_251),
.Y(n_4942)
);

AOI22xp5_ASAP7_75t_L g4943 ( 
.A1(n_4645),
.A2(n_253),
.B1(n_251),
.B2(n_252),
.Y(n_4943)
);

INVx1_ASAP7_75t_L g4944 ( 
.A(n_4675),
.Y(n_4944)
);

INVx2_ASAP7_75t_L g4945 ( 
.A(n_4777),
.Y(n_4945)
);

AND2x4_ASAP7_75t_L g4946 ( 
.A(n_4678),
.B(n_253),
.Y(n_4946)
);

BUFx12f_ASAP7_75t_L g4947 ( 
.A(n_4705),
.Y(n_4947)
);

BUFx12f_ASAP7_75t_L g4948 ( 
.A(n_4683),
.Y(n_4948)
);

NAND2xp33_ASAP7_75t_R g4949 ( 
.A(n_4683),
.B(n_254),
.Y(n_4949)
);

BUFx4f_ASAP7_75t_SL g4950 ( 
.A(n_4807),
.Y(n_4950)
);

AOI22xp5_ASAP7_75t_L g4951 ( 
.A1(n_4773),
.A2(n_256),
.B1(n_254),
.B2(n_255),
.Y(n_4951)
);

INVx1_ASAP7_75t_L g4952 ( 
.A(n_4747),
.Y(n_4952)
);

INVx4_ASAP7_75t_L g4953 ( 
.A(n_4748),
.Y(n_4953)
);

INVx1_ASAP7_75t_L g4954 ( 
.A(n_4747),
.Y(n_4954)
);

AND2x6_ASAP7_75t_L g4955 ( 
.A(n_4773),
.B(n_255),
.Y(n_4955)
);

CKINVDCx20_ASAP7_75t_R g4956 ( 
.A(n_4691),
.Y(n_4956)
);

NAND2xp5_ASAP7_75t_L g4957 ( 
.A(n_4653),
.B(n_256),
.Y(n_4957)
);

AND2x2_ASAP7_75t_L g4958 ( 
.A(n_4800),
.B(n_258),
.Y(n_4958)
);

BUFx2_ASAP7_75t_L g4959 ( 
.A(n_4795),
.Y(n_4959)
);

HB1xp67_ASAP7_75t_L g4960 ( 
.A(n_4644),
.Y(n_4960)
);

NAND2x1p5_ASAP7_75t_L g4961 ( 
.A(n_4752),
.B(n_258),
.Y(n_4961)
);

NAND2xp5_ASAP7_75t_L g4962 ( 
.A(n_4755),
.B(n_260),
.Y(n_4962)
);

OA21x2_ASAP7_75t_L g4963 ( 
.A1(n_4784),
.A2(n_260),
.B(n_261),
.Y(n_4963)
);

BUFx2_ASAP7_75t_SL g4964 ( 
.A(n_4752),
.Y(n_4964)
);

AOI22xp33_ASAP7_75t_SL g4965 ( 
.A1(n_4743),
.A2(n_4731),
.B1(n_4697),
.B2(n_4791),
.Y(n_4965)
);

OAI221xp5_ASAP7_75t_L g4966 ( 
.A1(n_4756),
.A2(n_265),
.B1(n_262),
.B2(n_263),
.C(n_266),
.Y(n_4966)
);

OAI22xp5_ASAP7_75t_L g4967 ( 
.A1(n_4785),
.A2(n_266),
.B1(n_262),
.B2(n_263),
.Y(n_4967)
);

INVx1_ASAP7_75t_L g4968 ( 
.A(n_4755),
.Y(n_4968)
);

AOI221xp5_ASAP7_75t_L g4969 ( 
.A1(n_4740),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.C(n_270),
.Y(n_4969)
);

AOI22xp33_ASAP7_75t_SL g4970 ( 
.A1(n_4731),
.A2(n_270),
.B1(n_267),
.B2(n_269),
.Y(n_4970)
);

CKINVDCx5p33_ASAP7_75t_R g4971 ( 
.A(n_4795),
.Y(n_4971)
);

AND2x4_ASAP7_75t_L g4972 ( 
.A(n_4678),
.B(n_271),
.Y(n_4972)
);

AND2x4_ASAP7_75t_L g4973 ( 
.A(n_4636),
.B(n_272),
.Y(n_4973)
);

AOI22xp33_ASAP7_75t_L g4974 ( 
.A1(n_4818),
.A2(n_276),
.B1(n_273),
.B2(n_274),
.Y(n_4974)
);

AOI221xp5_ASAP7_75t_L g4975 ( 
.A1(n_4762),
.A2(n_277),
.B1(n_273),
.B2(n_274),
.C(n_280),
.Y(n_4975)
);

OAI222xp33_ASAP7_75t_L g4976 ( 
.A1(n_4765),
.A2(n_281),
.B1(n_283),
.B2(n_277),
.C1(n_280),
.C2(n_282),
.Y(n_4976)
);

AOI22xp33_ASAP7_75t_L g4977 ( 
.A1(n_4818),
.A2(n_285),
.B1(n_282),
.B2(n_284),
.Y(n_4977)
);

INVx2_ASAP7_75t_L g4978 ( 
.A(n_4685),
.Y(n_4978)
);

INVx2_ASAP7_75t_L g4979 ( 
.A(n_4973),
.Y(n_4979)
);

OR2x2_ASAP7_75t_L g4980 ( 
.A(n_4891),
.B(n_4699),
.Y(n_4980)
);

BUFx3_ASAP7_75t_L g4981 ( 
.A(n_4869),
.Y(n_4981)
);

OA21x2_ASAP7_75t_L g4982 ( 
.A1(n_4854),
.A2(n_4792),
.B(n_4784),
.Y(n_4982)
);

AOI221xp5_ASAP7_75t_L g4983 ( 
.A1(n_4835),
.A2(n_4778),
.B1(n_4805),
.B2(n_4772),
.C(n_4794),
.Y(n_4983)
);

A2O1A1Ixp33_ASAP7_75t_L g4984 ( 
.A1(n_4847),
.A2(n_4688),
.B(n_4746),
.C(n_4815),
.Y(n_4984)
);

AOI22xp33_ASAP7_75t_L g4985 ( 
.A1(n_4844),
.A2(n_4636),
.B1(n_4672),
.B2(n_4660),
.Y(n_4985)
);

HB1xp67_ASAP7_75t_L g4986 ( 
.A(n_4934),
.Y(n_4986)
);

OAI22xp5_ASAP7_75t_L g4987 ( 
.A1(n_4848),
.A2(n_4965),
.B1(n_4925),
.B2(n_4940),
.Y(n_4987)
);

AOI221xp5_ASAP7_75t_L g4988 ( 
.A1(n_4912),
.A2(n_4709),
.B1(n_4695),
.B2(n_4727),
.C(n_4816),
.Y(n_4988)
);

INVx2_ASAP7_75t_L g4989 ( 
.A(n_4973),
.Y(n_4989)
);

NAND2xp5_ASAP7_75t_L g4990 ( 
.A(n_4843),
.B(n_4849),
.Y(n_4990)
);

AND2x4_ASAP7_75t_L g4991 ( 
.A(n_4867),
.B(n_4659),
.Y(n_4991)
);

HB1xp67_ASAP7_75t_L g4992 ( 
.A(n_4918),
.Y(n_4992)
);

OAI21xp5_ASAP7_75t_SL g4993 ( 
.A1(n_4879),
.A2(n_4880),
.B(n_4927),
.Y(n_4993)
);

OAI22xp5_ASAP7_75t_L g4994 ( 
.A1(n_4848),
.A2(n_4696),
.B1(n_4729),
.B2(n_4810),
.Y(n_4994)
);

NAND2xp5_ASAP7_75t_L g4995 ( 
.A(n_4893),
.B(n_4672),
.Y(n_4995)
);

AOI21xp5_ASAP7_75t_L g4996 ( 
.A1(n_4894),
.A2(n_4637),
.B(n_4644),
.Y(n_4996)
);

INVx5_ASAP7_75t_SL g4997 ( 
.A(n_4890),
.Y(n_4997)
);

HB1xp67_ASAP7_75t_L g4998 ( 
.A(n_4831),
.Y(n_4998)
);

OAI211xp5_ASAP7_75t_L g4999 ( 
.A1(n_4975),
.A2(n_4707),
.B(n_4710),
.C(n_4828),
.Y(n_4999)
);

OA21x2_ASAP7_75t_L g5000 ( 
.A1(n_4960),
.A2(n_4796),
.B(n_4700),
.Y(n_5000)
);

AOI22xp33_ASAP7_75t_L g5001 ( 
.A1(n_4895),
.A2(n_4660),
.B1(n_4713),
.B2(n_4734),
.Y(n_5001)
);

OAI221xp5_ASAP7_75t_L g5002 ( 
.A1(n_4838),
.A2(n_4771),
.B1(n_4779),
.B2(n_4796),
.C(n_4736),
.Y(n_5002)
);

INVx1_ASAP7_75t_L g5003 ( 
.A(n_4833),
.Y(n_5003)
);

NAND2xp5_ASAP7_75t_L g5004 ( 
.A(n_4930),
.B(n_4728),
.Y(n_5004)
);

INVx3_ASAP7_75t_L g5005 ( 
.A(n_4953),
.Y(n_5005)
);

OR2x6_ASAP7_75t_L g5006 ( 
.A(n_4890),
.B(n_4906),
.Y(n_5006)
);

INVx1_ASAP7_75t_L g5007 ( 
.A(n_4845),
.Y(n_5007)
);

INVx1_ASAP7_75t_L g5008 ( 
.A(n_4853),
.Y(n_5008)
);

OAI22xp33_ASAP7_75t_L g5009 ( 
.A1(n_4949),
.A2(n_4771),
.B1(n_4810),
.B2(n_4823),
.Y(n_5009)
);

BUFx3_ASAP7_75t_L g5010 ( 
.A(n_4956),
.Y(n_5010)
);

OAI22xp33_ASAP7_75t_L g5011 ( 
.A1(n_4832),
.A2(n_4771),
.B1(n_4823),
.B2(n_4725),
.Y(n_5011)
);

OAI221xp5_ASAP7_75t_L g5012 ( 
.A1(n_4865),
.A2(n_4737),
.B1(n_4714),
.B2(n_4823),
.C(n_4804),
.Y(n_5012)
);

AOI22xp33_ASAP7_75t_L g5013 ( 
.A1(n_4903),
.A2(n_4728),
.B1(n_4702),
.B2(n_4764),
.Y(n_5013)
);

INVx2_ASAP7_75t_SL g5014 ( 
.A(n_4839),
.Y(n_5014)
);

INVx1_ASAP7_75t_L g5015 ( 
.A(n_4855),
.Y(n_5015)
);

OR2x6_ASAP7_75t_L g5016 ( 
.A(n_4906),
.B(n_4739),
.Y(n_5016)
);

AND2x2_ASAP7_75t_L g5017 ( 
.A(n_4888),
.B(n_4728),
.Y(n_5017)
);

OAI21xp33_ASAP7_75t_SL g5018 ( 
.A1(n_4889),
.A2(n_4763),
.B(n_4760),
.Y(n_5018)
);

AOI221xp5_ASAP7_75t_L g5019 ( 
.A1(n_4915),
.A2(n_4797),
.B1(n_4803),
.B2(n_4817),
.C(n_4723),
.Y(n_5019)
);

OAI22xp33_ASAP7_75t_L g5020 ( 
.A1(n_4936),
.A2(n_4728),
.B1(n_4738),
.B2(n_4666),
.Y(n_5020)
);

OAI21x1_ASAP7_75t_L g5021 ( 
.A1(n_4945),
.A2(n_4875),
.B(n_4852),
.Y(n_5021)
);

AO21x2_ASAP7_75t_L g5022 ( 
.A1(n_4962),
.A2(n_4662),
.B(n_4735),
.Y(n_5022)
);

AOI22xp33_ASAP7_75t_L g5023 ( 
.A1(n_4908),
.A2(n_4728),
.B1(n_4825),
.B2(n_4811),
.Y(n_5023)
);

INVx2_ASAP7_75t_L g5024 ( 
.A(n_4901),
.Y(n_5024)
);

OAI211xp5_ASAP7_75t_L g5025 ( 
.A1(n_4969),
.A2(n_4786),
.B(n_4809),
.C(n_4819),
.Y(n_5025)
);

AND2x2_ASAP7_75t_L g5026 ( 
.A(n_4959),
.B(n_4775),
.Y(n_5026)
);

OAI211xp5_ASAP7_75t_L g5027 ( 
.A1(n_4913),
.A2(n_4821),
.B(n_4790),
.C(n_4718),
.Y(n_5027)
);

OAI22xp33_ASAP7_75t_L g5028 ( 
.A1(n_4963),
.A2(n_4738),
.B1(n_4814),
.B2(n_4686),
.Y(n_5028)
);

AOI22xp33_ASAP7_75t_L g5029 ( 
.A1(n_4863),
.A2(n_4824),
.B1(n_4788),
.B2(n_4802),
.Y(n_5029)
);

AOI22xp33_ASAP7_75t_L g5030 ( 
.A1(n_4842),
.A2(n_4717),
.B1(n_4766),
.B2(n_4703),
.Y(n_5030)
);

BUFx3_ASAP7_75t_L g5031 ( 
.A(n_4917),
.Y(n_5031)
);

AOI22xp33_ASAP7_75t_L g5032 ( 
.A1(n_4963),
.A2(n_4745),
.B1(n_4701),
.B2(n_4768),
.Y(n_5032)
);

OAI22xp5_ASAP7_75t_L g5033 ( 
.A1(n_4964),
.A2(n_4738),
.B1(n_4730),
.B2(n_4663),
.Y(n_5033)
);

CKINVDCx5p33_ASAP7_75t_R g5034 ( 
.A(n_4834),
.Y(n_5034)
);

INVx2_ASAP7_75t_L g5035 ( 
.A(n_4901),
.Y(n_5035)
);

OR2x2_ASAP7_75t_L g5036 ( 
.A(n_4876),
.B(n_286),
.Y(n_5036)
);

AOI21xp5_ASAP7_75t_L g5037 ( 
.A1(n_4858),
.A2(n_287),
.B(n_289),
.Y(n_5037)
);

NAND2xp5_ASAP7_75t_L g5038 ( 
.A(n_4939),
.B(n_287),
.Y(n_5038)
);

CKINVDCx6p67_ASAP7_75t_R g5039 ( 
.A(n_4883),
.Y(n_5039)
);

AOI21xp5_ASAP7_75t_L g5040 ( 
.A1(n_4928),
.A2(n_290),
.B(n_291),
.Y(n_5040)
);

AOI22xp33_ASAP7_75t_L g5041 ( 
.A1(n_4966),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_5041)
);

AOI21xp33_ASAP7_75t_L g5042 ( 
.A1(n_4837),
.A2(n_294),
.B(n_295),
.Y(n_5042)
);

INVxp67_ASAP7_75t_L g5043 ( 
.A(n_4941),
.Y(n_5043)
);

INVx2_ASAP7_75t_L g5044 ( 
.A(n_4901),
.Y(n_5044)
);

NOR2xp33_ASAP7_75t_L g5045 ( 
.A(n_4932),
.B(n_297),
.Y(n_5045)
);

AOI21x1_ASAP7_75t_L g5046 ( 
.A1(n_4905),
.A2(n_298),
.B(n_299),
.Y(n_5046)
);

OR2x2_ASAP7_75t_L g5047 ( 
.A(n_4860),
.B(n_298),
.Y(n_5047)
);

AOI221xp5_ASAP7_75t_L g5048 ( 
.A1(n_4967),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.C(n_304),
.Y(n_5048)
);

AO21x2_ASAP7_75t_L g5049 ( 
.A1(n_4886),
.A2(n_301),
.B(n_305),
.Y(n_5049)
);

OA21x2_ASAP7_75t_L g5050 ( 
.A1(n_4878),
.A2(n_305),
.B(n_306),
.Y(n_5050)
);

OR2x6_ASAP7_75t_L g5051 ( 
.A(n_4921),
.B(n_306),
.Y(n_5051)
);

BUFx2_ASAP7_75t_L g5052 ( 
.A(n_4948),
.Y(n_5052)
);

NAND2xp5_ASAP7_75t_L g5053 ( 
.A(n_4942),
.B(n_307),
.Y(n_5053)
);

NAND2xp5_ASAP7_75t_L g5054 ( 
.A(n_4864),
.B(n_308),
.Y(n_5054)
);

INVx1_ASAP7_75t_L g5055 ( 
.A(n_4866),
.Y(n_5055)
);

INVx1_ASAP7_75t_L g5056 ( 
.A(n_4872),
.Y(n_5056)
);

AOI221xp5_ASAP7_75t_L g5057 ( 
.A1(n_4882),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.C(n_312),
.Y(n_5057)
);

AND2x4_ASAP7_75t_L g5058 ( 
.A(n_4902),
.B(n_310),
.Y(n_5058)
);

O2A1O1Ixp33_ASAP7_75t_L g5059 ( 
.A1(n_4976),
.A2(n_314),
.B(n_311),
.C(n_313),
.Y(n_5059)
);

AND2x2_ASAP7_75t_L g5060 ( 
.A(n_4874),
.B(n_314),
.Y(n_5060)
);

INVx2_ASAP7_75t_L g5061 ( 
.A(n_4877),
.Y(n_5061)
);

INVx4_ASAP7_75t_L g5062 ( 
.A(n_4881),
.Y(n_5062)
);

OAI211xp5_ASAP7_75t_SL g5063 ( 
.A1(n_4870),
.A2(n_4840),
.B(n_4830),
.C(n_4857),
.Y(n_5063)
);

OAI21xp5_ASAP7_75t_L g5064 ( 
.A1(n_4970),
.A2(n_315),
.B(n_318),
.Y(n_5064)
);

AOI22xp33_ASAP7_75t_L g5065 ( 
.A1(n_4836),
.A2(n_319),
.B1(n_315),
.B2(n_318),
.Y(n_5065)
);

AND2x4_ASAP7_75t_L g5066 ( 
.A(n_4902),
.B(n_320),
.Y(n_5066)
);

OR2x6_ASAP7_75t_L g5067 ( 
.A(n_4921),
.B(n_322),
.Y(n_5067)
);

AOI221xp5_ASAP7_75t_L g5068 ( 
.A1(n_4933),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.C(n_325),
.Y(n_5068)
);

OR2x2_ASAP7_75t_L g5069 ( 
.A(n_4898),
.B(n_4919),
.Y(n_5069)
);

BUFx3_ASAP7_75t_L g5070 ( 
.A(n_4896),
.Y(n_5070)
);

OAI22x1_ASAP7_75t_L g5071 ( 
.A1(n_4961),
.A2(n_4931),
.B1(n_4904),
.B2(n_4897),
.Y(n_5071)
);

AND2x4_ASAP7_75t_SL g5072 ( 
.A(n_4862),
.B(n_4946),
.Y(n_5072)
);

HB1xp67_ASAP7_75t_L g5073 ( 
.A(n_4923),
.Y(n_5073)
);

O2A1O1Ixp33_ASAP7_75t_L g5074 ( 
.A1(n_4909),
.A2(n_327),
.B(n_324),
.C(n_326),
.Y(n_5074)
);

AOI221xp5_ASAP7_75t_L g5075 ( 
.A1(n_4935),
.A2(n_329),
.B1(n_327),
.B2(n_328),
.C(n_330),
.Y(n_5075)
);

INVx1_ASAP7_75t_L g5076 ( 
.A(n_4926),
.Y(n_5076)
);

INVx2_ASAP7_75t_SL g5077 ( 
.A(n_4896),
.Y(n_5077)
);

OAI22xp5_ASAP7_75t_L g5078 ( 
.A1(n_4951),
.A2(n_333),
.B1(n_330),
.B2(n_332),
.Y(n_5078)
);

INVx1_ASAP7_75t_L g5079 ( 
.A(n_4944),
.Y(n_5079)
);

AOI222xp33_ASAP7_75t_L g5080 ( 
.A1(n_4974),
.A2(n_332),
.B1(n_335),
.B2(n_336),
.C1(n_337),
.C2(n_340),
.Y(n_5080)
);

OAI221xp5_ASAP7_75t_L g5081 ( 
.A1(n_4977),
.A2(n_343),
.B1(n_337),
.B2(n_341),
.C(n_344),
.Y(n_5081)
);

OR2x2_ASAP7_75t_L g5082 ( 
.A(n_4952),
.B(n_341),
.Y(n_5082)
);

OAI22xp5_ASAP7_75t_L g5083 ( 
.A1(n_4905),
.A2(n_346),
.B1(n_344),
.B2(n_345),
.Y(n_5083)
);

INVx1_ASAP7_75t_L g5084 ( 
.A(n_4954),
.Y(n_5084)
);

AND2x2_ASAP7_75t_L g5085 ( 
.A(n_4929),
.B(n_347),
.Y(n_5085)
);

AOI322xp5_ASAP7_75t_L g5086 ( 
.A1(n_4943),
.A2(n_4892),
.A3(n_4910),
.B1(n_4920),
.B2(n_4958),
.C1(n_4868),
.C2(n_4957),
.Y(n_5086)
);

INVx3_ASAP7_75t_L g5087 ( 
.A(n_4841),
.Y(n_5087)
);

INVx1_ASAP7_75t_L g5088 ( 
.A(n_4968),
.Y(n_5088)
);

INVx1_ASAP7_75t_L g5089 ( 
.A(n_4911),
.Y(n_5089)
);

HB1xp67_ASAP7_75t_L g5090 ( 
.A(n_4922),
.Y(n_5090)
);

OAI21xp33_ASAP7_75t_L g5091 ( 
.A1(n_4841),
.A2(n_350),
.B(n_351),
.Y(n_5091)
);

OAI211xp5_ASAP7_75t_L g5092 ( 
.A1(n_4916),
.A2(n_353),
.B(n_351),
.C(n_352),
.Y(n_5092)
);

AOI211xp5_ASAP7_75t_L g5093 ( 
.A1(n_4851),
.A2(n_354),
.B(n_352),
.C(n_353),
.Y(n_5093)
);

INVx1_ASAP7_75t_L g5094 ( 
.A(n_4978),
.Y(n_5094)
);

BUFx6f_ASAP7_75t_L g5095 ( 
.A(n_4914),
.Y(n_5095)
);

AOI222xp33_ASAP7_75t_SL g5096 ( 
.A1(n_4907),
.A2(n_355),
.B1(n_356),
.B2(n_358),
.C1(n_360),
.C2(n_361),
.Y(n_5096)
);

NAND2xp5_ASAP7_75t_SL g5097 ( 
.A(n_4937),
.B(n_355),
.Y(n_5097)
);

AOI22xp33_ASAP7_75t_L g5098 ( 
.A1(n_4955),
.A2(n_360),
.B1(n_356),
.B2(n_358),
.Y(n_5098)
);

AOI22xp33_ASAP7_75t_L g5099 ( 
.A1(n_4955),
.A2(n_4873),
.B1(n_4856),
.B2(n_4846),
.Y(n_5099)
);

INVxp67_ASAP7_75t_SL g5100 ( 
.A(n_4846),
.Y(n_5100)
);

AOI22xp33_ASAP7_75t_L g5101 ( 
.A1(n_4955),
.A2(n_364),
.B1(n_362),
.B2(n_363),
.Y(n_5101)
);

AOI222xp33_ASAP7_75t_L g5102 ( 
.A1(n_4937),
.A2(n_363),
.B1(n_364),
.B2(n_365),
.C1(n_367),
.C2(n_368),
.Y(n_5102)
);

AOI22xp33_ASAP7_75t_SL g5103 ( 
.A1(n_4897),
.A2(n_368),
.B1(n_365),
.B2(n_367),
.Y(n_5103)
);

INVx2_ASAP7_75t_L g5104 ( 
.A(n_4924),
.Y(n_5104)
);

OR2x2_ASAP7_75t_L g5105 ( 
.A(n_4871),
.B(n_369),
.Y(n_5105)
);

OAI22xp5_ASAP7_75t_L g5106 ( 
.A1(n_4904),
.A2(n_372),
.B1(n_369),
.B2(n_371),
.Y(n_5106)
);

INVx3_ASAP7_75t_L g5107 ( 
.A(n_4850),
.Y(n_5107)
);

AOI21xp33_ASAP7_75t_L g5108 ( 
.A1(n_4871),
.A2(n_371),
.B(n_373),
.Y(n_5108)
);

AOI22xp33_ASAP7_75t_L g5109 ( 
.A1(n_4885),
.A2(n_375),
.B1(n_373),
.B2(n_374),
.Y(n_5109)
);

AOI21x1_ASAP7_75t_L g5110 ( 
.A1(n_4972),
.A2(n_4946),
.B(n_4900),
.Y(n_5110)
);

INVx2_ASAP7_75t_SL g5111 ( 
.A(n_4861),
.Y(n_5111)
);

AOI21xp5_ASAP7_75t_L g5112 ( 
.A1(n_4972),
.A2(n_4938),
.B(n_4859),
.Y(n_5112)
);

AOI22xp33_ASAP7_75t_L g5113 ( 
.A1(n_4947),
.A2(n_376),
.B1(n_374),
.B2(n_375),
.Y(n_5113)
);

INVx1_ASAP7_75t_L g5114 ( 
.A(n_4884),
.Y(n_5114)
);

AOI22xp33_ASAP7_75t_L g5115 ( 
.A1(n_4899),
.A2(n_378),
.B1(n_376),
.B2(n_377),
.Y(n_5115)
);

OAI221xp5_ASAP7_75t_L g5116 ( 
.A1(n_4971),
.A2(n_377),
.B1(n_378),
.B2(n_379),
.C(n_381),
.Y(n_5116)
);

INVx2_ASAP7_75t_L g5117 ( 
.A(n_4850),
.Y(n_5117)
);

OAI211xp5_ASAP7_75t_L g5118 ( 
.A1(n_4850),
.A2(n_383),
.B(n_381),
.C(n_382),
.Y(n_5118)
);

AND2x4_ASAP7_75t_L g5119 ( 
.A(n_4981),
.B(n_4859),
.Y(n_5119)
);

NAND2xp33_ASAP7_75t_R g5120 ( 
.A(n_5058),
.B(n_382),
.Y(n_5120)
);

NOR2xp33_ASAP7_75t_R g5121 ( 
.A(n_5034),
.B(n_4950),
.Y(n_5121)
);

NAND2xp5_ASAP7_75t_L g5122 ( 
.A(n_5090),
.B(n_4859),
.Y(n_5122)
);

NAND2xp33_ASAP7_75t_R g5123 ( 
.A(n_5058),
.B(n_383),
.Y(n_5123)
);

INVxp67_ASAP7_75t_L g5124 ( 
.A(n_5006),
.Y(n_5124)
);

NAND2xp5_ASAP7_75t_L g5125 ( 
.A(n_5009),
.B(n_4887),
.Y(n_5125)
);

NAND2xp5_ASAP7_75t_L g5126 ( 
.A(n_4984),
.B(n_4887),
.Y(n_5126)
);

CKINVDCx11_ASAP7_75t_R g5127 ( 
.A(n_5039),
.Y(n_5127)
);

AND2x4_ASAP7_75t_L g5128 ( 
.A(n_5005),
.B(n_384),
.Y(n_5128)
);

CKINVDCx12_ASAP7_75t_R g5129 ( 
.A(n_5051),
.Y(n_5129)
);

NAND2xp33_ASAP7_75t_R g5130 ( 
.A(n_5066),
.B(n_384),
.Y(n_5130)
);

NAND2xp33_ASAP7_75t_R g5131 ( 
.A(n_5066),
.B(n_386),
.Y(n_5131)
);

NAND2xp5_ASAP7_75t_L g5132 ( 
.A(n_4986),
.B(n_386),
.Y(n_5132)
);

NAND2xp33_ASAP7_75t_R g5133 ( 
.A(n_5006),
.B(n_387),
.Y(n_5133)
);

BUFx10_ASAP7_75t_L g5134 ( 
.A(n_5045),
.Y(n_5134)
);

NAND2xp33_ASAP7_75t_R g5135 ( 
.A(n_5051),
.B(n_387),
.Y(n_5135)
);

NOR2xp33_ASAP7_75t_R g5136 ( 
.A(n_5070),
.B(n_388),
.Y(n_5136)
);

XNOR2xp5_ASAP7_75t_L g5137 ( 
.A(n_5010),
.B(n_388),
.Y(n_5137)
);

NOR2xp33_ASAP7_75t_R g5138 ( 
.A(n_5077),
.B(n_389),
.Y(n_5138)
);

INVxp67_ASAP7_75t_L g5139 ( 
.A(n_5002),
.Y(n_5139)
);

AND2x2_ASAP7_75t_L g5140 ( 
.A(n_5005),
.B(n_390),
.Y(n_5140)
);

XNOR2xp5_ASAP7_75t_L g5141 ( 
.A(n_5071),
.B(n_390),
.Y(n_5141)
);

NAND2xp33_ASAP7_75t_R g5142 ( 
.A(n_5067),
.B(n_391),
.Y(n_5142)
);

NOR2xp33_ASAP7_75t_SL g5143 ( 
.A(n_5062),
.B(n_392),
.Y(n_5143)
);

AND2x4_ASAP7_75t_L g5144 ( 
.A(n_4979),
.B(n_4989),
.Y(n_5144)
);

NAND2xp33_ASAP7_75t_R g5145 ( 
.A(n_5067),
.B(n_392),
.Y(n_5145)
);

NOR2xp33_ASAP7_75t_R g5146 ( 
.A(n_5052),
.B(n_393),
.Y(n_5146)
);

BUFx12f_ASAP7_75t_L g5147 ( 
.A(n_5062),
.Y(n_5147)
);

CKINVDCx20_ASAP7_75t_R g5148 ( 
.A(n_5031),
.Y(n_5148)
);

BUFx3_ASAP7_75t_L g5149 ( 
.A(n_5072),
.Y(n_5149)
);

OR2x4_ASAP7_75t_L g5150 ( 
.A(n_4993),
.B(n_393),
.Y(n_5150)
);

NOR2xp33_ASAP7_75t_R g5151 ( 
.A(n_5014),
.B(n_394),
.Y(n_5151)
);

INVx2_ASAP7_75t_L g5152 ( 
.A(n_5095),
.Y(n_5152)
);

NAND2xp5_ASAP7_75t_SL g5153 ( 
.A(n_4996),
.B(n_5099),
.Y(n_5153)
);

INVx1_ASAP7_75t_L g5154 ( 
.A(n_4998),
.Y(n_5154)
);

AND2x4_ASAP7_75t_L g5155 ( 
.A(n_5110),
.B(n_395),
.Y(n_5155)
);

INVx2_ASAP7_75t_L g5156 ( 
.A(n_5095),
.Y(n_5156)
);

NAND2xp33_ASAP7_75t_R g5157 ( 
.A(n_5016),
.B(n_395),
.Y(n_5157)
);

NAND2xp33_ASAP7_75t_R g5158 ( 
.A(n_5016),
.B(n_396),
.Y(n_5158)
);

NOR2xp33_ASAP7_75t_R g5159 ( 
.A(n_5111),
.B(n_397),
.Y(n_5159)
);

AND2x4_ASAP7_75t_L g5160 ( 
.A(n_5112),
.B(n_4991),
.Y(n_5160)
);

OR2x6_ASAP7_75t_L g5161 ( 
.A(n_5040),
.B(n_397),
.Y(n_5161)
);

NAND2xp5_ASAP7_75t_L g5162 ( 
.A(n_5011),
.B(n_398),
.Y(n_5162)
);

NAND2xp5_ASAP7_75t_L g5163 ( 
.A(n_5022),
.B(n_399),
.Y(n_5163)
);

NOR2xp33_ASAP7_75t_R g5164 ( 
.A(n_5046),
.B(n_399),
.Y(n_5164)
);

AND2x4_ASAP7_75t_L g5165 ( 
.A(n_4991),
.B(n_400),
.Y(n_5165)
);

NOR2xp33_ASAP7_75t_R g5166 ( 
.A(n_5036),
.B(n_400),
.Y(n_5166)
);

XNOR2xp5_ASAP7_75t_L g5167 ( 
.A(n_4987),
.B(n_4994),
.Y(n_5167)
);

INVx2_ASAP7_75t_L g5168 ( 
.A(n_5095),
.Y(n_5168)
);

NOR2xp33_ASAP7_75t_R g5169 ( 
.A(n_5060),
.B(n_401),
.Y(n_5169)
);

NAND2xp33_ASAP7_75t_R g5170 ( 
.A(n_5050),
.B(n_402),
.Y(n_5170)
);

AND2x4_ASAP7_75t_L g5171 ( 
.A(n_5017),
.B(n_402),
.Y(n_5171)
);

NAND2xp33_ASAP7_75t_R g5172 ( 
.A(n_5050),
.B(n_403),
.Y(n_5172)
);

NOR2xp33_ASAP7_75t_R g5173 ( 
.A(n_5085),
.B(n_403),
.Y(n_5173)
);

AND2x4_ASAP7_75t_L g5174 ( 
.A(n_5100),
.B(n_404),
.Y(n_5174)
);

INVxp67_ASAP7_75t_L g5175 ( 
.A(n_5114),
.Y(n_5175)
);

NAND2xp33_ASAP7_75t_R g5176 ( 
.A(n_5105),
.B(n_404),
.Y(n_5176)
);

NAND2xp33_ASAP7_75t_R g5177 ( 
.A(n_5107),
.B(n_405),
.Y(n_5177)
);

AND2x4_ASAP7_75t_L g5178 ( 
.A(n_5087),
.B(n_405),
.Y(n_5178)
);

INVx2_ASAP7_75t_L g5179 ( 
.A(n_5022),
.Y(n_5179)
);

NAND2xp5_ASAP7_75t_SL g5180 ( 
.A(n_5020),
.B(n_406),
.Y(n_5180)
);

NAND2xp5_ASAP7_75t_L g5181 ( 
.A(n_5054),
.B(n_406),
.Y(n_5181)
);

AND2x4_ASAP7_75t_L g5182 ( 
.A(n_5087),
.B(n_407),
.Y(n_5182)
);

XNOR2xp5_ASAP7_75t_L g5183 ( 
.A(n_5093),
.B(n_407),
.Y(n_5183)
);

XOR2xp5_ASAP7_75t_L g5184 ( 
.A(n_5103),
.B(n_408),
.Y(n_5184)
);

OR2x6_ASAP7_75t_L g5185 ( 
.A(n_5037),
.B(n_409),
.Y(n_5185)
);

INVx2_ASAP7_75t_L g5186 ( 
.A(n_5000),
.Y(n_5186)
);

AND2x4_ASAP7_75t_L g5187 ( 
.A(n_5117),
.B(n_410),
.Y(n_5187)
);

AND2x4_ASAP7_75t_L g5188 ( 
.A(n_5107),
.B(n_413),
.Y(n_5188)
);

NAND2xp33_ASAP7_75t_R g5189 ( 
.A(n_5064),
.B(n_414),
.Y(n_5189)
);

BUFx8_ASAP7_75t_SL g5190 ( 
.A(n_5038),
.Y(n_5190)
);

NAND2xp33_ASAP7_75t_R g5191 ( 
.A(n_5114),
.B(n_415),
.Y(n_5191)
);

BUFx3_ASAP7_75t_L g5192 ( 
.A(n_5053),
.Y(n_5192)
);

BUFx2_ASAP7_75t_L g5193 ( 
.A(n_5018),
.Y(n_5193)
);

NOR2xp33_ASAP7_75t_R g5194 ( 
.A(n_5047),
.B(n_415),
.Y(n_5194)
);

INVx1_ASAP7_75t_L g5195 ( 
.A(n_5073),
.Y(n_5195)
);

INVx1_ASAP7_75t_L g5196 ( 
.A(n_5007),
.Y(n_5196)
);

NAND2xp33_ASAP7_75t_R g5197 ( 
.A(n_5026),
.B(n_416),
.Y(n_5197)
);

INVx1_ASAP7_75t_L g5198 ( 
.A(n_5007),
.Y(n_5198)
);

AND2x4_ASAP7_75t_L g5199 ( 
.A(n_5055),
.B(n_416),
.Y(n_5199)
);

NAND2xp33_ASAP7_75t_R g5200 ( 
.A(n_5082),
.B(n_4995),
.Y(n_5200)
);

NOR2xp33_ASAP7_75t_R g5201 ( 
.A(n_5113),
.B(n_417),
.Y(n_5201)
);

NAND2xp33_ASAP7_75t_R g5202 ( 
.A(n_4997),
.B(n_418),
.Y(n_5202)
);

NAND2xp5_ASAP7_75t_L g5203 ( 
.A(n_5019),
.B(n_418),
.Y(n_5203)
);

INVxp67_ASAP7_75t_L g5204 ( 
.A(n_5049),
.Y(n_5204)
);

OR2x6_ASAP7_75t_L g5205 ( 
.A(n_5097),
.B(n_420),
.Y(n_5205)
);

NAND2xp33_ASAP7_75t_R g5206 ( 
.A(n_4997),
.B(n_421),
.Y(n_5206)
);

XNOR2xp5_ASAP7_75t_L g5207 ( 
.A(n_5083),
.B(n_422),
.Y(n_5207)
);

CKINVDCx11_ASAP7_75t_R g5208 ( 
.A(n_5106),
.Y(n_5208)
);

NAND2xp33_ASAP7_75t_R g5209 ( 
.A(n_5000),
.B(n_424),
.Y(n_5209)
);

AND2x2_ASAP7_75t_L g5210 ( 
.A(n_5004),
.B(n_426),
.Y(n_5210)
);

INVxp67_ASAP7_75t_L g5211 ( 
.A(n_5049),
.Y(n_5211)
);

XNOR2xp5_ASAP7_75t_L g5212 ( 
.A(n_4988),
.B(n_427),
.Y(n_5212)
);

AND2x2_ASAP7_75t_L g5213 ( 
.A(n_4980),
.B(n_5061),
.Y(n_5213)
);

AND2x4_ASAP7_75t_L g5214 ( 
.A(n_5055),
.B(n_427),
.Y(n_5214)
);

NAND2xp33_ASAP7_75t_R g5215 ( 
.A(n_5063),
.B(n_428),
.Y(n_5215)
);

BUFx3_ASAP7_75t_L g5216 ( 
.A(n_5021),
.Y(n_5216)
);

AND2x2_ASAP7_75t_L g5217 ( 
.A(n_5003),
.B(n_428),
.Y(n_5217)
);

AND2x2_ASAP7_75t_L g5218 ( 
.A(n_5008),
.B(n_429),
.Y(n_5218)
);

NAND2xp33_ASAP7_75t_R g5219 ( 
.A(n_4990),
.B(n_430),
.Y(n_5219)
);

NOR2xp33_ASAP7_75t_R g5220 ( 
.A(n_5043),
.B(n_430),
.Y(n_5220)
);

AND2x4_ASAP7_75t_L g5221 ( 
.A(n_5015),
.B(n_431),
.Y(n_5221)
);

NAND2xp5_ASAP7_75t_L g5222 ( 
.A(n_5001),
.B(n_5056),
.Y(n_5222)
);

OR2x2_ASAP7_75t_L g5223 ( 
.A(n_5069),
.B(n_431),
.Y(n_5223)
);

INVx1_ASAP7_75t_L g5224 ( 
.A(n_5076),
.Y(n_5224)
);

NAND2xp5_ASAP7_75t_L g5225 ( 
.A(n_5079),
.B(n_432),
.Y(n_5225)
);

XNOR2xp5_ASAP7_75t_L g5226 ( 
.A(n_4983),
.B(n_433),
.Y(n_5226)
);

INVx2_ASAP7_75t_L g5227 ( 
.A(n_5186),
.Y(n_5227)
);

NAND2xp5_ASAP7_75t_L g5228 ( 
.A(n_5163),
.B(n_4992),
.Y(n_5228)
);

AND2x2_ASAP7_75t_L g5229 ( 
.A(n_5193),
.B(n_5084),
.Y(n_5229)
);

AND2x2_ASAP7_75t_L g5230 ( 
.A(n_5160),
.B(n_5088),
.Y(n_5230)
);

AO21x2_ASAP7_75t_L g5231 ( 
.A1(n_5126),
.A2(n_5035),
.B(n_5024),
.Y(n_5231)
);

AND2x2_ASAP7_75t_L g5232 ( 
.A(n_5175),
.B(n_5149),
.Y(n_5232)
);

INVx1_ASAP7_75t_L g5233 ( 
.A(n_5196),
.Y(n_5233)
);

INVx1_ASAP7_75t_L g5234 ( 
.A(n_5224),
.Y(n_5234)
);

INVx1_ASAP7_75t_L g5235 ( 
.A(n_5198),
.Y(n_5235)
);

AND2x2_ASAP7_75t_L g5236 ( 
.A(n_5119),
.B(n_5029),
.Y(n_5236)
);

OR2x2_ASAP7_75t_L g5237 ( 
.A(n_5154),
.B(n_5033),
.Y(n_5237)
);

INVx2_ASAP7_75t_L g5238 ( 
.A(n_5192),
.Y(n_5238)
);

INVx3_ASAP7_75t_L g5239 ( 
.A(n_5147),
.Y(n_5239)
);

OR2x2_ASAP7_75t_L g5240 ( 
.A(n_5195),
.B(n_5012),
.Y(n_5240)
);

HB1xp67_ASAP7_75t_L g5241 ( 
.A(n_5223),
.Y(n_5241)
);

HB1xp67_ASAP7_75t_L g5242 ( 
.A(n_5124),
.Y(n_5242)
);

INVx2_ASAP7_75t_L g5243 ( 
.A(n_5204),
.Y(n_5243)
);

INVx4_ASAP7_75t_L g5244 ( 
.A(n_5127),
.Y(n_5244)
);

NAND2xp5_ASAP7_75t_L g5245 ( 
.A(n_5211),
.B(n_5027),
.Y(n_5245)
);

NAND2xp5_ASAP7_75t_L g5246 ( 
.A(n_5199),
.B(n_5086),
.Y(n_5246)
);

INVx2_ASAP7_75t_L g5247 ( 
.A(n_5199),
.Y(n_5247)
);

BUFx3_ASAP7_75t_L g5248 ( 
.A(n_5148),
.Y(n_5248)
);

INVx1_ASAP7_75t_L g5249 ( 
.A(n_5132),
.Y(n_5249)
);

AND2x2_ASAP7_75t_L g5250 ( 
.A(n_5153),
.B(n_5023),
.Y(n_5250)
);

AND2x2_ASAP7_75t_L g5251 ( 
.A(n_5213),
.B(n_4985),
.Y(n_5251)
);

NAND2xp5_ASAP7_75t_L g5252 ( 
.A(n_5214),
.B(n_5091),
.Y(n_5252)
);

NAND2xp5_ASAP7_75t_L g5253 ( 
.A(n_5214),
.B(n_5030),
.Y(n_5253)
);

AND2x2_ASAP7_75t_L g5254 ( 
.A(n_5171),
.B(n_5032),
.Y(n_5254)
);

AND2x2_ASAP7_75t_L g5255 ( 
.A(n_5122),
.B(n_5013),
.Y(n_5255)
);

OR2x2_ASAP7_75t_L g5256 ( 
.A(n_5222),
.B(n_5089),
.Y(n_5256)
);

NAND3xp33_ASAP7_75t_L g5257 ( 
.A(n_5139),
.B(n_5096),
.C(n_5057),
.Y(n_5257)
);

OR2x2_ASAP7_75t_L g5258 ( 
.A(n_5125),
.B(n_5028),
.Y(n_5258)
);

INVx2_ASAP7_75t_L g5259 ( 
.A(n_5155),
.Y(n_5259)
);

INVx4_ASAP7_75t_L g5260 ( 
.A(n_5161),
.Y(n_5260)
);

OR2x2_ASAP7_75t_L g5261 ( 
.A(n_5162),
.B(n_5094),
.Y(n_5261)
);

INVx2_ASAP7_75t_L g5262 ( 
.A(n_5174),
.Y(n_5262)
);

INVx1_ASAP7_75t_L g5263 ( 
.A(n_5225),
.Y(n_5263)
);

INVx2_ASAP7_75t_L g5264 ( 
.A(n_5174),
.Y(n_5264)
);

INVx2_ASAP7_75t_L g5265 ( 
.A(n_5179),
.Y(n_5265)
);

BUFx2_ASAP7_75t_L g5266 ( 
.A(n_5150),
.Y(n_5266)
);

INVx1_ASAP7_75t_L g5267 ( 
.A(n_5217),
.Y(n_5267)
);

INVx1_ASAP7_75t_L g5268 ( 
.A(n_5218),
.Y(n_5268)
);

INVx2_ASAP7_75t_L g5269 ( 
.A(n_5144),
.Y(n_5269)
);

INVx1_ASAP7_75t_L g5270 ( 
.A(n_5203),
.Y(n_5270)
);

AND2x2_ASAP7_75t_L g5271 ( 
.A(n_5210),
.B(n_5108),
.Y(n_5271)
);

HB1xp67_ASAP7_75t_L g5272 ( 
.A(n_5152),
.Y(n_5272)
);

INVx2_ASAP7_75t_SL g5273 ( 
.A(n_5134),
.Y(n_5273)
);

OR2x2_ASAP7_75t_L g5274 ( 
.A(n_5156),
.B(n_4982),
.Y(n_5274)
);

AND2x2_ASAP7_75t_L g5275 ( 
.A(n_5221),
.B(n_4982),
.Y(n_5275)
);

AND2x2_ASAP7_75t_L g5276 ( 
.A(n_5140),
.B(n_5168),
.Y(n_5276)
);

AND2x2_ASAP7_75t_L g5277 ( 
.A(n_5178),
.B(n_5042),
.Y(n_5277)
);

BUFx2_ASAP7_75t_L g5278 ( 
.A(n_5121),
.Y(n_5278)
);

INVx1_ASAP7_75t_L g5279 ( 
.A(n_5181),
.Y(n_5279)
);

INVx1_ASAP7_75t_L g5280 ( 
.A(n_5129),
.Y(n_5280)
);

NAND2xp5_ASAP7_75t_L g5281 ( 
.A(n_5178),
.B(n_4999),
.Y(n_5281)
);

INVxp67_ASAP7_75t_SL g5282 ( 
.A(n_5157),
.Y(n_5282)
);

AND2x2_ASAP7_75t_L g5283 ( 
.A(n_5182),
.B(n_5104),
.Y(n_5283)
);

INVx1_ASAP7_75t_L g5284 ( 
.A(n_5182),
.Y(n_5284)
);

HB1xp67_ASAP7_75t_L g5285 ( 
.A(n_5141),
.Y(n_5285)
);

INVx2_ASAP7_75t_L g5286 ( 
.A(n_5161),
.Y(n_5286)
);

BUFx6f_ASAP7_75t_L g5287 ( 
.A(n_5185),
.Y(n_5287)
);

HB1xp67_ASAP7_75t_L g5288 ( 
.A(n_5200),
.Y(n_5288)
);

INVx2_ASAP7_75t_L g5289 ( 
.A(n_5185),
.Y(n_5289)
);

BUFx2_ASAP7_75t_L g5290 ( 
.A(n_5190),
.Y(n_5290)
);

INVx2_ASAP7_75t_L g5291 ( 
.A(n_5205),
.Y(n_5291)
);

INVx2_ASAP7_75t_SL g5292 ( 
.A(n_5165),
.Y(n_5292)
);

OR2x6_ASAP7_75t_L g5293 ( 
.A(n_5180),
.B(n_5074),
.Y(n_5293)
);

INVx1_ASAP7_75t_L g5294 ( 
.A(n_5187),
.Y(n_5294)
);

INVx1_ASAP7_75t_L g5295 ( 
.A(n_5216),
.Y(n_5295)
);

INVx1_ASAP7_75t_L g5296 ( 
.A(n_5188),
.Y(n_5296)
);

INVx2_ASAP7_75t_L g5297 ( 
.A(n_5205),
.Y(n_5297)
);

NAND2xp33_ASAP7_75t_SL g5298 ( 
.A(n_5158),
.B(n_5098),
.Y(n_5298)
);

AND2x4_ASAP7_75t_L g5299 ( 
.A(n_5128),
.B(n_5044),
.Y(n_5299)
);

INVx2_ASAP7_75t_L g5300 ( 
.A(n_5208),
.Y(n_5300)
);

CKINVDCx8_ASAP7_75t_R g5301 ( 
.A(n_5215),
.Y(n_5301)
);

AND2x2_ASAP7_75t_L g5302 ( 
.A(n_5167),
.B(n_5065),
.Y(n_5302)
);

NAND2xp5_ASAP7_75t_L g5303 ( 
.A(n_5164),
.B(n_5025),
.Y(n_5303)
);

NAND3xp33_ASAP7_75t_L g5304 ( 
.A(n_5288),
.B(n_5189),
.C(n_5197),
.Y(n_5304)
);

HB1xp67_ASAP7_75t_L g5305 ( 
.A(n_5242),
.Y(n_5305)
);

AOI22xp33_ASAP7_75t_L g5306 ( 
.A1(n_5250),
.A2(n_5183),
.B1(n_5201),
.B2(n_5226),
.Y(n_5306)
);

AND2x2_ASAP7_75t_SL g5307 ( 
.A(n_5266),
.B(n_5143),
.Y(n_5307)
);

AND2x2_ASAP7_75t_L g5308 ( 
.A(n_5290),
.B(n_5151),
.Y(n_5308)
);

OAI22xp5_ASAP7_75t_L g5309 ( 
.A1(n_5266),
.A2(n_5207),
.B1(n_5137),
.B2(n_5212),
.Y(n_5309)
);

NAND2xp5_ASAP7_75t_L g5310 ( 
.A(n_5241),
.B(n_5166),
.Y(n_5310)
);

NAND2xp5_ASAP7_75t_L g5311 ( 
.A(n_5267),
.B(n_5194),
.Y(n_5311)
);

AND2x2_ASAP7_75t_L g5312 ( 
.A(n_5232),
.B(n_5138),
.Y(n_5312)
);

NAND3xp33_ASAP7_75t_L g5313 ( 
.A(n_5257),
.B(n_5191),
.C(n_5209),
.Y(n_5313)
);

AND2x2_ASAP7_75t_L g5314 ( 
.A(n_5232),
.B(n_5159),
.Y(n_5314)
);

AND2x2_ASAP7_75t_L g5315 ( 
.A(n_5290),
.B(n_5146),
.Y(n_5315)
);

AND2x2_ASAP7_75t_L g5316 ( 
.A(n_5244),
.B(n_5136),
.Y(n_5316)
);

NAND2xp5_ASAP7_75t_L g5317 ( 
.A(n_5268),
.B(n_5173),
.Y(n_5317)
);

AOI22xp33_ASAP7_75t_L g5318 ( 
.A1(n_5250),
.A2(n_5184),
.B1(n_5220),
.B2(n_5116),
.Y(n_5318)
);

OA21x2_ASAP7_75t_L g5319 ( 
.A1(n_5245),
.A2(n_5075),
.B(n_5048),
.Y(n_5319)
);

AND2x2_ASAP7_75t_L g5320 ( 
.A(n_5230),
.B(n_5169),
.Y(n_5320)
);

NAND2xp5_ASAP7_75t_L g5321 ( 
.A(n_5238),
.B(n_5102),
.Y(n_5321)
);

AND2x2_ASAP7_75t_L g5322 ( 
.A(n_5244),
.B(n_5101),
.Y(n_5322)
);

NAND3xp33_ASAP7_75t_L g5323 ( 
.A(n_5293),
.B(n_5219),
.C(n_5142),
.Y(n_5323)
);

OA21x2_ASAP7_75t_L g5324 ( 
.A1(n_5243),
.A2(n_5303),
.B(n_5246),
.Y(n_5324)
);

NAND2xp5_ASAP7_75t_L g5325 ( 
.A(n_5238),
.B(n_5059),
.Y(n_5325)
);

AND2x2_ASAP7_75t_L g5326 ( 
.A(n_5244),
.B(n_5300),
.Y(n_5326)
);

OAI221xp5_ASAP7_75t_L g5327 ( 
.A1(n_5301),
.A2(n_5177),
.B1(n_5135),
.B2(n_5145),
.C(n_5172),
.Y(n_5327)
);

NAND2xp5_ASAP7_75t_L g5328 ( 
.A(n_5271),
.B(n_5078),
.Y(n_5328)
);

AND2x2_ASAP7_75t_L g5329 ( 
.A(n_5300),
.B(n_5041),
.Y(n_5329)
);

NOR2xp33_ASAP7_75t_L g5330 ( 
.A(n_5248),
.B(n_5092),
.Y(n_5330)
);

NAND2xp5_ASAP7_75t_L g5331 ( 
.A(n_5271),
.B(n_5080),
.Y(n_5331)
);

NAND2xp5_ASAP7_75t_L g5332 ( 
.A(n_5279),
.B(n_5068),
.Y(n_5332)
);

NAND2xp5_ASAP7_75t_L g5333 ( 
.A(n_5279),
.B(n_5270),
.Y(n_5333)
);

NAND3xp33_ASAP7_75t_L g5334 ( 
.A(n_5293),
.B(n_5170),
.C(n_5133),
.Y(n_5334)
);

NAND2x1_ASAP7_75t_L g5335 ( 
.A(n_5260),
.B(n_5120),
.Y(n_5335)
);

OAI22xp5_ASAP7_75t_L g5336 ( 
.A1(n_5258),
.A2(n_5109),
.B1(n_5115),
.B2(n_5081),
.Y(n_5336)
);

NAND2xp5_ASAP7_75t_L g5337 ( 
.A(n_5249),
.B(n_5118),
.Y(n_5337)
);

AOI22xp33_ASAP7_75t_SL g5338 ( 
.A1(n_5258),
.A2(n_5176),
.B1(n_5130),
.B2(n_5131),
.Y(n_5338)
);

NAND2xp5_ASAP7_75t_L g5339 ( 
.A(n_5249),
.B(n_5123),
.Y(n_5339)
);

NAND3xp33_ASAP7_75t_L g5340 ( 
.A(n_5293),
.B(n_5206),
.C(n_5202),
.Y(n_5340)
);

NAND3xp33_ASAP7_75t_L g5341 ( 
.A(n_5293),
.B(n_435),
.C(n_437),
.Y(n_5341)
);

AND2x2_ASAP7_75t_L g5342 ( 
.A(n_5230),
.B(n_435),
.Y(n_5342)
);

BUFx2_ASAP7_75t_L g5343 ( 
.A(n_5248),
.Y(n_5343)
);

NAND3xp33_ASAP7_75t_L g5344 ( 
.A(n_5298),
.B(n_438),
.C(n_439),
.Y(n_5344)
);

NAND3xp33_ASAP7_75t_L g5345 ( 
.A(n_5298),
.B(n_438),
.C(n_442),
.Y(n_5345)
);

NAND3xp33_ASAP7_75t_L g5346 ( 
.A(n_5301),
.B(n_443),
.C(n_444),
.Y(n_5346)
);

OAI21xp33_ASAP7_75t_L g5347 ( 
.A1(n_5240),
.A2(n_443),
.B(n_445),
.Y(n_5347)
);

NAND4xp25_ASAP7_75t_L g5348 ( 
.A(n_5278),
.B(n_448),
.C(n_446),
.D(n_447),
.Y(n_5348)
);

AND2x2_ASAP7_75t_L g5349 ( 
.A(n_5273),
.B(n_447),
.Y(n_5349)
);

AND2x2_ASAP7_75t_L g5350 ( 
.A(n_5273),
.B(n_450),
.Y(n_5350)
);

AND2x2_ASAP7_75t_L g5351 ( 
.A(n_5236),
.B(n_450),
.Y(n_5351)
);

NAND3xp33_ASAP7_75t_L g5352 ( 
.A(n_5240),
.B(n_451),
.C(n_452),
.Y(n_5352)
);

NAND2xp5_ASAP7_75t_L g5353 ( 
.A(n_5247),
.B(n_451),
.Y(n_5353)
);

NAND2xp5_ASAP7_75t_L g5354 ( 
.A(n_5247),
.B(n_453),
.Y(n_5354)
);

INVx2_ASAP7_75t_L g5355 ( 
.A(n_5343),
.Y(n_5355)
);

NAND2xp5_ASAP7_75t_L g5356 ( 
.A(n_5351),
.B(n_5262),
.Y(n_5356)
);

INVx1_ASAP7_75t_L g5357 ( 
.A(n_5305),
.Y(n_5357)
);

INVx2_ASAP7_75t_SL g5358 ( 
.A(n_5326),
.Y(n_5358)
);

INVx1_ASAP7_75t_L g5359 ( 
.A(n_5305),
.Y(n_5359)
);

INVx2_ASAP7_75t_L g5360 ( 
.A(n_5307),
.Y(n_5360)
);

OAI221xp5_ASAP7_75t_SL g5361 ( 
.A1(n_5323),
.A2(n_5281),
.B1(n_5282),
.B2(n_5302),
.C(n_5243),
.Y(n_5361)
);

OR2x2_ASAP7_75t_L g5362 ( 
.A(n_5333),
.B(n_5325),
.Y(n_5362)
);

BUFx3_ASAP7_75t_L g5363 ( 
.A(n_5316),
.Y(n_5363)
);

INVx4_ASAP7_75t_L g5364 ( 
.A(n_5349),
.Y(n_5364)
);

OR2x2_ASAP7_75t_L g5365 ( 
.A(n_5328),
.B(n_5263),
.Y(n_5365)
);

OR2x2_ASAP7_75t_SL g5366 ( 
.A(n_5304),
.B(n_5287),
.Y(n_5366)
);

AOI22xp5_ASAP7_75t_L g5367 ( 
.A1(n_5313),
.A2(n_5251),
.B1(n_5285),
.B2(n_5302),
.Y(n_5367)
);

AND2x2_ASAP7_75t_L g5368 ( 
.A(n_5315),
.B(n_5278),
.Y(n_5368)
);

OR2x2_ASAP7_75t_L g5369 ( 
.A(n_5310),
.B(n_5228),
.Y(n_5369)
);

NOR2xp67_ASAP7_75t_L g5370 ( 
.A(n_5340),
.B(n_5260),
.Y(n_5370)
);

AND2x2_ASAP7_75t_L g5371 ( 
.A(n_5308),
.B(n_5239),
.Y(n_5371)
);

INVx2_ASAP7_75t_L g5372 ( 
.A(n_5307),
.Y(n_5372)
);

NAND2xp5_ASAP7_75t_L g5373 ( 
.A(n_5347),
.B(n_5262),
.Y(n_5373)
);

OR2x2_ASAP7_75t_L g5374 ( 
.A(n_5311),
.B(n_5237),
.Y(n_5374)
);

AND2x4_ASAP7_75t_L g5375 ( 
.A(n_5312),
.B(n_5260),
.Y(n_5375)
);

AOI221xp5_ASAP7_75t_L g5376 ( 
.A1(n_5334),
.A2(n_5295),
.B1(n_5227),
.B2(n_5253),
.C(n_5287),
.Y(n_5376)
);

HB1xp67_ASAP7_75t_L g5377 ( 
.A(n_5319),
.Y(n_5377)
);

NAND3xp33_ASAP7_75t_L g5378 ( 
.A(n_5344),
.B(n_5345),
.C(n_5319),
.Y(n_5378)
);

AND2x2_ASAP7_75t_L g5379 ( 
.A(n_5312),
.B(n_5239),
.Y(n_5379)
);

INVx1_ASAP7_75t_L g5380 ( 
.A(n_5353),
.Y(n_5380)
);

INVx1_ASAP7_75t_L g5381 ( 
.A(n_5354),
.Y(n_5381)
);

NAND2xp5_ASAP7_75t_L g5382 ( 
.A(n_5330),
.B(n_5342),
.Y(n_5382)
);

INVx2_ASAP7_75t_L g5383 ( 
.A(n_5324),
.Y(n_5383)
);

AOI22xp33_ASAP7_75t_L g5384 ( 
.A1(n_5331),
.A2(n_5251),
.B1(n_5287),
.B2(n_5261),
.Y(n_5384)
);

INVx2_ASAP7_75t_L g5385 ( 
.A(n_5324),
.Y(n_5385)
);

INVx5_ASAP7_75t_L g5386 ( 
.A(n_5350),
.Y(n_5386)
);

HB1xp67_ASAP7_75t_L g5387 ( 
.A(n_5319),
.Y(n_5387)
);

OAI22xp5_ASAP7_75t_L g5388 ( 
.A1(n_5338),
.A2(n_5237),
.B1(n_5292),
.B2(n_5252),
.Y(n_5388)
);

AND2x4_ASAP7_75t_L g5389 ( 
.A(n_5363),
.B(n_5320),
.Y(n_5389)
);

HB1xp67_ASAP7_75t_L g5390 ( 
.A(n_5368),
.Y(n_5390)
);

AND2x2_ASAP7_75t_L g5391 ( 
.A(n_5371),
.B(n_5314),
.Y(n_5391)
);

INVx2_ASAP7_75t_L g5392 ( 
.A(n_5383),
.Y(n_5392)
);

AND2x2_ASAP7_75t_L g5393 ( 
.A(n_5379),
.B(n_5314),
.Y(n_5393)
);

AND2x2_ASAP7_75t_L g5394 ( 
.A(n_5363),
.B(n_5239),
.Y(n_5394)
);

NOR2xp67_ASAP7_75t_L g5395 ( 
.A(n_5386),
.B(n_5320),
.Y(n_5395)
);

AND2x2_ASAP7_75t_L g5396 ( 
.A(n_5386),
.B(n_5322),
.Y(n_5396)
);

AND2x2_ASAP7_75t_L g5397 ( 
.A(n_5386),
.B(n_5229),
.Y(n_5397)
);

AND2x2_ASAP7_75t_L g5398 ( 
.A(n_5386),
.B(n_5229),
.Y(n_5398)
);

INVx1_ASAP7_75t_L g5399 ( 
.A(n_5383),
.Y(n_5399)
);

INVx2_ASAP7_75t_L g5400 ( 
.A(n_5385),
.Y(n_5400)
);

INVx1_ASAP7_75t_L g5401 ( 
.A(n_5385),
.Y(n_5401)
);

NAND2xp5_ASAP7_75t_SL g5402 ( 
.A(n_5375),
.B(n_5338),
.Y(n_5402)
);

OR2x2_ASAP7_75t_L g5403 ( 
.A(n_5377),
.B(n_5387),
.Y(n_5403)
);

HB1xp67_ASAP7_75t_L g5404 ( 
.A(n_5355),
.Y(n_5404)
);

BUFx2_ASAP7_75t_L g5405 ( 
.A(n_5364),
.Y(n_5405)
);

INVx1_ASAP7_75t_L g5406 ( 
.A(n_5377),
.Y(n_5406)
);

NAND2xp5_ASAP7_75t_L g5407 ( 
.A(n_5355),
.B(n_5330),
.Y(n_5407)
);

NOR2xp67_ASAP7_75t_L g5408 ( 
.A(n_5364),
.B(n_5280),
.Y(n_5408)
);

INVx1_ASAP7_75t_L g5409 ( 
.A(n_5387),
.Y(n_5409)
);

INVx1_ASAP7_75t_L g5410 ( 
.A(n_5357),
.Y(n_5410)
);

INVx1_ASAP7_75t_L g5411 ( 
.A(n_5359),
.Y(n_5411)
);

AND2x2_ASAP7_75t_L g5412 ( 
.A(n_5375),
.B(n_5236),
.Y(n_5412)
);

INVx1_ASAP7_75t_L g5413 ( 
.A(n_5365),
.Y(n_5413)
);

OR2x2_ASAP7_75t_L g5414 ( 
.A(n_5362),
.B(n_5324),
.Y(n_5414)
);

AND2x2_ASAP7_75t_L g5415 ( 
.A(n_5358),
.B(n_5276),
.Y(n_5415)
);

INVx1_ASAP7_75t_L g5416 ( 
.A(n_5403),
.Y(n_5416)
);

INVx1_ASAP7_75t_L g5417 ( 
.A(n_5403),
.Y(n_5417)
);

INVx1_ASAP7_75t_L g5418 ( 
.A(n_5404),
.Y(n_5418)
);

INVx1_ASAP7_75t_L g5419 ( 
.A(n_5390),
.Y(n_5419)
);

OR2x2_ASAP7_75t_L g5420 ( 
.A(n_5414),
.B(n_5388),
.Y(n_5420)
);

HB1xp67_ASAP7_75t_L g5421 ( 
.A(n_5389),
.Y(n_5421)
);

AND2x4_ASAP7_75t_SL g5422 ( 
.A(n_5389),
.B(n_5280),
.Y(n_5422)
);

AND2x2_ASAP7_75t_L g5423 ( 
.A(n_5391),
.B(n_5370),
.Y(n_5423)
);

INVx1_ASAP7_75t_SL g5424 ( 
.A(n_5391),
.Y(n_5424)
);

AND2x2_ASAP7_75t_L g5425 ( 
.A(n_5393),
.B(n_5382),
.Y(n_5425)
);

BUFx2_ASAP7_75t_L g5426 ( 
.A(n_5389),
.Y(n_5426)
);

INVx2_ASAP7_75t_L g5427 ( 
.A(n_5406),
.Y(n_5427)
);

AND2x2_ASAP7_75t_L g5428 ( 
.A(n_5393),
.B(n_5360),
.Y(n_5428)
);

INVx2_ASAP7_75t_L g5429 ( 
.A(n_5409),
.Y(n_5429)
);

INVx2_ASAP7_75t_L g5430 ( 
.A(n_5414),
.Y(n_5430)
);

AND2x2_ASAP7_75t_L g5431 ( 
.A(n_5394),
.B(n_5360),
.Y(n_5431)
);

INVx1_ASAP7_75t_L g5432 ( 
.A(n_5392),
.Y(n_5432)
);

AND2x2_ASAP7_75t_L g5433 ( 
.A(n_5394),
.B(n_5372),
.Y(n_5433)
);

AND2x2_ASAP7_75t_L g5434 ( 
.A(n_5396),
.B(n_5397),
.Y(n_5434)
);

NAND2xp5_ASAP7_75t_L g5435 ( 
.A(n_5425),
.B(n_5396),
.Y(n_5435)
);

NAND2xp5_ASAP7_75t_L g5436 ( 
.A(n_5425),
.B(n_5397),
.Y(n_5436)
);

AOI22xp5_ASAP7_75t_L g5437 ( 
.A1(n_5420),
.A2(n_5378),
.B1(n_5367),
.B2(n_5335),
.Y(n_5437)
);

CKINVDCx5p33_ASAP7_75t_R g5438 ( 
.A(n_5422),
.Y(n_5438)
);

OAI221xp5_ASAP7_75t_L g5439 ( 
.A1(n_5420),
.A2(n_5361),
.B1(n_5376),
.B2(n_5384),
.C(n_5372),
.Y(n_5439)
);

NAND2xp33_ASAP7_75t_SL g5440 ( 
.A(n_5426),
.B(n_5398),
.Y(n_5440)
);

CKINVDCx5p33_ASAP7_75t_R g5441 ( 
.A(n_5422),
.Y(n_5441)
);

NOR2x1_ASAP7_75t_L g5442 ( 
.A(n_5434),
.B(n_5405),
.Y(n_5442)
);

NAND2xp5_ASAP7_75t_L g5443 ( 
.A(n_5424),
.B(n_5398),
.Y(n_5443)
);

OAI22xp5_ASAP7_75t_L g5444 ( 
.A1(n_5430),
.A2(n_5395),
.B1(n_5408),
.B2(n_5361),
.Y(n_5444)
);

NOR2xp33_ASAP7_75t_L g5445 ( 
.A(n_5421),
.B(n_5402),
.Y(n_5445)
);

NAND2xp5_ASAP7_75t_L g5446 ( 
.A(n_5434),
.B(n_5405),
.Y(n_5446)
);

INVx2_ASAP7_75t_SL g5447 ( 
.A(n_5431),
.Y(n_5447)
);

AO221x2_ASAP7_75t_L g5448 ( 
.A1(n_5419),
.A2(n_5407),
.B1(n_5410),
.B2(n_5411),
.C(n_5413),
.Y(n_5448)
);

NAND2xp5_ASAP7_75t_L g5449 ( 
.A(n_5447),
.B(n_5428),
.Y(n_5449)
);

INVx1_ASAP7_75t_SL g5450 ( 
.A(n_5435),
.Y(n_5450)
);

INVx2_ASAP7_75t_L g5451 ( 
.A(n_5442),
.Y(n_5451)
);

NOR2x1_ASAP7_75t_L g5452 ( 
.A(n_5446),
.B(n_5416),
.Y(n_5452)
);

AND2x2_ASAP7_75t_L g5453 ( 
.A(n_5445),
.B(n_5428),
.Y(n_5453)
);

INVx2_ASAP7_75t_L g5454 ( 
.A(n_5438),
.Y(n_5454)
);

OAI21xp33_ASAP7_75t_L g5455 ( 
.A1(n_5437),
.A2(n_5412),
.B(n_5423),
.Y(n_5455)
);

INVx1_ASAP7_75t_L g5456 ( 
.A(n_5436),
.Y(n_5456)
);

OR2x2_ASAP7_75t_L g5457 ( 
.A(n_5443),
.B(n_5418),
.Y(n_5457)
);

INVx1_ASAP7_75t_L g5458 ( 
.A(n_5448),
.Y(n_5458)
);

INVx1_ASAP7_75t_L g5459 ( 
.A(n_5448),
.Y(n_5459)
);

AND2x2_ASAP7_75t_L g5460 ( 
.A(n_5441),
.B(n_5423),
.Y(n_5460)
);

INVx1_ASAP7_75t_L g5461 ( 
.A(n_5440),
.Y(n_5461)
);

NOR2xp33_ASAP7_75t_L g5462 ( 
.A(n_5439),
.B(n_5412),
.Y(n_5462)
);

AND2x4_ASAP7_75t_L g5463 ( 
.A(n_5444),
.B(n_5431),
.Y(n_5463)
);

NOR2x1_ASAP7_75t_L g5464 ( 
.A(n_5442),
.B(n_5417),
.Y(n_5464)
);

AND2x2_ASAP7_75t_L g5465 ( 
.A(n_5453),
.B(n_5415),
.Y(n_5465)
);

AND2x2_ASAP7_75t_L g5466 ( 
.A(n_5460),
.B(n_5415),
.Y(n_5466)
);

INVx1_ASAP7_75t_L g5467 ( 
.A(n_5449),
.Y(n_5467)
);

INVx1_ASAP7_75t_L g5468 ( 
.A(n_5464),
.Y(n_5468)
);

NAND2xp5_ASAP7_75t_L g5469 ( 
.A(n_5450),
.B(n_5433),
.Y(n_5469)
);

AND2x4_ASAP7_75t_L g5470 ( 
.A(n_5452),
.B(n_5433),
.Y(n_5470)
);

NAND2xp5_ASAP7_75t_L g5471 ( 
.A(n_5463),
.B(n_5451),
.Y(n_5471)
);

INVx1_ASAP7_75t_L g5472 ( 
.A(n_5457),
.Y(n_5472)
);

OR2x2_ASAP7_75t_L g5473 ( 
.A(n_5459),
.B(n_5374),
.Y(n_5473)
);

AND2x2_ASAP7_75t_L g5474 ( 
.A(n_5463),
.B(n_5430),
.Y(n_5474)
);

NAND2xp5_ASAP7_75t_L g5475 ( 
.A(n_5461),
.B(n_5376),
.Y(n_5475)
);

NAND2xp5_ASAP7_75t_L g5476 ( 
.A(n_5459),
.B(n_5356),
.Y(n_5476)
);

OAI21xp5_ASAP7_75t_SL g5477 ( 
.A1(n_5470),
.A2(n_5462),
.B(n_5455),
.Y(n_5477)
);

OAI22xp33_ASAP7_75t_L g5478 ( 
.A1(n_5469),
.A2(n_5400),
.B1(n_5392),
.B2(n_5432),
.Y(n_5478)
);

OAI221xp5_ASAP7_75t_L g5479 ( 
.A1(n_5475),
.A2(n_5384),
.B1(n_5400),
.B2(n_5427),
.C(n_5429),
.Y(n_5479)
);

OAI32xp33_ASAP7_75t_L g5480 ( 
.A1(n_5468),
.A2(n_5458),
.A3(n_5427),
.B1(n_5429),
.B2(n_5401),
.Y(n_5480)
);

NAND2xp5_ASAP7_75t_L g5481 ( 
.A(n_5470),
.B(n_5465),
.Y(n_5481)
);

NAND2xp5_ASAP7_75t_L g5482 ( 
.A(n_5466),
.B(n_5456),
.Y(n_5482)
);

INVx1_ASAP7_75t_L g5483 ( 
.A(n_5474),
.Y(n_5483)
);

OAI21xp5_ASAP7_75t_L g5484 ( 
.A1(n_5471),
.A2(n_5401),
.B(n_5399),
.Y(n_5484)
);

OR2x2_ASAP7_75t_L g5485 ( 
.A(n_5473),
.B(n_5369),
.Y(n_5485)
);

OAI31xp33_ASAP7_75t_L g5486 ( 
.A1(n_5472),
.A2(n_5399),
.A3(n_5352),
.B(n_5341),
.Y(n_5486)
);

AOI22xp33_ASAP7_75t_L g5487 ( 
.A1(n_5479),
.A2(n_5227),
.B1(n_5265),
.B2(n_5476),
.Y(n_5487)
);

OAI21xp5_ASAP7_75t_L g5488 ( 
.A1(n_5481),
.A2(n_5467),
.B(n_5454),
.Y(n_5488)
);

INVxp67_ASAP7_75t_L g5489 ( 
.A(n_5485),
.Y(n_5489)
);

AOI31xp33_ASAP7_75t_L g5490 ( 
.A1(n_5483),
.A2(n_5381),
.A3(n_5380),
.B(n_5339),
.Y(n_5490)
);

INVx1_ASAP7_75t_L g5491 ( 
.A(n_5482),
.Y(n_5491)
);

AND2x2_ASAP7_75t_L g5492 ( 
.A(n_5484),
.B(n_5477),
.Y(n_5492)
);

AOI211xp5_ASAP7_75t_SL g5493 ( 
.A1(n_5478),
.A2(n_5366),
.B(n_5327),
.C(n_5373),
.Y(n_5493)
);

INVx1_ASAP7_75t_L g5494 ( 
.A(n_5480),
.Y(n_5494)
);

NOR2xp33_ASAP7_75t_L g5495 ( 
.A(n_5486),
.B(n_5317),
.Y(n_5495)
);

INVx1_ASAP7_75t_L g5496 ( 
.A(n_5489),
.Y(n_5496)
);

INVx1_ASAP7_75t_L g5497 ( 
.A(n_5492),
.Y(n_5497)
);

NAND2xp5_ASAP7_75t_L g5498 ( 
.A(n_5493),
.B(n_5329),
.Y(n_5498)
);

INVx2_ASAP7_75t_L g5499 ( 
.A(n_5491),
.Y(n_5499)
);

OAI22x1_ASAP7_75t_L g5500 ( 
.A1(n_5494),
.A2(n_5297),
.B1(n_5291),
.B2(n_5286),
.Y(n_5500)
);

INVx1_ASAP7_75t_L g5501 ( 
.A(n_5488),
.Y(n_5501)
);

XNOR2x1_ASAP7_75t_L g5502 ( 
.A(n_5490),
.B(n_5309),
.Y(n_5502)
);

INVx1_ASAP7_75t_L g5503 ( 
.A(n_5495),
.Y(n_5503)
);

AND2x2_ASAP7_75t_L g5504 ( 
.A(n_5487),
.B(n_5292),
.Y(n_5504)
);

NOR2xp33_ASAP7_75t_L g5505 ( 
.A(n_5489),
.B(n_5321),
.Y(n_5505)
);

AND2x2_ASAP7_75t_L g5506 ( 
.A(n_5492),
.B(n_5264),
.Y(n_5506)
);

O2A1O1Ixp33_ASAP7_75t_L g5507 ( 
.A1(n_5489),
.A2(n_5346),
.B(n_5332),
.C(n_5348),
.Y(n_5507)
);

NAND2xp5_ASAP7_75t_L g5508 ( 
.A(n_5489),
.B(n_5318),
.Y(n_5508)
);

INVx1_ASAP7_75t_L g5509 ( 
.A(n_5489),
.Y(n_5509)
);

INVx1_ASAP7_75t_L g5510 ( 
.A(n_5489),
.Y(n_5510)
);

NAND2xp5_ASAP7_75t_L g5511 ( 
.A(n_5489),
.B(n_5318),
.Y(n_5511)
);

INVx2_ASAP7_75t_L g5512 ( 
.A(n_5492),
.Y(n_5512)
);

INVx1_ASAP7_75t_L g5513 ( 
.A(n_5489),
.Y(n_5513)
);

INVx2_ASAP7_75t_L g5514 ( 
.A(n_5512),
.Y(n_5514)
);

INVx1_ASAP7_75t_L g5515 ( 
.A(n_5498),
.Y(n_5515)
);

INVx1_ASAP7_75t_SL g5516 ( 
.A(n_5501),
.Y(n_5516)
);

AND2x2_ASAP7_75t_L g5517 ( 
.A(n_5506),
.B(n_5497),
.Y(n_5517)
);

INVx2_ASAP7_75t_L g5518 ( 
.A(n_5499),
.Y(n_5518)
);

INVx1_ASAP7_75t_L g5519 ( 
.A(n_5508),
.Y(n_5519)
);

INVx1_ASAP7_75t_L g5520 ( 
.A(n_5511),
.Y(n_5520)
);

INVxp33_ASAP7_75t_L g5521 ( 
.A(n_5505),
.Y(n_5521)
);

INVx1_ASAP7_75t_L g5522 ( 
.A(n_5496),
.Y(n_5522)
);

HB1xp67_ASAP7_75t_L g5523 ( 
.A(n_5500),
.Y(n_5523)
);

XNOR2x1_ASAP7_75t_L g5524 ( 
.A(n_5502),
.B(n_5286),
.Y(n_5524)
);

INVxp33_ASAP7_75t_SL g5525 ( 
.A(n_5496),
.Y(n_5525)
);

BUFx2_ASAP7_75t_L g5526 ( 
.A(n_5509),
.Y(n_5526)
);

INVx1_ASAP7_75t_L g5527 ( 
.A(n_5504),
.Y(n_5527)
);

INVx1_ASAP7_75t_L g5528 ( 
.A(n_5510),
.Y(n_5528)
);

INVx2_ASAP7_75t_SL g5529 ( 
.A(n_5513),
.Y(n_5529)
);

INVx1_ASAP7_75t_SL g5530 ( 
.A(n_5503),
.Y(n_5530)
);

INVx1_ASAP7_75t_L g5531 ( 
.A(n_5507),
.Y(n_5531)
);

INVx1_ASAP7_75t_L g5532 ( 
.A(n_5498),
.Y(n_5532)
);

INVx1_ASAP7_75t_L g5533 ( 
.A(n_5498),
.Y(n_5533)
);

INVx1_ASAP7_75t_L g5534 ( 
.A(n_5498),
.Y(n_5534)
);

INVx1_ASAP7_75t_L g5535 ( 
.A(n_5498),
.Y(n_5535)
);

INVx1_ASAP7_75t_L g5536 ( 
.A(n_5498),
.Y(n_5536)
);

INVxp33_ASAP7_75t_SL g5537 ( 
.A(n_5505),
.Y(n_5537)
);

INVx1_ASAP7_75t_L g5538 ( 
.A(n_5498),
.Y(n_5538)
);

INVx1_ASAP7_75t_L g5539 ( 
.A(n_5498),
.Y(n_5539)
);

NOR2x1_ASAP7_75t_L g5540 ( 
.A(n_5518),
.B(n_5337),
.Y(n_5540)
);

INVx1_ASAP7_75t_L g5541 ( 
.A(n_5517),
.Y(n_5541)
);

AOI211xp5_ASAP7_75t_L g5542 ( 
.A1(n_5516),
.A2(n_5272),
.B(n_5297),
.C(n_5291),
.Y(n_5542)
);

INVx1_ASAP7_75t_SL g5543 ( 
.A(n_5516),
.Y(n_5543)
);

NAND4xp25_ASAP7_75t_L g5544 ( 
.A(n_5526),
.B(n_5306),
.C(n_5289),
.D(n_5277),
.Y(n_5544)
);

NAND2x1p5_ASAP7_75t_L g5545 ( 
.A(n_5514),
.B(n_5287),
.Y(n_5545)
);

INVx1_ASAP7_75t_L g5546 ( 
.A(n_5523),
.Y(n_5546)
);

OAI221xp5_ASAP7_75t_L g5547 ( 
.A1(n_5523),
.A2(n_5287),
.B1(n_5306),
.B2(n_5289),
.C(n_5265),
.Y(n_5547)
);

AOI221xp5_ASAP7_75t_L g5548 ( 
.A1(n_5525),
.A2(n_5336),
.B1(n_5274),
.B2(n_5275),
.C(n_5255),
.Y(n_5548)
);

AOI21xp5_ASAP7_75t_L g5549 ( 
.A1(n_5529),
.A2(n_5264),
.B(n_5276),
.Y(n_5549)
);

INVxp67_ASAP7_75t_L g5550 ( 
.A(n_5524),
.Y(n_5550)
);

OAI22xp33_ASAP7_75t_SL g5551 ( 
.A1(n_5537),
.A2(n_5274),
.B1(n_5256),
.B2(n_5259),
.Y(n_5551)
);

A2O1A1Ixp33_ASAP7_75t_L g5552 ( 
.A1(n_5528),
.A2(n_5233),
.B(n_5255),
.C(n_5275),
.Y(n_5552)
);

INVx1_ASAP7_75t_L g5553 ( 
.A(n_5522),
.Y(n_5553)
);

NAND3xp33_ASAP7_75t_L g5554 ( 
.A(n_5515),
.B(n_5256),
.C(n_5259),
.Y(n_5554)
);

AOI22xp33_ASAP7_75t_SL g5555 ( 
.A1(n_5532),
.A2(n_5277),
.B1(n_5254),
.B2(n_5231),
.Y(n_5555)
);

NAND2xp33_ASAP7_75t_L g5556 ( 
.A(n_5527),
.B(n_5284),
.Y(n_5556)
);

OAI211xp5_ASAP7_75t_L g5557 ( 
.A1(n_5533),
.A2(n_5535),
.B(n_5536),
.C(n_5534),
.Y(n_5557)
);

NOR2xp67_ASAP7_75t_L g5558 ( 
.A(n_5538),
.B(n_5284),
.Y(n_5558)
);

AOI221xp5_ASAP7_75t_L g5559 ( 
.A1(n_5539),
.A2(n_5254),
.B1(n_5231),
.B2(n_5233),
.C(n_5234),
.Y(n_5559)
);

NAND2xp5_ASAP7_75t_L g5560 ( 
.A(n_5530),
.B(n_5294),
.Y(n_5560)
);

AOI21xp5_ASAP7_75t_L g5561 ( 
.A1(n_5530),
.A2(n_5235),
.B(n_5296),
.Y(n_5561)
);

AOI221xp5_ASAP7_75t_L g5562 ( 
.A1(n_5531),
.A2(n_5231),
.B1(n_5261),
.B2(n_5299),
.C(n_5269),
.Y(n_5562)
);

AOI22xp5_ASAP7_75t_L g5563 ( 
.A1(n_5519),
.A2(n_5299),
.B1(n_5269),
.B2(n_5283),
.Y(n_5563)
);

INVx2_ASAP7_75t_L g5564 ( 
.A(n_5520),
.Y(n_5564)
);

NAND2xp5_ASAP7_75t_L g5565 ( 
.A(n_5521),
.B(n_5283),
.Y(n_5565)
);

AOI211xp5_ASAP7_75t_L g5566 ( 
.A1(n_5516),
.A2(n_5299),
.B(n_455),
.C(n_453),
.Y(n_5566)
);

OR2x2_ASAP7_75t_L g5567 ( 
.A(n_5523),
.B(n_454),
.Y(n_5567)
);

A2O1A1Ixp33_ASAP7_75t_L g5568 ( 
.A1(n_5529),
.A2(n_454),
.B(n_455),
.C(n_456),
.Y(n_5568)
);

OAI211xp5_ASAP7_75t_L g5569 ( 
.A1(n_5543),
.A2(n_456),
.B(n_457),
.C(n_458),
.Y(n_5569)
);

OAI22xp5_ASAP7_75t_L g5570 ( 
.A1(n_5546),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_5570)
);

NAND3xp33_ASAP7_75t_L g5571 ( 
.A(n_5550),
.B(n_459),
.C(n_460),
.Y(n_5571)
);

AOI221xp5_ASAP7_75t_L g5572 ( 
.A1(n_5541),
.A2(n_460),
.B1(n_461),
.B2(n_462),
.C(n_464),
.Y(n_5572)
);

XOR2xp5_ASAP7_75t_L g5573 ( 
.A(n_5545),
.B(n_5544),
.Y(n_5573)
);

OAI222xp33_ASAP7_75t_L g5574 ( 
.A1(n_5555),
.A2(n_462),
.B1(n_465),
.B2(n_467),
.C1(n_470),
.C2(n_471),
.Y(n_5574)
);

OAI222xp33_ASAP7_75t_L g5575 ( 
.A1(n_5547),
.A2(n_5540),
.B1(n_5567),
.B2(n_5553),
.C1(n_5549),
.C2(n_5560),
.Y(n_5575)
);

OAI211xp5_ASAP7_75t_SL g5576 ( 
.A1(n_5557),
.A2(n_5564),
.B(n_5556),
.C(n_5542),
.Y(n_5576)
);

O2A1O1Ixp5_ASAP7_75t_L g5577 ( 
.A1(n_5565),
.A2(n_470),
.B(n_472),
.C(n_473),
.Y(n_5577)
);

OAI221xp5_ASAP7_75t_L g5578 ( 
.A1(n_5559),
.A2(n_473),
.B1(n_474),
.B2(n_475),
.C(n_476),
.Y(n_5578)
);

O2A1O1Ixp33_ASAP7_75t_L g5579 ( 
.A1(n_5568),
.A2(n_476),
.B(n_477),
.C(n_481),
.Y(n_5579)
);

AOI222xp33_ASAP7_75t_L g5580 ( 
.A1(n_5558),
.A2(n_481),
.B1(n_482),
.B2(n_483),
.C1(n_484),
.C2(n_487),
.Y(n_5580)
);

OAI22xp5_ASAP7_75t_L g5581 ( 
.A1(n_5552),
.A2(n_482),
.B1(n_483),
.B2(n_484),
.Y(n_5581)
);

AOI321xp33_ASAP7_75t_L g5582 ( 
.A1(n_5551),
.A2(n_487),
.A3(n_488),
.B1(n_489),
.B2(n_490),
.C(n_491),
.Y(n_5582)
);

OAI211xp5_ASAP7_75t_SL g5583 ( 
.A1(n_5562),
.A2(n_488),
.B(n_490),
.C(n_493),
.Y(n_5583)
);

AOI22xp5_ASAP7_75t_L g5584 ( 
.A1(n_5554),
.A2(n_493),
.B1(n_494),
.B2(n_495),
.Y(n_5584)
);

AND4x1_ASAP7_75t_L g5585 ( 
.A(n_5566),
.B(n_494),
.C(n_496),
.D(n_497),
.Y(n_5585)
);

OAI222xp33_ASAP7_75t_L g5586 ( 
.A1(n_5561),
.A2(n_496),
.B1(n_497),
.B2(n_498),
.C1(n_499),
.C2(n_500),
.Y(n_5586)
);

NAND2xp5_ASAP7_75t_L g5587 ( 
.A(n_5563),
.B(n_499),
.Y(n_5587)
);

NOR3x1_ASAP7_75t_L g5588 ( 
.A(n_5548),
.B(n_500),
.C(n_501),
.Y(n_5588)
);

OAI211xp5_ASAP7_75t_L g5589 ( 
.A1(n_5543),
.A2(n_503),
.B(n_504),
.C(n_505),
.Y(n_5589)
);

AOI22xp5_ASAP7_75t_L g5590 ( 
.A1(n_5546),
.A2(n_503),
.B1(n_505),
.B2(n_508),
.Y(n_5590)
);

NOR2xp33_ASAP7_75t_L g5591 ( 
.A(n_5543),
.B(n_508),
.Y(n_5591)
);

INVx1_ASAP7_75t_L g5592 ( 
.A(n_5545),
.Y(n_5592)
);

INVx1_ASAP7_75t_L g5593 ( 
.A(n_5545),
.Y(n_5593)
);

NAND2xp5_ASAP7_75t_SL g5594 ( 
.A(n_5582),
.B(n_509),
.Y(n_5594)
);

INVx1_ASAP7_75t_SL g5595 ( 
.A(n_5573),
.Y(n_5595)
);

AOI221xp5_ASAP7_75t_L g5596 ( 
.A1(n_5576),
.A2(n_509),
.B1(n_510),
.B2(n_513),
.C(n_514),
.Y(n_5596)
);

NAND4xp25_ASAP7_75t_L g5597 ( 
.A(n_5588),
.B(n_513),
.C(n_514),
.D(n_515),
.Y(n_5597)
);

OAI22xp5_ASAP7_75t_L g5598 ( 
.A1(n_5592),
.A2(n_516),
.B1(n_517),
.B2(n_518),
.Y(n_5598)
);

XNOR2xp5_ASAP7_75t_L g5599 ( 
.A(n_5585),
.B(n_516),
.Y(n_5599)
);

OAI21xp5_ASAP7_75t_SL g5600 ( 
.A1(n_5575),
.A2(n_517),
.B(n_519),
.Y(n_5600)
);

AOI221xp5_ASAP7_75t_L g5601 ( 
.A1(n_5574),
.A2(n_520),
.B1(n_521),
.B2(n_522),
.C(n_523),
.Y(n_5601)
);

AOI221xp5_ASAP7_75t_SL g5602 ( 
.A1(n_5593),
.A2(n_520),
.B1(n_521),
.B2(n_523),
.C(n_525),
.Y(n_5602)
);

NAND2xp5_ASAP7_75t_L g5603 ( 
.A(n_5580),
.B(n_526),
.Y(n_5603)
);

AOI221xp5_ASAP7_75t_L g5604 ( 
.A1(n_5583),
.A2(n_526),
.B1(n_527),
.B2(n_528),
.C(n_529),
.Y(n_5604)
);

HB1xp67_ASAP7_75t_L g5605 ( 
.A(n_5591),
.Y(n_5605)
);

A2O1A1Ixp33_ASAP7_75t_L g5606 ( 
.A1(n_5579),
.A2(n_528),
.B(n_529),
.C(n_530),
.Y(n_5606)
);

OAI22xp5_ASAP7_75t_L g5607 ( 
.A1(n_5584),
.A2(n_530),
.B1(n_532),
.B2(n_534),
.Y(n_5607)
);

XNOR2xp5_ASAP7_75t_L g5608 ( 
.A(n_5571),
.B(n_535),
.Y(n_5608)
);

OAI211xp5_ASAP7_75t_SL g5609 ( 
.A1(n_5578),
.A2(n_538),
.B(n_539),
.C(n_540),
.Y(n_5609)
);

OAI311xp33_ASAP7_75t_L g5610 ( 
.A1(n_5587),
.A2(n_538),
.A3(n_541),
.B1(n_542),
.C1(n_543),
.Y(n_5610)
);

AO22x2_ASAP7_75t_L g5611 ( 
.A1(n_5581),
.A2(n_541),
.B1(n_542),
.B2(n_544),
.Y(n_5611)
);

AOI22xp5_ASAP7_75t_L g5612 ( 
.A1(n_5595),
.A2(n_5589),
.B1(n_5569),
.B2(n_5590),
.Y(n_5612)
);

OAI22xp33_ASAP7_75t_L g5613 ( 
.A1(n_5603),
.A2(n_5570),
.B1(n_5572),
.B2(n_5586),
.Y(n_5613)
);

INVx1_ASAP7_75t_L g5614 ( 
.A(n_5599),
.Y(n_5614)
);

OR2x2_ASAP7_75t_L g5615 ( 
.A(n_5597),
.B(n_5577),
.Y(n_5615)
);

OR2x2_ASAP7_75t_L g5616 ( 
.A(n_5594),
.B(n_545),
.Y(n_5616)
);

INVx1_ASAP7_75t_L g5617 ( 
.A(n_5605),
.Y(n_5617)
);

OR2x6_ASAP7_75t_L g5618 ( 
.A(n_5600),
.B(n_546),
.Y(n_5618)
);

NOR2x1_ASAP7_75t_L g5619 ( 
.A(n_5598),
.B(n_5609),
.Y(n_5619)
);

OAI211xp5_ASAP7_75t_L g5620 ( 
.A1(n_5596),
.A2(n_546),
.B(n_547),
.C(n_548),
.Y(n_5620)
);

INVx1_ASAP7_75t_L g5621 ( 
.A(n_5611),
.Y(n_5621)
);

AND2x4_ASAP7_75t_L g5622 ( 
.A(n_5606),
.B(n_547),
.Y(n_5622)
);

AOI22xp5_ASAP7_75t_L g5623 ( 
.A1(n_5601),
.A2(n_548),
.B1(n_549),
.B2(n_550),
.Y(n_5623)
);

AOI22xp5_ASAP7_75t_L g5624 ( 
.A1(n_5607),
.A2(n_5604),
.B1(n_5602),
.B2(n_5608),
.Y(n_5624)
);

NAND2xp5_ASAP7_75t_SL g5625 ( 
.A(n_5610),
.B(n_550),
.Y(n_5625)
);

NAND2xp5_ASAP7_75t_L g5626 ( 
.A(n_5611),
.B(n_551),
.Y(n_5626)
);

OAI221xp5_ASAP7_75t_L g5627 ( 
.A1(n_5617),
.A2(n_551),
.B1(n_552),
.B2(n_553),
.C(n_554),
.Y(n_5627)
);

NOR2xp67_ASAP7_75t_L g5628 ( 
.A(n_5626),
.B(n_5620),
.Y(n_5628)
);

INVx2_ASAP7_75t_L g5629 ( 
.A(n_5621),
.Y(n_5629)
);

OAI211xp5_ASAP7_75t_L g5630 ( 
.A1(n_5612),
.A2(n_552),
.B(n_553),
.C(n_554),
.Y(n_5630)
);

NAND4xp25_ASAP7_75t_L g5631 ( 
.A(n_5625),
.B(n_555),
.C(n_556),
.D(n_558),
.Y(n_5631)
);

NAND3xp33_ASAP7_75t_SL g5632 ( 
.A(n_5614),
.B(n_555),
.C(n_558),
.Y(n_5632)
);

A2O1A1Ixp33_ASAP7_75t_L g5633 ( 
.A1(n_5615),
.A2(n_5624),
.B(n_5623),
.C(n_5616),
.Y(n_5633)
);

INVx1_ASAP7_75t_L g5634 ( 
.A(n_5618),
.Y(n_5634)
);

OR2x2_ASAP7_75t_L g5635 ( 
.A(n_5618),
.B(n_559),
.Y(n_5635)
);

NOR4xp75_ASAP7_75t_L g5636 ( 
.A(n_5619),
.B(n_559),
.C(n_560),
.D(n_562),
.Y(n_5636)
);

AOI21xp5_ASAP7_75t_L g5637 ( 
.A1(n_5613),
.A2(n_5622),
.B(n_562),
.Y(n_5637)
);

OAI22xp5_ASAP7_75t_L g5638 ( 
.A1(n_5617),
.A2(n_560),
.B1(n_564),
.B2(n_567),
.Y(n_5638)
);

OAI321xp33_ASAP7_75t_L g5639 ( 
.A1(n_5617),
.A2(n_567),
.A3(n_568),
.B1(n_569),
.B2(n_570),
.C(n_571),
.Y(n_5639)
);

NOR2x1_ASAP7_75t_L g5640 ( 
.A(n_5617),
.B(n_568),
.Y(n_5640)
);

NAND2xp33_ASAP7_75t_SL g5641 ( 
.A(n_5635),
.B(n_570),
.Y(n_5641)
);

NOR2xp33_ASAP7_75t_L g5642 ( 
.A(n_5629),
.B(n_571),
.Y(n_5642)
);

NAND2xp5_ASAP7_75t_L g5643 ( 
.A(n_5628),
.B(n_573),
.Y(n_5643)
);

NOR2xp33_ASAP7_75t_R g5644 ( 
.A(n_5632),
.B(n_574),
.Y(n_5644)
);

NAND2xp5_ASAP7_75t_SL g5645 ( 
.A(n_5639),
.B(n_575),
.Y(n_5645)
);

NAND2xp5_ASAP7_75t_L g5646 ( 
.A(n_5634),
.B(n_575),
.Y(n_5646)
);

NAND2xp5_ASAP7_75t_L g5647 ( 
.A(n_5640),
.B(n_576),
.Y(n_5647)
);

NOR2xp33_ASAP7_75t_R g5648 ( 
.A(n_5631),
.B(n_576),
.Y(n_5648)
);

NAND2xp5_ASAP7_75t_L g5649 ( 
.A(n_5633),
.B(n_577),
.Y(n_5649)
);

NAND2xp33_ASAP7_75t_SL g5650 ( 
.A(n_5638),
.B(n_578),
.Y(n_5650)
);

NAND2xp5_ASAP7_75t_L g5651 ( 
.A(n_5637),
.B(n_578),
.Y(n_5651)
);

INVx3_ASAP7_75t_L g5652 ( 
.A(n_5647),
.Y(n_5652)
);

INVxp67_ASAP7_75t_SL g5653 ( 
.A(n_5643),
.Y(n_5653)
);

OR4x2_ASAP7_75t_L g5654 ( 
.A(n_5648),
.B(n_5636),
.C(n_5630),
.D(n_5627),
.Y(n_5654)
);

AOI22x1_ASAP7_75t_L g5655 ( 
.A1(n_5649),
.A2(n_580),
.B1(n_581),
.B2(n_582),
.Y(n_5655)
);

INVx1_ASAP7_75t_L g5656 ( 
.A(n_5646),
.Y(n_5656)
);

INVx1_ASAP7_75t_L g5657 ( 
.A(n_5641),
.Y(n_5657)
);

NAND5xp2_ASAP7_75t_L g5658 ( 
.A(n_5651),
.B(n_581),
.C(n_582),
.D(n_583),
.E(n_584),
.Y(n_5658)
);

CKINVDCx12_ASAP7_75t_R g5659 ( 
.A(n_5653),
.Y(n_5659)
);

AND2x2_ASAP7_75t_L g5660 ( 
.A(n_5657),
.B(n_5642),
.Y(n_5660)
);

CKINVDCx20_ASAP7_75t_R g5661 ( 
.A(n_5656),
.Y(n_5661)
);

INVx1_ASAP7_75t_L g5662 ( 
.A(n_5659),
.Y(n_5662)
);

INVx2_ASAP7_75t_SL g5663 ( 
.A(n_5661),
.Y(n_5663)
);

INVx1_ASAP7_75t_L g5664 ( 
.A(n_5663),
.Y(n_5664)
);

INVxp67_ASAP7_75t_L g5665 ( 
.A(n_5662),
.Y(n_5665)
);

OAI22xp33_ASAP7_75t_SL g5666 ( 
.A1(n_5664),
.A2(n_5652),
.B1(n_5655),
.B2(n_5645),
.Y(n_5666)
);

OAI22xp5_ASAP7_75t_L g5667 ( 
.A1(n_5665),
.A2(n_5660),
.B1(n_5654),
.B2(n_5658),
.Y(n_5667)
);

XOR2xp5_ASAP7_75t_L g5668 ( 
.A(n_5664),
.B(n_5644),
.Y(n_5668)
);

AOI22xp33_ASAP7_75t_L g5669 ( 
.A1(n_5667),
.A2(n_5650),
.B1(n_586),
.B2(n_587),
.Y(n_5669)
);

AOI22xp33_ASAP7_75t_L g5670 ( 
.A1(n_5668),
.A2(n_584),
.B1(n_587),
.B2(n_589),
.Y(n_5670)
);

O2A1O1Ixp33_ASAP7_75t_R g5671 ( 
.A1(n_5666),
.A2(n_589),
.B(n_590),
.C(n_591),
.Y(n_5671)
);

AOI31xp33_ASAP7_75t_L g5672 ( 
.A1(n_5667),
.A2(n_592),
.A3(n_593),
.B(n_594),
.Y(n_5672)
);

INVx2_ASAP7_75t_L g5673 ( 
.A(n_5671),
.Y(n_5673)
);

BUFx2_ASAP7_75t_L g5674 ( 
.A(n_5672),
.Y(n_5674)
);

OAI21xp5_ASAP7_75t_L g5675 ( 
.A1(n_5669),
.A2(n_592),
.B(n_593),
.Y(n_5675)
);

INVx1_ASAP7_75t_L g5676 ( 
.A(n_5670),
.Y(n_5676)
);

HB1xp67_ASAP7_75t_L g5677 ( 
.A(n_5669),
.Y(n_5677)
);

AOI21x1_ASAP7_75t_L g5678 ( 
.A1(n_5673),
.A2(n_595),
.B(n_596),
.Y(n_5678)
);

AOI22xp5_ASAP7_75t_L g5679 ( 
.A1(n_5674),
.A2(n_595),
.B1(n_596),
.B2(n_597),
.Y(n_5679)
);

OR2x2_ASAP7_75t_L g5680 ( 
.A(n_5677),
.B(n_598),
.Y(n_5680)
);

AOI22xp5_ASAP7_75t_L g5681 ( 
.A1(n_5676),
.A2(n_5675),
.B1(n_599),
.B2(n_600),
.Y(n_5681)
);

AOI222xp33_ASAP7_75t_L g5682 ( 
.A1(n_5673),
.A2(n_598),
.B1(n_599),
.B2(n_601),
.C1(n_602),
.C2(n_603),
.Y(n_5682)
);

OAI21x1_ASAP7_75t_L g5683 ( 
.A1(n_5673),
.A2(n_601),
.B(n_605),
.Y(n_5683)
);

OAI22x1_ASAP7_75t_L g5684 ( 
.A1(n_5673),
.A2(n_605),
.B1(n_606),
.B2(n_607),
.Y(n_5684)
);

AOI22xp33_ASAP7_75t_L g5685 ( 
.A1(n_5673),
.A2(n_607),
.B1(n_608),
.B2(n_609),
.Y(n_5685)
);

AOI22xp33_ASAP7_75t_L g5686 ( 
.A1(n_5673),
.A2(n_608),
.B1(n_609),
.B2(n_610),
.Y(n_5686)
);

OR2x6_ASAP7_75t_L g5687 ( 
.A(n_5674),
.B(n_610),
.Y(n_5687)
);

INVx1_ASAP7_75t_L g5688 ( 
.A(n_5673),
.Y(n_5688)
);

OAI22x1_ASAP7_75t_L g5689 ( 
.A1(n_5688),
.A2(n_611),
.B1(n_612),
.B2(n_614),
.Y(n_5689)
);

AOI21xp5_ASAP7_75t_L g5690 ( 
.A1(n_5680),
.A2(n_611),
.B(n_612),
.Y(n_5690)
);

AOI22xp33_ASAP7_75t_L g5691 ( 
.A1(n_5687),
.A2(n_614),
.B1(n_615),
.B2(n_616),
.Y(n_5691)
);

AOI22xp5_ASAP7_75t_L g5692 ( 
.A1(n_5687),
.A2(n_617),
.B1(n_618),
.B2(n_620),
.Y(n_5692)
);

INVx1_ASAP7_75t_L g5693 ( 
.A(n_5681),
.Y(n_5693)
);

INVx1_ASAP7_75t_L g5694 ( 
.A(n_5678),
.Y(n_5694)
);

AOI222xp33_ASAP7_75t_L g5695 ( 
.A1(n_5684),
.A2(n_618),
.B1(n_620),
.B2(n_622),
.C1(n_623),
.C2(n_624),
.Y(n_5695)
);

AOI221x1_ASAP7_75t_L g5696 ( 
.A1(n_5683),
.A2(n_622),
.B1(n_623),
.B2(n_625),
.C(n_627),
.Y(n_5696)
);

INVxp67_ASAP7_75t_L g5697 ( 
.A(n_5682),
.Y(n_5697)
);

XNOR2xp5_ASAP7_75t_L g5698 ( 
.A(n_5694),
.B(n_5679),
.Y(n_5698)
);

INVx1_ASAP7_75t_L g5699 ( 
.A(n_5697),
.Y(n_5699)
);

INVx1_ASAP7_75t_L g5700 ( 
.A(n_5693),
.Y(n_5700)
);

OAI222xp33_ASAP7_75t_L g5701 ( 
.A1(n_5692),
.A2(n_5686),
.B1(n_5685),
.B2(n_631),
.C1(n_632),
.C2(n_633),
.Y(n_5701)
);

INVx1_ASAP7_75t_L g5702 ( 
.A(n_5690),
.Y(n_5702)
);

NAND2xp5_ASAP7_75t_L g5703 ( 
.A(n_5696),
.B(n_628),
.Y(n_5703)
);

INVxp67_ASAP7_75t_L g5704 ( 
.A(n_5700),
.Y(n_5704)
);

AO221x2_ASAP7_75t_L g5705 ( 
.A1(n_5699),
.A2(n_5689),
.B1(n_5695),
.B2(n_5691),
.C(n_634),
.Y(n_5705)
);

OAI321xp33_ASAP7_75t_L g5706 ( 
.A1(n_5702),
.A2(n_629),
.A3(n_631),
.B1(n_633),
.B2(n_634),
.C(n_635),
.Y(n_5706)
);

OAI221xp5_ASAP7_75t_R g5707 ( 
.A1(n_5704),
.A2(n_5698),
.B1(n_5701),
.B2(n_5703),
.C(n_640),
.Y(n_5707)
);

AOI221xp5_ASAP7_75t_L g5708 ( 
.A1(n_5707),
.A2(n_5706),
.B1(n_5705),
.B2(n_639),
.C(n_640),
.Y(n_5708)
);

AOI211xp5_ASAP7_75t_L g5709 ( 
.A1(n_5708),
.A2(n_635),
.B(n_637),
.C(n_639),
.Y(n_5709)
);


endmodule