module fake_jpeg_255_n_398 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_398);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_398;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx16_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_11),
.B(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_2),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx10_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

BUFx6f_ASAP7_75t_SL g39 ( 
.A(n_2),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_8),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_2),
.Y(n_43)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_SL g46 ( 
.A(n_3),
.Y(n_46)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_11),
.B(n_5),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_14),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_54),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_29),
.Y(n_55)
);

INVx5_ASAP7_75t_L g172 ( 
.A(n_55),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_56),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_15),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_57),
.B(n_58),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_26),
.B(n_15),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_25),
.Y(n_59)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_59),
.Y(n_165)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_60),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_61),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_20),
.B(n_14),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_62),
.B(n_68),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_12),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_63),
.B(n_81),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_65),
.Y(n_124)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_17),
.Y(n_66)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_66),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_67),
.B(n_94),
.Y(n_112)
);

AND2x2_ASAP7_75t_SL g68 ( 
.A(n_35),
.B(n_1),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_70),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_24),
.Y(n_71)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_71),
.Y(n_117)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_24),
.Y(n_73)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_73),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_24),
.Y(n_74)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_74),
.Y(n_136)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_36),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g146 ( 
.A(n_75),
.Y(n_146)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_49),
.Y(n_76)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_77),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_78),
.Y(n_138)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx3_ASAP7_75t_SL g80 ( 
.A(n_36),
.Y(n_80)
);

CKINVDCx6p67_ASAP7_75t_R g130 ( 
.A(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_18),
.B(n_1),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_82),
.Y(n_159)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_29),
.Y(n_84)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_22),
.Y(n_86)
);

INVxp67_ASAP7_75t_SL g156 ( 
.A(n_86),
.Y(n_156)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_28),
.Y(n_87)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_87),
.Y(n_135)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_38),
.Y(n_88)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_88),
.Y(n_161)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_38),
.Y(n_89)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_89),
.Y(n_147)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_27),
.Y(n_90)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_90),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_46),
.Y(n_92)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_92),
.Y(n_168)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

CKINVDCx16_ASAP7_75t_R g128 ( 
.A(n_93),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_17),
.B(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_29),
.Y(n_95)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_95),
.Y(n_154)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_96),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_18),
.B(n_2),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_97),
.B(n_98),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_37),
.Y(n_98)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_37),
.Y(n_99)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_99),
.Y(n_111)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_42),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_100),
.B(n_102),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_101),
.B(n_105),
.Y(n_120)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_103),
.B(n_106),
.Y(n_133)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_21),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_104),
.B(n_107),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_37),
.Y(n_105)
);

BUFx2_ASAP7_75t_L g106 ( 
.A(n_36),
.Y(n_106)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_39),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_108),
.B(n_109),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_110),
.B(n_23),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_32),
.B1(n_21),
.B2(n_43),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_116),
.A2(n_126),
.B1(n_129),
.B2(n_131),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_86),
.A2(n_39),
.B1(n_47),
.B2(n_32),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_39),
.B1(n_51),
.B2(n_50),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_94),
.A2(n_47),
.B1(n_51),
.B2(n_50),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_57),
.B(n_58),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g184 ( 
.A(n_142),
.B(n_160),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_56),
.A2(n_52),
.B1(n_41),
.B2(n_34),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_145),
.A2(n_108),
.B1(n_169),
.B2(n_158),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_106),
.A2(n_52),
.B1(n_41),
.B2(n_34),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_148),
.A2(n_158),
.B1(n_169),
.B2(n_173),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_149),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_62),
.B(n_23),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_150),
.B(n_152),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_68),
.B(n_45),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_19),
.B1(n_43),
.B2(n_40),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_155),
.A2(n_167),
.B1(n_128),
.B2(n_135),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_75),
.A2(n_19),
.B1(n_40),
.B2(n_33),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_45),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_55),
.B(n_33),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_177),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_73),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_61),
.A2(n_31),
.B1(n_30),
.B2(n_36),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_64),
.A2(n_36),
.B1(n_4),
.B2(n_5),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_69),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_174),
.A2(n_179),
.B1(n_98),
.B2(n_84),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_74),
.B(n_3),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_175),
.B(n_178),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_70),
.B(n_11),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_77),
.B(n_4),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_99),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_179)
);

OA22x2_ASAP7_75t_SL g180 ( 
.A1(n_80),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_180)
);

O2A1O1Ixp33_ASAP7_75t_SL g199 ( 
.A1(n_180),
.A2(n_145),
.B(n_167),
.C(n_173),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_131),
.A2(n_78),
.B(n_8),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_181),
.A2(n_200),
.B(n_220),
.Y(n_250)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_137),
.Y(n_182)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_182),
.Y(n_262)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_130),
.Y(n_185)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_185),
.Y(n_259)
);

BUFx8_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_186),
.Y(n_279)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_130),
.Y(n_188)
);

INVx3_ASAP7_75t_L g241 ( 
.A(n_188),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_189),
.A2(n_236),
.B(n_181),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_170),
.B(n_85),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_190),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_119),
.A2(n_95),
.B1(n_101),
.B2(n_105),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_191),
.A2(n_185),
.B1(n_188),
.B2(n_197),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_139),
.B(n_11),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_192),
.B(n_215),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_193),
.A2(n_220),
.B1(n_234),
.B2(n_181),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_112),
.B(n_113),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_194),
.B(n_210),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_139),
.B(n_151),
.Y(n_195)
);

OAI21xp33_ASAP7_75t_L g247 ( 
.A1(n_195),
.A2(n_199),
.B(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_130),
.Y(n_196)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_197),
.Y(n_258)
);

O2A1O1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_180),
.A2(n_156),
.B(n_120),
.C(n_148),
.Y(n_200)
);

INVx3_ASAP7_75t_L g201 ( 
.A(n_165),
.Y(n_201)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_201),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_180),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_202),
.B(n_205),
.Y(n_264)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_147),
.Y(n_203)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_203),
.Y(n_266)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_134),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_204),
.B(n_217),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_157),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g206 ( 
.A(n_125),
.B(n_133),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_206),
.B(n_207),
.Y(n_268)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_121),
.B(n_124),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_159),
.B(n_161),
.C(n_115),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_209),
.B(n_223),
.C(n_222),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_114),
.B(n_168),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_146),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_211),
.B(n_213),
.Y(n_275)
);

AOI32xp33_ASAP7_75t_L g213 ( 
.A1(n_143),
.A2(n_153),
.A3(n_154),
.B1(n_138),
.B2(n_162),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_156),
.B(n_132),
.Y(n_215)
);

OAI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_216),
.A2(n_231),
.B1(n_205),
.B2(n_196),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_172),
.Y(n_217)
);

NOR2x1_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_117),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_218),
.B(n_219),
.Y(n_265)
);

INVx3_ASAP7_75t_SL g219 ( 
.A(n_117),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_174),
.A2(n_127),
.B1(n_126),
.B2(n_179),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_221),
.B(n_222),
.Y(n_277)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_146),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g223 ( 
.A(n_138),
.B(n_122),
.Y(n_223)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_143),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_224),
.A2(n_229),
.B1(n_233),
.B2(n_237),
.Y(n_278)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_118),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_SL g254 ( 
.A(n_225),
.B(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_122),
.B(n_153),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_227),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_118),
.B(n_136),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_140),
.B(n_136),
.Y(n_228)
);

MAJx2_ASAP7_75t_L g272 ( 
.A(n_228),
.B(n_230),
.C(n_238),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_141),
.B(n_123),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_140),
.B(n_157),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g231 ( 
.A1(n_164),
.A2(n_171),
.B1(n_141),
.B2(n_176),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_164),
.Y(n_232)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_171),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_176),
.B(n_113),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_235),
.A2(n_223),
.B(n_186),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_112),
.A2(n_139),
.B1(n_63),
.B2(n_167),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_144),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_170),
.B(n_112),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_242),
.A2(n_250),
.B(n_269),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_202),
.A2(n_182),
.B1(n_236),
.B2(n_214),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_244),
.B1(n_248),
.B2(n_249),
.Y(n_290)
);

A2O1A1Ixp33_ASAP7_75t_L g246 ( 
.A1(n_192),
.A2(n_200),
.B(n_183),
.C(n_199),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_246),
.B(n_247),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_234),
.A2(n_204),
.B1(n_216),
.B2(n_199),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_189),
.A2(n_198),
.B1(n_184),
.B2(n_230),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_193),
.A2(n_228),
.B1(n_212),
.B2(n_187),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g252 ( 
.A1(n_212),
.A2(n_198),
.B1(n_221),
.B2(n_225),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_184),
.A2(n_232),
.B1(n_219),
.B2(n_203),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_206),
.A2(n_209),
.B1(n_235),
.B2(n_201),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_260),
.B(n_263),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_219),
.A2(n_218),
.B1(n_237),
.B2(n_207),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_261),
.A2(n_270),
.B1(n_273),
.B2(n_274),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g289 ( 
.A1(n_267),
.A2(n_271),
.B1(n_265),
.B2(n_275),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g291 ( 
.A(n_269),
.B(n_265),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_224),
.A2(n_223),
.B1(n_217),
.B2(n_186),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_186),
.A2(n_202),
.B1(n_182),
.B2(n_236),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_202),
.A2(n_182),
.B1(n_236),
.B2(n_214),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_202),
.A2(n_182),
.B1(n_236),
.B2(n_214),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_242),
.Y(n_286)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_281),
.A2(n_286),
.B(n_301),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_272),
.B(n_273),
.CI(n_274),
.CON(n_282),
.SN(n_282)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_287),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_271),
.A2(n_250),
.B1(n_248),
.B2(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_283),
.A2(n_289),
.B1(n_307),
.B2(n_259),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_253),
.B(n_251),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_284),
.B(n_285),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_262),
.B(n_240),
.Y(n_285)
);

NOR3xp33_ASAP7_75t_SL g287 ( 
.A(n_275),
.B(n_264),
.C(n_246),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_266),
.Y(n_288)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_288),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_291),
.A2(n_303),
.B(n_309),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_268),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_292),
.B(n_293),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_277),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_266),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_294),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_262),
.B(n_240),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_295),
.B(n_296),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_272),
.B(n_268),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_297),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_260),
.B(n_280),
.C(n_243),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_304),
.C(n_305),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_249),
.B(n_256),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_302),
.B(n_306),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_265),
.A2(n_254),
.B(n_278),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_239),
.B(n_263),
.C(n_252),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_255),
.B(n_239),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_257),
.B1(n_261),
.B2(n_276),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_276),
.B(n_241),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_308),
.B(n_311),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_254),
.A2(n_270),
.B(n_241),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_277),
.Y(n_310)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_310),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_279),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_315),
.A2(n_331),
.B1(n_307),
.B2(n_289),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_292),
.B(n_245),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_318),
.B(n_322),
.C(n_324),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_300),
.B(n_258),
.C(n_259),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_300),
.B(n_258),
.C(n_279),
.Y(n_324)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_328),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_296),
.B(n_279),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_329),
.B(n_333),
.C(n_303),
.Y(n_338)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_330),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_283),
.A2(n_298),
.B1(n_290),
.B2(n_302),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_284),
.C(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_317),
.B(n_295),
.Y(n_335)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_335),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_321),
.A2(n_301),
.B(n_286),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_337),
.B(n_343),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_338),
.B(n_347),
.Y(n_356)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_312),
.Y(n_340)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_340),
.Y(n_358)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_341),
.A2(n_331),
.B1(n_315),
.B2(n_325),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_316),
.B(n_305),
.C(n_285),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_342),
.B(n_318),
.C(n_322),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_SL g343 ( 
.A(n_314),
.B(n_287),
.C(n_306),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g344 ( 
.A1(n_321),
.A2(n_291),
.B(n_309),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_344),
.B(n_349),
.Y(n_354)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_312),
.Y(n_345)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_345),
.Y(n_362)
);

NOR3xp33_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_287),
.C(n_282),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_346),
.B(n_350),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_316),
.B(n_305),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_319),
.A2(n_290),
.B(n_298),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_348),
.B(n_319),
.Y(n_357)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g350 ( 
.A(n_332),
.B(n_293),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_351),
.B(n_341),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_359),
.C(n_360),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_357),
.A2(n_337),
.B(n_348),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_324),
.C(n_333),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_334),
.B(n_329),
.C(n_320),
.Y(n_360)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_334),
.B(n_320),
.C(n_327),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_363),
.B(n_356),
.Y(n_366)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_358),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_366),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_367),
.A2(n_372),
.B1(n_373),
.B2(n_351),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g368 ( 
.A(n_353),
.B(n_323),
.Y(n_368)
);

AOI322xp5_ASAP7_75t_L g380 ( 
.A1(n_368),
.A2(n_323),
.A3(n_335),
.B1(n_327),
.B2(n_317),
.C1(n_326),
.C2(n_308),
.Y(n_380)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_362),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g374 ( 
.A1(n_369),
.A2(n_370),
.B1(n_371),
.B2(n_350),
.Y(n_374)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_352),
.Y(n_370)
);

AOI31xp67_ASAP7_75t_L g371 ( 
.A1(n_361),
.A2(n_344),
.A3(n_343),
.B(n_346),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_SL g372 ( 
.A(n_356),
.B(n_363),
.Y(n_372)
);

OR2x2_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_379),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_377),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_367),
.A2(n_373),
.B1(n_325),
.B2(n_354),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_371),
.A2(n_354),
.B1(n_357),
.B2(n_299),
.Y(n_378)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_378),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_366),
.A2(n_326),
.B(n_332),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_380),
.B(n_336),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_375),
.B(n_365),
.C(n_372),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_355),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_376),
.A2(n_374),
.B(n_378),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_377),
.B(n_379),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_385),
.B(n_376),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_387),
.B(n_388),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_382),
.B(n_365),
.C(n_359),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_389),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_390),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_392),
.A2(n_386),
.B(n_381),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_394),
.A2(n_395),
.B(n_391),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_393),
.B(n_389),
.C(n_386),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g397 ( 
.A1(n_396),
.A2(n_384),
.B1(n_349),
.B2(n_345),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_397),
.B(n_339),
.Y(n_398)
);


endmodule