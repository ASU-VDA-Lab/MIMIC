module fake_jpeg_13096_n_62 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_18),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_25),
.A2(n_26),
.B(n_1),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_0),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_12),
.B1(n_20),
.B2(n_19),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_31),
.A2(n_33),
.B1(n_28),
.B2(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_32),
.Y(n_36)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_22),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_24),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_35),
.B(n_37),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_34),
.B(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_R g50 ( 
.A(n_39),
.B(n_3),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g41 ( 
.A(n_34),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_42),
.A2(n_28),
.B1(n_23),
.B2(n_4),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_43),
.A2(n_45),
.B1(n_21),
.B2(n_9),
.Y(n_51)
);

BUFx24_ASAP7_75t_SL g44 ( 
.A(n_39),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_46),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_36),
.B1(n_23),
.B2(n_40),
.Y(n_45)
);

OAI32xp33_ASAP7_75t_L g46 ( 
.A1(n_36),
.A2(n_2),
.A3(n_3),
.B1(n_4),
.B2(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_47),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_50),
.B(n_14),
.Y(n_54)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_49),
.A2(n_7),
.B1(n_10),
.B2(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_54),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_56),
.B(n_55),
.Y(n_58)
);

OAI221xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_53),
.B1(n_57),
.B2(n_52),
.C(n_51),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_59),
.B(n_48),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_60),
.B(n_48),
.C(n_16),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_15),
.Y(n_62)
);


endmodule