module fake_jpeg_23284_n_205 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_205);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_205;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_11),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx24_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx16f_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_5),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_15),
.B(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_29),
.B(n_34),
.Y(n_54)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_30),
.Y(n_53)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_32),
.Y(n_39)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_19),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_23),
.Y(n_55)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g40 ( 
.A1(n_34),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_44),
.B1(n_45),
.B2(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_29),
.B(n_21),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_41),
.B(n_14),
.Y(n_61)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_37),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_37),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_37),
.A2(n_19),
.B1(n_26),
.B2(n_21),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_34),
.A2(n_26),
.B(n_16),
.C(n_15),
.Y(n_46)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_46),
.A2(n_35),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_36),
.A2(n_26),
.B1(n_20),
.B2(n_16),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_31),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_31),
.B(n_27),
.Y(n_52)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_55),
.B(n_35),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_53),
.A2(n_31),
.B1(n_30),
.B2(n_27),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_67),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_61),
.B(n_70),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_23),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_49),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_46),
.B(n_32),
.Y(n_65)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_62),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_53),
.A2(n_30),
.B1(n_14),
.B2(n_22),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_38),
.B1(n_36),
.B2(n_30),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_53),
.A2(n_22),
.B1(n_36),
.B2(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_71),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_33),
.B(n_16),
.C(n_38),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_72),
.B(n_73),
.Y(n_78)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_74),
.B(n_76),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_75),
.A2(n_39),
.B(n_68),
.Y(n_105)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_60),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_81),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_79),
.B(n_88),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_65),
.B(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_54),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_70),
.Y(n_83)
);

NOR3xp33_ASAP7_75t_SL g106 ( 
.A(n_83),
.B(n_66),
.C(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_70),
.Y(n_85)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

AO22x2_ASAP7_75t_L g87 ( 
.A1(n_64),
.A2(n_40),
.B1(n_45),
.B2(n_33),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_87),
.A2(n_71),
.B1(n_63),
.B2(n_67),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_55),
.C(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_61),
.B(n_28),
.Y(n_91)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_91),
.Y(n_109)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_78),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_92),
.B(n_102),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g94 ( 
.A1(n_80),
.A2(n_65),
.B(n_72),
.Y(n_94)
);

A2O1A1O1Ixp25_ASAP7_75t_L g119 ( 
.A1(n_94),
.A2(n_87),
.B(n_105),
.C(n_93),
.D(n_101),
.Y(n_119)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_96),
.A2(n_106),
.B1(n_32),
.B2(n_35),
.Y(n_122)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_74),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_58),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_79),
.Y(n_112)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_86),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_69),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_89),
.A2(n_58),
.B1(n_63),
.B2(n_68),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_104),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_105),
.A2(n_87),
.B(n_88),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_77),
.Y(n_108)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_108),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_103),
.A2(n_87),
.B1(n_85),
.B2(n_81),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_110),
.A2(n_50),
.B1(n_56),
.B2(n_33),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_116),
.B(n_121),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_112),
.B(n_119),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_92),
.B(n_84),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_113),
.B(n_115),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_109),
.B(n_84),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_75),
.C(n_87),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_127),
.C(n_99),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_76),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_120),
.B(n_126),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_96),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_125),
.B1(n_48),
.B2(n_104),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_95),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_94),
.B(n_47),
.C(n_39),
.Y(n_127)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_124),
.Y(n_128)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_129),
.A2(n_135),
.B1(n_136),
.B2(n_144),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_133),
.C(n_139),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_117),
.B(n_97),
.C(n_98),
.Y(n_133)
);

XNOR2x1_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_97),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_134),
.B(n_140),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_125),
.A2(n_100),
.B1(n_106),
.B2(n_91),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_123),
.A2(n_43),
.B1(n_51),
.B2(n_18),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_43),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_114),
.C(n_126),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_50),
.C(n_51),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_123),
.A2(n_28),
.B(n_25),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_127),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_139),
.B(n_115),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_145),
.B(n_153),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_142),
.B(n_112),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_121),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_141),
.B(n_118),
.Y(n_148)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_148),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_110),
.Y(n_149)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_149),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_137),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_132),
.B(n_113),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_154),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_130),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_157),
.A2(n_158),
.B1(n_25),
.B2(n_18),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g158 ( 
.A(n_144),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_159),
.B(n_166),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_133),
.C(n_131),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_161),
.B(n_165),
.C(n_167),
.Y(n_172)
);

XNOR2x1_ASAP7_75t_SL g162 ( 
.A(n_146),
.B(n_134),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_162),
.A2(n_147),
.B1(n_23),
.B2(n_2),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_150),
.B(n_130),
.C(n_140),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_146),
.B(n_121),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_155),
.B(n_143),
.C(n_56),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_169),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_163),
.A2(n_152),
.B1(n_158),
.B2(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_171),
.B(n_176),
.Y(n_181)
);

XOR2x1_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_166),
.Y(n_173)
);

OAI21x1_ASAP7_75t_L g182 ( 
.A1(n_173),
.A2(n_170),
.B(n_1),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_168),
.A2(n_152),
.B1(n_160),
.B2(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_175),
.B(n_7),
.Y(n_185)
);

AND2x2_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_156),
.Y(n_176)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_9),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_164),
.B(n_151),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

AOI21x1_ASAP7_75t_L g190 ( 
.A1(n_182),
.A2(n_12),
.B(n_3),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_174),
.B(n_0),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_183),
.A2(n_184),
.B(n_185),
.Y(n_191)
);

NAND4xp25_ASAP7_75t_L g184 ( 
.A(n_173),
.B(n_56),
.C(n_1),
.D(n_2),
.Y(n_184)
);

OAI221xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_7),
.B1(n_3),
.B2(n_4),
.C(n_5),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_12),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_9),
.C(n_3),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_189),
.A2(n_193),
.B(n_6),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_190),
.A2(n_183),
.B(n_4),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_181),
.A2(n_176),
.B1(n_172),
.B2(n_177),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_192),
.B(n_194),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_188),
.A2(n_172),
.B(n_177),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_195),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_189),
.A2(n_56),
.B(n_6),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_196),
.B(n_197),
.C(n_10),
.Y(n_201)
);

AOI321xp33_ASAP7_75t_L g199 ( 
.A1(n_198),
.A2(n_191),
.A3(n_9),
.B1(n_10),
.B2(n_13),
.C(n_0),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_199),
.B(n_201),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_200),
.B(n_10),
.C(n_13),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_203),
.B(n_13),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_204),
.B(n_202),
.Y(n_205)
);


endmodule