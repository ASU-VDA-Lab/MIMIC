module fake_jpeg_128_n_697 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_697);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_697;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_417;
wire n_362;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx11_ASAP7_75t_SL g22 ( 
.A(n_19),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_10),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_2),
.Y(n_37)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_4),
.Y(n_38)
);

BUFx8_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

BUFx5_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_1),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_3),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_11),
.Y(n_53)
);

HB1xp67_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_3),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_11),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_19),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_63),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_20),
.B(n_19),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_64),
.B(n_78),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_65),
.Y(n_150)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx4_ASAP7_75t_SL g170 ( 
.A(n_66),
.Y(n_170)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_52),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g187 ( 
.A(n_67),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_68),
.Y(n_207)
);

INVx13_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVxp67_ASAP7_75t_SL g142 ( 
.A(n_69),
.Y(n_142)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_71),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g200 ( 
.A(n_72),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

INVx6_ASAP7_75t_L g165 ( 
.A(n_73),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_75),
.Y(n_178)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx5_ASAP7_75t_L g147 ( 
.A(n_76),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_77),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_20),
.B(n_18),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_36),
.Y(n_79)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_79),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_36),
.Y(n_80)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_80),
.Y(n_223)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_81),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_18),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_82),
.B(n_54),
.Y(n_136)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_83),
.Y(n_162)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_37),
.Y(n_85)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_85),
.Y(n_168)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_58),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_86),
.Y(n_212)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_40),
.Y(n_87)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_87),
.Y(n_152)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_22),
.Y(n_88)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_89),
.Y(n_153)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_90),
.Y(n_157)
);

BUFx24_ASAP7_75t_L g91 ( 
.A(n_39),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_36),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_92),
.Y(n_155)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_58),
.Y(n_93)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_93),
.Y(n_174)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_94),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_36),
.Y(n_95)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_95),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_23),
.B(n_17),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_96),
.B(n_24),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_97),
.Y(n_184)
);

INVx4_ASAP7_75t_SL g98 ( 
.A(n_39),
.Y(n_98)
);

BUFx3_ASAP7_75t_L g222 ( 
.A(n_98),
.Y(n_222)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_26),
.Y(n_99)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_99),
.Y(n_149)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_38),
.Y(n_100)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_37),
.Y(n_101)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_26),
.Y(n_102)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_102),
.Y(n_166)
);

INVx5_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_104),
.Y(n_159)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_28),
.Y(n_105)
);

INVx5_ASAP7_75t_L g191 ( 
.A(n_105),
.Y(n_191)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_43),
.Y(n_106)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_106),
.Y(n_210)
);

INVx8_ASAP7_75t_L g107 ( 
.A(n_41),
.Y(n_107)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_107),
.Y(n_214)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_38),
.Y(n_108)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_108),
.Y(n_203)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_109),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_39),
.Y(n_110)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_110),
.Y(n_219)
);

INVx2_ASAP7_75t_SL g111 ( 
.A(n_39),
.Y(n_111)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_43),
.Y(n_112)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

BUFx12f_ASAP7_75t_SL g226 ( 
.A(n_113),
.Y(n_226)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_50),
.Y(n_114)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_114),
.Y(n_164)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_38),
.Y(n_115)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_43),
.Y(n_116)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_116),
.Y(n_201)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_117),
.Y(n_202)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_37),
.Y(n_118)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_118),
.Y(n_211)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_53),
.Y(n_119)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_121),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_53),
.Y(n_122)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_34),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_126),
.Y(n_145)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_41),
.Y(n_124)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_124),
.Y(n_217)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_31),
.Y(n_125)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_125),
.Y(n_221)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_41),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_31),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_132),
.Y(n_144)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_55),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_128),
.B(n_129),
.Y(n_224)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_130),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_56),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_131),
.Y(n_171)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_55),
.Y(n_132)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_45),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g176 ( 
.A(n_133),
.B(n_44),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_136),
.B(n_148),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_68),
.B(n_60),
.C(n_61),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_137),
.B(n_140),
.C(n_190),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_86),
.B(n_60),
.C(n_61),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_64),
.A2(n_96),
.B1(n_78),
.B2(n_130),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_141),
.A2(n_172),
.B1(n_185),
.B2(n_208),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_98),
.B(n_27),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_106),
.A2(n_56),
.B1(n_57),
.B2(n_48),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_151),
.A2(n_161),
.B1(n_169),
.B2(n_215),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_111),
.B(n_27),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_154),
.B(n_182),
.Y(n_250)
);

HAxp5_ASAP7_75t_SL g156 ( 
.A(n_69),
.B(n_50),
.CON(n_156),
.SN(n_156)
);

OR2x2_ASAP7_75t_L g244 ( 
.A(n_156),
.B(n_220),
.Y(n_244)
);

OAI22xp33_ASAP7_75t_L g161 ( 
.A1(n_119),
.A2(n_57),
.B1(n_48),
.B2(n_47),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_62),
.A2(n_72),
.B1(n_131),
.B2(n_122),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_65),
.A2(n_56),
.B1(n_57),
.B2(n_48),
.Y(n_172)
);

CKINVDCx14_ASAP7_75t_R g306 ( 
.A(n_176),
.Y(n_306)
);

INVx6_ASAP7_75t_SL g177 ( 
.A(n_91),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_177),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_71),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_197),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_110),
.B(n_23),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_73),
.A2(n_56),
.B1(n_57),
.B2(n_48),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_44),
.C(n_49),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_110),
.B(n_24),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_196),
.B(n_204),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_132),
.B(n_30),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_74),
.B(n_30),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_205),
.B(n_209),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_75),
.A2(n_47),
.B1(n_35),
.B2(n_42),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_77),
.B(n_51),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_76),
.A2(n_29),
.B1(n_34),
.B2(n_55),
.Y(n_213)
);

AOI21xp5_ASAP7_75t_L g298 ( 
.A1(n_213),
.A2(n_0),
.B(n_2),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_79),
.A2(n_35),
.B1(n_42),
.B2(n_47),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_51),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_218),
.B(n_225),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_80),
.B(n_46),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_107),
.B(n_49),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_193),
.A2(n_46),
.B(n_55),
.C(n_45),
.Y(n_227)
);

AOI21xp33_ASAP7_75t_L g358 ( 
.A1(n_227),
.A2(n_281),
.B(n_297),
.Y(n_358)
);

BUFx12f_ASAP7_75t_L g228 ( 
.A(n_219),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g317 ( 
.A(n_228),
.Y(n_317)
);

AND2x4_ASAP7_75t_SL g229 ( 
.A(n_138),
.B(n_35),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g367 ( 
.A(n_229),
.B(n_4),
.Y(n_367)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_134),
.Y(n_230)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_230),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_156),
.A2(n_29),
.B1(n_34),
.B2(n_47),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_231),
.A2(n_240),
.B1(n_246),
.B2(n_251),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_35),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_SL g309 ( 
.A(n_232),
.B(n_283),
.Y(n_309)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_234),
.Y(n_323)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_146),
.Y(n_237)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_237),
.Y(n_319)
);

INVx6_ASAP7_75t_L g238 ( 
.A(n_143),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_238),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_208),
.A2(n_120),
.B1(n_116),
.B2(n_112),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_239),
.A2(n_272),
.B1(n_287),
.B2(n_187),
.Y(n_328)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_145),
.A2(n_29),
.B1(n_42),
.B2(n_92),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_149),
.Y(n_241)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_241),
.Y(n_332)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_166),
.Y(n_242)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_242),
.Y(n_335)
);

INVx6_ASAP7_75t_L g243 ( 
.A(n_143),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

INVx4_ASAP7_75t_L g245 ( 
.A(n_158),
.Y(n_245)
);

INVx4_ASAP7_75t_L g308 ( 
.A(n_245),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_145),
.A2(n_142),
.B1(n_158),
.B2(n_206),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx2_ASAP7_75t_L g340 ( 
.A(n_247),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_150),
.Y(n_248)
);

INVx5_ASAP7_75t_L g343 ( 
.A(n_248),
.Y(n_343)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_174),
.Y(n_249)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_249),
.Y(n_348)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_142),
.A2(n_42),
.B1(n_95),
.B2(n_97),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_144),
.Y(n_252)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_252),
.Y(n_330)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_167),
.Y(n_254)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_254),
.Y(n_365)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_222),
.Y(n_255)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_222),
.Y(n_256)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_256),
.Y(n_314)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_174),
.Y(n_257)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_257),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_164),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_258),
.B(n_271),
.Y(n_315)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_158),
.Y(n_259)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_259),
.Y(n_345)
);

INVx5_ASAP7_75t_L g262 ( 
.A(n_219),
.Y(n_262)
);

INVx3_ASAP7_75t_L g316 ( 
.A(n_262),
.Y(n_316)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_216),
.Y(n_263)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

AO22x2_ASAP7_75t_L g264 ( 
.A1(n_161),
.A2(n_45),
.B1(n_2),
.B2(n_3),
.Y(n_264)
);

AO22x1_ASAP7_75t_SL g363 ( 
.A1(n_264),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_169),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_265),
.A2(n_178),
.B1(n_173),
.B2(n_180),
.Y(n_321)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_189),
.Y(n_266)
);

INVx3_ASAP7_75t_L g352 ( 
.A(n_266),
.Y(n_352)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_207),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_267),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_226),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_SL g324 ( 
.A1(n_270),
.A2(n_286),
.B1(n_298),
.B2(n_300),
.Y(n_324)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_160),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_213),
.A2(n_16),
.B1(n_14),
.B2(n_13),
.Y(n_272)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_147),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_273),
.B(n_274),
.Y(n_342)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_201),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_188),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_275),
.B(n_277),
.Y(n_351)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_198),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_188),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_278),
.B(n_279),
.Y(n_356)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_217),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_150),
.Y(n_280)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

A2O1A1Ixp33_ASAP7_75t_L g281 ( 
.A1(n_159),
.A2(n_16),
.B(n_14),
.C(n_13),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_282),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_153),
.B(n_13),
.Y(n_283)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_157),
.B(n_152),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_284),
.B(n_299),
.C(n_175),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g285 ( 
.A(n_195),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_285),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_200),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_139),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_207),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_288),
.B(n_290),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g289 ( 
.A1(n_226),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_289),
.A2(n_224),
.B(n_194),
.Y(n_336)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_192),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_147),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_292),
.Y(n_360)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_203),
.Y(n_292)
);

BUFx2_ASAP7_75t_L g293 ( 
.A(n_191),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_293),
.B(n_294),
.Y(n_364)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_212),
.Y(n_294)
);

INVx4_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_295),
.B(n_296),
.Y(n_337)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_200),
.Y(n_296)
);

AND2x2_ASAP7_75t_L g297 ( 
.A(n_224),
.B(n_10),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_202),
.B(n_203),
.C(n_211),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_199),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_165),
.Y(n_301)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_301),
.A2(n_302),
.B1(n_303),
.B2(n_305),
.Y(n_333)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_170),
.Y(n_302)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_212),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_155),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_304),
.B(n_187),
.Y(n_307)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_170),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_307),
.Y(n_385)
);

AOI22xp33_ASAP7_75t_L g310 ( 
.A1(n_235),
.A2(n_171),
.B1(n_163),
.B2(n_155),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g401 ( 
.A1(n_310),
.A2(n_328),
.B1(n_341),
.B2(n_5),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_236),
.A2(n_244),
.B1(n_269),
.B2(n_306),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_313),
.A2(n_320),
.B1(n_321),
.B2(n_329),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_260),
.B(n_210),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_318),
.B(n_322),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_244),
.A2(n_165),
.B1(n_180),
.B2(n_178),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_233),
.B(n_210),
.Y(n_322)
);

OAI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_227),
.A2(n_206),
.B1(n_194),
.B2(n_168),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_276),
.B(n_191),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_331),
.B(n_344),
.Y(n_376)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_336),
.Y(n_415)
);

AOI22xp33_ASAP7_75t_SL g338 ( 
.A1(n_270),
.A2(n_186),
.B1(n_168),
.B2(n_214),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_338),
.A2(n_366),
.B1(n_259),
.B2(n_355),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g341 ( 
.A1(n_264),
.A2(n_184),
.B1(n_181),
.B2(n_186),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_232),
.B(n_181),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g386 ( 
.A(n_347),
.B(n_363),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_231),
.A2(n_175),
.B1(n_162),
.B2(n_223),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_349),
.A2(n_350),
.B1(n_355),
.B2(n_366),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_264),
.A2(n_173),
.B1(n_184),
.B2(n_135),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_253),
.B(n_0),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_353),
.B(n_367),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g355 ( 
.A1(n_240),
.A2(n_223),
.B1(n_135),
.B2(n_162),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_250),
.B(n_10),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_357),
.B(n_261),
.C(n_297),
.Y(n_370)
);

O2A1O1Ixp33_ASAP7_75t_SL g361 ( 
.A1(n_264),
.A2(n_4),
.B(n_5),
.C(n_6),
.Y(n_361)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_281),
.B(n_289),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_251),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_367),
.B(n_363),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_369),
.B(n_400),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_370),
.B(n_354),
.Y(n_425)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_311),
.Y(n_371)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_371),
.Y(n_428)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_374),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_328),
.A2(n_268),
.B1(n_229),
.B2(n_296),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_375),
.A2(n_378),
.B1(n_390),
.B2(n_395),
.Y(n_419)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_319),
.Y(n_377)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_377),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_322),
.A2(n_229),
.B1(n_284),
.B2(n_301),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g379 ( 
.A1(n_321),
.A2(n_291),
.B1(n_273),
.B2(n_282),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g444 ( 
.A1(n_379),
.A2(n_404),
.B1(n_339),
.B2(n_316),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_330),
.B(n_258),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_380),
.B(n_387),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_381),
.B(n_392),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g382 ( 
.A(n_318),
.B(n_246),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_354),
.Y(n_435)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_383),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_SL g384 ( 
.A1(n_350),
.A2(n_320),
.B1(n_312),
.B2(n_313),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g429 ( 
.A1(n_384),
.A2(n_416),
.B(n_343),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_309),
.B(n_295),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_347),
.B(n_255),
.C(n_293),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_388),
.B(n_406),
.C(n_409),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_330),
.B(n_262),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_SL g451 ( 
.A(n_389),
.B(n_396),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_336),
.A2(n_243),
.B1(n_238),
.B2(n_285),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_351),
.Y(n_392)
);

AOI32xp33_ASAP7_75t_L g393 ( 
.A1(n_358),
.A2(n_245),
.A3(n_294),
.B1(n_267),
.B2(n_303),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_393),
.B(n_407),
.Y(n_443)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_319),
.Y(n_394)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_394),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_324),
.A2(n_286),
.B1(n_280),
.B2(n_248),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_309),
.B(n_256),
.Y(n_396)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_344),
.A2(n_288),
.B1(n_228),
.B2(n_7),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g421 ( 
.A1(n_397),
.A2(n_401),
.B1(n_405),
.B2(n_317),
.Y(n_421)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_365),
.Y(n_398)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_398),
.Y(n_440)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_365),
.Y(n_399)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_399),
.Y(n_455)
);

AO22x1_ASAP7_75t_SL g400 ( 
.A1(n_361),
.A2(n_228),
.B1(n_6),
.B2(n_7),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_353),
.B(n_9),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_402),
.B(n_403),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_331),
.B(n_9),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_363),
.A2(n_8),
.B1(n_367),
.B2(n_357),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_359),
.B(n_8),
.C(n_307),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_337),
.Y(n_407)
);

CKINVDCx14_ASAP7_75t_R g439 ( 
.A(n_408),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_342),
.B(n_360),
.C(n_315),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_410),
.B(n_385),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_332),
.B(n_335),
.C(n_340),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_411),
.B(n_314),
.C(n_382),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_327),
.B(n_364),
.Y(n_412)
);

CKINVDCx14_ASAP7_75t_R g450 ( 
.A(n_412),
.Y(n_450)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_334),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_413),
.B(n_417),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_325),
.B(n_352),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_414),
.B(n_348),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_SL g416 ( 
.A1(n_327),
.A2(n_368),
.B1(n_362),
.B2(n_326),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_334),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_415),
.A2(n_333),
.B(n_317),
.Y(n_418)
);

AOI21xp5_ASAP7_75t_L g488 ( 
.A1(n_418),
.A2(n_432),
.B(n_383),
.Y(n_488)
);

AOI22xp33_ASAP7_75t_L g420 ( 
.A1(n_375),
.A2(n_368),
.B1(n_362),
.B2(n_334),
.Y(n_420)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_420),
.A2(n_417),
.B1(n_413),
.B2(n_374),
.Y(n_486)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_421),
.B(n_444),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_425),
.B(n_382),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_373),
.B(n_323),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_426),
.B(n_435),
.C(n_457),
.Y(n_459)
);

INVx4_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_427),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_429),
.A2(n_441),
.B(n_452),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_393),
.A2(n_326),
.B(n_308),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_SL g467 ( 
.A(n_434),
.B(n_454),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_SL g441 ( 
.A1(n_386),
.A2(n_316),
.B(n_325),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_391),
.A2(n_346),
.B1(n_343),
.B2(n_339),
.Y(n_442)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_442),
.A2(n_445),
.B1(n_449),
.B2(n_453),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_384),
.A2(n_346),
.B1(n_352),
.B2(n_348),
.Y(n_445)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_412),
.Y(n_446)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_446),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_447),
.B(n_456),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_391),
.A2(n_346),
.B1(n_323),
.B2(n_335),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_386),
.A2(n_332),
.B(n_340),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_372),
.A2(n_345),
.B1(n_314),
.B2(n_308),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_414),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_376),
.B(n_345),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g458 ( 
.A1(n_385),
.A2(n_387),
.B1(n_390),
.B2(n_407),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g463 ( 
.A1(n_458),
.A2(n_386),
.B(n_408),
.Y(n_463)
);

INVxp67_ASAP7_75t_L g509 ( 
.A(n_463),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_424),
.B(n_392),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g503 ( 
.A(n_465),
.B(n_480),
.Y(n_503)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_428),
.Y(n_466)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_466),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_443),
.A2(n_373),
.B(n_386),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_SL g512 ( 
.A(n_468),
.B(n_496),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_419),
.A2(n_372),
.B1(n_376),
.B2(n_378),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_469),
.A2(n_471),
.B1(n_479),
.B2(n_481),
.Y(n_499)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_428),
.Y(n_470)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_470),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_419),
.A2(n_408),
.B1(n_395),
.B2(n_369),
.Y(n_471)
);

XOR2xp5_ASAP7_75t_L g516 ( 
.A(n_472),
.B(n_484),
.Y(n_516)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_431),
.Y(n_473)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_473),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_448),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_474),
.B(n_475),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_454),
.B(n_412),
.Y(n_475)
);

OR2x2_ASAP7_75t_L g476 ( 
.A(n_427),
.B(n_408),
.Y(n_476)
);

CKINVDCx20_ASAP7_75t_R g498 ( 
.A(n_476),
.Y(n_498)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_431),
.Y(n_477)
);

INVx2_ASAP7_75t_SL g526 ( 
.A(n_477),
.Y(n_526)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_448),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_478),
.B(n_487),
.Y(n_513)
);

AOI22xp5_ASAP7_75t_L g479 ( 
.A1(n_443),
.A2(n_432),
.B1(n_445),
.B2(n_456),
.Y(n_479)
);

BUFx24_ASAP7_75t_SL g480 ( 
.A(n_424),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g481 ( 
.A(n_434),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g484 ( 
.A(n_425),
.B(n_388),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g485 ( 
.A(n_423),
.B(n_409),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_485),
.B(n_495),
.C(n_435),
.Y(n_501)
);

OAI22xp5_ASAP7_75t_L g518 ( 
.A1(n_486),
.A2(n_488),
.B1(n_492),
.B2(n_418),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_403),
.Y(n_487)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_429),
.A2(n_416),
.B(n_396),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_489),
.B(n_490),
.Y(n_521)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_436),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_436),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_491),
.B(n_493),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_433),
.A2(n_405),
.B1(n_381),
.B2(n_410),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_447),
.Y(n_493)
);

OAI21x1_ASAP7_75t_SL g494 ( 
.A1(n_433),
.A2(n_400),
.B(n_404),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_494),
.B(n_400),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_423),
.B(n_370),
.Y(n_495)
);

OAI21xp5_ASAP7_75t_L g496 ( 
.A1(n_439),
.A2(n_406),
.B(n_389),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g497 ( 
.A(n_495),
.B(n_423),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_497),
.B(n_525),
.Y(n_557)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_469),
.A2(n_433),
.B1(n_430),
.B2(n_439),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g564 ( 
.A1(n_500),
.A2(n_522),
.B1(n_476),
.B2(n_460),
.Y(n_564)
);

XNOR2xp5_ASAP7_75t_L g565 ( 
.A(n_501),
.B(n_502),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_484),
.B(n_435),
.C(n_457),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_485),
.B(n_380),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g549 ( 
.A(n_504),
.B(n_517),
.Y(n_549)
);

CKINVDCx16_ASAP7_75t_R g506 ( 
.A(n_475),
.Y(n_506)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_506),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_457),
.C(n_441),
.Y(n_507)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g510 ( 
.A1(n_468),
.A2(n_467),
.B(n_496),
.Y(n_510)
);

INVxp67_ASAP7_75t_L g562 ( 
.A(n_510),
.Y(n_562)
);

OAI22xp5_ASAP7_75t_SL g511 ( 
.A1(n_479),
.A2(n_458),
.B1(n_433),
.B2(n_421),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_511),
.A2(n_519),
.B1(n_520),
.B2(n_530),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_467),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_SL g544 ( 
.A1(n_518),
.A2(n_483),
.B1(n_461),
.B2(n_464),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g519 ( 
.A1(n_471),
.A2(n_420),
.B1(n_442),
.B2(n_449),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g520 ( 
.A1(n_492),
.A2(n_450),
.B1(n_453),
.B2(n_446),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_483),
.A2(n_450),
.B1(n_444),
.B2(n_427),
.Y(n_522)
);

AOI22xp5_ASAP7_75t_SL g523 ( 
.A1(n_474),
.A2(n_422),
.B1(n_451),
.B2(n_437),
.Y(n_523)
);

AO21x1_ASAP7_75t_L g535 ( 
.A1(n_523),
.A2(n_531),
.B(n_534),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_462),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_524),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_459),
.B(n_452),
.C(n_455),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g527 ( 
.A(n_462),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_527),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_472),
.B(n_455),
.C(n_440),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_529),
.B(n_533),
.Y(n_554)
);

OAI22xp5_ASAP7_75t_SL g530 ( 
.A1(n_488),
.A2(n_440),
.B1(n_438),
.B2(n_379),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_463),
.B(n_422),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_532),
.B(n_478),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_464),
.B(n_438),
.C(n_377),
.Y(n_533)
);

XOR2x2_ASAP7_75t_SL g534 ( 
.A(n_487),
.B(n_476),
.Y(n_534)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_508),
.Y(n_537)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_537),
.Y(n_571)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_508),
.Y(n_540)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_540),
.Y(n_572)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_542),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_513),
.B(n_493),
.Y(n_543)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_543),
.Y(n_578)
);

OAI22xp5_ASAP7_75t_L g581 ( 
.A1(n_544),
.A2(n_548),
.B1(n_559),
.B2(n_560),
.Y(n_581)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_521),
.A2(n_482),
.B(n_489),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_545),
.B(n_553),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_461),
.Y(n_546)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_546),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_528),
.B(n_466),
.Y(n_547)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

AOI22xp5_ASAP7_75t_L g548 ( 
.A1(n_499),
.A2(n_483),
.B1(n_494),
.B2(n_460),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_528),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_550),
.B(n_555),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g551 ( 
.A(n_526),
.B(n_491),
.Y(n_551)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_551),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_526),
.B(n_490),
.Y(n_552)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_552),
.Y(n_586)
);

BUFx12f_ASAP7_75t_SL g553 ( 
.A(n_509),
.Y(n_553)
);

CKINVDCx16_ASAP7_75t_R g555 ( 
.A(n_523),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_526),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_556),
.B(n_558),
.Y(n_595)
);

NAND3xp33_ASAP7_75t_SL g558 ( 
.A(n_513),
.B(n_437),
.C(n_482),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_505),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_505),
.Y(n_560)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_514),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g592 ( 
.A1(n_563),
.A2(n_566),
.B1(n_567),
.B2(n_515),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_SL g574 ( 
.A1(n_564),
.A2(n_511),
.B1(n_520),
.B2(n_519),
.Y(n_574)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_514),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_515),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_503),
.B(n_451),
.Y(n_568)
);

CKINVDCx16_ASAP7_75t_R g587 ( 
.A(n_568),
.Y(n_587)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_565),
.B(n_502),
.Y(n_569)
);

MAJx2_ASAP7_75t_L g619 ( 
.A(n_569),
.B(n_575),
.C(n_579),
.Y(n_619)
);

FAx1_ASAP7_75t_SL g573 ( 
.A(n_535),
.B(n_534),
.CI(n_512),
.CON(n_573),
.SN(n_573)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_573),
.B(n_535),
.Y(n_598)
);

OAI22xp5_ASAP7_75t_SL g605 ( 
.A1(n_574),
.A2(n_580),
.B1(n_541),
.B2(n_544),
.Y(n_605)
);

XOR2x2_ASAP7_75t_L g575 ( 
.A(n_542),
.B(n_532),
.Y(n_575)
);

XNOR2xp5_ASAP7_75t_L g577 ( 
.A(n_557),
.B(n_525),
.Y(n_577)
);

XNOR2xp5_ASAP7_75t_L g620 ( 
.A(n_577),
.B(n_596),
.Y(n_620)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_565),
.B(n_507),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g580 ( 
.A1(n_550),
.A2(n_564),
.B1(n_555),
.B2(n_537),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_557),
.B(n_516),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g607 ( 
.A(n_582),
.B(n_588),
.Y(n_607)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_561),
.B(n_497),
.C(n_501),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_583),
.B(n_585),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_554),
.B(n_516),
.C(n_529),
.Y(n_585)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_554),
.B(n_512),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_SL g589 ( 
.A1(n_548),
.A2(n_500),
.B1(n_522),
.B2(n_498),
.Y(n_589)
);

AOI22xp5_ASAP7_75t_L g608 ( 
.A1(n_589),
.A2(n_498),
.B1(n_547),
.B2(n_539),
.Y(n_608)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_592),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g593 ( 
.A(n_543),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_593),
.B(n_549),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_546),
.B(n_509),
.C(n_521),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_594),
.B(n_536),
.C(n_556),
.Y(n_599)
);

XNOR2xp5_ASAP7_75t_L g596 ( 
.A(n_535),
.B(n_531),
.Y(n_596)
);

XOR2xp5_ASAP7_75t_SL g635 ( 
.A(n_598),
.B(n_570),
.Y(n_635)
);

NOR2xp67_ASAP7_75t_SL g622 ( 
.A(n_599),
.B(n_604),
.Y(n_622)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_578),
.Y(n_601)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_601),
.Y(n_628)
);

INVxp67_ASAP7_75t_L g602 ( 
.A(n_594),
.Y(n_602)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_602),
.Y(n_637)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_597),
.Y(n_603)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_603),
.Y(n_642)
);

MAJIxp5_ASAP7_75t_L g604 ( 
.A(n_579),
.B(n_562),
.C(n_545),
.Y(n_604)
);

AOI22xp5_ASAP7_75t_L g639 ( 
.A1(n_605),
.A2(n_530),
.B1(n_573),
.B2(n_553),
.Y(n_639)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_569),
.B(n_541),
.C(n_540),
.Y(n_606)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_606),
.B(n_610),
.C(n_575),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_SL g627 ( 
.A1(n_608),
.A2(n_613),
.B1(n_584),
.B2(n_586),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_588),
.B(n_582),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_SL g638 ( 
.A(n_609),
.B(n_589),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_577),
.B(n_551),
.C(n_552),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_595),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g630 ( 
.A(n_611),
.B(n_616),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g613 ( 
.A1(n_581),
.A2(n_538),
.B1(n_539),
.B2(n_549),
.Y(n_613)
);

OAI21xp5_ASAP7_75t_L g614 ( 
.A1(n_570),
.A2(n_553),
.B(n_538),
.Y(n_614)
);

MAJx2_ASAP7_75t_L g634 ( 
.A(n_614),
.B(n_590),
.C(n_591),
.Y(n_634)
);

BUFx2_ASAP7_75t_L g631 ( 
.A(n_615),
.Y(n_631)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_587),
.B(n_568),
.Y(n_616)
);

CKINVDCx20_ASAP7_75t_R g617 ( 
.A(n_595),
.Y(n_617)
);

NOR2xp33_ASAP7_75t_L g625 ( 
.A(n_617),
.B(n_618),
.Y(n_625)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_586),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_585),
.B(n_536),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_621),
.B(n_572),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_623),
.B(n_626),
.Y(n_650)
);

XNOR2x1_ASAP7_75t_L g624 ( 
.A(n_604),
.B(n_590),
.Y(n_624)
);

XOR2xp5_ASAP7_75t_L g648 ( 
.A(n_624),
.B(n_638),
.Y(n_648)
);

MAJIxp5_ASAP7_75t_L g626 ( 
.A(n_606),
.B(n_583),
.C(n_576),
.Y(n_626)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_627),
.Y(n_652)
);

OAI22xp5_ASAP7_75t_SL g629 ( 
.A1(n_613),
.A2(n_580),
.B1(n_574),
.B2(n_571),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_629),
.B(n_641),
.Y(n_647)
);

FAx1_ASAP7_75t_SL g632 ( 
.A(n_598),
.B(n_573),
.CI(n_596),
.CON(n_632),
.SN(n_632)
);

OAI21xp5_ASAP7_75t_L g654 ( 
.A1(n_632),
.A2(n_620),
.B(n_607),
.Y(n_654)
);

MAJIxp5_ASAP7_75t_L g633 ( 
.A(n_612),
.B(n_576),
.C(n_590),
.Y(n_633)
);

HB1xp67_ASAP7_75t_L g658 ( 
.A(n_633),
.Y(n_658)
);

INVxp67_ASAP7_75t_L g645 ( 
.A(n_634),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_635),
.B(n_602),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g644 ( 
.A(n_636),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g656 ( 
.A1(n_639),
.A2(n_640),
.B1(n_559),
.B2(n_605),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_614),
.A2(n_567),
.B1(n_566),
.B2(n_563),
.Y(n_640)
);

XNOR2xp5_ASAP7_75t_L g641 ( 
.A(n_610),
.B(n_560),
.Y(n_641)
);

OAI22xp5_ASAP7_75t_L g643 ( 
.A1(n_631),
.A2(n_608),
.B1(n_601),
.B2(n_600),
.Y(n_643)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_643),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_L g646 ( 
.A1(n_625),
.A2(n_600),
.B1(n_603),
.B2(n_618),
.Y(n_646)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_646),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_649),
.B(n_651),
.Y(n_671)
);

MAJIxp5_ASAP7_75t_L g651 ( 
.A(n_626),
.B(n_599),
.C(n_619),
.Y(n_651)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_631),
.B(n_620),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g664 ( 
.A(n_653),
.Y(n_664)
);

XOR2xp5_ASAP7_75t_L g660 ( 
.A(n_654),
.B(n_655),
.Y(n_660)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_641),
.B(n_619),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_SL g672 ( 
.A1(n_656),
.A2(n_642),
.B1(n_628),
.B2(n_632),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g657 ( 
.A(n_630),
.B(n_371),
.Y(n_657)
);

XNOR2xp5_ASAP7_75t_L g661 ( 
.A(n_657),
.B(n_659),
.Y(n_661)
);

XOR2xp5_ASAP7_75t_L g659 ( 
.A(n_624),
.B(n_607),
.Y(n_659)
);

MAJIxp5_ASAP7_75t_L g662 ( 
.A(n_658),
.B(n_637),
.C(n_622),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_662),
.B(n_663),
.Y(n_680)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_655),
.B(n_633),
.Y(n_663)
);

A2O1A1Ixp33_ASAP7_75t_SL g665 ( 
.A1(n_649),
.A2(n_634),
.B(n_639),
.C(n_635),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_665),
.B(n_645),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_644),
.B(n_623),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_SL g675 ( 
.A(n_667),
.B(n_647),
.Y(n_675)
);

MAJIxp5_ASAP7_75t_L g669 ( 
.A(n_651),
.B(n_638),
.C(n_609),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_669),
.B(n_670),
.Y(n_681)
);

XNOR2xp5_ASAP7_75t_L g670 ( 
.A(n_648),
.B(n_640),
.Y(n_670)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_672),
.Y(n_679)
);

OAI21x1_ASAP7_75t_SL g685 ( 
.A1(n_673),
.A2(n_676),
.B(n_654),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_671),
.B(n_650),
.Y(n_674)
);

CKINVDCx20_ASAP7_75t_R g686 ( 
.A(n_674),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_675),
.B(n_677),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_662),
.B(n_648),
.Y(n_676)
);

MAJIxp5_ASAP7_75t_L g677 ( 
.A(n_664),
.B(n_652),
.C(n_645),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_SL g678 ( 
.A(n_661),
.B(n_649),
.Y(n_678)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_678),
.B(n_669),
.Y(n_683)
);

OAI22xp33_ASAP7_75t_L g682 ( 
.A1(n_679),
.A2(n_666),
.B1(n_668),
.B2(n_646),
.Y(n_682)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_682),
.A2(n_685),
.B(n_681),
.Y(n_689)
);

O2A1O1Ixp33_ASAP7_75t_SL g690 ( 
.A1(n_683),
.A2(n_684),
.B(n_665),
.C(n_660),
.Y(n_690)
);

AOI22xp33_ASAP7_75t_L g684 ( 
.A1(n_673),
.A2(n_665),
.B1(n_470),
.B2(n_473),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_687),
.B(n_680),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_688),
.B(n_689),
.Y(n_692)
);

OAI311xp33_ASAP7_75t_L g691 ( 
.A1(n_690),
.A2(n_665),
.A3(n_686),
.B1(n_660),
.C1(n_632),
.Y(n_691)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_691),
.B(n_659),
.C(n_477),
.Y(n_693)
);

OAI21xp5_ASAP7_75t_SL g694 ( 
.A1(n_693),
.A2(n_692),
.B(n_394),
.Y(n_694)
);

MAJIxp5_ASAP7_75t_L g695 ( 
.A(n_694),
.B(n_398),
.C(n_399),
.Y(n_695)
);

MAJIxp5_ASAP7_75t_L g696 ( 
.A(n_695),
.B(n_411),
.C(n_397),
.Y(n_696)
);

MAJx2_ASAP7_75t_L g697 ( 
.A(n_696),
.B(n_400),
.C(n_402),
.Y(n_697)
);


endmodule