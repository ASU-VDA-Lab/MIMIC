module fake_jpeg_11260_n_534 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_534);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_534;

wire n_529;
wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_16),
.B(n_18),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx4f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_8),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_8),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_9),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_12),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_53),
.Y(n_107)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_55),
.Y(n_162)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx4f_ASAP7_75t_SL g111 ( 
.A(n_56),
.Y(n_111)
);

AOI21xp33_ASAP7_75t_L g57 ( 
.A1(n_22),
.A2(n_18),
.B(n_16),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_57),
.B(n_1),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_22),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_58),
.B(n_99),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_59),
.Y(n_129)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx5_ASAP7_75t_L g112 ( 
.A(n_60),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_34),
.B(n_15),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_66),
.Y(n_106)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_30),
.Y(n_63)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_63),
.Y(n_126)
);

HB1xp67_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_64),
.Y(n_133)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_30),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_46),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_69),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

BUFx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

INVx4_ASAP7_75t_SL g72 ( 
.A(n_21),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g146 ( 
.A(n_72),
.Y(n_146)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_26),
.Y(n_73)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_74),
.Y(n_149)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_75),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_76),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx8_ASAP7_75t_L g144 ( 
.A(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_40),
.Y(n_80)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_80),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_81),
.Y(n_154)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_83),
.Y(n_139)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_84),
.Y(n_124)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

BUFx12f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_51),
.Y(n_88)
);

INVx4_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_89),
.B(n_91),
.Y(n_108)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_28),
.Y(n_90)
);

BUFx10_ASAP7_75t_L g158 ( 
.A(n_90),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_25),
.B(n_15),
.Y(n_91)
);

BUFx16f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_98),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_93),
.B(n_94),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_25),
.B(n_15),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_33),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_95),
.B(n_96),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_20),
.Y(n_96)
);

INVx13_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_97),
.Y(n_125)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_28),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_37),
.B(n_0),
.Y(n_99)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_101),
.Y(n_114)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_26),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_20),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_102),
.B(n_104),
.Y(n_127)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_43),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_103),
.B(n_48),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_24),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_53),
.A2(n_43),
.B1(n_50),
.B2(n_29),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_105),
.A2(n_45),
.B1(n_47),
.B2(n_42),
.Y(n_164)
);

NOR2xp67_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_27),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_117),
.B(n_145),
.Y(n_181)
);

NOR4xp25_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_1),
.C(n_2),
.D(n_3),
.Y(n_118)
);

NAND3xp33_ASAP7_75t_L g173 ( 
.A(n_118),
.B(n_1),
.C(n_2),
.Y(n_173)
);

OAI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_43),
.B1(n_39),
.B2(n_24),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_120),
.A2(n_122),
.B1(n_123),
.B2(n_31),
.Y(n_196)
);

OAI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_102),
.A2(n_39),
.B1(n_50),
.B2(n_29),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_85),
.A2(n_39),
.B1(n_49),
.B2(n_32),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_92),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_130),
.B(n_132),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_61),
.B(n_45),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_64),
.A2(n_49),
.B1(n_32),
.B2(n_19),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_134),
.A2(n_124),
.B(n_146),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_60),
.A2(n_49),
.B1(n_32),
.B2(n_19),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_141),
.A2(n_147),
.B1(n_159),
.B2(n_98),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_143),
.B(n_150),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_56),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_90),
.A2(n_49),
.B1(n_32),
.B2(n_23),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_100),
.B(n_41),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_56),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_155),
.B(n_111),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_157),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_103),
.A2(n_86),
.B1(n_80),
.B2(n_81),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_164),
.A2(n_174),
.B1(n_179),
.B2(n_185),
.Y(n_233)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_133),
.Y(n_165)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_126),
.Y(n_166)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_166),
.Y(n_253)
);

AOI22xp33_ASAP7_75t_SL g248 ( 
.A1(n_167),
.A2(n_187),
.B1(n_221),
.B2(n_201),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_108),
.B(n_104),
.C(n_83),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_168),
.B(n_128),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_114),
.Y(n_169)
);

INVx4_ASAP7_75t_SL g267 ( 
.A(n_169),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g170 ( 
.A(n_107),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g171 ( 
.A(n_144),
.Y(n_171)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_171),
.Y(n_268)
);

BUFx2_ASAP7_75t_SL g172 ( 
.A(n_146),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_172),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_173),
.B(n_184),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_156),
.A2(n_74),
.B1(n_67),
.B2(n_68),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_115),
.B(n_23),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_175),
.B(n_176),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_48),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_133),
.Y(n_177)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_177),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_72),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_178),
.B(n_206),
.Y(n_237)
);

OAI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_157),
.A2(n_93),
.B1(n_88),
.B2(n_59),
.Y(n_179)
);

A2O1A1Ixp33_ASAP7_75t_L g180 ( 
.A1(n_106),
.A2(n_27),
.B(n_47),
.C(n_42),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g264 ( 
.A(n_180),
.B(n_208),
.Y(n_264)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_126),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_135),
.Y(n_183)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_183),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_159),
.A2(n_77),
.B1(n_76),
.B2(n_69),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_135),
.Y(n_186)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_186),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_123),
.A2(n_49),
.B1(n_41),
.B2(n_35),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_148),
.Y(n_188)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_188),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_189),
.B(n_190),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_158),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_191),
.B(n_192),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_124),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_131),
.A2(n_100),
.B1(n_35),
.B2(n_31),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g243 ( 
.A1(n_193),
.A2(n_137),
.B(n_154),
.Y(n_243)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_148),
.Y(n_194)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_194),
.Y(n_263)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_196),
.Y(n_240)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_105),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_197),
.A2(n_199),
.B1(n_201),
.B2(n_205),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_160),
.A2(n_134),
.B1(n_127),
.B2(n_147),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_121),
.B(n_3),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_202),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_141),
.A2(n_13),
.B1(n_4),
.B2(n_5),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_3),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_149),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_163),
.B1(n_136),
.B2(n_129),
.Y(n_224)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_151),
.Y(n_204)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_131),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_125),
.B(n_10),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_207),
.B(n_209),
.Y(n_258)
);

A2O1A1Ixp33_ASAP7_75t_L g208 ( 
.A1(n_146),
.A2(n_10),
.B(n_11),
.C(n_12),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_113),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_111),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g229 ( 
.A(n_210),
.B(n_212),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_211),
.Y(n_223)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_113),
.Y(n_212)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVx4_ASAP7_75t_L g265 ( 
.A(n_214),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_144),
.B(n_153),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_215),
.B(n_139),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_111),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_216),
.B(n_217),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_137),
.B(n_10),
.Y(n_217)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_107),
.Y(n_219)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_219),
.Y(n_254)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_109),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_220),
.B(n_191),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_119),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_196),
.A2(n_109),
.B1(n_153),
.B2(n_149),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_222),
.A2(n_224),
.B1(n_242),
.B2(n_260),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_199),
.A2(n_163),
.B1(n_152),
.B2(n_129),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_225),
.A2(n_226),
.B1(n_262),
.B2(n_171),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g226 ( 
.A1(n_198),
.A2(n_152),
.B1(n_136),
.B2(n_119),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_175),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_238),
.B(n_184),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_170),
.Y(n_239)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_239),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_128),
.B1(n_154),
.B2(n_112),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_243),
.B(n_214),
.Y(n_310)
);

O2A1O1Ixp33_ASAP7_75t_L g244 ( 
.A1(n_208),
.A2(n_112),
.B(n_116),
.C(n_138),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_206),
.B(n_216),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_245),
.B(n_178),
.Y(n_282)
);

BUFx5_ASAP7_75t_L g247 ( 
.A(n_220),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_247),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_248),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_178),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_250),
.B(n_271),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_255),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_202),
.B(n_13),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_176),
.A2(n_139),
.B1(n_161),
.B2(n_116),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_L g261 ( 
.A1(n_168),
.A2(n_161),
.B1(n_138),
.B2(n_13),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_272),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_174),
.A2(n_138),
.B1(n_161),
.B2(n_164),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_266),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_215),
.A2(n_193),
.B1(n_181),
.B2(n_213),
.Y(n_270)
);

AOI22xp33_ASAP7_75t_L g312 ( 
.A1(n_270),
.A2(n_204),
.B1(n_205),
.B2(n_192),
.Y(n_312)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_213),
.B(n_207),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_206),
.B(n_200),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_257),
.Y(n_273)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_273),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_229),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_275),
.B(n_277),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g277 ( 
.A(n_269),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_245),
.B(n_169),
.C(n_218),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_278),
.B(n_282),
.C(n_290),
.Y(n_347)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_227),
.Y(n_280)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_280),
.Y(n_352)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_283),
.B(n_304),
.Y(n_338)
);

AO22x2_ASAP7_75t_L g284 ( 
.A1(n_243),
.A2(n_171),
.B1(n_195),
.B2(n_209),
.Y(n_284)
);

A2O1A1Ixp33_ASAP7_75t_SL g343 ( 
.A1(n_284),
.A2(n_240),
.B(n_267),
.C(n_249),
.Y(n_343)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_227),
.Y(n_285)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_285),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_286),
.B(n_294),
.Y(n_345)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_230),
.Y(n_287)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_287),
.Y(n_323)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_288),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_237),
.B(n_194),
.C(n_188),
.Y(n_290)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_254),
.Y(n_291)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_291),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_217),
.B(n_180),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_292),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_212),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_263),
.Y(n_295)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_295),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_237),
.B(n_165),
.C(n_177),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_296),
.B(n_300),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_190),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_297),
.B(n_305),
.Y(n_348)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_298),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_238),
.B(n_166),
.C(n_186),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_228),
.B(n_189),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_301),
.B(n_234),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_246),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_302),
.B(n_303),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_258),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_231),
.B(n_264),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_230),
.Y(n_306)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_306),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_228),
.B(n_236),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_313),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_182),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_311),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_310),
.A2(n_251),
.B(n_244),
.Y(n_326)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_312),
.A2(n_233),
.B1(n_256),
.B2(n_268),
.Y(n_341)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_258),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g314 ( 
.A(n_258),
.Y(n_314)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_314),
.Y(n_333)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_232),
.Y(n_315)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_315),
.Y(n_358)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_232),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_319),
.Y(n_344)
);

INVx13_ASAP7_75t_L g317 ( 
.A(n_251),
.Y(n_317)
);

BUFx12f_ASAP7_75t_L g320 ( 
.A(n_317),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_252),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g322 ( 
.A(n_318),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_255),
.B(n_183),
.Y(n_319)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_325),
.B(n_329),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g373 ( 
.A(n_326),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_273),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_288),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_331),
.B(n_360),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_307),
.A2(n_240),
.B1(n_222),
.B2(n_264),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g392 ( 
.A1(n_332),
.A2(n_342),
.B1(n_254),
.B2(n_281),
.Y(n_392)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_292),
.Y(n_336)
);

INVxp67_ASAP7_75t_L g378 ( 
.A(n_336),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_307),
.A2(n_256),
.B1(n_233),
.B2(n_262),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_340),
.A2(n_349),
.B1(n_350),
.B2(n_289),
.Y(n_370)
);

CKINVDCx14_ASAP7_75t_R g368 ( 
.A(n_341),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_304),
.A2(n_240),
.B1(n_224),
.B2(n_261),
.Y(n_342)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_343),
.A2(n_354),
.B(n_359),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_SL g349 ( 
.A1(n_294),
.A2(n_299),
.B1(n_314),
.B2(n_313),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_299),
.A2(n_272),
.B1(n_203),
.B2(n_241),
.Y(n_350)
);

A2O1A1O1Ixp25_ASAP7_75t_L g354 ( 
.A1(n_293),
.A2(n_267),
.B(n_249),
.C(n_234),
.D(n_247),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g375 ( 
.A(n_356),
.B(n_290),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_283),
.A2(n_267),
.B(n_265),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_357),
.A2(n_279),
.B(n_282),
.Y(n_366)
);

OAI22x1_ASAP7_75t_L g359 ( 
.A1(n_279),
.A2(n_268),
.B1(n_265),
.B2(n_219),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_295),
.Y(n_360)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_310),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_361),
.B(n_298),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_321),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_363),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_322),
.B(n_309),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_344),
.B(n_335),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_369),
.Y(n_419)
);

OAI21xp5_ASAP7_75t_SL g414 ( 
.A1(n_366),
.A2(n_386),
.B(n_387),
.Y(n_414)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_328),
.Y(n_367)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_367),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_344),
.B(n_276),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g428 ( 
.A1(n_370),
.A2(n_376),
.B1(n_334),
.B2(n_352),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_278),
.C(n_301),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_372),
.B(n_347),
.C(n_355),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g374 ( 
.A1(n_357),
.A2(n_284),
.B(n_274),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_L g426 ( 
.A1(n_374),
.A2(n_388),
.B(n_396),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g411 ( 
.A(n_375),
.B(n_350),
.Y(n_411)
);

OAI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_342),
.A2(n_289),
.B1(n_284),
.B2(n_302),
.Y(n_376)
);

CKINVDCx20_ASAP7_75t_R g377 ( 
.A(n_335),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_384),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_327),
.B(n_276),
.Y(n_380)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_380),
.Y(n_416)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_328),
.Y(n_381)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_381),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g383 ( 
.A(n_338),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_339),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_345),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g385 ( 
.A1(n_346),
.A2(n_284),
.B(n_296),
.Y(n_385)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_385),
.Y(n_415)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_338),
.A2(n_326),
.B(n_343),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_346),
.A2(n_284),
.B(n_300),
.Y(n_387)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_338),
.A2(n_354),
.B(n_333),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_358),
.B(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_389),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_348),
.B(n_316),
.Y(n_390)
);

NAND3xp33_ASAP7_75t_L g402 ( 
.A(n_390),
.B(n_394),
.C(n_353),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g391 ( 
.A1(n_332),
.A2(n_280),
.B1(n_287),
.B2(n_291),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_391),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g417 ( 
.A(n_392),
.B(n_395),
.Y(n_417)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_337),
.Y(n_393)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_393),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_351),
.B(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_337),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g396 ( 
.A1(n_349),
.A2(n_274),
.B(n_317),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_358),
.B(n_281),
.Y(n_397)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_397),
.Y(n_399)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_400),
.B(n_409),
.C(n_412),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g401 ( 
.A1(n_370),
.A2(n_340),
.B1(n_343),
.B2(n_324),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g435 ( 
.A1(n_401),
.A2(n_428),
.B1(n_392),
.B2(n_391),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_402),
.B(n_407),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_375),
.B(n_355),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_376),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_362),
.Y(n_406)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_371),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_408),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_356),
.C(n_343),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_411),
.B(n_364),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_372),
.B(n_375),
.C(n_366),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_366),
.B(n_343),
.C(n_330),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_413),
.B(n_423),
.C(n_386),
.Y(n_444)
);

OAI21xp33_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_339),
.B(n_353),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_371),
.Y(n_440)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_422),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_323),
.C(n_334),
.Y(n_423)
);

FAx1_ASAP7_75t_SL g425 ( 
.A(n_369),
.B(n_359),
.CI(n_323),
.CON(n_425),
.SN(n_425)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_425),
.B(n_379),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_404),
.B(n_388),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_430),
.B(n_433),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_416),
.A2(n_370),
.B1(n_380),
.B2(n_390),
.Y(n_431)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_431),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_405),
.A2(n_363),
.B1(n_396),
.B2(n_365),
.Y(n_432)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_432),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_400),
.B(n_387),
.Y(n_433)
);

XOR2xp5_ASAP7_75t_L g462 ( 
.A(n_434),
.B(n_444),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_435),
.A2(n_427),
.B1(n_396),
.B2(n_421),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_406),
.B(n_378),
.Y(n_438)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_438),
.B(n_443),
.Y(n_458)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_440),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_409),
.B(n_386),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_441),
.B(n_449),
.Y(n_464)
);

NAND3xp33_ASAP7_75t_SL g461 ( 
.A(n_442),
.B(n_379),
.C(n_399),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_424),
.B(n_365),
.Y(n_443)
);

XNOR2x1_ASAP7_75t_L g445 ( 
.A(n_423),
.B(n_383),
.Y(n_445)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_445),
.B(n_448),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_424),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_447),
.B(n_452),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_411),
.Y(n_449)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_415),
.B(n_373),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_450),
.B(n_426),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_415),
.B(n_414),
.C(n_413),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_451),
.B(n_453),
.C(n_426),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_419),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_414),
.B(n_382),
.C(n_391),
.Y(n_453)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_410),
.A2(n_389),
.B(n_397),
.Y(n_454)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_454),
.Y(n_468)
);

MAJx2_ASAP7_75t_L g491 ( 
.A(n_456),
.B(n_465),
.C(n_474),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_439),
.B(n_410),
.Y(n_460)
);

NAND3xp33_ASAP7_75t_L g490 ( 
.A(n_460),
.B(n_471),
.C(n_474),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_461),
.A2(n_394),
.B(n_352),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_467),
.A2(n_469),
.B1(n_368),
.B2(n_446),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g469 ( 
.A1(n_453),
.A2(n_377),
.B1(n_374),
.B2(n_401),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g470 ( 
.A(n_429),
.B(n_417),
.C(n_374),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g480 ( 
.A(n_470),
.B(n_475),
.C(n_449),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_440),
.B(n_425),
.Y(n_471)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_434),
.A2(n_417),
.B1(n_368),
.B2(n_425),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g476 ( 
.A1(n_472),
.A2(n_444),
.B1(n_451),
.B2(n_445),
.Y(n_476)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_433),
.B(n_417),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_429),
.B(n_403),
.C(n_418),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_477),
.Y(n_495)
);

A2O1A1O1Ixp25_ASAP7_75t_L g478 ( 
.A1(n_468),
.A2(n_448),
.B(n_430),
.C(n_441),
.D(n_446),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_478),
.B(n_480),
.Y(n_496)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_466),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_479),
.A2(n_482),
.B1(n_486),
.B2(n_488),
.Y(n_493)
);

NOR2xp33_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_436),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_SL g497 ( 
.A(n_481),
.B(n_492),
.Y(n_497)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_475),
.B(n_450),
.C(n_437),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_483),
.B(n_462),
.C(n_464),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_467),
.B(n_408),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_484),
.B(n_485),
.Y(n_494)
);

OA21x2_ASAP7_75t_L g485 ( 
.A1(n_469),
.A2(n_398),
.B(n_395),
.Y(n_485)
);

OAI21x1_ASAP7_75t_SL g486 ( 
.A1(n_459),
.A2(n_393),
.B(n_381),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_487),
.A2(n_472),
.B1(n_465),
.B2(n_473),
.Y(n_499)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_455),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_456),
.A2(n_320),
.B(n_253),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_490),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_470),
.B(n_320),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_498),
.B(n_499),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_483),
.B(n_462),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_505),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g501 ( 
.A(n_480),
.B(n_464),
.Y(n_501)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_501),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_457),
.Y(n_503)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_503),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_485),
.B(n_457),
.Y(n_504)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_504),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_477),
.A2(n_473),
.B1(n_235),
.B2(n_239),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_484),
.B(n_320),
.Y(n_506)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_506),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_496),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g521 ( 
.A(n_509),
.B(n_516),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g511 ( 
.A(n_498),
.B(n_478),
.Y(n_511)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_511),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_SL g513 ( 
.A1(n_502),
.A2(n_491),
.B(n_487),
.Y(n_513)
);

OAI21xp5_ASAP7_75t_SL g520 ( 
.A1(n_513),
.A2(n_517),
.B(n_504),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_497),
.B(n_484),
.Y(n_516)
);

NOR2xp67_ASAP7_75t_SL g517 ( 
.A(n_502),
.B(n_476),
.Y(n_517)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_512),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_519),
.B(n_522),
.Y(n_526)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_520),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_SL g522 ( 
.A1(n_507),
.A2(n_503),
.B1(n_494),
.B2(n_506),
.Y(n_522)
);

FAx1_ASAP7_75t_SL g523 ( 
.A(n_508),
.B(n_494),
.CI(n_493),
.CON(n_523),
.SN(n_523)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_523),
.B(n_524),
.Y(n_527)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_510),
.A2(n_495),
.B1(n_489),
.B2(n_491),
.Y(n_524)
);

INVxp67_ASAP7_75t_L g525 ( 
.A(n_521),
.Y(n_525)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_525),
.Y(n_530)
);

OAI311xp33_ASAP7_75t_L g529 ( 
.A1(n_526),
.A2(n_523),
.A3(n_515),
.B1(n_495),
.C1(n_514),
.Y(n_529)
);

AOI21xp33_ASAP7_75t_L g532 ( 
.A1(n_529),
.A2(n_235),
.B(n_259),
.Y(n_532)
);

AOI322xp5_ASAP7_75t_L g531 ( 
.A1(n_530),
.A2(n_528),
.A3(n_519),
.B1(n_518),
.B2(n_516),
.C1(n_527),
.C2(n_320),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_531),
.B(n_532),
.C(n_170),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_533),
.B(n_259),
.Y(n_534)
);


endmodule