module fake_netlist_5_1490_n_2157 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_223, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_222, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2157);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_223;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_222;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2157;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_2022;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_677;
wire n_293;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_604;
wire n_433;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1400;
wire n_1342;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_1115;
wire n_980;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1996;
wire n_597;
wire n_1879;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g224 ( 
.A(n_155),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_20),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_65),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_13),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_161),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_66),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_6),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_222),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_104),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_187),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_24),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_159),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

BUFx10_ASAP7_75t_L g238 ( 
.A(n_23),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_31),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

CKINVDCx14_ASAP7_75t_R g241 ( 
.A(n_57),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_71),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_79),
.Y(n_243)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_70),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_101),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_192),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_184),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_124),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_59),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_219),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_19),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_47),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_5),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_129),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_151),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_158),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_29),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_70),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_200),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_152),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_107),
.Y(n_263)
);

HB1xp67_ASAP7_75t_L g264 ( 
.A(n_93),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_24),
.Y(n_265)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_77),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_135),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_143),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_7),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_52),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_19),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_59),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_45),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_204),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_132),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_168),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_94),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_213),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_17),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_99),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_193),
.Y(n_281)
);

CKINVDCx14_ASAP7_75t_R g282 ( 
.A(n_54),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_206),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_78),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_174),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_140),
.Y(n_286)
);

BUFx10_ASAP7_75t_L g287 ( 
.A(n_22),
.Y(n_287)
);

BUFx10_ASAP7_75t_L g288 ( 
.A(n_57),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_115),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_51),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_123),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_51),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_172),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_66),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_160),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_139),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_191),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_178),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_167),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_2),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_202),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_52),
.Y(n_302)
);

BUFx2_ASAP7_75t_L g303 ( 
.A(n_95),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_11),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_48),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_56),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_162),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_119),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_46),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_61),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_218),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_0),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_73),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_5),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_31),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_86),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_89),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_212),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_23),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g320 ( 
.A(n_12),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_54),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_41),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_69),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_68),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_190),
.Y(n_325)
);

BUFx2_ASAP7_75t_SL g326 ( 
.A(n_196),
.Y(n_326)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_125),
.Y(n_327)
);

BUFx3_ASAP7_75t_L g328 ( 
.A(n_199),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_157),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_34),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_147),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_18),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_40),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_28),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_102),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_75),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_189),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_114),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_91),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_153),
.Y(n_342)
);

BUFx10_ASAP7_75t_L g343 ( 
.A(n_138),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_164),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_98),
.Y(n_345)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_183),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_180),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_131),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_118),
.Y(n_349)
);

CKINVDCx14_ASAP7_75t_R g350 ( 
.A(n_173),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_154),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_10),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_142),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_150),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_127),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_75),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_113),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_40),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_74),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_67),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g361 ( 
.A(n_16),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_194),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_111),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_16),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_121),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_148),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_39),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_67),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_26),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_71),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_48),
.Y(n_371)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_84),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_117),
.Y(n_373)
);

BUFx3_ASAP7_75t_L g374 ( 
.A(n_76),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_34),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_198),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_76),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_69),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_9),
.Y(n_379)
);

INVx2_ASAP7_75t_L g380 ( 
.A(n_43),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_96),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_217),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_90),
.Y(n_383)
);

BUFx10_ASAP7_75t_L g384 ( 
.A(n_10),
.Y(n_384)
);

BUFx10_ASAP7_75t_L g385 ( 
.A(n_85),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_110),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_42),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_106),
.Y(n_388)
);

BUFx5_ASAP7_75t_L g389 ( 
.A(n_1),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_188),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_137),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_223),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_122),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_136),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_100),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_92),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_25),
.Y(n_397)
);

INVxp67_ASAP7_75t_R g398 ( 
.A(n_203),
.Y(n_398)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_33),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_13),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_15),
.Y(n_401)
);

BUFx10_ASAP7_75t_L g402 ( 
.A(n_3),
.Y(n_402)
);

BUFx10_ASAP7_75t_L g403 ( 
.A(n_108),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_185),
.Y(n_404)
);

BUFx3_ASAP7_75t_L g405 ( 
.A(n_68),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_64),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_175),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_82),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_65),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_41),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_30),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_61),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_7),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_30),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_103),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_17),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_37),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_221),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_3),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_35),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_216),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_50),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_27),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_145),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_109),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_182),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_72),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_208),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_134),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_177),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_80),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_201),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_81),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_88),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_171),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_112),
.Y(n_436)
);

INVx1_ASAP7_75t_SL g437 ( 
.A(n_1),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_105),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_20),
.Y(n_439)
);

INVx2_ASAP7_75t_SL g440 ( 
.A(n_83),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_389),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_231),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_389),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_389),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_389),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_389),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_265),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_389),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_389),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_241),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_233),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_244),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_234),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_244),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_315),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_296),
.Y(n_457)
);

BUFx6f_ASAP7_75t_SL g458 ( 
.A(n_240),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_282),
.Y(n_459)
);

INVx2_ASAP7_75t_L g460 ( 
.A(n_244),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_370),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_299),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_315),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_315),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_315),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_252),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_320),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_315),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_301),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_252),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g471 ( 
.A(n_357),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_252),
.Y(n_472)
);

BUFx6f_ASAP7_75t_SL g473 ( 
.A(n_240),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_401),
.B(n_0),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_333),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_308),
.Y(n_476)
);

INVxp67_ASAP7_75t_SL g477 ( 
.A(n_264),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_290),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_333),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_294),
.Y(n_480)
);

CKINVDCx20_ASAP7_75t_R g481 ( 
.A(n_372),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_350),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_253),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_275),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_253),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_302),
.Y(n_486)
);

INVxp67_ASAP7_75t_L g487 ( 
.A(n_306),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_276),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_332),
.Y(n_489)
);

BUFx2_ASAP7_75t_L g490 ( 
.A(n_332),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_304),
.Y(n_491)
);

CKINVDCx20_ASAP7_75t_R g492 ( 
.A(n_277),
.Y(n_492)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_283),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_374),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_374),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_225),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_405),
.Y(n_497)
);

INVxp67_ASAP7_75t_L g498 ( 
.A(n_238),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_405),
.Y(n_499)
);

INVxp67_ASAP7_75t_SL g500 ( 
.A(n_254),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_333),
.Y(n_501)
);

BUFx2_ASAP7_75t_L g502 ( 
.A(n_225),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_309),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_333),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_333),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_310),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_284),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_361),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_361),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_361),
.Y(n_510)
);

CKINVDCx20_ASAP7_75t_R g511 ( 
.A(n_286),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_361),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_229),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_361),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_313),
.Y(n_515)
);

BUFx2_ASAP7_75t_L g516 ( 
.A(n_226),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

CKINVDCx20_ASAP7_75t_R g518 ( 
.A(n_289),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_399),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_295),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_298),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_399),
.Y(n_522)
);

HB1xp67_ASAP7_75t_L g523 ( 
.A(n_226),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_399),
.Y(n_524)
);

OR2x2_ASAP7_75t_L g525 ( 
.A(n_227),
.B(n_2),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_314),
.Y(n_526)
);

INVxp67_ASAP7_75t_L g527 ( 
.A(n_238),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_316),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_303),
.B(n_4),
.Y(n_529)
);

INVxp67_ASAP7_75t_SL g530 ( 
.A(n_308),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_230),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_399),
.Y(n_532)
);

HB1xp67_ASAP7_75t_L g533 ( 
.A(n_230),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_322),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_232),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_235),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_323),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_237),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_273),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g540 ( 
.A(n_328),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_237),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_239),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_324),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_280),
.B(n_4),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_330),
.Y(n_545)
);

INVxp67_ASAP7_75t_SL g546 ( 
.A(n_328),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_273),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_292),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_280),
.B(n_318),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_336),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_292),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_339),
.Y(n_552)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_317),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_335),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_318),
.B(n_6),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_259),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_380),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_354),
.B(n_8),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_444),
.Y(n_559)
);

BUFx8_ASAP7_75t_L g560 ( 
.A(n_458),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_456),
.Y(n_561)
);

AND2x2_ASAP7_75t_SL g562 ( 
.A(n_555),
.B(n_266),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_456),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_451),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_463),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_463),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_460),
.B(n_354),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_464),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_464),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g570 ( 
.A(n_453),
.B(n_440),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_444),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_446),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_549),
.B(n_440),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_465),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_496),
.Y(n_575)
);

BUFx6f_ASAP7_75t_L g576 ( 
.A(n_446),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_530),
.B(n_228),
.Y(n_577)
);

BUFx6f_ASAP7_75t_L g578 ( 
.A(n_447),
.Y(n_578)
);

INVx6_ASAP7_75t_L g579 ( 
.A(n_476),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_465),
.Y(n_580)
);

INVx3_ASAP7_75t_L g581 ( 
.A(n_447),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_450),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_450),
.Y(n_583)
);

INVxp67_ASAP7_75t_L g584 ( 
.A(n_523),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_445),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_441),
.Y(n_586)
);

AND2x4_ASAP7_75t_L g587 ( 
.A(n_460),
.B(n_266),
.Y(n_587)
);

AND2x2_ASAP7_75t_SL g588 ( 
.A(n_529),
.B(n_278),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_449),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_468),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_540),
.B(n_228),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_468),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_544),
.B(n_558),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_441),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_443),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_475),
.Y(n_596)
);

OA21x2_ASAP7_75t_L g597 ( 
.A1(n_443),
.A2(n_387),
.B(n_380),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_475),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_479),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_510),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_546),
.B(n_236),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_510),
.Y(n_603)
);

NOR2xp33_ASAP7_75t_L g604 ( 
.A(n_500),
.B(n_477),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_512),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_455),
.B(n_278),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_476),
.B(n_325),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_512),
.Y(n_608)
);

HB1xp67_ASAP7_75t_L g609 ( 
.A(n_531),
.Y(n_609)
);

INVx3_ASAP7_75t_L g610 ( 
.A(n_514),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_514),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_517),
.Y(n_612)
);

INVx3_ASAP7_75t_L g613 ( 
.A(n_517),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_519),
.Y(n_614)
);

AND2x4_ASAP7_75t_L g615 ( 
.A(n_466),
.B(n_325),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_501),
.B(n_236),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_519),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_522),
.Y(n_618)
);

INVx3_ASAP7_75t_L g619 ( 
.A(n_522),
.Y(n_619)
);

AND2x4_ASAP7_75t_L g620 ( 
.A(n_466),
.B(n_327),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_524),
.Y(n_621)
);

CKINVDCx20_ASAP7_75t_R g622 ( 
.A(n_442),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_524),
.Y(n_623)
);

AND2x4_ASAP7_75t_L g624 ( 
.A(n_470),
.B(n_327),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_532),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_532),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_470),
.B(n_329),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_472),
.Y(n_628)
);

HB1xp67_ASAP7_75t_L g629 ( 
.A(n_533),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_504),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_505),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_508),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_509),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_472),
.B(n_483),
.Y(n_634)
);

NAND2xp5_ASAP7_75t_L g635 ( 
.A(n_485),
.B(n_243),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_539),
.Y(n_636)
);

AND2x4_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_329),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_547),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_547),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_548),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_548),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_551),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_489),
.B(n_243),
.Y(n_643)
);

BUFx6f_ASAP7_75t_L g644 ( 
.A(n_551),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_451),
.B(n_240),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_484),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_494),
.B(n_245),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_459),
.B(n_343),
.Y(n_648)
);

INVxp67_ASAP7_75t_L g649 ( 
.A(n_538),
.Y(n_649)
);

NOR2xp33_ASAP7_75t_L g650 ( 
.A(n_487),
.B(n_274),
.Y(n_650)
);

NOR2x1p5_ASAP7_75t_L g651 ( 
.A(n_573),
.B(n_459),
.Y(n_651)
);

AO22x2_ASAP7_75t_L g652 ( 
.A1(n_593),
.A2(n_461),
.B1(n_525),
.B2(n_387),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_588),
.B(n_467),
.Y(n_653)
);

HB1xp67_ASAP7_75t_L g654 ( 
.A(n_609),
.Y(n_654)
);

BUFx3_ASAP7_75t_L g655 ( 
.A(n_579),
.Y(n_655)
);

INVx4_ASAP7_75t_L g656 ( 
.A(n_586),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_586),
.Y(n_657)
);

INVx3_ASAP7_75t_L g658 ( 
.A(n_576),
.Y(n_658)
);

NAND2xp5_ASAP7_75t_SL g659 ( 
.A(n_562),
.B(n_337),
.Y(n_659)
);

BUFx3_ASAP7_75t_L g660 ( 
.A(n_579),
.Y(n_660)
);

INVx2_ASAP7_75t_SL g661 ( 
.A(n_579),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_588),
.B(n_467),
.Y(n_663)
);

INVx8_ASAP7_75t_L g664 ( 
.A(n_567),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_576),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_585),
.Y(n_666)
);

BUFx2_ASAP7_75t_L g667 ( 
.A(n_564),
.Y(n_667)
);

NAND3xp33_ASAP7_75t_L g668 ( 
.A(n_650),
.B(n_480),
.C(n_478),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_585),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_585),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_559),
.Y(n_671)
);

BUFx6f_ASAP7_75t_SL g672 ( 
.A(n_588),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_585),
.Y(n_673)
);

INVx4_ASAP7_75t_L g674 ( 
.A(n_586),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_589),
.Y(n_675)
);

AOI22xp5_ASAP7_75t_L g676 ( 
.A1(n_604),
.A2(n_488),
.B1(n_493),
.B2(n_492),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx3_ASAP7_75t_L g678 ( 
.A(n_576),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_646),
.Y(n_679)
);

NOR2xp33_ASAP7_75t_L g680 ( 
.A(n_593),
.B(n_507),
.Y(n_680)
);

AND2x4_ASAP7_75t_L g681 ( 
.A(n_607),
.B(n_535),
.Y(n_681)
);

INVx1_ASAP7_75t_SL g682 ( 
.A(n_622),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_646),
.Y(n_683)
);

AND3x2_ASAP7_75t_L g684 ( 
.A(n_564),
.B(n_347),
.C(n_337),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_589),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_589),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_559),
.Y(n_687)
);

BUFx10_ASAP7_75t_L g688 ( 
.A(n_650),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_559),
.Y(n_689)
);

OR2x6_ASAP7_75t_L g690 ( 
.A(n_645),
.B(n_525),
.Y(n_690)
);

OAI22xp33_ASAP7_75t_L g691 ( 
.A1(n_575),
.A2(n_437),
.B1(n_279),
.B2(n_474),
.Y(n_691)
);

INVx3_ASAP7_75t_L g692 ( 
.A(n_576),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_582),
.Y(n_693)
);

HB1xp67_ASAP7_75t_L g694 ( 
.A(n_609),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_588),
.B(n_478),
.Y(n_695)
);

AOI22xp5_ASAP7_75t_L g696 ( 
.A1(n_604),
.A2(n_562),
.B1(n_648),
.B2(n_645),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_579),
.Y(n_697)
);

NAND3xp33_ASAP7_75t_L g698 ( 
.A(n_635),
.B(n_647),
.C(n_643),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_589),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_562),
.B(n_480),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_582),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_SL g702 ( 
.A(n_562),
.B(n_347),
.Y(n_702)
);

INVx3_ASAP7_75t_L g703 ( 
.A(n_576),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_622),
.Y(n_704)
);

INVx3_ASAP7_75t_L g705 ( 
.A(n_576),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_582),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_577),
.B(n_511),
.Y(n_707)
);

AND2x4_ASAP7_75t_SL g708 ( 
.A(n_629),
.B(n_452),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_595),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_595),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_582),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_577),
.B(n_365),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_627),
.B(n_365),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_591),
.B(n_518),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_583),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_SL g716 ( 
.A(n_591),
.B(n_602),
.Y(n_716)
);

AND2x2_ASAP7_75t_L g717 ( 
.A(n_607),
.B(n_495),
.Y(n_717)
);

OR2x6_ASAP7_75t_L g718 ( 
.A(n_648),
.B(n_635),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_583),
.Y(n_719)
);

INVx3_ASAP7_75t_L g720 ( 
.A(n_576),
.Y(n_720)
);

INVx2_ASAP7_75t_SL g721 ( 
.A(n_579),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_595),
.Y(n_722)
);

AOI22xp5_ASAP7_75t_L g723 ( 
.A1(n_575),
.A2(n_520),
.B1(n_528),
.B2(n_521),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_602),
.B(n_553),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_583),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_L g726 ( 
.A(n_573),
.B(n_263),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_583),
.Y(n_727)
);

INVx1_ASAP7_75t_SL g728 ( 
.A(n_564),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_595),
.Y(n_729)
);

BUFx6f_ASAP7_75t_L g730 ( 
.A(n_597),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_597),
.Y(n_731)
);

OAI22xp33_ASAP7_75t_SL g732 ( 
.A1(n_579),
.A2(n_398),
.B1(n_527),
.B2(n_498),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_630),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_630),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_616),
.B(n_486),
.Y(n_735)
);

BUFx10_ASAP7_75t_L g736 ( 
.A(n_629),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_587),
.B(n_263),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_576),
.Y(n_738)
);

NAND3xp33_ASAP7_75t_L g739 ( 
.A(n_643),
.B(n_491),
.C(n_486),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_L g740 ( 
.A(n_584),
.B(n_554),
.Y(n_740)
);

INVx2_ASAP7_75t_SL g741 ( 
.A(n_607),
.Y(n_741)
);

AND2x6_ASAP7_75t_L g742 ( 
.A(n_627),
.B(n_263),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_SL g743 ( 
.A(n_587),
.B(n_263),
.Y(n_743)
);

OAI22xp5_ASAP7_75t_L g744 ( 
.A1(n_584),
.A2(n_649),
.B1(n_482),
.B2(n_503),
.Y(n_744)
);

INVx2_ASAP7_75t_L g745 ( 
.A(n_630),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_570),
.B(n_497),
.Y(n_746)
);

BUFx4f_ASAP7_75t_L g747 ( 
.A(n_597),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_567),
.B(n_627),
.Y(n_748)
);

BUFx10_ASAP7_75t_L g749 ( 
.A(n_567),
.Y(n_749)
);

NOR2xp33_ASAP7_75t_L g750 ( 
.A(n_649),
.B(n_491),
.Y(n_750)
);

BUFx10_ASAP7_75t_L g751 ( 
.A(n_567),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_616),
.B(n_570),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_SL g753 ( 
.A(n_587),
.B(n_263),
.Y(n_753)
);

NAND2xp33_ASAP7_75t_SL g754 ( 
.A(n_647),
.B(n_334),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_570),
.B(n_499),
.Y(n_755)
);

AND2x6_ASAP7_75t_L g756 ( 
.A(n_587),
.B(n_224),
.Y(n_756)
);

INVx3_ASAP7_75t_L g757 ( 
.A(n_578),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_634),
.B(n_503),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_606),
.B(n_490),
.Y(n_759)
);

AND3x1_ASAP7_75t_L g760 ( 
.A(n_606),
.B(n_448),
.C(n_312),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_597),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_586),
.B(n_506),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_630),
.Y(n_763)
);

AOI22xp5_ASAP7_75t_L g764 ( 
.A1(n_567),
.A2(n_515),
.B1(n_526),
.B2(n_506),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_606),
.B(n_567),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_597),
.A2(n_516),
.B1(n_541),
.B2(n_502),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_632),
.Y(n_767)
);

OAI22xp33_ASAP7_75t_SL g768 ( 
.A1(n_634),
.A2(n_526),
.B1(n_534),
.B2(n_515),
.Y(n_768)
);

OR2x2_ASAP7_75t_L g769 ( 
.A(n_631),
.B(n_513),
.Y(n_769)
);

NAND2x1p5_ASAP7_75t_L g770 ( 
.A(n_587),
.B(n_355),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_632),
.Y(n_771)
);

OAI22xp33_ASAP7_75t_L g772 ( 
.A1(n_639),
.A2(n_356),
.B1(n_358),
.B2(n_352),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_631),
.B(n_534),
.Y(n_773)
);

OR2x6_ASAP7_75t_L g774 ( 
.A(n_587),
.B(n_326),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_615),
.B(n_537),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_586),
.B(n_537),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_586),
.B(n_543),
.Y(n_777)
);

INVx3_ASAP7_75t_L g778 ( 
.A(n_578),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_586),
.B(n_543),
.Y(n_779)
);

AND3x2_ASAP7_75t_L g780 ( 
.A(n_615),
.B(n_516),
.C(n_502),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_561),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_639),
.B(n_490),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_615),
.B(n_545),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_561),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_578),
.Y(n_785)
);

INVxp67_ASAP7_75t_SL g786 ( 
.A(n_578),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_642),
.B(n_545),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_563),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_632),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_632),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_563),
.Y(n_791)
);

INVx3_ASAP7_75t_L g792 ( 
.A(n_578),
.Y(n_792)
);

INVx2_ASAP7_75t_L g793 ( 
.A(n_633),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_565),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_586),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_594),
.B(n_550),
.Y(n_796)
);

NAND2xp33_ASAP7_75t_L g797 ( 
.A(n_594),
.B(n_246),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_565),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_633),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_633),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_633),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_566),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_568),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_578),
.Y(n_804)
);

INVx1_ASAP7_75t_SL g805 ( 
.A(n_637),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_598),
.Y(n_806)
);

INVx4_ASAP7_75t_L g807 ( 
.A(n_594),
.Y(n_807)
);

O2A1O1Ixp33_ASAP7_75t_L g808 ( 
.A1(n_659),
.A2(n_300),
.B(n_321),
.C(n_319),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_659),
.A2(n_371),
.B1(n_377),
.B2(n_360),
.Y(n_809)
);

AND2x2_ASAP7_75t_L g810 ( 
.A(n_759),
.B(n_550),
.Y(n_810)
);

BUFx6f_ASAP7_75t_SL g811 ( 
.A(n_736),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_716),
.B(n_594),
.Y(n_812)
);

INVx3_ASAP7_75t_L g813 ( 
.A(n_748),
.Y(n_813)
);

INVx3_ASAP7_75t_L g814 ( 
.A(n_748),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_716),
.B(n_594),
.Y(n_815)
);

NOR2x1p5_ASAP7_75t_L g816 ( 
.A(n_769),
.B(n_735),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_752),
.B(n_594),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_SL g818 ( 
.A(n_662),
.B(n_247),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_750),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_741),
.B(n_594),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_696),
.A2(n_454),
.B1(n_462),
.B2(n_457),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_741),
.B(n_594),
.Y(n_822)
);

OR2x6_ASAP7_75t_L g823 ( 
.A(n_667),
.B(n_541),
.Y(n_823)
);

INVx8_ASAP7_75t_L g824 ( 
.A(n_672),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_698),
.B(n_578),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_805),
.B(n_578),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_695),
.B(n_552),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_759),
.B(n_552),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_688),
.B(n_469),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_700),
.B(n_560),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_653),
.B(n_245),
.Y(n_831)
);

AOI22xp33_ASAP7_75t_L g832 ( 
.A1(n_702),
.A2(n_378),
.B1(n_414),
.B2(n_406),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_747),
.B(n_560),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_748),
.B(n_615),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_758),
.B(n_615),
.Y(n_835)
);

NOR2xp67_ASAP7_75t_L g836 ( 
.A(n_668),
.B(n_642),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_671),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_765),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_713),
.B(n_338),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_677),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_765),
.Y(n_841)
);

BUFx3_ASAP7_75t_L g842 ( 
.A(n_681),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_766),
.B(n_560),
.C(n_397),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_SL g844 ( 
.A(n_747),
.B(n_662),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_740),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_762),
.B(n_615),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_672),
.A2(n_471),
.B1(n_481),
.B2(n_285),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_687),
.Y(n_848)
);

INVx3_ASAP7_75t_L g849 ( 
.A(n_749),
.Y(n_849)
);

AOI22xp5_ASAP7_75t_L g850 ( 
.A1(n_672),
.A2(n_341),
.B1(n_342),
.B2(n_340),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_776),
.B(n_777),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_SL g852 ( 
.A(n_747),
.B(n_560),
.Y(n_852)
);

AND2x6_ASAP7_75t_SL g853 ( 
.A(n_680),
.B(n_416),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_662),
.B(n_730),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_688),
.B(n_238),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_717),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_718),
.A2(n_345),
.B1(n_348),
.B2(n_344),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_654),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_688),
.B(n_782),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_779),
.B(n_620),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_702),
.A2(n_419),
.B1(n_439),
.B2(n_417),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_796),
.B(n_620),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_717),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_662),
.B(n_620),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_689),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_662),
.B(n_620),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_730),
.B(n_731),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_730),
.B(n_620),
.Y(n_868)
);

OAI22xp5_ASAP7_75t_L g869 ( 
.A1(n_663),
.A2(n_268),
.B1(n_281),
.B2(n_257),
.Y(n_869)
);

NOR2xp67_ASAP7_75t_L g870 ( 
.A(n_676),
.B(n_640),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_781),
.Y(n_871)
);

NOR2xp33_ASAP7_75t_L g872 ( 
.A(n_707),
.B(n_248),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_718),
.A2(n_353),
.B1(n_386),
.B2(n_351),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_SL g874 ( 
.A(n_730),
.B(n_560),
.Y(n_874)
);

CKINVDCx5p33_ASAP7_75t_R g875 ( 
.A(n_679),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_784),
.Y(n_876)
);

NAND2xp33_ASAP7_75t_L g877 ( 
.A(n_713),
.B(n_394),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_730),
.B(n_620),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_788),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_693),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_714),
.B(n_560),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_724),
.B(n_628),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_749),
.B(n_628),
.Y(n_883)
);

AOI22xp33_ASAP7_75t_L g884 ( 
.A1(n_652),
.A2(n_761),
.B1(n_712),
.B2(n_690),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_791),
.B(n_624),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_794),
.B(n_624),
.Y(n_886)
);

NAND2xp5_ASAP7_75t_SL g887 ( 
.A(n_749),
.B(n_628),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_798),
.B(n_624),
.Y(n_888)
);

AOI22xp5_ASAP7_75t_L g889 ( 
.A1(n_718),
.A2(n_783),
.B1(n_775),
.B2(n_754),
.Y(n_889)
);

AOI22xp5_ASAP7_75t_L g890 ( 
.A1(n_718),
.A2(n_783),
.B1(n_775),
.B2(n_754),
.Y(n_890)
);

A2O1A1Ixp33_ASAP7_75t_L g891 ( 
.A1(n_712),
.A2(n_624),
.B(n_542),
.C(n_556),
.Y(n_891)
);

OAI22xp5_ASAP7_75t_L g892 ( 
.A1(n_690),
.A2(n_362),
.B1(n_388),
.B2(n_395),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_802),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_787),
.A2(n_624),
.B(n_536),
.C(n_637),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_803),
.B(n_624),
.Y(n_895)
);

BUFx3_ASAP7_75t_L g896 ( 
.A(n_681),
.Y(n_896)
);

BUFx6f_ASAP7_75t_L g897 ( 
.A(n_664),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_681),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_751),
.B(n_770),
.Y(n_899)
);

INVx2_ASAP7_75t_L g900 ( 
.A(n_701),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_769),
.B(n_248),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_786),
.B(n_637),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_706),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_773),
.B(n_637),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_770),
.B(n_637),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_713),
.B(n_637),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_736),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_746),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_664),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_751),
.B(n_628),
.Y(n_910)
);

NAND3xp33_ASAP7_75t_L g911 ( 
.A(n_739),
.B(n_409),
.C(n_359),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_713),
.B(n_571),
.Y(n_912)
);

NOR2xp33_ASAP7_75t_L g913 ( 
.A(n_690),
.B(n_250),
.Y(n_913)
);

NAND2xp33_ASAP7_75t_L g914 ( 
.A(n_713),
.B(n_407),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_713),
.B(n_571),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_746),
.B(n_571),
.Y(n_916)
);

A2O1A1Ixp33_ASAP7_75t_L g917 ( 
.A1(n_755),
.A2(n_782),
.B(n_764),
.C(n_726),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_736),
.Y(n_918)
);

OAI22xp33_ASAP7_75t_L g919 ( 
.A1(n_690),
.A2(n_375),
.B1(n_400),
.B2(n_260),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_755),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_694),
.Y(n_921)
);

INVx3_ASAP7_75t_L g922 ( 
.A(n_751),
.Y(n_922)
);

AO221x1_ASAP7_75t_L g923 ( 
.A1(n_652),
.A2(n_691),
.B1(n_772),
.B2(n_744),
.C(n_291),
.Y(n_923)
);

AND2x6_ASAP7_75t_L g924 ( 
.A(n_658),
.B(n_293),
.Y(n_924)
);

NAND3xp33_ASAP7_75t_L g925 ( 
.A(n_760),
.B(n_411),
.C(n_410),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_706),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_733),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_664),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_733),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_768),
.B(n_628),
.Y(n_930)
);

INVxp67_ASAP7_75t_L g931 ( 
.A(n_728),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_658),
.B(n_571),
.Y(n_932)
);

AOI22xp33_ASAP7_75t_L g933 ( 
.A1(n_652),
.A2(n_331),
.B1(n_297),
.B2(n_438),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_734),
.Y(n_934)
);

BUFx5_ASAP7_75t_L g935 ( 
.A(n_756),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_732),
.B(n_628),
.Y(n_936)
);

INVx5_ASAP7_75t_L g937 ( 
.A(n_742),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_658),
.B(n_571),
.Y(n_938)
);

NOR3xp33_ASAP7_75t_L g939 ( 
.A(n_682),
.B(n_704),
.C(n_723),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_734),
.Y(n_940)
);

NOR2xp33_ASAP7_75t_L g941 ( 
.A(n_780),
.B(n_250),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_665),
.B(n_572),
.Y(n_942)
);

OAI22xp5_ASAP7_75t_SL g943 ( 
.A1(n_679),
.A2(n_249),
.B1(n_242),
.B2(n_305),
.Y(n_943)
);

INVxp67_ASAP7_75t_L g944 ( 
.A(n_651),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_745),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_665),
.B(n_572),
.Y(n_946)
);

AOI22xp5_ASAP7_75t_L g947 ( 
.A1(n_652),
.A2(n_425),
.B1(n_408),
.B2(n_418),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_785),
.B(n_628),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_664),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_SL g950 ( 
.A(n_785),
.B(n_628),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_665),
.B(n_572),
.Y(n_951)
);

INVx2_ASAP7_75t_L g952 ( 
.A(n_711),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_711),
.Y(n_953)
);

NOR2xp33_ASAP7_75t_L g954 ( 
.A(n_684),
.B(n_251),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_745),
.Y(n_955)
);

BUFx2_ASAP7_75t_L g956 ( 
.A(n_683),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_763),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_678),
.B(n_572),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_785),
.B(n_307),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_678),
.B(n_572),
.Y(n_960)
);

AND2x2_ASAP7_75t_L g961 ( 
.A(n_708),
.B(n_287),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_785),
.B(n_311),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_774),
.B(n_709),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_L g964 ( 
.A(n_774),
.B(n_710),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_678),
.B(n_581),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_763),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_767),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_692),
.B(n_581),
.Y(n_968)
);

BUFx3_ASAP7_75t_L g969 ( 
.A(n_655),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_SL g970 ( 
.A(n_785),
.B(n_346),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_774),
.B(n_251),
.Y(n_971)
);

INVx8_ASAP7_75t_L g972 ( 
.A(n_774),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_692),
.B(n_581),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_872),
.B(n_692),
.Y(n_974)
);

INVx1_ASAP7_75t_SL g975 ( 
.A(n_858),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_872),
.B(n_703),
.Y(n_976)
);

AOI22xp5_ASAP7_75t_L g977 ( 
.A1(n_827),
.A2(n_756),
.B1(n_721),
.B2(n_661),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_837),
.Y(n_978)
);

AOI21x1_ASAP7_75t_L g979 ( 
.A1(n_818),
.A2(n_882),
.B(n_883),
.Y(n_979)
);

AND2x4_ASAP7_75t_L g980 ( 
.A(n_842),
.B(n_655),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_827),
.B(n_831),
.Y(n_981)
);

OAI22xp5_ASAP7_75t_L g982 ( 
.A1(n_889),
.A2(n_661),
.B1(n_721),
.B2(n_697),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_864),
.A2(n_729),
.B(n_722),
.Y(n_983)
);

HB1xp67_ASAP7_75t_L g984 ( 
.A(n_931),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_866),
.A2(n_697),
.B(n_660),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_L g986 ( 
.A1(n_890),
.A2(n_756),
.B1(n_742),
.B2(n_660),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_868),
.A2(n_743),
.B(n_737),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_831),
.B(n_835),
.Y(n_988)
);

O2A1O1Ixp5_ASAP7_75t_L g989 ( 
.A1(n_930),
.A2(n_743),
.B(n_753),
.C(n_737),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_878),
.A2(n_753),
.B(n_657),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_867),
.B(n_703),
.Y(n_991)
);

OAI22xp5_ASAP7_75t_L g992 ( 
.A1(n_884),
.A2(n_705),
.B1(n_720),
.B2(n_703),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_904),
.B(n_705),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_L g994 ( 
.A(n_819),
.B(n_683),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_838),
.B(n_705),
.Y(n_995)
);

NOR2xp67_ASAP7_75t_L g996 ( 
.A(n_845),
.B(n_666),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_841),
.B(n_720),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_898),
.Y(n_998)
);

O2A1O1Ixp33_ASAP7_75t_L g999 ( 
.A1(n_917),
.A2(n_726),
.B(n_797),
.C(n_670),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_817),
.B(n_720),
.Y(n_1000)
);

NOR2x2_ASAP7_75t_L g1001 ( 
.A(n_823),
.B(n_708),
.Y(n_1001)
);

NAND2x1p5_ASAP7_75t_L g1002 ( 
.A(n_928),
.B(n_738),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_851),
.B(n_738),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_859),
.B(n_256),
.Y(n_1004)
);

INVx1_ASAP7_75t_SL g1005 ( 
.A(n_921),
.Y(n_1005)
);

OAI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_812),
.A2(n_673),
.B(n_669),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_SL g1007 ( 
.A(n_813),
.B(n_256),
.Y(n_1007)
);

AND2x2_ASAP7_75t_SL g1008 ( 
.A(n_956),
.B(n_829),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_916),
.B(n_738),
.Y(n_1009)
);

NOR2xp67_ASAP7_75t_L g1010 ( 
.A(n_907),
.B(n_675),
.Y(n_1010)
);

AOI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_902),
.A2(n_657),
.B(n_656),
.Y(n_1011)
);

NOR2xp33_ASAP7_75t_L g1012 ( 
.A(n_901),
.B(n_458),
.Y(n_1012)
);

AOI21x1_ASAP7_75t_L g1013 ( 
.A1(n_882),
.A2(n_686),
.B(n_685),
.Y(n_1013)
);

INVx1_ASAP7_75t_L g1014 ( 
.A(n_871),
.Y(n_1014)
);

NOR3xp33_ASAP7_75t_L g1015 ( 
.A(n_919),
.B(n_901),
.C(n_939),
.Y(n_1015)
);

BUFx6f_ASAP7_75t_L g1016 ( 
.A(n_969),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_810),
.B(n_458),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_846),
.A2(n_657),
.B(n_656),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_876),
.B(n_757),
.Y(n_1019)
);

INVx2_ASAP7_75t_L g1020 ( 
.A(n_840),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_879),
.Y(n_1021)
);

AOI22xp5_ASAP7_75t_L g1022 ( 
.A1(n_813),
.A2(n_756),
.B1(n_742),
.B2(n_792),
.Y(n_1022)
);

AOI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_860),
.A2(n_674),
.B(n_656),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_854),
.A2(n_795),
.B(n_674),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_854),
.A2(n_795),
.B(n_674),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_862),
.A2(n_807),
.B(n_795),
.Y(n_1026)
);

AND2x2_ASAP7_75t_L g1027 ( 
.A(n_828),
.B(n_287),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_893),
.B(n_757),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_826),
.A2(n_807),
.B(n_778),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_834),
.Y(n_1030)
);

HB1xp67_ASAP7_75t_L g1031 ( 
.A(n_823),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_814),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_844),
.A2(n_807),
.B(n_778),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_844),
.A2(n_905),
.B(n_906),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_884),
.A2(n_757),
.B1(n_804),
.B2(n_778),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_928),
.B(n_792),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_883),
.A2(n_804),
.B(n_792),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_887),
.A2(n_804),
.B(n_797),
.Y(n_1038)
);

O2A1O1Ixp5_ASAP7_75t_L g1039 ( 
.A1(n_930),
.A2(n_699),
.B(n_806),
.C(n_800),
.Y(n_1039)
);

O2A1O1Ixp33_ASAP7_75t_SL g1040 ( 
.A1(n_894),
.A2(n_349),
.B(n_373),
.C(n_396),
.Y(n_1040)
);

BUFx3_ASAP7_75t_L g1041 ( 
.A(n_875),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_917),
.B(n_715),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_887),
.A2(n_719),
.B(n_715),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_910),
.A2(n_725),
.B(n_719),
.Y(n_1044)
);

NAND2x1p5_ASAP7_75t_L g1045 ( 
.A(n_949),
.B(n_725),
.Y(n_1045)
);

NOR2xp33_ASAP7_75t_L g1046 ( 
.A(n_855),
.B(n_473),
.Y(n_1046)
);

OAI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_815),
.A2(n_727),
.B(n_806),
.Y(n_1047)
);

INVxp67_ASAP7_75t_L g1048 ( 
.A(n_961),
.Y(n_1048)
);

INVxp67_ASAP7_75t_L g1049 ( 
.A(n_823),
.Y(n_1049)
);

A2O1A1Ixp33_ASAP7_75t_L g1050 ( 
.A1(n_913),
.A2(n_432),
.B(n_424),
.C(n_415),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_814),
.B(n_727),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_885),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_910),
.A2(n_581),
.B(n_767),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_825),
.A2(n_581),
.B(n_771),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_820),
.A2(n_789),
.B(n_771),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_886),
.Y(n_1056)
);

NAND2xp33_ASAP7_75t_SL g1057 ( 
.A(n_816),
.B(n_473),
.Y(n_1057)
);

BUFx12f_ASAP7_75t_L g1058 ( 
.A(n_918),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_856),
.B(n_756),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_822),
.A2(n_790),
.B(n_789),
.Y(n_1060)
);

NOR3xp33_ASAP7_75t_L g1061 ( 
.A(n_919),
.B(n_261),
.C(n_258),
.Y(n_1061)
);

O2A1O1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_908),
.A2(n_404),
.B(n_612),
.C(n_568),
.Y(n_1062)
);

AOI21xp33_ASAP7_75t_L g1063 ( 
.A1(n_913),
.A2(n_413),
.B(n_412),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_863),
.B(n_756),
.Y(n_1064)
);

OAI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_933),
.A2(n_430),
.B1(n_261),
.B2(n_262),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_920),
.B(n_742),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_888),
.Y(n_1067)
);

INVx8_ASAP7_75t_L g1068 ( 
.A(n_972),
.Y(n_1068)
);

OAI21xp33_ASAP7_75t_L g1069 ( 
.A1(n_809),
.A2(n_249),
.B(n_242),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_L g1070 ( 
.A(n_809),
.B(n_742),
.Y(n_1070)
);

BUFx2_ASAP7_75t_L g1071 ( 
.A(n_896),
.Y(n_1071)
);

BUFx6f_ASAP7_75t_L g1072 ( 
.A(n_969),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_912),
.A2(n_915),
.B(n_899),
.Y(n_1073)
);

NAND2xp5_ASAP7_75t_L g1074 ( 
.A(n_832),
.B(n_742),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_869),
.A2(n_580),
.B(n_612),
.C(n_601),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_899),
.A2(n_793),
.B(n_790),
.Y(n_1076)
);

BUFx4f_ASAP7_75t_L g1077 ( 
.A(n_824),
.Y(n_1077)
);

O2A1O1Ixp33_ASAP7_75t_L g1078 ( 
.A1(n_891),
.A2(n_892),
.B(n_881),
.C(n_894),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_832),
.B(n_793),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_895),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_861),
.B(n_799),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_861),
.B(n_799),
.Y(n_1082)
);

NAND3xp33_ASAP7_75t_SL g1083 ( 
.A(n_821),
.B(n_260),
.C(n_255),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_836),
.B(n_800),
.Y(n_1084)
);

A2O1A1Ixp33_ASAP7_75t_L g1085 ( 
.A1(n_971),
.A2(n_640),
.B(n_801),
.C(n_433),
.Y(n_1085)
);

INVxp67_ASAP7_75t_L g1086 ( 
.A(n_954),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_932),
.A2(n_801),
.B(n_599),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_SL g1088 ( 
.A(n_870),
.B(n_258),
.Y(n_1088)
);

NAND2xp5_ASAP7_75t_L g1089 ( 
.A(n_849),
.B(n_640),
.Y(n_1089)
);

OAI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_933),
.A2(n_428),
.B1(n_262),
.B2(n_435),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_938),
.A2(n_599),
.B(n_598),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_942),
.A2(n_599),
.B(n_598),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_L g1093 ( 
.A(n_849),
.B(n_640),
.Y(n_1093)
);

BUFx2_ASAP7_75t_L g1094 ( 
.A(n_944),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_SL g1095 ( 
.A(n_897),
.B(n_267),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_946),
.A2(n_599),
.B(n_598),
.Y(n_1096)
);

INVx5_ASAP7_75t_L g1097 ( 
.A(n_897),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_L g1098 ( 
.A(n_911),
.B(n_473),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_824),
.Y(n_1099)
);

OAI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_881),
.A2(n_428),
.B1(n_267),
.B2(n_435),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_927),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_922),
.B(n_640),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_891),
.A2(n_936),
.B(n_808),
.C(n_830),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_951),
.A2(n_608),
.B(n_605),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_922),
.B(n_569),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_958),
.A2(n_608),
.B(n_605),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_SL g1107 ( 
.A(n_897),
.B(n_363),
.Y(n_1107)
);

OAI22xp5_ASAP7_75t_L g1108 ( 
.A1(n_830),
.A2(n_363),
.B1(n_366),
.B2(n_376),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_963),
.B(n_569),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_847),
.B(n_366),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_963),
.B(n_574),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_960),
.A2(n_608),
.B(n_605),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_964),
.B(n_929),
.Y(n_1113)
);

NOR3xp33_ASAP7_75t_L g1114 ( 
.A(n_941),
.B(n_381),
.C(n_376),
.Y(n_1114)
);

AND2x4_ASAP7_75t_L g1115 ( 
.A(n_949),
.B(n_557),
.Y(n_1115)
);

OAI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_964),
.A2(n_580),
.B(n_574),
.Y(n_1116)
);

AND2x4_ASAP7_75t_L g1117 ( 
.A(n_897),
.B(n_557),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_SL g1118 ( 
.A(n_909),
.B(n_381),
.Y(n_1118)
);

NOR2xp33_ASAP7_75t_L g1119 ( 
.A(n_943),
.B(n_382),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_934),
.B(n_590),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_909),
.B(n_382),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_909),
.B(n_383),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_848),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_824),
.Y(n_1124)
);

O2A1O1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_936),
.A2(n_596),
.B(n_592),
.C(n_625),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_940),
.B(n_590),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_972),
.Y(n_1127)
);

OAI21xp33_ASAP7_75t_L g1128 ( 
.A1(n_925),
.A2(n_427),
.B(n_269),
.Y(n_1128)
);

INVx4_ASAP7_75t_L g1129 ( 
.A(n_909),
.Y(n_1129)
);

INVx2_ASAP7_75t_L g1130 ( 
.A(n_865),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_965),
.A2(n_617),
.B(n_605),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_941),
.B(n_287),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_968),
.A2(n_614),
.B(n_608),
.Y(n_1133)
);

AND2x2_ASAP7_75t_SL g1134 ( 
.A(n_971),
.B(n_343),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_973),
.A2(n_614),
.B(n_621),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_948),
.A2(n_614),
.B(n_621),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_839),
.A2(n_914),
.B(n_877),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_945),
.B(n_592),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_948),
.A2(n_617),
.B(n_614),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_955),
.B(n_596),
.Y(n_1140)
);

BUFx2_ASAP7_75t_L g1141 ( 
.A(n_853),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_950),
.A2(n_617),
.B(n_621),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_950),
.A2(n_621),
.B(n_617),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_L g1144 ( 
.A1(n_959),
.A2(n_601),
.B(n_618),
.C(n_625),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_957),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_966),
.B(n_618),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_967),
.B(n_600),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_937),
.A2(n_623),
.B(n_626),
.Y(n_1148)
);

O2A1O1Ixp33_ASAP7_75t_SL g1149 ( 
.A1(n_959),
.A2(n_636),
.B(n_600),
.C(n_619),
.Y(n_1149)
);

OAI22xp5_ASAP7_75t_L g1150 ( 
.A1(n_874),
.A2(n_431),
.B1(n_383),
.B2(n_390),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_923),
.B(n_600),
.Y(n_1151)
);

CKINVDCx8_ASAP7_75t_R g1152 ( 
.A(n_972),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_937),
.A2(n_623),
.B(n_626),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_880),
.Y(n_1154)
);

OR2x6_ASAP7_75t_L g1155 ( 
.A(n_843),
.B(n_636),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_937),
.A2(n_874),
.B(n_852),
.Y(n_1156)
);

AOI22xp5_ASAP7_75t_L g1157 ( 
.A1(n_947),
.A2(n_873),
.B1(n_857),
.B2(n_850),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_937),
.B(n_390),
.Y(n_1158)
);

OAI21xp33_ASAP7_75t_L g1159 ( 
.A1(n_954),
.A2(n_255),
.B(n_269),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_900),
.B(n_600),
.Y(n_1160)
);

HB1xp67_ASAP7_75t_L g1161 ( 
.A(n_975),
.Y(n_1161)
);

O2A1O1Ixp33_ASAP7_75t_L g1162 ( 
.A1(n_981),
.A2(n_852),
.B(n_833),
.C(n_970),
.Y(n_1162)
);

AOI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1137),
.A2(n_833),
.B(n_962),
.Y(n_1163)
);

NOR2xp33_ASAP7_75t_L g1164 ( 
.A(n_994),
.B(n_811),
.Y(n_1164)
);

OAI21xp5_ASAP7_75t_L g1165 ( 
.A1(n_988),
.A2(n_953),
.B(n_952),
.Y(n_1165)
);

NAND2xp5_ASAP7_75t_L g1166 ( 
.A(n_1030),
.B(n_903),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_1041),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_1129),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1052),
.B(n_926),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_L g1170 ( 
.A(n_1056),
.B(n_924),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1067),
.B(n_924),
.Y(n_1171)
);

BUFx2_ASAP7_75t_SL g1172 ( 
.A(n_1005),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1154),
.Y(n_1173)
);

AOI22xp33_ASAP7_75t_L g1174 ( 
.A1(n_1015),
.A2(n_924),
.B1(n_962),
.B2(n_970),
.Y(n_1174)
);

A2O1A1Ixp33_ASAP7_75t_SL g1175 ( 
.A1(n_1012),
.A2(n_619),
.B(n_611),
.C(n_600),
.Y(n_1175)
);

HB1xp67_ASAP7_75t_L g1176 ( 
.A(n_984),
.Y(n_1176)
);

AOI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1034),
.A2(n_935),
.B(n_603),
.Y(n_1177)
);

INVx3_ASAP7_75t_L g1178 ( 
.A(n_1129),
.Y(n_1178)
);

OR2x2_ASAP7_75t_SL g1179 ( 
.A(n_1083),
.B(n_811),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1003),
.A2(n_935),
.B(n_603),
.Y(n_1180)
);

BUFx3_ASAP7_75t_L g1181 ( 
.A(n_1058),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_1094),
.Y(n_1182)
);

NOR2xp33_ASAP7_75t_R g1183 ( 
.A(n_1077),
.B(n_924),
.Y(n_1183)
);

AO32x1_ASAP7_75t_L g1184 ( 
.A1(n_992),
.A2(n_641),
.A3(n_638),
.B1(n_626),
.B2(n_623),
.Y(n_1184)
);

BUFx6f_ASAP7_75t_L g1185 ( 
.A(n_1016),
.Y(n_1185)
);

AOI21x1_ASAP7_75t_L g1186 ( 
.A1(n_979),
.A2(n_976),
.B(n_974),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1080),
.B(n_924),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_L g1188 ( 
.A(n_996),
.B(n_935),
.Y(n_1188)
);

AOI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1013),
.A2(n_623),
.B(n_626),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1014),
.B(n_935),
.Y(n_1190)
);

BUFx6f_ASAP7_75t_L g1191 ( 
.A(n_1016),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1031),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_SL g1193 ( 
.A(n_1134),
.B(n_1016),
.Y(n_1193)
);

INVx4_ASAP7_75t_L g1194 ( 
.A(n_1097),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1086),
.B(n_420),
.Y(n_1195)
);

NOR2xp67_ASAP7_75t_SL g1196 ( 
.A(n_1097),
.B(n_391),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_L g1197 ( 
.A1(n_1061),
.A2(n_935),
.B1(n_343),
.B2(n_385),
.Y(n_1197)
);

AND3x4_ASAP7_75t_L g1198 ( 
.A(n_1114),
.B(n_402),
.C(n_384),
.Y(n_1198)
);

NAND2xp5_ASAP7_75t_L g1199 ( 
.A(n_1021),
.B(n_935),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1072),
.B(n_391),
.Y(n_1200)
);

NOR2xp67_ASAP7_75t_L g1201 ( 
.A(n_1048),
.B(n_421),
.Y(n_1201)
);

INVxp67_ASAP7_75t_L g1202 ( 
.A(n_1027),
.Y(n_1202)
);

OAI22x1_ASAP7_75t_L g1203 ( 
.A1(n_1157),
.A2(n_305),
.B1(n_427),
.B2(n_272),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1072),
.B(n_392),
.Y(n_1204)
);

NOR3xp33_ASAP7_75t_L g1205 ( 
.A(n_1110),
.B(n_422),
.C(n_423),
.Y(n_1205)
);

NOR2xp33_ASAP7_75t_SL g1206 ( 
.A(n_1152),
.B(n_385),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_993),
.A2(n_613),
.B(n_619),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_983),
.A2(n_613),
.B(n_619),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_998),
.Y(n_1209)
);

CKINVDCx5p33_ASAP7_75t_R g1210 ( 
.A(n_1099),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1004),
.B(n_270),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_SL g1212 ( 
.A(n_1072),
.B(n_392),
.Y(n_1212)
);

OA22x2_ASAP7_75t_L g1213 ( 
.A1(n_1159),
.A2(n_1049),
.B1(n_1132),
.B2(n_1069),
.Y(n_1213)
);

AOI22xp33_ASAP7_75t_L g1214 ( 
.A1(n_1063),
.A2(n_403),
.B1(n_385),
.B2(n_393),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1008),
.B(n_393),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1026),
.A2(n_613),
.B(n_619),
.Y(n_1216)
);

AOI21x1_ASAP7_75t_L g1217 ( 
.A1(n_1073),
.A2(n_641),
.B(n_638),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1026),
.A2(n_611),
.B(n_613),
.Y(n_1218)
);

BUFx2_ASAP7_75t_L g1219 ( 
.A(n_1071),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_1000),
.A2(n_611),
.B(n_613),
.Y(n_1220)
);

AND2x2_ASAP7_75t_SL g1221 ( 
.A(n_1077),
.B(n_403),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1101),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_978),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1124),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1097),
.B(n_429),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_1113),
.B(n_429),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1042),
.A2(n_641),
.B(n_638),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1141),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1119),
.A2(n_384),
.B1(n_402),
.B2(n_288),
.Y(n_1229)
);

OAI22xp5_ASAP7_75t_SL g1230 ( 
.A1(n_1017),
.A2(n_1046),
.B1(n_271),
.B2(n_272),
.Y(n_1230)
);

HB1xp67_ASAP7_75t_L g1231 ( 
.A(n_1115),
.Y(n_1231)
);

NAND2xp5_ASAP7_75t_L g1232 ( 
.A(n_1109),
.B(n_1111),
.Y(n_1232)
);

NOR2xp33_ASAP7_75t_L g1233 ( 
.A(n_1128),
.B(n_270),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_SL g1234 ( 
.A1(n_1098),
.A2(n_611),
.B(n_610),
.C(n_603),
.Y(n_1234)
);

AND2x4_ASAP7_75t_L g1235 ( 
.A(n_1115),
.B(n_980),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1151),
.A2(n_641),
.B(n_638),
.C(n_610),
.Y(n_1236)
);

O2A1O1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_1050),
.A2(n_611),
.B(n_610),
.C(n_603),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1145),
.B(n_991),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_980),
.B(n_87),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_990),
.A2(n_610),
.B(n_603),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_1097),
.B(n_430),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1032),
.B(n_431),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1020),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1120),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_990),
.A2(n_610),
.B(n_426),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1117),
.B(n_433),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_1126),
.Y(n_1247)
);

OAI21xp33_ASAP7_75t_L g1248 ( 
.A1(n_1065),
.A2(n_379),
.B(n_364),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_R g1249 ( 
.A(n_1057),
.B(n_434),
.Y(n_1249)
);

INVx4_ASAP7_75t_L g1250 ( 
.A(n_1068),
.Y(n_1250)
);

INVx3_ASAP7_75t_SL g1251 ( 
.A(n_1001),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1138),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_987),
.A2(n_644),
.B(n_436),
.Y(n_1253)
);

O2A1O1Ixp5_ASAP7_75t_SL g1254 ( 
.A1(n_1088),
.A2(n_403),
.B(n_288),
.C(n_402),
.Y(n_1254)
);

NOR2xp33_ASAP7_75t_L g1255 ( 
.A(n_1007),
.B(n_271),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1117),
.B(n_434),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1140),
.Y(n_1257)
);

AOI21xp5_ASAP7_75t_L g1258 ( 
.A1(n_987),
.A2(n_644),
.B(n_436),
.Y(n_1258)
);

OR2x6_ASAP7_75t_L g1259 ( 
.A(n_1068),
.B(n_1155),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1146),
.Y(n_1260)
);

OAI22xp5_ASAP7_75t_L g1261 ( 
.A1(n_986),
.A2(n_379),
.B1(n_369),
.B2(n_368),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1018),
.A2(n_1023),
.B(n_985),
.Y(n_1262)
);

O2A1O1Ixp33_ASAP7_75t_L g1263 ( 
.A1(n_1085),
.A2(n_384),
.B(n_288),
.C(n_644),
.Y(n_1263)
);

INVx11_ASAP7_75t_L g1264 ( 
.A(n_1127),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1127),
.B(n_364),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_L g1266 ( 
.A(n_1009),
.B(n_644),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_R g1267 ( 
.A(n_1068),
.B(n_367),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_977),
.A2(n_369),
.B1(n_368),
.B2(n_367),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_SL g1269 ( 
.A(n_1010),
.B(n_644),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1116),
.B(n_644),
.Y(n_1270)
);

BUFx6f_ASAP7_75t_L g1271 ( 
.A(n_1002),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1123),
.Y(n_1272)
);

AO21x1_ASAP7_75t_L g1273 ( 
.A1(n_1078),
.A2(n_1103),
.B(n_1156),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_1155),
.Y(n_1274)
);

NOR2x1_ASAP7_75t_L g1275 ( 
.A(n_1095),
.B(n_644),
.Y(n_1275)
);

NAND2x1_ASAP7_75t_L g1276 ( 
.A(n_1130),
.B(n_644),
.Y(n_1276)
);

NOR2xp33_ASAP7_75t_L g1277 ( 
.A(n_1100),
.B(n_8),
.Y(n_1277)
);

AO21x1_ASAP7_75t_L g1278 ( 
.A1(n_999),
.A2(n_9),
.B(n_11),
.Y(n_1278)
);

O2A1O1Ixp33_ASAP7_75t_SL g1279 ( 
.A1(n_1059),
.A2(n_215),
.B(n_214),
.C(n_211),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1033),
.A2(n_209),
.B(n_207),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_995),
.B(n_14),
.Y(n_1281)
);

OAI22xp5_ASAP7_75t_L g1282 ( 
.A1(n_1064),
.A2(n_205),
.B1(n_197),
.B2(n_195),
.Y(n_1282)
);

INVx1_ASAP7_75t_SL g1283 ( 
.A(n_1155),
.Y(n_1283)
);

OR2x6_ASAP7_75t_SL g1284 ( 
.A(n_1090),
.B(n_14),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_985),
.A2(n_186),
.B(n_181),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_989),
.A2(n_15),
.B(n_18),
.C(n_21),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1107),
.B(n_21),
.Y(n_1287)
);

BUFx6f_ASAP7_75t_L g1288 ( 
.A(n_1002),
.Y(n_1288)
);

A2O1A1Ixp33_ASAP7_75t_SL g1289 ( 
.A1(n_1062),
.A2(n_179),
.B(n_176),
.C(n_170),
.Y(n_1289)
);

NAND2xp5_ASAP7_75t_SL g1290 ( 
.A(n_1118),
.B(n_1121),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1122),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1108),
.B(n_25),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_997),
.B(n_26),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1150),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1105),
.B(n_27),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1084),
.B(n_28),
.Y(n_1296)
);

OAI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1066),
.A2(n_169),
.B1(n_166),
.B2(n_165),
.Y(n_1297)
);

HB1xp67_ASAP7_75t_L g1298 ( 
.A(n_1019),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1022),
.A2(n_163),
.B1(n_156),
.B2(n_149),
.Y(n_1299)
);

BUFx4f_ASAP7_75t_SL g1300 ( 
.A(n_1158),
.Y(n_1300)
);

INVx2_ASAP7_75t_L g1301 ( 
.A(n_1051),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_SL g1302 ( 
.A(n_1028),
.B(n_146),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1070),
.B(n_1074),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1011),
.A2(n_133),
.B(n_130),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1079),
.B(n_29),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1081),
.Y(n_1306)
);

A2O1A1Ixp33_ASAP7_75t_L g1307 ( 
.A1(n_1038),
.A2(n_32),
.B(n_33),
.C(n_35),
.Y(n_1307)
);

A2O1A1Ixp33_ASAP7_75t_L g1308 ( 
.A1(n_1039),
.A2(n_32),
.B(n_36),
.C(n_37),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1125),
.Y(n_1309)
);

INVxp67_ASAP7_75t_L g1310 ( 
.A(n_1082),
.Y(n_1310)
);

OAI22xp5_ASAP7_75t_L g1311 ( 
.A1(n_1045),
.A2(n_141),
.B1(n_126),
.B2(n_120),
.Y(n_1311)
);

NAND2xp5_ASAP7_75t_L g1312 ( 
.A(n_1089),
.B(n_36),
.Y(n_1312)
);

AOI22xp5_ASAP7_75t_L g1313 ( 
.A1(n_982),
.A2(n_116),
.B1(n_97),
.B2(n_42),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1093),
.B(n_38),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1147),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1102),
.B(n_38),
.Y(n_1316)
);

A2O1A1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1006),
.A2(n_39),
.B(n_43),
.C(n_44),
.Y(n_1317)
);

HB1xp67_ASAP7_75t_L g1318 ( 
.A(n_1035),
.Y(n_1318)
);

CKINVDCx8_ASAP7_75t_R g1319 ( 
.A(n_1036),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1232),
.B(n_1054),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1185),
.Y(n_1321)
);

AOI21xp5_ASAP7_75t_SL g1322 ( 
.A1(n_1162),
.A2(n_1045),
.B(n_1036),
.Y(n_1322)
);

AO31x2_ASAP7_75t_L g1323 ( 
.A1(n_1273),
.A2(n_1076),
.A3(n_1029),
.B(n_1025),
.Y(n_1323)
);

OAI21x1_ASAP7_75t_L g1324 ( 
.A1(n_1189),
.A2(n_1055),
.B(n_1060),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_L g1325 ( 
.A1(n_1163),
.A2(n_1024),
.B(n_1025),
.Y(n_1325)
);

AOI21xp5_ASAP7_75t_L g1326 ( 
.A1(n_1163),
.A2(n_1162),
.B(n_1262),
.Y(n_1326)
);

HB1xp67_ASAP7_75t_L g1327 ( 
.A(n_1161),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1169),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1231),
.B(n_1047),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1278),
.A2(n_1024),
.A3(n_1087),
.B(n_1096),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1262),
.A2(n_1037),
.B(n_1087),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1229),
.A2(n_1075),
.B(n_1053),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1202),
.B(n_1160),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1303),
.A2(n_1044),
.B(n_1043),
.Y(n_1334)
);

AOI21xp5_ASAP7_75t_L g1335 ( 
.A1(n_1270),
.A2(n_1040),
.B(n_1091),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1188),
.A2(n_1091),
.B(n_1092),
.Y(n_1336)
);

AOI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1177),
.A2(n_1092),
.B(n_1096),
.Y(n_1337)
);

INVx2_ASAP7_75t_L g1338 ( 
.A(n_1222),
.Y(n_1338)
);

BUFx4f_ASAP7_75t_L g1339 ( 
.A(n_1185),
.Y(n_1339)
);

OAI22xp5_ASAP7_75t_L g1340 ( 
.A1(n_1318),
.A2(n_1136),
.B1(n_1142),
.B2(n_1104),
.Y(n_1340)
);

AOI211x1_ASAP7_75t_L g1341 ( 
.A1(n_1248),
.A2(n_1209),
.B(n_1193),
.C(n_1290),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1294),
.B(n_1149),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_SL g1343 ( 
.A(n_1167),
.B(n_1144),
.Y(n_1343)
);

NAND2xp5_ASAP7_75t_L g1344 ( 
.A(n_1244),
.B(n_1247),
.Y(n_1344)
);

NOR2xp33_ASAP7_75t_L g1345 ( 
.A(n_1176),
.B(n_1135),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1177),
.A2(n_1135),
.B(n_1106),
.Y(n_1346)
);

AOI21x1_ASAP7_75t_L g1347 ( 
.A1(n_1186),
.A2(n_1104),
.B(n_1106),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1166),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1217),
.A2(n_1227),
.B(n_1218),
.Y(n_1349)
);

NAND3x1_ASAP7_75t_L g1350 ( 
.A(n_1205),
.B(n_44),
.C(n_45),
.Y(n_1350)
);

NAND2xp5_ASAP7_75t_SL g1351 ( 
.A(n_1235),
.B(n_1112),
.Y(n_1351)
);

AOI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1291),
.A2(n_1153),
.B1(n_1148),
.B2(n_1112),
.Y(n_1352)
);

NOR2xp33_ASAP7_75t_L g1353 ( 
.A(n_1195),
.B(n_1133),
.Y(n_1353)
);

AOI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1305),
.A2(n_1133),
.B(n_1131),
.Y(n_1354)
);

AOI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1266),
.A2(n_1131),
.B(n_1139),
.Y(n_1355)
);

AO31x2_ASAP7_75t_L g1356 ( 
.A1(n_1286),
.A2(n_1308),
.A3(n_1258),
.B(n_1253),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1306),
.A2(n_1142),
.B(n_1136),
.Y(n_1357)
);

AOI21xp5_ASAP7_75t_L g1358 ( 
.A1(n_1170),
.A2(n_1143),
.B(n_49),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_L g1359 ( 
.A1(n_1171),
.A2(n_47),
.B(n_49),
.Y(n_1359)
);

NAND2xp5_ASAP7_75t_L g1360 ( 
.A(n_1252),
.B(n_50),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1223),
.Y(n_1361)
);

NAND2xp33_ASAP7_75t_L g1362 ( 
.A(n_1183),
.B(n_53),
.Y(n_1362)
);

NAND2xp5_ASAP7_75t_L g1363 ( 
.A(n_1257),
.B(n_74),
.Y(n_1363)
);

OA21x2_ASAP7_75t_L g1364 ( 
.A1(n_1253),
.A2(n_1258),
.B(n_1306),
.Y(n_1364)
);

INVx1_ASAP7_75t_SL g1365 ( 
.A(n_1172),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1216),
.A2(n_53),
.B(n_55),
.Y(n_1366)
);

AO32x2_ASAP7_75t_L g1367 ( 
.A1(n_1261),
.A2(n_55),
.A3(n_56),
.B1(n_58),
.B2(n_60),
.Y(n_1367)
);

AO21x2_ASAP7_75t_L g1368 ( 
.A1(n_1175),
.A2(n_58),
.B(n_60),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1216),
.A2(n_62),
.B(n_63),
.Y(n_1369)
);

AND2x4_ASAP7_75t_L g1370 ( 
.A(n_1235),
.B(n_62),
.Y(n_1370)
);

AO21x1_ASAP7_75t_L g1371 ( 
.A1(n_1263),
.A2(n_63),
.B(n_64),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1221),
.B(n_72),
.Y(n_1372)
);

AOI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1187),
.A2(n_73),
.B(n_1238),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1226),
.B(n_1192),
.Y(n_1374)
);

BUFx10_ASAP7_75t_L g1375 ( 
.A(n_1164),
.Y(n_1375)
);

BUFx3_ASAP7_75t_L g1376 ( 
.A(n_1182),
.Y(n_1376)
);

NOR2x1_ASAP7_75t_L g1377 ( 
.A(n_1250),
.B(n_1194),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1234),
.A2(n_1236),
.B(n_1245),
.Y(n_1378)
);

AO32x2_ASAP7_75t_L g1379 ( 
.A1(n_1230),
.A2(n_1268),
.A3(n_1299),
.B1(n_1297),
.B2(n_1282),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_L g1380 ( 
.A1(n_1218),
.A2(n_1240),
.B(n_1180),
.Y(n_1380)
);

A2O1A1Ixp33_ASAP7_75t_L g1381 ( 
.A1(n_1233),
.A2(n_1277),
.B(n_1292),
.C(n_1255),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1260),
.B(n_1301),
.Y(n_1382)
);

AND2x4_ASAP7_75t_L g1383 ( 
.A(n_1250),
.B(n_1259),
.Y(n_1383)
);

AOI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1180),
.A2(n_1165),
.B(n_1199),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1310),
.B(n_1298),
.Y(n_1385)
);

INVx5_ASAP7_75t_L g1386 ( 
.A(n_1185),
.Y(n_1386)
);

OAI21xp5_ASAP7_75t_L g1387 ( 
.A1(n_1310),
.A2(n_1312),
.B(n_1314),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1243),
.Y(n_1388)
);

OAI21x1_ASAP7_75t_SL g1389 ( 
.A1(n_1285),
.A2(n_1304),
.B(n_1236),
.Y(n_1389)
);

AOI21xp5_ASAP7_75t_L g1390 ( 
.A1(n_1190),
.A2(n_1309),
.B(n_1304),
.Y(n_1390)
);

AOI21xp5_ASAP7_75t_L g1391 ( 
.A1(n_1302),
.A2(n_1245),
.B(n_1315),
.Y(n_1391)
);

AOI21xp5_ASAP7_75t_L g1392 ( 
.A1(n_1208),
.A2(n_1174),
.B(n_1184),
.Y(n_1392)
);

AO21x2_ASAP7_75t_L g1393 ( 
.A1(n_1208),
.A2(n_1240),
.B(n_1285),
.Y(n_1393)
);

O2A1O1Ixp5_ASAP7_75t_L g1394 ( 
.A1(n_1316),
.A2(n_1296),
.B(n_1295),
.C(n_1196),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1291),
.B(n_1274),
.Y(n_1395)
);

AO31x2_ASAP7_75t_L g1396 ( 
.A1(n_1307),
.A2(n_1317),
.A3(n_1207),
.B(n_1220),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1272),
.Y(n_1397)
);

AO31x2_ASAP7_75t_L g1398 ( 
.A1(n_1207),
.A2(n_1220),
.A3(n_1293),
.B(n_1281),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1184),
.A2(n_1269),
.B(n_1263),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1198),
.A2(n_1215),
.B1(n_1283),
.B2(n_1214),
.Y(n_1400)
);

NOR2x1_ASAP7_75t_SL g1401 ( 
.A(n_1259),
.B(n_1271),
.Y(n_1401)
);

INVx2_ASAP7_75t_SL g1402 ( 
.A(n_1219),
.Y(n_1402)
);

AND2x4_ASAP7_75t_L g1403 ( 
.A(n_1259),
.B(n_1239),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1246),
.B(n_1256),
.Y(n_1404)
);

A2O1A1Ixp33_ASAP7_75t_L g1405 ( 
.A1(n_1313),
.A2(n_1197),
.B(n_1229),
.C(n_1287),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1173),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1210),
.Y(n_1407)
);

OAI22x1_ASAP7_75t_L g1408 ( 
.A1(n_1251),
.A2(n_1284),
.B1(n_1265),
.B2(n_1212),
.Y(n_1408)
);

AND2x4_ASAP7_75t_L g1409 ( 
.A(n_1239),
.B(n_1191),
.Y(n_1409)
);

AOI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1184),
.A2(n_1280),
.B(n_1275),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1242),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1168),
.A2(n_1178),
.B(n_1279),
.Y(n_1412)
);

INVx2_ASAP7_75t_SL g1413 ( 
.A(n_1191),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1213),
.A2(n_1254),
.B(n_1237),
.Y(n_1414)
);

OAI21xp5_ASAP7_75t_SL g1415 ( 
.A1(n_1211),
.A2(n_1204),
.B(n_1200),
.Y(n_1415)
);

OR2x2_ASAP7_75t_L g1416 ( 
.A(n_1203),
.B(n_1191),
.Y(n_1416)
);

HB1xp67_ASAP7_75t_L g1417 ( 
.A(n_1224),
.Y(n_1417)
);

OR2x2_ASAP7_75t_L g1418 ( 
.A(n_1228),
.B(n_1179),
.Y(n_1418)
);

OAI22x1_ASAP7_75t_L g1419 ( 
.A1(n_1213),
.A2(n_1225),
.B1(n_1241),
.B2(n_1168),
.Y(n_1419)
);

INVx4_ASAP7_75t_L g1420 ( 
.A(n_1264),
.Y(n_1420)
);

AOI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1178),
.A2(n_1289),
.B(n_1311),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_SL g1422 ( 
.A1(n_1276),
.A2(n_1237),
.B(n_1319),
.C(n_1300),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1271),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1201),
.A2(n_1271),
.B(n_1288),
.Y(n_1424)
);

A2O1A1Ixp33_ASAP7_75t_L g1425 ( 
.A1(n_1206),
.A2(n_1288),
.B(n_1181),
.C(n_1249),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1288),
.A2(n_1137),
.B(n_851),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_L g1427 ( 
.A1(n_1267),
.A2(n_981),
.B(n_988),
.Y(n_1427)
);

AOI22xp5_ASAP7_75t_L g1428 ( 
.A1(n_1294),
.A2(n_872),
.B1(n_740),
.B2(n_452),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1169),
.Y(n_1429)
);

AOI22xp5_ASAP7_75t_L g1430 ( 
.A1(n_1294),
.A2(n_872),
.B1(n_740),
.B2(n_452),
.Y(n_1430)
);

INVx3_ASAP7_75t_L g1431 ( 
.A(n_1194),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1167),
.Y(n_1432)
);

AO31x2_ASAP7_75t_L g1433 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1433)
);

AO31x2_ASAP7_75t_L g1434 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1434)
);

O2A1O1Ixp33_ASAP7_75t_L g1435 ( 
.A1(n_1277),
.A2(n_981),
.B(n_872),
.C(n_1015),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1294),
.B(n_845),
.Y(n_1436)
);

AOI21xp5_ASAP7_75t_L g1437 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1437)
);

OAI21xp33_ASAP7_75t_L g1438 ( 
.A1(n_1229),
.A2(n_872),
.B(n_901),
.Y(n_1438)
);

O2A1O1Ixp33_ASAP7_75t_L g1439 ( 
.A1(n_1277),
.A2(n_981),
.B(n_872),
.C(n_1015),
.Y(n_1439)
);

OAI21xp5_ASAP7_75t_L g1440 ( 
.A1(n_1232),
.A2(n_981),
.B(n_988),
.Y(n_1440)
);

OAI21xp5_ASAP7_75t_L g1441 ( 
.A1(n_1232),
.A2(n_981),
.B(n_988),
.Y(n_1441)
);

NAND2xp5_ASAP7_75t_L g1442 ( 
.A(n_1232),
.B(n_981),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1189),
.A2(n_1262),
.B(n_1217),
.Y(n_1443)
);

AOI21xp5_ASAP7_75t_L g1444 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1189),
.A2(n_1262),
.B(n_1217),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1232),
.B(n_981),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1189),
.A2(n_1262),
.B(n_1217),
.Y(n_1447)
);

CKINVDCx20_ASAP7_75t_R g1448 ( 
.A(n_1167),
.Y(n_1448)
);

AOI21xp5_ASAP7_75t_L g1449 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_SL g1450 ( 
.A(n_1181),
.Y(n_1450)
);

AO31x2_ASAP7_75t_L g1451 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1262),
.A2(n_1273),
.B(n_1163),
.Y(n_1452)
);

AOI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1231),
.B(n_859),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1455)
);

NOR2xp33_ASAP7_75t_L g1456 ( 
.A(n_1294),
.B(n_845),
.Y(n_1456)
);

AND2x4_ASAP7_75t_L g1457 ( 
.A(n_1235),
.B(n_1250),
.Y(n_1457)
);

AOI21xp5_ASAP7_75t_SL g1458 ( 
.A1(n_1162),
.A2(n_909),
.B(n_897),
.Y(n_1458)
);

CKINVDCx6p67_ASAP7_75t_R g1459 ( 
.A(n_1172),
.Y(n_1459)
);

AO31x2_ASAP7_75t_L g1460 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1460)
);

AOI21xp5_ASAP7_75t_L g1461 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1461)
);

AOI21xp5_ASAP7_75t_L g1462 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1462)
);

AND2x4_ASAP7_75t_L g1463 ( 
.A(n_1235),
.B(n_1250),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1232),
.A2(n_981),
.B1(n_672),
.B2(n_696),
.Y(n_1464)
);

AO31x2_ASAP7_75t_L g1465 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1465)
);

AO21x2_ASAP7_75t_L g1466 ( 
.A1(n_1163),
.A2(n_1262),
.B(n_1273),
.Y(n_1466)
);

A2O1A1Ixp33_ASAP7_75t_L g1467 ( 
.A1(n_1162),
.A2(n_981),
.B(n_696),
.C(n_872),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1169),
.Y(n_1468)
);

A2O1A1Ixp33_ASAP7_75t_L g1469 ( 
.A1(n_1162),
.A2(n_981),
.B(n_696),
.C(n_872),
.Y(n_1469)
);

AO31x2_ASAP7_75t_L g1470 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1470)
);

AOI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1203),
.A2(n_1015),
.B1(n_919),
.B2(n_1063),
.C(n_691),
.Y(n_1471)
);

AOI21xp5_ASAP7_75t_L g1472 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1472)
);

AO31x2_ASAP7_75t_L g1473 ( 
.A1(n_1273),
.A2(n_1278),
.A3(n_1262),
.B(n_1163),
.Y(n_1473)
);

OR2x2_ASAP7_75t_L g1474 ( 
.A(n_1161),
.B(n_682),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1232),
.B(n_981),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1189),
.A2(n_1262),
.B(n_1217),
.Y(n_1476)
);

NAND2xp33_ASAP7_75t_L g1477 ( 
.A(n_1183),
.B(n_981),
.Y(n_1477)
);

INVx5_ASAP7_75t_SL g1478 ( 
.A(n_1264),
.Y(n_1478)
);

NOR2xp67_ASAP7_75t_L g1479 ( 
.A(n_1202),
.B(n_931),
.Y(n_1479)
);

AOI221xp5_ASAP7_75t_L g1480 ( 
.A1(n_1203),
.A2(n_1015),
.B1(n_919),
.B2(n_1063),
.C(n_691),
.Y(n_1480)
);

NAND2xp5_ASAP7_75t_SL g1481 ( 
.A(n_1294),
.B(n_994),
.Y(n_1481)
);

NOR2xp33_ASAP7_75t_SL g1482 ( 
.A(n_1167),
.B(n_875),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_SL g1483 ( 
.A1(n_1203),
.A2(n_919),
.B1(n_1277),
.B2(n_1292),
.C(n_1248),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_1167),
.Y(n_1484)
);

NOR2xp67_ASAP7_75t_L g1485 ( 
.A(n_1202),
.B(n_931),
.Y(n_1485)
);

AOI21xp5_ASAP7_75t_L g1486 ( 
.A1(n_1163),
.A2(n_1137),
.B(n_851),
.Y(n_1486)
);

NOR4xp25_ASAP7_75t_L g1487 ( 
.A(n_1317),
.B(n_981),
.C(n_919),
.D(n_872),
.Y(n_1487)
);

BUFx2_ASAP7_75t_L g1488 ( 
.A(n_1376),
.Y(n_1488)
);

CKINVDCx11_ASAP7_75t_R g1489 ( 
.A(n_1432),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_SL g1490 ( 
.A1(n_1362),
.A2(n_1427),
.B1(n_1436),
.B2(n_1456),
.Y(n_1490)
);

BUFx4f_ASAP7_75t_SL g1491 ( 
.A(n_1448),
.Y(n_1491)
);

BUFx4f_ASAP7_75t_SL g1492 ( 
.A(n_1459),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_L g1493 ( 
.A1(n_1438),
.A2(n_1471),
.B1(n_1480),
.B2(n_1430),
.Y(n_1493)
);

BUFx8_ASAP7_75t_L g1494 ( 
.A(n_1450),
.Y(n_1494)
);

AOI22xp33_ASAP7_75t_L g1495 ( 
.A1(n_1428),
.A2(n_1372),
.B1(n_1481),
.B2(n_1464),
.Y(n_1495)
);

OAI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1400),
.A2(n_1343),
.B1(n_1475),
.B2(n_1442),
.Y(n_1496)
);

OAI22xp5_ASAP7_75t_L g1497 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1344),
.B2(n_1405),
.Y(n_1497)
);

CKINVDCx20_ASAP7_75t_R g1498 ( 
.A(n_1484),
.Y(n_1498)
);

AOI22xp33_ASAP7_75t_L g1499 ( 
.A1(n_1411),
.A2(n_1353),
.B1(n_1408),
.B2(n_1371),
.Y(n_1499)
);

CKINVDCx20_ASAP7_75t_R g1500 ( 
.A(n_1407),
.Y(n_1500)
);

OAI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1482),
.A2(n_1415),
.B1(n_1374),
.B2(n_1365),
.Y(n_1501)
);

BUFx2_ASAP7_75t_L g1502 ( 
.A(n_1402),
.Y(n_1502)
);

BUFx10_ASAP7_75t_L g1503 ( 
.A(n_1450),
.Y(n_1503)
);

NAND2x1p5_ASAP7_75t_L g1504 ( 
.A(n_1383),
.B(n_1386),
.Y(n_1504)
);

BUFx12f_ASAP7_75t_L g1505 ( 
.A(n_1420),
.Y(n_1505)
);

BUFx6f_ASAP7_75t_L g1506 ( 
.A(n_1339),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1375),
.Y(n_1507)
);

CKINVDCx16_ASAP7_75t_R g1508 ( 
.A(n_1420),
.Y(n_1508)
);

BUFx6f_ASAP7_75t_L g1509 ( 
.A(n_1339),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_L g1510 ( 
.A1(n_1404),
.A2(n_1342),
.B1(n_1345),
.B2(n_1419),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1375),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1361),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_L g1513 ( 
.A1(n_1387),
.A2(n_1440),
.B1(n_1441),
.B2(n_1351),
.Y(n_1513)
);

BUFx10_ASAP7_75t_L g1514 ( 
.A(n_1370),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1328),
.B(n_1348),
.Y(n_1515)
);

OAI22xp33_ASAP7_75t_L g1516 ( 
.A1(n_1416),
.A2(n_1363),
.B1(n_1360),
.B2(n_1385),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_L g1517 ( 
.A(n_1328),
.B(n_1348),
.Y(n_1517)
);

INVx6_ASAP7_75t_L g1518 ( 
.A(n_1386),
.Y(n_1518)
);

AOI22xp33_ASAP7_75t_L g1519 ( 
.A1(n_1454),
.A2(n_1403),
.B1(n_1329),
.B2(n_1370),
.Y(n_1519)
);

INVx1_ASAP7_75t_SL g1520 ( 
.A(n_1474),
.Y(n_1520)
);

BUFx2_ASAP7_75t_SL g1521 ( 
.A(n_1386),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_SL g1522 ( 
.A1(n_1403),
.A2(n_1401),
.B1(n_1477),
.B2(n_1483),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1395),
.Y(n_1523)
);

INVxp67_ASAP7_75t_L g1524 ( 
.A(n_1417),
.Y(n_1524)
);

CKINVDCx11_ASAP7_75t_R g1525 ( 
.A(n_1321),
.Y(n_1525)
);

OAI22xp33_ASAP7_75t_L g1526 ( 
.A1(n_1382),
.A2(n_1418),
.B1(n_1479),
.B2(n_1485),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1333),
.A2(n_1468),
.B1(n_1429),
.B2(n_1373),
.Y(n_1527)
);

CKINVDCx11_ASAP7_75t_R g1528 ( 
.A(n_1321),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1429),
.A2(n_1468),
.B1(n_1414),
.B2(n_1359),
.Y(n_1529)
);

BUFx4f_ASAP7_75t_L g1530 ( 
.A(n_1457),
.Y(n_1530)
);

CKINVDCx6p67_ASAP7_75t_R g1531 ( 
.A(n_1321),
.Y(n_1531)
);

AOI22xp5_ASAP7_75t_L g1532 ( 
.A1(n_1350),
.A2(n_1409),
.B1(n_1383),
.B2(n_1332),
.Y(n_1532)
);

BUFx10_ASAP7_75t_L g1533 ( 
.A(n_1457),
.Y(n_1533)
);

BUFx6f_ASAP7_75t_L g1534 ( 
.A(n_1463),
.Y(n_1534)
);

BUFx6f_ASAP7_75t_L g1535 ( 
.A(n_1463),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1364),
.A2(n_1397),
.B1(n_1388),
.B2(n_1409),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1406),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1413),
.Y(n_1538)
);

AOI22xp33_ASAP7_75t_SL g1539 ( 
.A1(n_1389),
.A2(n_1435),
.B1(n_1439),
.B2(n_1379),
.Y(n_1539)
);

CKINVDCx20_ASAP7_75t_R g1540 ( 
.A(n_1478),
.Y(n_1540)
);

BUFx12f_ASAP7_75t_L g1541 ( 
.A(n_1478),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1364),
.A2(n_1391),
.B1(n_1320),
.B2(n_1358),
.Y(n_1542)
);

AOI22xp33_ASAP7_75t_SL g1543 ( 
.A1(n_1379),
.A2(n_1487),
.B1(n_1366),
.B2(n_1369),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1423),
.Y(n_1544)
);

BUFx12f_ASAP7_75t_L g1545 ( 
.A(n_1425),
.Y(n_1545)
);

OAI22xp5_ASAP7_75t_L g1546 ( 
.A1(n_1467),
.A2(n_1469),
.B1(n_1341),
.B2(n_1392),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1424),
.Y(n_1547)
);

INVx2_ASAP7_75t_SL g1548 ( 
.A(n_1377),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1368),
.A2(n_1466),
.B1(n_1326),
.B2(n_1393),
.Y(n_1549)
);

BUFx10_ASAP7_75t_L g1550 ( 
.A(n_1394),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1352),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1368),
.A2(n_1466),
.B1(n_1393),
.B2(n_1378),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1367),
.Y(n_1553)
);

INVx6_ASAP7_75t_L g1554 ( 
.A(n_1431),
.Y(n_1554)
);

INVx3_ASAP7_75t_L g1555 ( 
.A(n_1396),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_SL g1556 ( 
.A1(n_1379),
.A2(n_1421),
.B1(n_1452),
.B2(n_1367),
.Y(n_1556)
);

INVx1_ASAP7_75t_SL g1557 ( 
.A(n_1452),
.Y(n_1557)
);

INVx1_ASAP7_75t_SL g1558 ( 
.A(n_1412),
.Y(n_1558)
);

AOI22xp33_ASAP7_75t_L g1559 ( 
.A1(n_1378),
.A2(n_1426),
.B1(n_1390),
.B2(n_1340),
.Y(n_1559)
);

INVx2_ASAP7_75t_SL g1560 ( 
.A(n_1396),
.Y(n_1560)
);

AOI22xp33_ASAP7_75t_L g1561 ( 
.A1(n_1357),
.A2(n_1334),
.B1(n_1384),
.B2(n_1399),
.Y(n_1561)
);

OAI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1437),
.A2(n_1449),
.B1(n_1472),
.B2(n_1462),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_SL g1563 ( 
.A1(n_1367),
.A2(n_1486),
.B1(n_1461),
.B2(n_1444),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1433),
.B(n_1470),
.Y(n_1564)
);

AOI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1422),
.A2(n_1455),
.B1(n_1453),
.B2(n_1335),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_L g1566 ( 
.A1(n_1325),
.A2(n_1336),
.B1(n_1337),
.B2(n_1346),
.Y(n_1566)
);

CKINVDCx5p33_ASAP7_75t_R g1567 ( 
.A(n_1322),
.Y(n_1567)
);

BUFx2_ASAP7_75t_SL g1568 ( 
.A(n_1410),
.Y(n_1568)
);

INVx1_ASAP7_75t_L g1569 ( 
.A(n_1434),
.Y(n_1569)
);

OAI22x1_ASAP7_75t_L g1570 ( 
.A1(n_1354),
.A2(n_1347),
.B1(n_1458),
.B2(n_1356),
.Y(n_1570)
);

BUFx12f_ASAP7_75t_L g1571 ( 
.A(n_1398),
.Y(n_1571)
);

BUFx4f_ASAP7_75t_SL g1572 ( 
.A(n_1356),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1355),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1356),
.B(n_1451),
.Y(n_1574)
);

BUFx6f_ASAP7_75t_L g1575 ( 
.A(n_1380),
.Y(n_1575)
);

AOI22xp33_ASAP7_75t_SL g1576 ( 
.A1(n_1331),
.A2(n_1445),
.B1(n_1447),
.B2(n_1443),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1460),
.B(n_1473),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1460),
.Y(n_1578)
);

OAI22x1_ASAP7_75t_L g1579 ( 
.A1(n_1460),
.A2(n_1473),
.B1(n_1470),
.B2(n_1465),
.Y(n_1579)
);

INVx1_ASAP7_75t_SL g1580 ( 
.A(n_1349),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1465),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_SL g1582 ( 
.A1(n_1476),
.A2(n_1465),
.B1(n_1470),
.B2(n_1473),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1398),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1398),
.Y(n_1584)
);

BUFx8_ASAP7_75t_L g1585 ( 
.A(n_1330),
.Y(n_1585)
);

INVxp33_ASAP7_75t_SL g1586 ( 
.A(n_1324),
.Y(n_1586)
);

INVx4_ASAP7_75t_L g1587 ( 
.A(n_1330),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1330),
.A2(n_1438),
.B1(n_1134),
.B2(n_1015),
.Y(n_1588)
);

BUFx3_ASAP7_75t_L g1589 ( 
.A(n_1323),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1323),
.Y(n_1590)
);

CKINVDCx6p67_ASAP7_75t_R g1591 ( 
.A(n_1432),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1593)
);

INVx6_ASAP7_75t_L g1594 ( 
.A(n_1386),
.Y(n_1594)
);

INVx6_ASAP7_75t_L g1595 ( 
.A(n_1386),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_SL g1597 ( 
.A(n_1381),
.B(n_1427),
.Y(n_1597)
);

BUFx2_ASAP7_75t_R g1598 ( 
.A(n_1484),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1338),
.Y(n_1599)
);

OAI22xp5_ASAP7_75t_L g1600 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1475),
.B2(n_1442),
.Y(n_1600)
);

AOI22xp33_ASAP7_75t_SL g1601 ( 
.A1(n_1362),
.A2(n_1134),
.B1(n_452),
.B2(n_454),
.Y(n_1601)
);

INVx6_ASAP7_75t_L g1602 ( 
.A(n_1386),
.Y(n_1602)
);

AOI22xp33_ASAP7_75t_L g1603 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1338),
.Y(n_1604)
);

AOI22xp33_ASAP7_75t_L g1605 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1605)
);

INVx8_ASAP7_75t_L g1606 ( 
.A(n_1386),
.Y(n_1606)
);

AOI22xp33_ASAP7_75t_SL g1607 ( 
.A1(n_1362),
.A2(n_1134),
.B1(n_1221),
.B2(n_981),
.Y(n_1607)
);

AOI22xp33_ASAP7_75t_L g1608 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_1438),
.B2(n_1381),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1407),
.Y(n_1610)
);

OAI21xp33_ASAP7_75t_L g1611 ( 
.A1(n_1381),
.A2(n_1438),
.B(n_872),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1338),
.Y(n_1612)
);

BUFx3_ASAP7_75t_L g1613 ( 
.A(n_1376),
.Y(n_1613)
);

AOI22xp33_ASAP7_75t_L g1614 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1614)
);

AOI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_1438),
.B2(n_1381),
.Y(n_1615)
);

OAI22xp5_ASAP7_75t_L g1616 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1475),
.B2(n_1442),
.Y(n_1616)
);

AOI22xp33_ASAP7_75t_SL g1617 ( 
.A1(n_1362),
.A2(n_1134),
.B1(n_1221),
.B2(n_981),
.Y(n_1617)
);

AOI22xp33_ASAP7_75t_L g1618 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1618)
);

INVx6_ASAP7_75t_L g1619 ( 
.A(n_1386),
.Y(n_1619)
);

OAI22xp5_ASAP7_75t_L g1620 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1475),
.B2(n_1442),
.Y(n_1620)
);

INVx1_ASAP7_75t_SL g1621 ( 
.A(n_1327),
.Y(n_1621)
);

OAI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_696),
.B2(n_981),
.Y(n_1622)
);

AOI22xp33_ASAP7_75t_SL g1623 ( 
.A1(n_1362),
.A2(n_1134),
.B1(n_1221),
.B2(n_981),
.Y(n_1623)
);

INVx6_ASAP7_75t_L g1624 ( 
.A(n_1386),
.Y(n_1624)
);

AOI22xp33_ASAP7_75t_L g1625 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1625)
);

INVx2_ASAP7_75t_SL g1626 ( 
.A(n_1407),
.Y(n_1626)
);

AOI22xp33_ASAP7_75t_L g1627 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1627)
);

AOI22xp33_ASAP7_75t_L g1628 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1338),
.Y(n_1631)
);

INVx1_ASAP7_75t_SL g1632 ( 
.A(n_1327),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1475),
.B2(n_1442),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1381),
.A2(n_1446),
.B1(n_1475),
.B2(n_1442),
.Y(n_1634)
);

OAI22xp33_ASAP7_75t_L g1635 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_696),
.B2(n_981),
.Y(n_1635)
);

AOI22xp33_ASAP7_75t_SL g1636 ( 
.A1(n_1362),
.A2(n_1134),
.B1(n_1221),
.B2(n_981),
.Y(n_1636)
);

CKINVDCx11_ASAP7_75t_R g1637 ( 
.A(n_1432),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1338),
.Y(n_1638)
);

OAI22xp33_ASAP7_75t_L g1639 ( 
.A1(n_1428),
.A2(n_1430),
.B1(n_696),
.B2(n_981),
.Y(n_1639)
);

AOI22xp33_ASAP7_75t_L g1640 ( 
.A1(n_1438),
.A2(n_1134),
.B1(n_1015),
.B2(n_1471),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1440),
.B(n_1441),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1338),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1338),
.Y(n_1643)
);

CKINVDCx11_ASAP7_75t_R g1644 ( 
.A(n_1432),
.Y(n_1644)
);

OR2x2_ASAP7_75t_L g1645 ( 
.A(n_1374),
.B(n_1385),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1569),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1578),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1523),
.Y(n_1648)
);

OAI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1493),
.A2(n_1609),
.B1(n_1615),
.B2(n_1614),
.C(n_1640),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1600),
.B(n_1616),
.Y(n_1650)
);

AOI21x1_ASAP7_75t_L g1651 ( 
.A1(n_1570),
.A2(n_1597),
.B(n_1546),
.Y(n_1651)
);

OAI21x1_ASAP7_75t_L g1652 ( 
.A1(n_1559),
.A2(n_1566),
.B(n_1565),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1504),
.Y(n_1653)
);

INVx2_ASAP7_75t_SL g1654 ( 
.A(n_1554),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1622),
.A2(n_1635),
.B1(n_1639),
.B2(n_1611),
.Y(n_1655)
);

NAND2xp5_ASAP7_75t_L g1656 ( 
.A(n_1600),
.B(n_1616),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1583),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1584),
.Y(n_1658)
);

HB1xp67_ASAP7_75t_L g1659 ( 
.A(n_1621),
.Y(n_1659)
);

HB1xp67_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1556),
.B(n_1574),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1554),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1590),
.Y(n_1663)
);

AO21x2_ASAP7_75t_L g1664 ( 
.A1(n_1562),
.A2(n_1577),
.B(n_1564),
.Y(n_1664)
);

OAI21x1_ASAP7_75t_L g1665 ( 
.A1(n_1542),
.A2(n_1549),
.B(n_1561),
.Y(n_1665)
);

AOI21x1_ASAP7_75t_L g1666 ( 
.A1(n_1546),
.A2(n_1497),
.B(n_1579),
.Y(n_1666)
);

AND2x2_ASAP7_75t_L g1667 ( 
.A(n_1574),
.B(n_1539),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1581),
.Y(n_1668)
);

INVxp67_ASAP7_75t_L g1669 ( 
.A(n_1645),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1551),
.B(n_1588),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1557),
.Y(n_1671)
);

OA21x2_ASAP7_75t_L g1672 ( 
.A1(n_1552),
.A2(n_1536),
.B(n_1557),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1555),
.Y(n_1673)
);

INVx4_ASAP7_75t_L g1674 ( 
.A(n_1606),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1560),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1553),
.B(n_1589),
.Y(n_1676)
);

INVx3_ASAP7_75t_L g1677 ( 
.A(n_1575),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1572),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1543),
.B(n_1587),
.Y(n_1679)
);

BUFx2_ASAP7_75t_L g1680 ( 
.A(n_1571),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1547),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1585),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1585),
.Y(n_1683)
);

AOI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1497),
.A2(n_1630),
.B(n_1629),
.Y(n_1684)
);

OAI21x1_ASAP7_75t_L g1685 ( 
.A1(n_1529),
.A2(n_1513),
.B(n_1596),
.Y(n_1685)
);

INVx2_ASAP7_75t_L g1686 ( 
.A(n_1580),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1580),
.Y(n_1687)
);

INVx2_ASAP7_75t_L g1688 ( 
.A(n_1558),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1515),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1515),
.Y(n_1690)
);

INVx6_ASAP7_75t_L g1691 ( 
.A(n_1533),
.Y(n_1691)
);

BUFx3_ASAP7_75t_L g1692 ( 
.A(n_1504),
.Y(n_1692)
);

BUFx6f_ASAP7_75t_L g1693 ( 
.A(n_1567),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1517),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1558),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1568),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1592),
.A2(n_1629),
.B(n_1596),
.Y(n_1697)
);

BUFx3_ASAP7_75t_L g1698 ( 
.A(n_1606),
.Y(n_1698)
);

AOI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1630),
.A2(n_1641),
.B(n_1633),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1632),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1641),
.Y(n_1701)
);

BUFx3_ASAP7_75t_L g1702 ( 
.A(n_1606),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1537),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1573),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1582),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1620),
.B(n_1633),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1599),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1604),
.Y(n_1708)
);

INVx1_ASAP7_75t_L g1709 ( 
.A(n_1612),
.Y(n_1709)
);

INVx3_ASAP7_75t_L g1710 ( 
.A(n_1550),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1631),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1638),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1642),
.Y(n_1713)
);

HB1xp67_ASAP7_75t_L g1714 ( 
.A(n_1632),
.Y(n_1714)
);

OAI21x1_ASAP7_75t_L g1715 ( 
.A1(n_1527),
.A2(n_1510),
.B(n_1618),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1643),
.Y(n_1716)
);

AOI21xp5_ASAP7_75t_L g1717 ( 
.A1(n_1620),
.A2(n_1634),
.B(n_1563),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1532),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1520),
.Y(n_1719)
);

OAI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1593),
.A2(n_1603),
.B(n_1627),
.Y(n_1720)
);

CKINVDCx20_ASAP7_75t_R g1721 ( 
.A(n_1489),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1550),
.Y(n_1722)
);

OA21x2_ASAP7_75t_L g1723 ( 
.A1(n_1605),
.A2(n_1608),
.B(n_1625),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1628),
.B(n_1512),
.Y(n_1724)
);

OR2x2_ASAP7_75t_L g1725 ( 
.A(n_1634),
.B(n_1520),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1586),
.Y(n_1726)
);

INVx4_ASAP7_75t_L g1727 ( 
.A(n_1518),
.Y(n_1727)
);

AOI22xp33_ASAP7_75t_SL g1728 ( 
.A1(n_1545),
.A2(n_1601),
.B1(n_1636),
.B2(n_1617),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1544),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1576),
.Y(n_1730)
);

BUFx3_ASAP7_75t_L g1731 ( 
.A(n_1518),
.Y(n_1731)
);

INVx2_ASAP7_75t_SL g1732 ( 
.A(n_1554),
.Y(n_1732)
);

HB1xp67_ASAP7_75t_L g1733 ( 
.A(n_1502),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1524),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1516),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1496),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1526),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1495),
.B(n_1499),
.Y(n_1738)
);

INVx2_ASAP7_75t_L g1739 ( 
.A(n_1548),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1601),
.A2(n_1607),
.B1(n_1623),
.B2(n_1490),
.Y(n_1740)
);

BUFx3_ASAP7_75t_L g1741 ( 
.A(n_1594),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1522),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1594),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1595),
.Y(n_1744)
);

BUFx6f_ASAP7_75t_L g1745 ( 
.A(n_1530),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1519),
.B(n_1535),
.Y(n_1746)
);

INVx2_ASAP7_75t_L g1747 ( 
.A(n_1602),
.Y(n_1747)
);

OR2x2_ASAP7_75t_L g1748 ( 
.A(n_1501),
.B(n_1488),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1619),
.Y(n_1749)
);

INVx1_ASAP7_75t_SL g1750 ( 
.A(n_1491),
.Y(n_1750)
);

CKINVDCx20_ASAP7_75t_R g1751 ( 
.A(n_1637),
.Y(n_1751)
);

INVxp67_ASAP7_75t_SL g1752 ( 
.A(n_1534),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1624),
.Y(n_1753)
);

INVx4_ASAP7_75t_L g1754 ( 
.A(n_1530),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1521),
.Y(n_1755)
);

AO31x2_ASAP7_75t_L g1756 ( 
.A1(n_1531),
.A2(n_1514),
.A3(n_1525),
.B(n_1528),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1538),
.Y(n_1757)
);

INVx2_ASAP7_75t_SL g1758 ( 
.A(n_1514),
.Y(n_1758)
);

INVx3_ASAP7_75t_L g1759 ( 
.A(n_1503),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1538),
.Y(n_1760)
);

A2O1A1Ixp33_ASAP7_75t_L g1761 ( 
.A1(n_1610),
.A2(n_1626),
.B(n_1509),
.C(n_1506),
.Y(n_1761)
);

OR2x6_ASAP7_75t_L g1762 ( 
.A(n_1717),
.B(n_1650),
.Y(n_1762)
);

AND2x2_ASAP7_75t_L g1763 ( 
.A(n_1667),
.B(n_1591),
.Y(n_1763)
);

AO21x2_ASAP7_75t_L g1764 ( 
.A1(n_1656),
.A2(n_1507),
.B(n_1511),
.Y(n_1764)
);

AOI22xp33_ASAP7_75t_L g1765 ( 
.A1(n_1649),
.A2(n_1494),
.B1(n_1613),
.B2(n_1541),
.Y(n_1765)
);

AND2x4_ASAP7_75t_L g1766 ( 
.A(n_1678),
.B(n_1506),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_L g1767 ( 
.A(n_1704),
.B(n_1644),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_L g1768 ( 
.A1(n_1740),
.A2(n_1598),
.B1(n_1492),
.B2(n_1508),
.Y(n_1768)
);

INVxp67_ASAP7_75t_L g1769 ( 
.A(n_1719),
.Y(n_1769)
);

AND2x4_ASAP7_75t_L g1770 ( 
.A(n_1678),
.B(n_1506),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1670),
.B(n_1598),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1655),
.A2(n_1706),
.B(n_1720),
.Y(n_1772)
);

OA21x2_ASAP7_75t_L g1773 ( 
.A1(n_1685),
.A2(n_1503),
.B(n_1509),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1682),
.B(n_1500),
.Y(n_1774)
);

AOI22xp33_ASAP7_75t_L g1775 ( 
.A1(n_1723),
.A2(n_1728),
.B1(n_1737),
.B2(n_1736),
.Y(n_1775)
);

INVx4_ASAP7_75t_L g1776 ( 
.A(n_1727),
.Y(n_1776)
);

OR2x2_ASAP7_75t_L g1777 ( 
.A(n_1725),
.B(n_1494),
.Y(n_1777)
);

A2O1A1Ixp33_ASAP7_75t_L g1778 ( 
.A1(n_1715),
.A2(n_1540),
.B(n_1498),
.C(n_1505),
.Y(n_1778)
);

HB1xp67_ASAP7_75t_L g1779 ( 
.A(n_1648),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1685),
.A2(n_1665),
.B(n_1652),
.Y(n_1780)
);

AOI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1738),
.A2(n_1723),
.B1(n_1736),
.B2(n_1742),
.Y(n_1781)
);

AOI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1723),
.A2(n_1742),
.B1(n_1737),
.B2(n_1718),
.Y(n_1782)
);

AOI221xp5_ASAP7_75t_L g1783 ( 
.A1(n_1735),
.A2(n_1670),
.B1(n_1669),
.B2(n_1714),
.C(n_1659),
.Y(n_1783)
);

HB1xp67_ASAP7_75t_SL g1784 ( 
.A(n_1704),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1750),
.B(n_1748),
.Y(n_1785)
);

INVx2_ASAP7_75t_SL g1786 ( 
.A(n_1733),
.Y(n_1786)
);

CKINVDCx5p33_ASAP7_75t_R g1787 ( 
.A(n_1721),
.Y(n_1787)
);

CKINVDCx20_ASAP7_75t_R g1788 ( 
.A(n_1751),
.Y(n_1788)
);

NAND3xp33_ASAP7_75t_L g1789 ( 
.A(n_1735),
.B(n_1723),
.C(n_1748),
.Y(n_1789)
);

AOI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1718),
.A2(n_1715),
.B1(n_1724),
.B2(n_1746),
.Y(n_1790)
);

AOI21xp5_ASAP7_75t_L g1791 ( 
.A1(n_1688),
.A2(n_1695),
.B(n_1664),
.Y(n_1791)
);

OAI22xp5_ASAP7_75t_SL g1792 ( 
.A1(n_1734),
.A2(n_1693),
.B1(n_1722),
.B2(n_1683),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1703),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1722),
.A2(n_1710),
.B(n_1761),
.C(n_1726),
.Y(n_1794)
);

AOI22xp5_ASAP7_75t_L g1795 ( 
.A1(n_1724),
.A2(n_1746),
.B1(n_1660),
.B2(n_1700),
.Y(n_1795)
);

OAI22xp5_ASAP7_75t_L g1796 ( 
.A1(n_1688),
.A2(n_1695),
.B1(n_1689),
.B2(n_1694),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1701),
.B(n_1689),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_SL g1798 ( 
.A1(n_1682),
.A2(n_1683),
.B(n_1755),
.C(n_1758),
.Y(n_1798)
);

OA21x2_ASAP7_75t_L g1799 ( 
.A1(n_1730),
.A2(n_1651),
.B(n_1666),
.Y(n_1799)
);

AND2x2_ASAP7_75t_L g1800 ( 
.A(n_1661),
.B(n_1680),
.Y(n_1800)
);

AO22x1_ASAP7_75t_L g1801 ( 
.A1(n_1693),
.A2(n_1759),
.B1(n_1755),
.B2(n_1752),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1661),
.B(n_1680),
.Y(n_1802)
);

A2O1A1Ixp33_ASAP7_75t_L g1803 ( 
.A1(n_1710),
.A2(n_1726),
.B(n_1759),
.C(n_1758),
.Y(n_1803)
);

AO32x2_ASAP7_75t_L g1804 ( 
.A1(n_1727),
.A2(n_1654),
.A3(n_1662),
.B1(n_1732),
.B2(n_1676),
.Y(n_1804)
);

AND2x4_ASAP7_75t_L g1805 ( 
.A(n_1653),
.B(n_1692),
.Y(n_1805)
);

OAI21x1_ASAP7_75t_SL g1806 ( 
.A1(n_1651),
.A2(n_1666),
.B(n_1684),
.Y(n_1806)
);

NOR2x1_ASAP7_75t_L g1807 ( 
.A(n_1759),
.B(n_1710),
.Y(n_1807)
);

AOI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1701),
.A2(n_1693),
.B1(n_1754),
.B2(n_1759),
.Y(n_1808)
);

OAI21xp5_ASAP7_75t_L g1809 ( 
.A1(n_1684),
.A2(n_1699),
.B(n_1695),
.Y(n_1809)
);

OAI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1699),
.A2(n_1688),
.B(n_1697),
.Y(n_1810)
);

NAND4xp25_ASAP7_75t_L g1811 ( 
.A(n_1707),
.B(n_1708),
.C(n_1709),
.D(n_1711),
.Y(n_1811)
);

O2A1O1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1739),
.A2(n_1760),
.B(n_1757),
.C(n_1696),
.Y(n_1812)
);

O2A1O1Ixp33_ASAP7_75t_SL g1813 ( 
.A1(n_1654),
.A2(n_1662),
.B(n_1732),
.C(n_1744),
.Y(n_1813)
);

AND2x4_ASAP7_75t_L g1814 ( 
.A(n_1653),
.B(n_1692),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1815)
);

AOI22xp5_ASAP7_75t_L g1816 ( 
.A1(n_1754),
.A2(n_1705),
.B1(n_1745),
.B2(n_1679),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1697),
.A2(n_1696),
.B(n_1705),
.Y(n_1817)
);

AO32x2_ASAP7_75t_L g1818 ( 
.A1(n_1727),
.A2(n_1674),
.A3(n_1668),
.B1(n_1671),
.B2(n_1646),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1729),
.B(n_1712),
.Y(n_1819)
);

AOI21xp5_ASAP7_75t_L g1820 ( 
.A1(n_1696),
.A2(n_1690),
.B(n_1694),
.Y(n_1820)
);

BUFx3_ASAP7_75t_L g1821 ( 
.A(n_1756),
.Y(n_1821)
);

AOI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1679),
.A2(n_1716),
.B1(n_1713),
.B2(n_1711),
.C(n_1709),
.Y(n_1822)
);

AO21x2_ASAP7_75t_L g1823 ( 
.A1(n_1675),
.A2(n_1657),
.B(n_1658),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_SL g1824 ( 
.A(n_1754),
.B(n_1745),
.Y(n_1824)
);

AOI22xp5_ASAP7_75t_L g1825 ( 
.A1(n_1754),
.A2(n_1745),
.B1(n_1739),
.B2(n_1690),
.Y(n_1825)
);

BUFx3_ASAP7_75t_L g1826 ( 
.A(n_1821),
.Y(n_1826)
);

AND2x2_ASAP7_75t_L g1827 ( 
.A(n_1804),
.B(n_1686),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1793),
.Y(n_1828)
);

NOR2x1_ASAP7_75t_L g1829 ( 
.A(n_1807),
.B(n_1739),
.Y(n_1829)
);

BUFx2_ASAP7_75t_L g1830 ( 
.A(n_1804),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1804),
.B(n_1686),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1817),
.B(n_1687),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1777),
.B(n_1749),
.Y(n_1833)
);

INVx4_ASAP7_75t_L g1834 ( 
.A(n_1776),
.Y(n_1834)
);

INVx3_ASAP7_75t_L g1835 ( 
.A(n_1819),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1817),
.B(n_1687),
.Y(n_1836)
);

INVxp67_ASAP7_75t_SL g1837 ( 
.A(n_1815),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1820),
.B(n_1658),
.Y(n_1838)
);

INVx2_ASAP7_75t_L g1839 ( 
.A(n_1823),
.Y(n_1839)
);

AND2x2_ASAP7_75t_L g1840 ( 
.A(n_1800),
.B(n_1672),
.Y(n_1840)
);

BUFx2_ASAP7_75t_L g1841 ( 
.A(n_1818),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1823),
.Y(n_1842)
);

AOI22xp33_ASAP7_75t_L g1843 ( 
.A1(n_1772),
.A2(n_1745),
.B1(n_1747),
.B2(n_1743),
.Y(n_1843)
);

INVxp67_ASAP7_75t_L g1844 ( 
.A(n_1811),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1802),
.B(n_1672),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1791),
.B(n_1810),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1818),
.B(n_1673),
.Y(n_1847)
);

BUFx3_ASAP7_75t_L g1848 ( 
.A(n_1773),
.Y(n_1848)
);

CKINVDCx20_ASAP7_75t_R g1849 ( 
.A(n_1788),
.Y(n_1849)
);

NOR2x1_ASAP7_75t_SL g1850 ( 
.A(n_1762),
.B(n_1796),
.Y(n_1850)
);

HB1xp67_ASAP7_75t_L g1851 ( 
.A(n_1779),
.Y(n_1851)
);

AOI22xp33_ASAP7_75t_SL g1852 ( 
.A1(n_1772),
.A2(n_1731),
.B1(n_1741),
.B2(n_1691),
.Y(n_1852)
);

AOI22xp33_ASAP7_75t_L g1853 ( 
.A1(n_1762),
.A2(n_1747),
.B1(n_1743),
.B2(n_1753),
.Y(n_1853)
);

INVxp67_ASAP7_75t_SL g1854 ( 
.A(n_1796),
.Y(n_1854)
);

AND2x4_ASAP7_75t_L g1855 ( 
.A(n_1805),
.B(n_1677),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1773),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1810),
.B(n_1663),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1811),
.Y(n_1858)
);

AND2x2_ASAP7_75t_L g1859 ( 
.A(n_1790),
.B(n_1681),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1790),
.B(n_1795),
.Y(n_1860)
);

INVx1_ASAP7_75t_L g1861 ( 
.A(n_1797),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1812),
.Y(n_1862)
);

INVx2_ASAP7_75t_L g1863 ( 
.A(n_1780),
.Y(n_1863)
);

BUFx2_ASAP7_75t_L g1864 ( 
.A(n_1848),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1830),
.B(n_1841),
.Y(n_1865)
);

INVx1_ASAP7_75t_SL g1866 ( 
.A(n_1846),
.Y(n_1866)
);

INVx3_ASAP7_75t_L g1867 ( 
.A(n_1835),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1828),
.Y(n_1868)
);

NAND3xp33_ASAP7_75t_L g1869 ( 
.A(n_1844),
.B(n_1783),
.C(n_1775),
.Y(n_1869)
);

AND2x4_ASAP7_75t_SL g1870 ( 
.A(n_1834),
.B(n_1808),
.Y(n_1870)
);

CKINVDCx5p33_ASAP7_75t_R g1871 ( 
.A(n_1849),
.Y(n_1871)
);

OR2x2_ASAP7_75t_L g1872 ( 
.A(n_1830),
.B(n_1780),
.Y(n_1872)
);

AO21x2_ASAP7_75t_L g1873 ( 
.A1(n_1839),
.A2(n_1806),
.B(n_1809),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1841),
.B(n_1809),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1827),
.B(n_1799),
.Y(n_1875)
);

INVx2_ASAP7_75t_L g1876 ( 
.A(n_1839),
.Y(n_1876)
);

AOI322xp5_ASAP7_75t_L g1877 ( 
.A1(n_1860),
.A2(n_1782),
.A3(n_1765),
.B1(n_1771),
.B2(n_1781),
.C1(n_1785),
.C2(n_1767),
.Y(n_1877)
);

HB1xp67_ASAP7_75t_L g1878 ( 
.A(n_1831),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1831),
.B(n_1795),
.Y(n_1879)
);

AOI22xp33_ASAP7_75t_L g1880 ( 
.A1(n_1860),
.A2(n_1762),
.B1(n_1768),
.B2(n_1789),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1854),
.B(n_1769),
.Y(n_1881)
);

AOI22xp33_ASAP7_75t_L g1882 ( 
.A1(n_1852),
.A2(n_1789),
.B1(n_1764),
.B2(n_1782),
.Y(n_1882)
);

AO21x2_ASAP7_75t_L g1883 ( 
.A1(n_1839),
.A2(n_1646),
.B(n_1647),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1862),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1816),
.Y(n_1885)
);

AND2x2_ASAP7_75t_L g1886 ( 
.A(n_1840),
.B(n_1816),
.Y(n_1886)
);

INVxp67_ASAP7_75t_L g1887 ( 
.A(n_1862),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1842),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1889)
);

HB1xp67_ASAP7_75t_L g1890 ( 
.A(n_1847),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_L g1891 ( 
.A(n_1854),
.B(n_1822),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1848),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_SL g1893 ( 
.A1(n_1850),
.A2(n_1778),
.B(n_1794),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1847),
.Y(n_1894)
);

AOI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1838),
.A2(n_1801),
.B(n_1813),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1837),
.B(n_1786),
.Y(n_1896)
);

AND2x2_ASAP7_75t_L g1897 ( 
.A(n_1845),
.B(n_1825),
.Y(n_1897)
);

INVx5_ASAP7_75t_SL g1898 ( 
.A(n_1855),
.Y(n_1898)
);

OAI211xp5_ASAP7_75t_L g1899 ( 
.A1(n_1844),
.A2(n_1781),
.B(n_1808),
.C(n_1803),
.Y(n_1899)
);

AND2x4_ASAP7_75t_L g1900 ( 
.A(n_1856),
.B(n_1814),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1861),
.B(n_1764),
.Y(n_1901)
);

HB1xp67_ASAP7_75t_L g1902 ( 
.A(n_1838),
.Y(n_1902)
);

BUFx2_ASAP7_75t_L g1903 ( 
.A(n_1829),
.Y(n_1903)
);

HB1xp67_ASAP7_75t_L g1904 ( 
.A(n_1902),
.Y(n_1904)
);

NOR2xp33_ASAP7_75t_L g1905 ( 
.A(n_1869),
.B(n_1858),
.Y(n_1905)
);

NAND2xp5_ASAP7_75t_L g1906 ( 
.A(n_1884),
.B(n_1887),
.Y(n_1906)
);

NOR2xp33_ASAP7_75t_L g1907 ( 
.A(n_1869),
.B(n_1858),
.Y(n_1907)
);

AND2x2_ASAP7_75t_L g1908 ( 
.A(n_1878),
.B(n_1850),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1883),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1878),
.B(n_1856),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1892),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1867),
.B(n_1856),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1890),
.B(n_1856),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1868),
.Y(n_1914)
);

AND2x2_ASAP7_75t_L g1915 ( 
.A(n_1890),
.B(n_1846),
.Y(n_1915)
);

NAND2x1_ASAP7_75t_L g1916 ( 
.A(n_1903),
.B(n_1829),
.Y(n_1916)
);

BUFx3_ASAP7_75t_L g1917 ( 
.A(n_1892),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1883),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1868),
.Y(n_1919)
);

HB1xp67_ASAP7_75t_L g1920 ( 
.A(n_1902),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1894),
.B(n_1832),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1884),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1883),
.Y(n_1923)
);

AND2x2_ASAP7_75t_L g1924 ( 
.A(n_1894),
.B(n_1832),
.Y(n_1924)
);

OR2x2_ASAP7_75t_L g1925 ( 
.A(n_1865),
.B(n_1857),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1875),
.B(n_1836),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1883),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1865),
.B(n_1857),
.Y(n_1928)
);

AND2x2_ASAP7_75t_L g1929 ( 
.A(n_1875),
.B(n_1836),
.Y(n_1929)
);

INVx2_ASAP7_75t_L g1930 ( 
.A(n_1876),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1876),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1887),
.B(n_1866),
.Y(n_1932)
);

AND2x2_ASAP7_75t_L g1933 ( 
.A(n_1875),
.B(n_1859),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1866),
.B(n_1861),
.Y(n_1934)
);

BUFx2_ASAP7_75t_L g1935 ( 
.A(n_1892),
.Y(n_1935)
);

INVx2_ASAP7_75t_L g1936 ( 
.A(n_1876),
.Y(n_1936)
);

NAND2x1p5_ASAP7_75t_L g1937 ( 
.A(n_1903),
.B(n_1863),
.Y(n_1937)
);

INVxp67_ASAP7_75t_L g1938 ( 
.A(n_1901),
.Y(n_1938)
);

NAND4xp25_ASAP7_75t_L g1939 ( 
.A(n_1877),
.B(n_1852),
.C(n_1853),
.D(n_1843),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_SL g1940 ( 
.A(n_1877),
.B(n_1792),
.Y(n_1940)
);

NOR2x1_ASAP7_75t_L g1941 ( 
.A(n_1893),
.B(n_1842),
.Y(n_1941)
);

INVx2_ASAP7_75t_L g1942 ( 
.A(n_1888),
.Y(n_1942)
);

AND2x2_ASAP7_75t_L g1943 ( 
.A(n_1933),
.B(n_1900),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1922),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1905),
.B(n_1891),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1905),
.B(n_1891),
.Y(n_1946)
);

INVx3_ASAP7_75t_L g1947 ( 
.A(n_1937),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1922),
.Y(n_1948)
);

OAI21xp33_ASAP7_75t_L g1949 ( 
.A1(n_1907),
.A2(n_1882),
.B(n_1880),
.Y(n_1949)
);

INVx1_ASAP7_75t_L g1950 ( 
.A(n_1904),
.Y(n_1950)
);

NOR2xp67_ASAP7_75t_L g1951 ( 
.A(n_1911),
.B(n_1895),
.Y(n_1951)
);

AND2x2_ASAP7_75t_L g1952 ( 
.A(n_1933),
.B(n_1900),
.Y(n_1952)
);

INVx2_ASAP7_75t_SL g1953 ( 
.A(n_1917),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1932),
.B(n_1874),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1937),
.Y(n_1955)
);

AND2x2_ASAP7_75t_L g1956 ( 
.A(n_1933),
.B(n_1908),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1904),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1908),
.B(n_1921),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1907),
.B(n_1885),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1937),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1932),
.B(n_1885),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1908),
.B(n_1900),
.Y(n_1962)
);

AND2x2_ASAP7_75t_L g1963 ( 
.A(n_1921),
.B(n_1900),
.Y(n_1963)
);

BUFx3_ASAP7_75t_L g1964 ( 
.A(n_1935),
.Y(n_1964)
);

OR2x6_ASAP7_75t_L g1965 ( 
.A(n_1941),
.B(n_1911),
.Y(n_1965)
);

AND2x4_ASAP7_75t_L g1966 ( 
.A(n_1917),
.B(n_1864),
.Y(n_1966)
);

NOR2xp33_ASAP7_75t_L g1967 ( 
.A(n_1940),
.B(n_1787),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1906),
.Y(n_1968)
);

INVx1_ASAP7_75t_SL g1969 ( 
.A(n_1917),
.Y(n_1969)
);

NAND2xp5_ASAP7_75t_L g1970 ( 
.A(n_1934),
.B(n_1885),
.Y(n_1970)
);

OR2x2_ASAP7_75t_L g1971 ( 
.A(n_1925),
.B(n_1874),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1940),
.A2(n_1899),
.B(n_1895),
.Y(n_1972)
);

INVxp67_ASAP7_75t_L g1973 ( 
.A(n_1906),
.Y(n_1973)
);

AND2x2_ASAP7_75t_L g1974 ( 
.A(n_1921),
.B(n_1900),
.Y(n_1974)
);

INVx1_ASAP7_75t_SL g1975 ( 
.A(n_1917),
.Y(n_1975)
);

INVxp67_ASAP7_75t_SL g1976 ( 
.A(n_1941),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1924),
.B(n_1898),
.Y(n_1977)
);

INVx2_ASAP7_75t_L g1978 ( 
.A(n_1937),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1924),
.B(n_1898),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1920),
.Y(n_1980)
);

INVx1_ASAP7_75t_L g1981 ( 
.A(n_1920),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1914),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1934),
.B(n_1886),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1938),
.B(n_1886),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1914),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1914),
.Y(n_1986)
);

AOI21xp33_ASAP7_75t_L g1987 ( 
.A1(n_1941),
.A2(n_1899),
.B(n_1901),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1938),
.B(n_1886),
.Y(n_1988)
);

INVx2_ASAP7_75t_L g1989 ( 
.A(n_1937),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1919),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1919),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1919),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1925),
.B(n_1874),
.Y(n_1993)
);

AND2x2_ASAP7_75t_L g1994 ( 
.A(n_1924),
.B(n_1898),
.Y(n_1994)
);

INVxp67_ASAP7_75t_SL g1995 ( 
.A(n_1916),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1915),
.B(n_1889),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1996),
.B(n_1925),
.Y(n_1997)
);

OR2x2_ASAP7_75t_L g1998 ( 
.A(n_1961),
.B(n_1928),
.Y(n_1998)
);

NAND2x1p5_ASAP7_75t_L g1999 ( 
.A(n_1951),
.B(n_1916),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1977),
.B(n_1935),
.Y(n_2000)
);

NOR2xp33_ASAP7_75t_L g2001 ( 
.A(n_1967),
.B(n_1871),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1977),
.B(n_1935),
.Y(n_2002)
);

AND2x2_ASAP7_75t_L g2003 ( 
.A(n_1979),
.B(n_1911),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1944),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1979),
.B(n_1911),
.Y(n_2005)
);

INVx2_ASAP7_75t_SL g2006 ( 
.A(n_1964),
.Y(n_2006)
);

AND2x2_ASAP7_75t_L g2007 ( 
.A(n_1994),
.B(n_1915),
.Y(n_2007)
);

AND2x2_ASAP7_75t_L g2008 ( 
.A(n_1994),
.B(n_1915),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1964),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1972),
.B(n_1889),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1982),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_L g2012 ( 
.A(n_1945),
.B(n_1889),
.Y(n_2012)
);

NAND2x1_ASAP7_75t_L g2013 ( 
.A(n_1965),
.B(n_1864),
.Y(n_2013)
);

INVx1_ASAP7_75t_L g2014 ( 
.A(n_1982),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1956),
.Y(n_2015)
);

INVx2_ASAP7_75t_SL g2016 ( 
.A(n_1965),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1956),
.B(n_1926),
.Y(n_2017)
);

NAND4xp25_ASAP7_75t_L g2018 ( 
.A(n_1946),
.B(n_1939),
.C(n_1881),
.D(n_1833),
.Y(n_2018)
);

INVx2_ASAP7_75t_L g2019 ( 
.A(n_1958),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1958),
.B(n_1926),
.Y(n_2020)
);

INVx1_ASAP7_75t_L g2021 ( 
.A(n_1944),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1965),
.B(n_1913),
.Y(n_2022)
);

INVx1_ASAP7_75t_L g2023 ( 
.A(n_1985),
.Y(n_2023)
);

OR2x2_ASAP7_75t_L g2024 ( 
.A(n_1984),
.B(n_1928),
.Y(n_2024)
);

NAND2xp5_ASAP7_75t_L g2025 ( 
.A(n_1949),
.B(n_1959),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1948),
.Y(n_2026)
);

AND2x4_ASAP7_75t_L g2027 ( 
.A(n_1965),
.B(n_1913),
.Y(n_2027)
);

INVx1_ASAP7_75t_L g2028 ( 
.A(n_1985),
.Y(n_2028)
);

HB1xp67_ASAP7_75t_L g2029 ( 
.A(n_1950),
.Y(n_2029)
);

INVx1_ASAP7_75t_L g2030 ( 
.A(n_1986),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1986),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_L g2032 ( 
.A(n_1973),
.B(n_1897),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1990),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1966),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_L g2035 ( 
.A(n_1968),
.B(n_1897),
.Y(n_2035)
);

NOR2xp33_ASAP7_75t_L g2036 ( 
.A(n_1987),
.B(n_1774),
.Y(n_2036)
);

OAI22xp33_ASAP7_75t_L g2037 ( 
.A1(n_2010),
.A2(n_1939),
.B1(n_1976),
.B2(n_1865),
.Y(n_2037)
);

AOI32xp33_ASAP7_75t_L g2038 ( 
.A1(n_2025),
.A2(n_1975),
.A3(n_1969),
.B1(n_1948),
.B2(n_1995),
.Y(n_2038)
);

AOI32xp33_ASAP7_75t_L g2039 ( 
.A1(n_2036),
.A2(n_1966),
.A3(n_1953),
.B1(n_1988),
.B2(n_1943),
.Y(n_2039)
);

INVx1_ASAP7_75t_SL g2040 ( 
.A(n_2000),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_2034),
.Y(n_2041)
);

AND2x2_ASAP7_75t_L g2042 ( 
.A(n_2000),
.B(n_1966),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_2009),
.B(n_1953),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_2009),
.B(n_1970),
.Y(n_2044)
);

INVx1_ASAP7_75t_L g2045 ( 
.A(n_2011),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_2011),
.Y(n_2046)
);

INVx1_ASAP7_75t_SL g2047 ( 
.A(n_2002),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_2006),
.B(n_1983),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_2006),
.B(n_1980),
.Y(n_2049)
);

OAI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2018),
.A2(n_2013),
.B1(n_1999),
.B2(n_2012),
.Y(n_2050)
);

OAI21xp5_ASAP7_75t_L g2051 ( 
.A1(n_2013),
.A2(n_1981),
.B(n_1957),
.Y(n_2051)
);

NOR2xp67_ASAP7_75t_L g2052 ( 
.A(n_2034),
.B(n_1947),
.Y(n_2052)
);

AOI22xp5_ASAP7_75t_L g2053 ( 
.A1(n_2002),
.A2(n_1792),
.B1(n_1950),
.B2(n_1957),
.Y(n_2053)
);

NAND3xp33_ASAP7_75t_L g2054 ( 
.A(n_2029),
.B(n_2016),
.C(n_2004),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_2022),
.Y(n_2055)
);

AOI22xp5_ASAP7_75t_SL g2056 ( 
.A1(n_2016),
.A2(n_1955),
.B1(n_1947),
.B2(n_1774),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_2014),
.Y(n_2057)
);

INVx1_ASAP7_75t_SL g2058 ( 
.A(n_2003),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_2001),
.A2(n_1916),
.B(n_1881),
.Y(n_2059)
);

AND2x2_ASAP7_75t_L g2060 ( 
.A(n_2003),
.B(n_1943),
.Y(n_2060)
);

INVx1_ASAP7_75t_SL g2061 ( 
.A(n_2005),
.Y(n_2061)
);

AOI21xp5_ASAP7_75t_L g2062 ( 
.A1(n_1999),
.A2(n_1954),
.B(n_1947),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_2014),
.Y(n_2063)
);

AND2x2_ASAP7_75t_L g2064 ( 
.A(n_2005),
.B(n_1952),
.Y(n_2064)
);

OR2x2_ASAP7_75t_L g2065 ( 
.A(n_2032),
.B(n_1954),
.Y(n_2065)
);

OAI322xp33_ASAP7_75t_L g2066 ( 
.A1(n_2037),
.A2(n_2021),
.A3(n_2026),
.B1(n_1999),
.B2(n_2019),
.C1(n_2015),
.C2(n_2024),
.Y(n_2066)
);

OAI21xp5_ASAP7_75t_L g2067 ( 
.A1(n_2037),
.A2(n_2027),
.B(n_2022),
.Y(n_2067)
);

INVx1_ASAP7_75t_L g2068 ( 
.A(n_2045),
.Y(n_2068)
);

INVxp33_ASAP7_75t_L g2069 ( 
.A(n_2056),
.Y(n_2069)
);

AO22x1_ASAP7_75t_L g2070 ( 
.A1(n_2051),
.A2(n_2027),
.B1(n_2022),
.B2(n_2007),
.Y(n_2070)
);

AOI22xp5_ASAP7_75t_L g2071 ( 
.A1(n_2050),
.A2(n_2008),
.B1(n_2007),
.B2(n_2019),
.Y(n_2071)
);

OAI211xp5_ASAP7_75t_L g2072 ( 
.A1(n_2038),
.A2(n_2008),
.B(n_2015),
.C(n_2024),
.Y(n_2072)
);

AOI22xp5_ASAP7_75t_L g2073 ( 
.A1(n_2050),
.A2(n_2035),
.B1(n_2027),
.B2(n_2020),
.Y(n_2073)
);

AND2x2_ASAP7_75t_L g2074 ( 
.A(n_2042),
.B(n_2020),
.Y(n_2074)
);

INVx1_ASAP7_75t_L g2075 ( 
.A(n_2046),
.Y(n_2075)
);

INVx2_ASAP7_75t_L g2076 ( 
.A(n_2042),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2057),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_L g2078 ( 
.A(n_2040),
.B(n_2017),
.Y(n_2078)
);

BUFx2_ASAP7_75t_L g2079 ( 
.A(n_2041),
.Y(n_2079)
);

AOI222xp33_ASAP7_75t_L g2080 ( 
.A1(n_2054),
.A2(n_2017),
.B1(n_1879),
.B2(n_2030),
.C1(n_2028),
.C2(n_2023),
.Y(n_2080)
);

NOR3xp33_ASAP7_75t_L g2081 ( 
.A(n_2043),
.B(n_1955),
.C(n_2023),
.Y(n_2081)
);

INVx2_ASAP7_75t_L g2082 ( 
.A(n_2060),
.Y(n_2082)
);

INVx1_ASAP7_75t_L g2083 ( 
.A(n_2063),
.Y(n_2083)
);

OAI22xp33_ASAP7_75t_L g2084 ( 
.A1(n_2053),
.A2(n_2047),
.B1(n_2061),
.B2(n_2058),
.Y(n_2084)
);

O2A1O1Ixp33_ASAP7_75t_L g2085 ( 
.A1(n_2049),
.A2(n_1955),
.B(n_2031),
.C(n_2030),
.Y(n_2085)
);

OAI22xp33_ASAP7_75t_SL g2086 ( 
.A1(n_2055),
.A2(n_1784),
.B1(n_1997),
.B2(n_1998),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_L g2087 ( 
.A(n_2041),
.B(n_1997),
.Y(n_2087)
);

INVxp33_ASAP7_75t_L g2088 ( 
.A(n_2052),
.Y(n_2088)
);

OAI31xp33_ASAP7_75t_L g2089 ( 
.A1(n_2084),
.A2(n_2059),
.A3(n_2062),
.B(n_2055),
.Y(n_2089)
);

O2A1O1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_2066),
.A2(n_2084),
.B(n_2067),
.C(n_2069),
.Y(n_2090)
);

AND2x2_ASAP7_75t_L g2091 ( 
.A(n_2074),
.B(n_2060),
.Y(n_2091)
);

NAND3xp33_ASAP7_75t_L g2092 ( 
.A(n_2080),
.B(n_2039),
.C(n_2048),
.Y(n_2092)
);

AOI21xp33_ASAP7_75t_L g2093 ( 
.A1(n_2069),
.A2(n_2044),
.B(n_2065),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_L g2094 ( 
.A(n_2076),
.B(n_2064),
.Y(n_2094)
);

NAND2xp5_ASAP7_75t_L g2095 ( 
.A(n_2079),
.B(n_2064),
.Y(n_2095)
);

AOI22xp5_ASAP7_75t_L g2096 ( 
.A1(n_2071),
.A2(n_2073),
.B1(n_2072),
.B2(n_2082),
.Y(n_2096)
);

OAI21xp33_ASAP7_75t_L g2097 ( 
.A1(n_2086),
.A2(n_1998),
.B(n_2033),
.Y(n_2097)
);

INVxp67_ASAP7_75t_L g2098 ( 
.A(n_2087),
.Y(n_2098)
);

AOI22xp5_ASAP7_75t_L g2099 ( 
.A1(n_2078),
.A2(n_2033),
.B1(n_2031),
.B2(n_2028),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2068),
.Y(n_2100)
);

INVx1_ASAP7_75t_L g2101 ( 
.A(n_2075),
.Y(n_2101)
);

OR2x2_ASAP7_75t_L g2102 ( 
.A(n_2070),
.B(n_1971),
.Y(n_2102)
);

INVx1_ASAP7_75t_L g2103 ( 
.A(n_2077),
.Y(n_2103)
);

OAI21xp5_ASAP7_75t_SL g2104 ( 
.A1(n_2088),
.A2(n_1763),
.B(n_1971),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_2089),
.B(n_2088),
.Y(n_2105)
);

OAI211xp5_ASAP7_75t_SL g2106 ( 
.A1(n_2090),
.A2(n_2085),
.B(n_2083),
.C(n_2081),
.Y(n_2106)
);

NAND2xp33_ASAP7_75t_R g2107 ( 
.A(n_2095),
.B(n_1993),
.Y(n_2107)
);

NOR3x1_ASAP7_75t_L g2108 ( 
.A(n_2092),
.B(n_1993),
.C(n_1991),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2094),
.Y(n_2109)
);

NOR3xp33_ASAP7_75t_L g2110 ( 
.A(n_2098),
.B(n_2081),
.C(n_1978),
.Y(n_2110)
);

NOR2x1_ASAP7_75t_L g2111 ( 
.A(n_2100),
.B(n_1960),
.Y(n_2111)
);

AOI221xp5_ASAP7_75t_L g2112 ( 
.A1(n_2093),
.A2(n_1989),
.B1(n_1978),
.B2(n_1960),
.C(n_1992),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_2102),
.B(n_1989),
.Y(n_2113)
);

OR2x2_ASAP7_75t_L g2114 ( 
.A(n_2091),
.B(n_1928),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_2101),
.Y(n_2115)
);

NOR3xp33_ASAP7_75t_L g2116 ( 
.A(n_2097),
.B(n_2104),
.C(n_2103),
.Y(n_2116)
);

INVx1_ASAP7_75t_L g2117 ( 
.A(n_2099),
.Y(n_2117)
);

AOI322xp5_ASAP7_75t_L g2118 ( 
.A1(n_2116),
.A2(n_2096),
.A3(n_1879),
.B1(n_2104),
.B2(n_1929),
.C1(n_1926),
.C2(n_1913),
.Y(n_2118)
);

AOI211xp5_ASAP7_75t_L g2119 ( 
.A1(n_2106),
.A2(n_1962),
.B(n_1798),
.C(n_1952),
.Y(n_2119)
);

INVx2_ASAP7_75t_L g2120 ( 
.A(n_2114),
.Y(n_2120)
);

NOR4xp25_ASAP7_75t_L g2121 ( 
.A(n_2105),
.B(n_1992),
.C(n_1991),
.D(n_1990),
.Y(n_2121)
);

AOI221xp5_ASAP7_75t_L g2122 ( 
.A1(n_2117),
.A2(n_1963),
.B1(n_1974),
.B2(n_1927),
.C(n_1923),
.Y(n_2122)
);

OAI21xp33_ASAP7_75t_L g2123 ( 
.A1(n_2113),
.A2(n_1962),
.B(n_1963),
.Y(n_2123)
);

AOI221xp5_ASAP7_75t_L g2124 ( 
.A1(n_2110),
.A2(n_1974),
.B1(n_1918),
.B2(n_1909),
.C(n_1923),
.Y(n_2124)
);

O2A1O1Ixp33_ASAP7_75t_L g2125 ( 
.A1(n_2115),
.A2(n_1872),
.B(n_1910),
.C(n_1909),
.Y(n_2125)
);

AOI22xp33_ASAP7_75t_L g2126 ( 
.A1(n_2120),
.A2(n_2109),
.B1(n_2112),
.B2(n_2111),
.Y(n_2126)
);

OAI22xp5_ASAP7_75t_L g2127 ( 
.A1(n_2119),
.A2(n_2108),
.B1(n_2107),
.B2(n_1912),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2121),
.A2(n_1918),
.B1(n_1909),
.B2(n_1923),
.C(n_1927),
.Y(n_2128)
);

AOI21xp5_ASAP7_75t_L g2129 ( 
.A1(n_2125),
.A2(n_1912),
.B(n_1910),
.Y(n_2129)
);

AOI22xp33_ASAP7_75t_L g2130 ( 
.A1(n_2123),
.A2(n_1873),
.B1(n_1826),
.B2(n_1870),
.Y(n_2130)
);

O2A1O1Ixp33_ASAP7_75t_L g2131 ( 
.A1(n_2122),
.A2(n_2124),
.B(n_2118),
.C(n_1910),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_2120),
.A2(n_1912),
.B1(n_1851),
.B2(n_1896),
.Y(n_2132)
);

HB1xp67_ASAP7_75t_L g2133 ( 
.A(n_2120),
.Y(n_2133)
);

NAND2xp5_ASAP7_75t_L g2134 ( 
.A(n_2133),
.B(n_1929),
.Y(n_2134)
);

XOR2xp5_ASAP7_75t_L g2135 ( 
.A(n_2126),
.B(n_1766),
.Y(n_2135)
);

OR2x2_ASAP7_75t_L g2136 ( 
.A(n_2127),
.B(n_1929),
.Y(n_2136)
);

XNOR2xp5_ASAP7_75t_L g2137 ( 
.A(n_2132),
.B(n_2130),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_2129),
.Y(n_2138)
);

NOR2x1_ASAP7_75t_L g2139 ( 
.A(n_2131),
.B(n_1912),
.Y(n_2139)
);

OAI211xp5_ASAP7_75t_SL g2140 ( 
.A1(n_2138),
.A2(n_2128),
.B(n_1824),
.C(n_1896),
.Y(n_2140)
);

OR3x2_ASAP7_75t_L g2141 ( 
.A(n_2136),
.B(n_1756),
.C(n_1872),
.Y(n_2141)
);

INVxp67_ASAP7_75t_L g2142 ( 
.A(n_2135),
.Y(n_2142)
);

NOR2xp67_ASAP7_75t_L g2143 ( 
.A(n_2134),
.B(n_1912),
.Y(n_2143)
);

OR2x2_ASAP7_75t_L g2144 ( 
.A(n_2142),
.B(n_2137),
.Y(n_2144)
);

AND2x4_ASAP7_75t_L g2145 ( 
.A(n_2143),
.B(n_2139),
.Y(n_2145)
);

OAI22xp33_ASAP7_75t_SL g2146 ( 
.A1(n_2144),
.A2(n_2141),
.B1(n_2140),
.B2(n_1912),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2146),
.A2(n_2145),
.B1(n_1931),
.B2(n_1942),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2146),
.B(n_1930),
.Y(n_2148)
);

INVx1_ASAP7_75t_L g2149 ( 
.A(n_2148),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2147),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_SL g2151 ( 
.A1(n_2150),
.A2(n_1702),
.B1(n_1698),
.B2(n_1674),
.Y(n_2151)
);

INVxp67_ASAP7_75t_SL g2152 ( 
.A(n_2149),
.Y(n_2152)
);

OAI21xp5_ASAP7_75t_L g2153 ( 
.A1(n_2152),
.A2(n_1770),
.B(n_1766),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_2153),
.B(n_2151),
.Y(n_2154)
);

OAI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_2154),
.A2(n_1936),
.B1(n_1942),
.B2(n_1931),
.Y(n_2155)
);

AOI221xp5_ASAP7_75t_L g2156 ( 
.A1(n_2155),
.A2(n_1936),
.B1(n_1942),
.B2(n_1931),
.C(n_1930),
.Y(n_2156)
);

AOI211xp5_ASAP7_75t_L g2157 ( 
.A1(n_2156),
.A2(n_1702),
.B(n_1698),
.C(n_1770),
.Y(n_2157)
);


endmodule