module fake_jpeg_12192_n_193 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_193);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_193;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx6_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_3),
.B(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_15),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_7),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx13_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_25),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_47),
.Y(n_60)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_41),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_25),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_42),
.B(n_43),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_23),
.B(n_14),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

OR2x2_ASAP7_75t_L g45 ( 
.A(n_27),
.B(n_31),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_45),
.B(n_49),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_21),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_17),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_21),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_42),
.A2(n_16),
.B1(n_19),
.B2(n_21),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_53),
.A2(n_16),
.B1(n_18),
.B2(n_32),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_62),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_30),
.Y(n_63)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_26),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_67),
.B(n_71),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g68 ( 
.A(n_35),
.B(n_29),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_31),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_69),
.B(n_0),
.Y(n_90)
);

A2O1A1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_37),
.A2(n_34),
.B(n_24),
.C(n_29),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_52),
.A2(n_18),
.B1(n_16),
.B2(n_32),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_72),
.A2(n_20),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_44),
.B(n_30),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_50),
.A2(n_46),
.B1(n_39),
.B2(n_51),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_78),
.A2(n_20),
.B1(n_1),
.B2(n_2),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_26),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_58),
.Y(n_104)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_58),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_80),
.Y(n_121)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_82),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_83),
.B(n_87),
.Y(n_115)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_66),
.A2(n_41),
.B1(n_40),
.B2(n_34),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_84),
.A2(n_94),
.B1(n_70),
.B2(n_61),
.Y(n_107)
);

INVx5_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_69),
.A2(n_24),
.B1(n_20),
.B2(n_17),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_88),
.B(n_100),
.Y(n_119)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_90),
.B(n_105),
.Y(n_110)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

AOI21xp33_ASAP7_75t_L g93 ( 
.A1(n_56),
.A2(n_1),
.B(n_4),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_93),
.B(n_77),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_75),
.A2(n_20),
.B1(n_5),
.B2(n_6),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_96),
.A2(n_97),
.B(n_103),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_68),
.A2(n_4),
.B(n_5),
.Y(n_97)
);

BUFx6f_ASAP7_75t_SL g98 ( 
.A(n_64),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_98),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_60),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_99),
.B(n_77),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_55),
.A2(n_6),
.B1(n_9),
.B2(n_11),
.Y(n_100)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_104),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_59),
.A2(n_12),
.B(n_13),
.Y(n_103)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_61),
.C(n_73),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g142 ( 
.A(n_106),
.B(n_105),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_107),
.A2(n_100),
.B1(n_92),
.B2(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_81),
.B(n_73),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_111),
.B(n_113),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_71),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_116),
.B(n_87),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g122 ( 
.A(n_95),
.B(n_64),
.C(n_54),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_122),
.B(n_123),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_95),
.A2(n_54),
.B(n_76),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_126),
.A2(n_96),
.B(n_80),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_103),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_127),
.B(n_131),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_128),
.B(n_138),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_101),
.Y(n_131)
);

FAx1_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_83),
.CI(n_98),
.CON(n_132),
.SN(n_132)
);

A2O1A1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_132),
.A2(n_115),
.B(n_119),
.C(n_117),
.Y(n_154)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_109),
.Y(n_133)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_133),
.Y(n_156)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_112),
.Y(n_134)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_134),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_137),
.B(n_143),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_110),
.B(n_99),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_82),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_140),
.Y(n_146)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_106),
.C(n_126),
.Y(n_149)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_118),
.Y(n_143)
);

A2O1A1O1Ixp25_ASAP7_75t_L g147 ( 
.A1(n_139),
.A2(n_129),
.B(n_128),
.C(n_136),
.D(n_138),
.Y(n_147)
);

AOI21xp33_ASAP7_75t_L g159 ( 
.A1(n_147),
.A2(n_151),
.B(n_132),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_149),
.B(n_152),
.C(n_143),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_114),
.B(n_124),
.C(n_123),
.D(n_115),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_142),
.B(n_124),
.C(n_118),
.Y(n_152)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_154),
.Y(n_160)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_153),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_158),
.A2(n_162),
.B1(n_163),
.B2(n_164),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_159),
.B(n_161),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_147),
.B(n_137),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_150),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_145),
.A2(n_132),
.A3(n_130),
.B1(n_134),
.B2(n_135),
.C(n_119),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_155),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_117),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_166),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_145),
.B(n_146),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_168),
.C(n_152),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_149),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_170),
.C(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_148),
.C(n_146),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_167),
.B(n_148),
.C(n_157),
.Y(n_171)
);

AOI321xp33_ASAP7_75t_L g172 ( 
.A1(n_160),
.A2(n_151),
.A3(n_154),
.B1(n_115),
.B2(n_120),
.C(n_119),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_172),
.B(n_133),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_160),
.B(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_162),
.C(n_156),
.Y(n_180)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_175),
.Y(n_177)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_177),
.Y(n_184)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_174),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_179),
.A2(n_102),
.B1(n_125),
.B2(n_86),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_181),
.B(n_182),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_170),
.A2(n_156),
.B(n_109),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_178),
.A2(n_173),
.B(n_176),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_185),
.B(n_178),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_186),
.A2(n_182),
.B1(n_180),
.B2(n_179),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_187),
.B(n_188),
.Y(n_190)
);

AOI321xp33_ASAP7_75t_L g189 ( 
.A1(n_184),
.A2(n_85),
.A3(n_89),
.B1(n_125),
.B2(n_177),
.C(n_183),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_189),
.B(n_85),
.C(n_121),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_191),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_190),
.Y(n_193)
);


endmodule