module fake_aes_5369_n_825 (n_52, n_50, n_7, n_3, n_34, n_25, n_9, n_96, n_72, n_77, n_90, n_99, n_43, n_73, n_62, n_97, n_33, n_4, n_59, n_76, n_6, n_74, n_8, n_61, n_44, n_66, n_88, n_46, n_37, n_18, n_65, n_87, n_5, n_81, n_85, n_47, n_1, n_16, n_78, n_95, n_40, n_68, n_36, n_11, n_15, n_71, n_70, n_94, n_2, n_17, n_58, n_20, n_84, n_12, n_56, n_80, n_67, n_22, n_19, n_26, n_39, n_98, n_38, n_100, n_24, n_35, n_91, n_32, n_93, n_48, n_63, n_54, n_41, n_55, n_29, n_60, n_10, n_30, n_13, n_92, n_75, n_82, n_53, n_64, n_69, n_83, n_23, n_0, n_57, n_51, n_45, n_42, n_21, n_86, n_27, n_89, n_28, n_79, n_49, n_14, n_31, n_825, n_804);
input n_52;
input n_50;
input n_7;
input n_3;
input n_34;
input n_25;
input n_9;
input n_96;
input n_72;
input n_77;
input n_90;
input n_99;
input n_43;
input n_73;
input n_62;
input n_97;
input n_33;
input n_4;
input n_59;
input n_76;
input n_6;
input n_74;
input n_8;
input n_61;
input n_44;
input n_66;
input n_88;
input n_46;
input n_37;
input n_18;
input n_65;
input n_87;
input n_5;
input n_81;
input n_85;
input n_47;
input n_1;
input n_16;
input n_78;
input n_95;
input n_40;
input n_68;
input n_36;
input n_11;
input n_15;
input n_71;
input n_70;
input n_94;
input n_2;
input n_17;
input n_58;
input n_20;
input n_84;
input n_12;
input n_56;
input n_80;
input n_67;
input n_22;
input n_19;
input n_26;
input n_39;
input n_98;
input n_38;
input n_100;
input n_24;
input n_35;
input n_91;
input n_32;
input n_93;
input n_48;
input n_63;
input n_54;
input n_41;
input n_55;
input n_29;
input n_60;
input n_10;
input n_30;
input n_13;
input n_92;
input n_75;
input n_82;
input n_53;
input n_64;
input n_69;
input n_83;
input n_23;
input n_0;
input n_57;
input n_51;
input n_45;
input n_42;
input n_21;
input n_86;
input n_27;
input n_89;
input n_28;
input n_79;
input n_49;
input n_14;
input n_31;
output n_825;
output n_804;
wire n_107;
wire n_646;
wire n_759;
wire n_658;
wire n_673;
wire n_156;
wire n_154;
wire n_239;
wire n_7;
wire n_309;
wire n_356;
wire n_327;
wire n_25;
wire n_204;
wire n_592;
wire n_769;
wire n_169;
wire n_370;
wire n_384;
wire n_439;
wire n_545;
wire n_180;
wire n_604;
wire n_99;
wire n_43;
wire n_73;
wire n_440;
wire n_199;
wire n_279;
wire n_786;
wire n_357;
wire n_74;
wire n_729;
wire n_308;
wire n_518;
wire n_394;
wire n_44;
wire n_189;
wire n_681;
wire n_226;
wire n_352;
wire n_447;
wire n_66;
wire n_379;
wire n_535;
wire n_689;
wire n_595;
wire n_626;
wire n_316;
wire n_285;
wire n_564;
wire n_586;
wire n_471;
wire n_47;
wire n_766;
wire n_475;
wire n_744;
wire n_281;
wire n_645;
wire n_497;
wire n_399;
wire n_11;
wire n_295;
wire n_371;
wire n_579;
wire n_516;
wire n_608;
wire n_368;
wire n_805;
wire n_373;
wire n_139;
wire n_342;
wire n_151;
wire n_71;
wire n_288;
wire n_557;
wire n_176;
wire n_753;
wire n_436;
wire n_438;
wire n_359;
wire n_195;
wire n_300;
wire n_487;
wire n_461;
wire n_723;
wire n_223;
wire n_405;
wire n_562;
wire n_19;
wire n_409;
wire n_482;
wire n_534;
wire n_569;
wire n_707;
wire n_526;
wire n_261;
wire n_483;
wire n_423;
wire n_220;
wire n_353;
wire n_410;
wire n_104;
wire n_709;
wire n_303;
wire n_502;
wire n_821;
wire n_468;
wire n_159;
wire n_566;
wire n_91;
wire n_301;
wire n_340;
wire n_148;
wire n_149;
wire n_567;
wire n_378;
wire n_752;
wire n_246;
wire n_676;
wire n_823;
wire n_191;
wire n_143;
wire n_780;
wire n_629;
wire n_446;
wire n_63;
wire n_402;
wire n_54;
wire n_387;
wire n_125;
wire n_145;
wire n_166;
wire n_558;
wire n_596;
wire n_492;
wire n_181;
wire n_123;
wire n_219;
wire n_343;
wire n_494;
wire n_553;
wire n_555;
wire n_135;
wire n_481;
wire n_621;
wire n_817;
wire n_776;
wire n_315;
wire n_397;
wire n_53;
wire n_213;
wire n_196;
wire n_293;
wire n_797;
wire n_127;
wire n_312;
wire n_742;
wire n_424;
wire n_23;
wire n_110;
wire n_182;
wire n_269;
wire n_663;
wire n_529;
wire n_656;
wire n_751;
wire n_186;
wire n_137;
wire n_507;
wire n_334;
wire n_164;
wire n_433;
wire n_660;
wire n_120;
wire n_392;
wire n_650;
wire n_806;
wire n_155;
wire n_162;
wire n_114;
wire n_772;
wire n_50;
wire n_789;
wire n_816;
wire n_3;
wire n_331;
wire n_651;
wire n_574;
wire n_636;
wire n_330;
wire n_614;
wire n_231;
wire n_9;
wire n_737;
wire n_428;
wire n_178;
wire n_478;
wire n_814;
wire n_652;
wire n_678;
wire n_708;
wire n_229;
wire n_97;
wire n_133;
wire n_324;
wire n_442;
wire n_422;
wire n_192;
wire n_699;
wire n_329;
wire n_6;
wire n_8;
wire n_578;
wire n_187;
wire n_548;
wire n_188;
wire n_443;
wire n_304;
wire n_18;
wire n_682;
wire n_801;
wire n_441;
wire n_628;
wire n_425;
wire n_314;
wire n_824;
wire n_601;
wire n_307;
wire n_517;
wire n_215;
wire n_736;
wire n_172;
wire n_109;
wire n_332;
wire n_198;
wire n_386;
wire n_653;
wire n_351;
wire n_1;
wire n_16;
wire n_670;
wire n_95;
wire n_40;
wire n_210;
wire n_426;
wire n_755;
wire n_716;
wire n_228;
wire n_671;
wire n_278;
wire n_115;
wire n_270;
wire n_476;
wire n_765;
wire n_599;
wire n_715;
wire n_179;
wire n_289;
wire n_404;
wire n_366;
wire n_721;
wire n_362;
wire n_617;
wire n_688;
wire n_485;
wire n_396;
wire n_549;
wire n_354;
wire n_720;
wire n_152;
wire n_70;
wire n_588;
wire n_458;
wire n_375;
wire n_17;
wire n_322;
wire n_317;
wire n_221;
wire n_328;
wire n_506;
wire n_711;
wire n_491;
wire n_800;
wire n_388;
wire n_773;
wire n_266;
wire n_763;
wire n_80;
wire n_632;
wire n_793;
wire n_679;
wire n_522;
wire n_546;
wire n_684;
wire n_615;
wire n_701;
wire n_326;
wire n_532;
wire n_756;
wire n_635;
wire n_544;
wire n_576;
wire n_275;
wire n_691;
wire n_661;
wire n_622;
wire n_493;
wire n_274;
wire n_150;
wire n_235;
wire n_690;
wire n_38;
wire n_533;
wire n_272;
wire n_686;
wire n_299;
wire n_100;
wire n_561;
wire n_581;
wire n_280;
wire n_141;
wire n_509;
wire n_160;
wire n_499;
wire n_377;
wire n_263;
wire n_757;
wire n_695;
wire n_193;
wire n_232;
wire n_344;
wire n_783;
wire n_812;
wire n_147;
wire n_185;
wire n_367;
wire n_795;
wire n_267;
wire n_687;
wire n_171;
wire n_638;
wire n_450;
wire n_585;
wire n_140;
wire n_644;
wire n_111;
wire n_746;
wire n_212;
wire n_779;
wire n_30;
wire n_634;
wire n_13;
wire n_254;
wire n_559;
wire n_704;
wire n_435;
wire n_728;
wire n_583;
wire n_64;
wire n_69;
wire n_248;
wire n_407;
wire n_527;
wire n_83;
wire n_200;
wire n_603;
wire n_262;
wire n_119;
wire n_667;
wire n_503;
wire n_339;
wire n_347;
wire n_124;
wire n_696;
wire n_748;
wire n_79;
wire n_129;
wire n_611;
wire n_521;
wire n_157;
wire n_774;
wire n_103;
wire n_808;
wire n_421;
wire n_52;
wire n_253;
wire n_434;
wire n_677;
wire n_624;
wire n_273;
wire n_325;
wire n_571;
wire n_524;
wire n_692;
wire n_530;
wire n_743;
wire n_163;
wire n_348;
wire n_96;
wire n_669;
wire n_685;
wire n_72;
wire n_77;
wire n_762;
wire n_594;
wire n_787;
wire n_214;
wire n_90;
wire n_770;
wire n_167;
wire n_809;
wire n_364;
wire n_33;
wire n_464;
wire n_76;
wire n_470;
wire n_590;
wire n_61;
wire n_463;
wire n_216;
wire n_153;
wire n_355;
wire n_609;
wire n_121;
wire n_286;
wire n_408;
wire n_247;
wire n_431;
wire n_161;
wire n_224;
wire n_484;
wire n_165;
wire n_413;
wire n_65;
wire n_537;
wire n_710;
wire n_525;
wire n_560;
wire n_5;
wire n_496;
wire n_393;
wire n_211;
wire n_85;
wire n_320;
wire n_264;
wire n_102;
wire n_283;
wire n_733;
wire n_290;
wire n_217;
wire n_201;
wire n_791;
wire n_277;
wire n_259;
wire n_612;
wire n_244;
wire n_666;
wire n_771;
wire n_276;
wire n_297;
wire n_225;
wire n_631;
wire n_350;
wire n_747;
wire n_208;
wire n_616;
wire n_815;
wire n_523;
wire n_528;
wire n_419;
wire n_252;
wire n_519;
wire n_168;
wire n_271;
wire n_693;
wire n_785;
wire n_739;
wire n_94;
wire n_194;
wire n_758;
wire n_282;
wire n_58;
wire n_775;
wire n_113;
wire n_242;
wire n_498;
wire n_501;
wire n_284;
wire n_321;
wire n_302;
wire n_538;
wire n_703;
wire n_811;
wire n_116;
wire n_734;
wire n_292;
wire n_547;
wire n_593;
wire n_118;
wire n_587;
wire n_233;
wire n_554;
wire n_597;
wire n_698;
wire n_705;
wire n_257;
wire n_741;
wire n_722;
wire n_203;
wire n_26;
wire n_477;
wire n_460;
wire n_243;
wire n_318;
wire n_346;
wire n_98;
wire n_345;
wire n_230;
wire n_452;
wire n_714;
wire n_146;
wire n_337;
wire n_32;
wire n_637;
wire n_641;
wire n_726;
wire n_531;
wire n_539;
wire n_93;
wire n_406;
wire n_372;
wire n_820;
wire n_713;
wire n_467;
wire n_702;
wire n_41;
wire n_760;
wire n_623;
wire n_417;
wire n_451;
wire n_665;
wire n_647;
wire n_445;
wire n_500;
wire n_732;
wire n_575;
wire n_10;
wire n_390;
wire n_600;
wire n_818;
wire n_75;
wire n_82;
wire n_183;
wire n_731;
wire n_550;
wire n_132;
wire n_643;
wire n_761;
wire n_778;
wire n_582;
wire n_784;
wire n_170;
wire n_205;
wire n_158;
wire n_126;
wire n_473;
wire n_249;
wire n_389;
wire n_510;
wire n_360;
wire n_363;
wire n_749;
wire n_427;
wire n_724;
wire n_106;
wire n_296;
wire n_605;
wire n_42;
wire n_21;
wire n_437;
wire n_620;
wire n_89;
wire n_480;
wire n_130;
wire n_341;
wire n_310;
wire n_700;
wire n_640;
wire n_14;
wire n_236;
wire n_639;
wire n_727;
wire n_136;
wire n_260;
wire n_580;
wire n_610;
wire n_222;
wire n_657;
wire n_822;
wire n_381;
wire n_34;
wire n_142;
wire n_754;
wire n_385;
wire n_798;
wire n_227;
wire n_395;
wire n_454;
wire n_453;
wire n_250;
wire n_551;
wire n_268;
wire n_190;
wire n_606;
wire n_62;
wire n_712;
wire n_777;
wire n_4;
wire n_59;
wire n_323;
wire n_565;
wire n_781;
wire n_376;
wire n_694;
wire n_240;
wire n_459;
wire n_768;
wire n_568;
wire n_807;
wire n_46;
wire n_174;
wire n_717;
wire n_88;
wire n_108;
wire n_335;
wire n_37;
wire n_122;
wire n_374;
wire n_613;
wire n_380;
wire n_515;
wire n_802;
wire n_672;
wire n_466;
wire n_87;
wire n_207;
wire n_197;
wire n_81;
wire n_541;
wire n_572;
wire n_298;
wire n_112;
wire n_630;
wire n_735;
wire n_649;
wire n_602;
wire n_78;
wire n_552;
wire n_68;
wire n_444;
wire n_105;
wire n_251;
wire n_598;
wire n_810;
wire n_416;
wire n_36;
wire n_432;
wire n_465;
wire n_414;
wire n_680;
wire n_730;
wire n_369;
wire n_469;
wire n_361;
wire n_767;
wire n_237;
wire n_654;
wire n_15;
wire n_520;
wire n_633;
wire n_429;
wire n_803;
wire n_256;
wire n_398;
wire n_668;
wire n_117;
wire n_238;
wire n_365;
wire n_577;
wire n_804;
wire n_796;
wire n_294;
wire n_2;
wire n_338;
wire n_662;
wire n_591;
wire n_391;
wire n_241;
wire n_209;
wire n_20;
wire n_84;
wire n_782;
wire n_449;
wire n_12;
wire n_56;
wire n_412;
wire n_455;
wire n_67;
wire n_504;
wire n_618;
wire n_790;
wire n_456;
wire n_22;
wire n_683;
wire n_479;
wire n_584;
wire n_311;
wire n_401;
wire n_383;
wire n_813;
wire n_202;
wire n_319;
wire n_542;
wire n_725;
wire n_819;
wire n_39;
wire n_101;
wire n_291;
wire n_489;
wire n_245;
wire n_664;
wire n_508;
wire n_764;
wire n_719;
wire n_486;
wire n_788;
wire n_24;
wire n_35;
wire n_655;
wire n_490;
wire n_472;
wire n_540;
wire n_400;
wire n_794;
wire n_457;
wire n_659;
wire n_134;
wire n_48;
wire n_255;
wire n_563;
wire n_513;
wire n_55;
wire n_718;
wire n_543;
wire n_336;
wire n_29;
wire n_218;
wire n_173;
wire n_488;
wire n_556;
wire n_648;
wire n_382;
wire n_799;
wire n_138;
wire n_60;
wire n_462;
wire n_536;
wire n_573;
wire n_474;
wire n_745;
wire n_305;
wire n_495;
wire n_430;
wire n_418;
wire n_505;
wire n_92;
wire n_313;
wire n_358;
wire n_333;
wire n_627;
wire n_706;
wire n_740;
wire n_589;
wire n_750;
wire n_175;
wire n_128;
wire n_306;
wire n_31;
wire n_415;
wire n_697;
wire n_0;
wire n_512;
wire n_258;
wire n_619;
wire n_675;
wire n_642;
wire n_234;
wire n_607;
wire n_184;
wire n_265;
wire n_57;
wire n_674;
wire n_51;
wire n_570;
wire n_411;
wire n_514;
wire n_287;
wire n_144;
wire n_403;
wire n_625;
wire n_45;
wire n_131;
wire n_420;
wire n_86;
wire n_27;
wire n_738;
wire n_177;
wire n_28;
wire n_511;
wire n_448;
wire n_49;
wire n_206;
wire n_349;
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_33), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_68), .Y(n_102) );
CKINVDCx5p33_ASAP7_75t_R g103 ( .A(n_55), .Y(n_103) );
INVx1_ASAP7_75t_SL g104 ( .A(n_20), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_22), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_98), .Y(n_106) );
BUFx6f_ASAP7_75t_L g107 ( .A(n_70), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_12), .Y(n_108) );
OR2x2_ASAP7_75t_L g109 ( .A(n_92), .B(n_19), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_41), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_67), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_15), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_40), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_81), .Y(n_114) );
INVxp67_ASAP7_75t_L g115 ( .A(n_15), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_51), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_23), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_12), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_34), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g120 ( .A(n_83), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_76), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_59), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_86), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_91), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_65), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_96), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_58), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_3), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_73), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_32), .Y(n_130) );
BUFx10_ASAP7_75t_L g131 ( .A(n_47), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_31), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_56), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_2), .Y(n_134) );
CKINVDCx5p33_ASAP7_75t_R g135 ( .A(n_71), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_48), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_49), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_10), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_117), .Y(n_139) );
AOI22xp5_ASAP7_75t_SL g140 ( .A1(n_138), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_140) );
AND2x4_ASAP7_75t_L g141 ( .A(n_117), .B(n_0), .Y(n_141) );
AND2x6_ASAP7_75t_L g142 ( .A(n_102), .B(n_18), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_107), .Y(n_143) );
INVx6_ASAP7_75t_L g144 ( .A(n_131), .Y(n_144) );
INVx6_ASAP7_75t_L g145 ( .A(n_131), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_108), .B(n_1), .Y(n_146) );
AND2x2_ASAP7_75t_L g147 ( .A(n_120), .B(n_3), .Y(n_147) );
AOI22xp5_ASAP7_75t_L g148 ( .A1(n_138), .A2(n_4), .B1(n_5), .B2(n_6), .Y(n_148) );
BUFx12f_ASAP7_75t_L g149 ( .A(n_131), .Y(n_149) );
INVx2_ASAP7_75t_L g150 ( .A(n_106), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_110), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_114), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_107), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_107), .Y(n_154) );
BUFx6f_ASAP7_75t_L g155 ( .A(n_107), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_119), .B(n_121), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_124), .Y(n_157) );
OA21x2_ASAP7_75t_L g158 ( .A1(n_125), .A2(n_52), .B(n_99), .Y(n_158) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_126), .A2(n_50), .B(n_97), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
CKINVDCx16_ASAP7_75t_R g161 ( .A(n_116), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_161), .Y(n_162) );
INVx6_ASAP7_75t_L g163 ( .A(n_141), .Y(n_163) );
AND2x6_ASAP7_75t_L g164 ( .A(n_141), .B(n_136), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
INVx4_ASAP7_75t_L g166 ( .A(n_142), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_142), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_141), .Y(n_168) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_149), .B(n_103), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g170 ( .A(n_144), .B(n_103), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_143), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
INVx2_ASAP7_75t_L g174 ( .A(n_143), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_141), .Y(n_175) );
INVx3_ASAP7_75t_L g176 ( .A(n_146), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g178 ( .A1(n_146), .A2(n_118), .B1(n_115), .B2(n_134), .Y(n_178) );
OAI22xp5_ASAP7_75t_L g179 ( .A1(n_144), .A2(n_116), .B1(n_112), .B2(n_128), .Y(n_179) );
INVx3_ASAP7_75t_L g180 ( .A(n_146), .Y(n_180) );
NAND2xp5_ASAP7_75t_SL g181 ( .A(n_149), .B(n_105), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_153), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g183 ( .A(n_144), .B(n_105), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_139), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_139), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_153), .Y(n_186) );
AOI22xp5_ASAP7_75t_L g187 ( .A1(n_146), .A2(n_137), .B1(n_135), .B2(n_133), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_144), .B(n_137), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
OR2x6_ASAP7_75t_L g190 ( .A(n_145), .B(n_109), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_145), .B(n_101), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_145), .B(n_111), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_157), .B(n_113), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_150), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_153), .Y(n_195) );
BUFx3_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
BUFx3_ASAP7_75t_L g197 ( .A(n_142), .Y(n_197) );
NOR2x1p5_ASAP7_75t_L g198 ( .A(n_147), .B(n_122), .Y(n_198) );
INVx3_ASAP7_75t_L g199 ( .A(n_154), .Y(n_199) );
INVx1_ASAP7_75t_L g200 ( .A(n_150), .Y(n_200) );
INVx2_ASAP7_75t_SL g201 ( .A(n_145), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_184), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_170), .B(n_147), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_194), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_183), .B(n_157), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_188), .B(n_156), .Y(n_207) );
OR2x6_ASAP7_75t_L g208 ( .A(n_190), .B(n_161), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_164), .B(n_151), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_184), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_185), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_176), .A2(n_159), .B(n_158), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_193), .B(n_160), .Y(n_213) );
NOR3xp33_ASAP7_75t_L g214 ( .A(n_179), .B(n_148), .C(n_152), .Y(n_214) );
BUFx4_ASAP7_75t_L g215 ( .A(n_162), .Y(n_215) );
AND2x2_ASAP7_75t_L g216 ( .A(n_190), .B(n_151), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_190), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_164), .B(n_152), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g219 ( .A(n_166), .B(n_160), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g220 ( .A(n_164), .B(n_142), .Y(n_220) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_164), .A2(n_142), .B1(n_158), .B2(n_159), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_191), .B(n_104), .Y(n_222) );
HB1xp67_ASAP7_75t_L g223 ( .A(n_190), .Y(n_223) );
INVx2_ASAP7_75t_L g224 ( .A(n_185), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_164), .B(n_142), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g226 ( .A(n_192), .B(n_123), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_164), .B(n_127), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_187), .Y(n_228) );
AOI22xp33_ASAP7_75t_L g229 ( .A1(n_164), .A2(n_158), .B1(n_159), .B2(n_155), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_187), .B(n_129), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_194), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_200), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_168), .B(n_130), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_178), .B(n_140), .Y(n_234) );
NAND2xp5_ASAP7_75t_SL g235 ( .A(n_166), .B(n_155), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_201), .B(n_159), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_198), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_169), .B(n_4), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_200), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_181), .B(n_5), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g241 ( .A(n_166), .B(n_155), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_168), .B(n_158), .Y(n_242) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_176), .A2(n_155), .B(n_154), .C(n_8), .Y(n_243) );
AOI22x1_ASAP7_75t_L g244 ( .A1(n_166), .A2(n_155), .B1(n_154), .B2(n_54), .Y(n_244) );
OR2x6_ASAP7_75t_L g245 ( .A(n_190), .B(n_154), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_175), .B(n_6), .Y(n_246) );
INVxp67_ASAP7_75t_L g247 ( .A(n_198), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_163), .Y(n_248) );
AOI22xp5_ASAP7_75t_L g249 ( .A1(n_163), .A2(n_7), .B1(n_8), .B2(n_9), .Y(n_249) );
BUFx5_ASAP7_75t_L g250 ( .A(n_167), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_201), .B(n_53), .Y(n_251) );
AND2x2_ASAP7_75t_L g252 ( .A(n_217), .B(n_176), .Y(n_252) );
AOI21x1_ASAP7_75t_L g253 ( .A1(n_212), .A2(n_175), .B(n_173), .Y(n_253) );
CKINVDCx11_ASAP7_75t_R g254 ( .A(n_208), .Y(n_254) );
CKINVDCx20_ASAP7_75t_R g255 ( .A(n_208), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_216), .B(n_176), .Y(n_256) );
O2A1O1Ixp33_ASAP7_75t_SL g257 ( .A1(n_242), .A2(n_202), .B(n_165), .C(n_171), .Y(n_257) );
AOI21xp5_ASAP7_75t_L g258 ( .A1(n_220), .A2(n_167), .B(n_197), .Y(n_258) );
INVx11_ASAP7_75t_L g259 ( .A(n_215), .Y(n_259) );
AOI22x1_ASAP7_75t_L g260 ( .A1(n_232), .A2(n_180), .B1(n_202), .B2(n_182), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_204), .B(n_180), .Y(n_261) );
AOI21xp5_ASAP7_75t_L g262 ( .A1(n_225), .A2(n_167), .B(n_197), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_236), .A2(n_196), .B(n_197), .Y(n_263) );
AO21x1_ASAP7_75t_L g264 ( .A1(n_236), .A2(n_202), .B(n_165), .Y(n_264) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_241), .A2(n_177), .B(n_174), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_208), .B(n_180), .Y(n_266) );
INVx4_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
AND2x2_ASAP7_75t_L g268 ( .A(n_228), .B(n_180), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_207), .B(n_163), .Y(n_269) );
NOR2xp33_ASAP7_75t_L g270 ( .A(n_230), .B(n_163), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_214), .B(n_196), .Y(n_271) );
AND2x2_ASAP7_75t_L g272 ( .A(n_234), .B(n_196), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_248), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_214), .B(n_7), .Y(n_274) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
AOI21x1_ASAP7_75t_L g276 ( .A1(n_241), .A2(n_177), .B(n_173), .Y(n_276) );
BUFx6f_ASAP7_75t_L g277 ( .A(n_245), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_206), .B(n_9), .Y(n_278) );
NOR2xp33_ASAP7_75t_L g279 ( .A(n_247), .B(n_10), .Y(n_279) );
NOR2xp67_ASAP7_75t_L g280 ( .A(n_237), .B(n_11), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_213), .B(n_11), .Y(n_281) );
O2A1O1Ixp33_ASAP7_75t_SL g282 ( .A1(n_243), .A2(n_182), .B(n_195), .C(n_171), .Y(n_282) );
AOI21xp5_ASAP7_75t_L g283 ( .A1(n_219), .A2(n_174), .B(n_186), .Y(n_283) );
OAI22xp5_ASAP7_75t_L g284 ( .A1(n_217), .A2(n_199), .B1(n_195), .B2(n_182), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_213), .B(n_13), .Y(n_285) );
O2A1O1Ixp33_ASAP7_75t_L g286 ( .A1(n_246), .A2(n_199), .B(n_189), .C(n_186), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_219), .A2(n_189), .B(n_195), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_222), .B(n_13), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_222), .B(n_14), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_203), .Y(n_290) );
BUFx3_ASAP7_75t_L g291 ( .A(n_254), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_263), .A2(n_235), .B(n_221), .Y(n_292) );
BUFx5_ASAP7_75t_L g293 ( .A(n_252), .Y(n_293) );
AO31x2_ASAP7_75t_L g294 ( .A1(n_264), .A2(n_251), .A3(n_205), .B(n_231), .Y(n_294) );
BUFx2_ASAP7_75t_L g295 ( .A(n_255), .Y(n_295) );
INVx5_ASAP7_75t_L g296 ( .A(n_277), .Y(n_296) );
AOI21xp5_ASAP7_75t_L g297 ( .A1(n_257), .A2(n_221), .B(n_229), .Y(n_297) );
AOI21xp5_ASAP7_75t_L g298 ( .A1(n_257), .A2(n_258), .B(n_262), .Y(n_298) );
NAND3x1_ASAP7_75t_L g299 ( .A(n_259), .B(n_249), .C(n_16), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_271), .A2(n_229), .B(n_233), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_256), .Y(n_301) );
OAI21x1_ASAP7_75t_L g302 ( .A1(n_253), .A2(n_276), .B(n_265), .Y(n_302) );
AO32x2_ASAP7_75t_L g303 ( .A1(n_267), .A2(n_251), .A3(n_223), .B1(n_240), .B2(n_238), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_277), .Y(n_304) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_270), .A2(n_218), .B(n_209), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_269), .A2(n_223), .B(n_227), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_274), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_261), .A2(n_211), .B(n_224), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_277), .Y(n_309) );
BUFx12f_ASAP7_75t_L g310 ( .A(n_254), .Y(n_310) );
OAI21x1_ASAP7_75t_SL g311 ( .A1(n_267), .A2(n_210), .B(n_239), .Y(n_311) );
OAI21x1_ASAP7_75t_SL g312 ( .A1(n_267), .A2(n_244), .B(n_250), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_272), .B(n_226), .Y(n_313) );
O2A1O1Ixp5_ASAP7_75t_SL g314 ( .A1(n_273), .A2(n_199), .B(n_172), .C(n_165), .Y(n_314) );
NAND2xp5_ASAP7_75t_SL g315 ( .A(n_277), .B(n_250), .Y(n_315) );
BUFx2_ASAP7_75t_L g316 ( .A(n_293), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_301), .Y(n_317) );
NOR2x1_ASAP7_75t_SL g318 ( .A(n_296), .B(n_290), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_310), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_302), .A2(n_286), .B(n_260), .Y(n_320) );
AOI21xp33_ASAP7_75t_L g321 ( .A1(n_307), .A2(n_288), .B(n_289), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_301), .Y(n_322) );
OAI21x1_ASAP7_75t_L g323 ( .A1(n_297), .A2(n_285), .B(n_281), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_308), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_313), .B(n_268), .Y(n_325) );
INVx3_ASAP7_75t_L g326 ( .A(n_309), .Y(n_326) );
OA21x2_ASAP7_75t_L g327 ( .A1(n_298), .A2(n_278), .B(n_287), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_293), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_293), .B(n_270), .Y(n_329) );
NOR2x1_ASAP7_75t_SL g330 ( .A(n_296), .B(n_290), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_293), .Y(n_331) );
OAI21xp5_ASAP7_75t_L g332 ( .A1(n_300), .A2(n_282), .B(n_252), .Y(n_332) );
OAI21x1_ASAP7_75t_L g333 ( .A1(n_314), .A2(n_283), .B(n_284), .Y(n_333) );
AO31x2_ASAP7_75t_L g334 ( .A1(n_292), .A2(n_279), .A3(n_282), .B(n_226), .Y(n_334) );
CKINVDCx5p33_ASAP7_75t_R g335 ( .A(n_291), .Y(n_335) );
AND2x4_ASAP7_75t_L g336 ( .A(n_296), .B(n_266), .Y(n_336) );
HB1xp67_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
AOI21xp5_ASAP7_75t_L g339 ( .A1(n_306), .A2(n_290), .B(n_275), .Y(n_339) );
OAI21x1_ASAP7_75t_L g340 ( .A1(n_312), .A2(n_280), .B(n_171), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_309), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_324), .Y(n_342) );
OAI21x1_ASAP7_75t_L g343 ( .A1(n_320), .A2(n_311), .B(n_315), .Y(n_343) );
BUFx3_ASAP7_75t_L g344 ( .A(n_316), .Y(n_344) );
INVx2_ASAP7_75t_L g345 ( .A(n_324), .Y(n_345) );
INVx2_ASAP7_75t_L g346 ( .A(n_322), .Y(n_346) );
NAND2xp33_ASAP7_75t_R g347 ( .A(n_335), .B(n_304), .Y(n_347) );
BUFx2_ASAP7_75t_R g348 ( .A(n_325), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_322), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_322), .Y(n_350) );
OAI21x1_ASAP7_75t_L g351 ( .A1(n_320), .A2(n_305), .B(n_304), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_317), .Y(n_352) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_325), .A2(n_255), .B1(n_279), .B2(n_290), .Y(n_353) );
OR2x2_ASAP7_75t_L g354 ( .A(n_317), .B(n_294), .Y(n_354) );
OAI21x1_ASAP7_75t_L g355 ( .A1(n_320), .A2(n_294), .B(n_299), .Y(n_355) );
BUFx3_ASAP7_75t_L g356 ( .A(n_316), .Y(n_356) );
BUFx2_ASAP7_75t_L g357 ( .A(n_328), .Y(n_357) );
BUFx2_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_331), .Y(n_359) );
INVx2_ASAP7_75t_L g360 ( .A(n_327), .Y(n_360) );
OA21x2_ASAP7_75t_L g361 ( .A1(n_323), .A2(n_294), .B(n_303), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_336), .B(n_303), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_338), .Y(n_364) );
BUFx10_ASAP7_75t_L g365 ( .A(n_336), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_327), .Y(n_366) );
INVx2_ASAP7_75t_L g367 ( .A(n_327), .Y(n_367) );
CKINVDCx11_ASAP7_75t_R g368 ( .A(n_319), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_327), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_338), .Y(n_370) );
AO21x2_ASAP7_75t_L g371 ( .A1(n_332), .A2(n_303), .B(n_172), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_338), .Y(n_372) );
BUFx3_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
AND2x6_ASAP7_75t_L g374 ( .A(n_341), .B(n_250), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_341), .Y(n_375) );
BUFx6f_ASAP7_75t_L g376 ( .A(n_326), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_341), .Y(n_377) );
INVx2_ASAP7_75t_L g378 ( .A(n_323), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_334), .B(n_14), .Y(n_379) );
OR2x2_ASAP7_75t_L g380 ( .A(n_337), .B(n_16), .Y(n_380) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_326), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_323), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_346), .B(n_334), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_379), .A2(n_321), .B1(n_329), .B2(n_336), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_360), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_342), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_342), .Y(n_388) );
AND2x2_ASAP7_75t_L g389 ( .A(n_346), .B(n_334), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_354), .B(n_329), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_346), .Y(n_391) );
AND2x2_ASAP7_75t_L g392 ( .A(n_349), .B(n_334), .Y(n_392) );
OR2x2_ASAP7_75t_L g393 ( .A(n_354), .B(n_334), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_352), .B(n_321), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_349), .B(n_334), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_349), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_350), .B(n_332), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_350), .B(n_379), .Y(n_398) );
OR2x2_ASAP7_75t_L g399 ( .A(n_357), .B(n_326), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_376), .Y(n_400) );
AND2x2_ASAP7_75t_L g401 ( .A(n_379), .B(n_326), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_352), .B(n_330), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_380), .B(n_353), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_380), .B(n_330), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_363), .B(n_318), .Y(n_405) );
INVx3_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
INVx2_ASAP7_75t_L g407 ( .A(n_360), .Y(n_407) );
AOI22xp33_ASAP7_75t_SL g408 ( .A1(n_365), .A2(n_318), .B1(n_340), .B2(n_339), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_360), .Y(n_409) );
BUFx2_ASAP7_75t_L g410 ( .A(n_344), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_359), .B(n_17), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_357), .B(n_358), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_365), .Y(n_413) );
BUFx2_ASAP7_75t_L g414 ( .A(n_344), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_359), .B(n_17), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_345), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_366), .Y(n_417) );
AND2x2_ASAP7_75t_L g418 ( .A(n_363), .B(n_340), .Y(n_418) );
AO21x2_ASAP7_75t_L g419 ( .A1(n_355), .A2(n_333), .B(n_340), .Y(n_419) );
BUFx6f_ASAP7_75t_L g420 ( .A(n_376), .Y(n_420) );
BUFx6f_ASAP7_75t_L g421 ( .A(n_376), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_366), .Y(n_422) );
INVx3_ASAP7_75t_L g423 ( .A(n_376), .Y(n_423) );
AND2x4_ASAP7_75t_L g424 ( .A(n_345), .B(n_333), .Y(n_424) );
BUFx2_ASAP7_75t_L g425 ( .A(n_344), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_366), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_345), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_364), .B(n_333), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_364), .B(n_21), .Y(n_429) );
NOR2x1_ASAP7_75t_R g430 ( .A(n_368), .B(n_250), .Y(n_430) );
BUFx2_ASAP7_75t_L g431 ( .A(n_356), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_362), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_362), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_367), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_358), .B(n_24), .Y(n_435) );
INVxp67_ASAP7_75t_L g436 ( .A(n_347), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_356), .B(n_25), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_367), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_367), .Y(n_439) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_356), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
AND2x2_ASAP7_75t_L g442 ( .A(n_370), .B(n_26), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_370), .B(n_27), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_369), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_369), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_372), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_375), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_377), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_375), .B(n_28), .Y(n_449) );
AND2x2_ASAP7_75t_L g450 ( .A(n_377), .B(n_29), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_382), .Y(n_451) );
AND2x4_ASAP7_75t_SL g452 ( .A(n_365), .B(n_172), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_372), .B(n_30), .Y(n_453) );
NOR2xp67_ASAP7_75t_SL g454 ( .A(n_437), .B(n_348), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_398), .B(n_373), .Y(n_455) );
NAND2x1p5_ASAP7_75t_L g456 ( .A(n_437), .B(n_373), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_386), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_398), .B(n_371), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_432), .B(n_373), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_386), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_432), .Y(n_461) );
NOR2xp67_ASAP7_75t_L g462 ( .A(n_436), .B(n_381), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_405), .B(n_365), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_433), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_390), .B(n_381), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_433), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_447), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_405), .B(n_377), .Y(n_468) );
HB1xp67_ASAP7_75t_L g469 ( .A(n_434), .Y(n_469) );
BUFx2_ASAP7_75t_L g470 ( .A(n_440), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_447), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g472 ( .A(n_394), .B(n_361), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_402), .B(n_361), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_418), .B(n_371), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_402), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_386), .Y(n_476) );
OR2x2_ASAP7_75t_L g477 ( .A(n_390), .B(n_361), .Y(n_477) );
OR2x2_ASAP7_75t_L g478 ( .A(n_412), .B(n_361), .Y(n_478) );
INVx2_ASAP7_75t_L g479 ( .A(n_407), .Y(n_479) );
AND2x2_ASAP7_75t_SL g480 ( .A(n_412), .B(n_361), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_418), .B(n_371), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_397), .B(n_371), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_397), .B(n_355), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_401), .B(n_355), .Y(n_484) );
INVx2_ASAP7_75t_SL g485 ( .A(n_410), .Y(n_485) );
AND2x4_ASAP7_75t_L g486 ( .A(n_401), .B(n_382), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_403), .B(n_376), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_434), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_384), .Y(n_489) );
AND2x4_ASAP7_75t_L g490 ( .A(n_410), .B(n_382), .Y(n_490) );
OR2x2_ASAP7_75t_L g491 ( .A(n_414), .B(n_378), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_407), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_384), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_407), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_404), .B(n_378), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_387), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_414), .B(n_348), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_409), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_425), .B(n_351), .Y(n_499) );
AND2x4_ASAP7_75t_L g500 ( .A(n_425), .B(n_378), .Y(n_500) );
OR2x2_ASAP7_75t_L g501 ( .A(n_431), .B(n_351), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_431), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_387), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_388), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_388), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_409), .Y(n_506) );
INVx2_ASAP7_75t_SL g507 ( .A(n_446), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_416), .Y(n_508) );
AND2x4_ASAP7_75t_L g509 ( .A(n_416), .B(n_343), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_427), .Y(n_510) );
AND2x2_ASAP7_75t_L g511 ( .A(n_383), .B(n_351), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_452), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_383), .B(n_343), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_385), .B(n_413), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_427), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g516 ( .A(n_413), .B(n_374), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_389), .B(n_392), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_389), .B(n_374), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_399), .B(n_343), .Y(n_519) );
INVx3_ASAP7_75t_L g520 ( .A(n_417), .Y(n_520) );
HB1xp67_ASAP7_75t_L g521 ( .A(n_438), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_393), .A2(n_415), .B1(n_411), .B2(n_395), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_399), .B(n_374), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_429), .B(n_374), .Y(n_524) );
OAI22xp5_ASAP7_75t_L g525 ( .A1(n_453), .A2(n_374), .B1(n_36), .B2(n_37), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_392), .B(n_374), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_395), .B(n_374), .Y(n_527) );
INVx2_ASAP7_75t_SL g528 ( .A(n_452), .Y(n_528) );
INVx2_ASAP7_75t_L g529 ( .A(n_417), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_391), .B(n_35), .Y(n_530) );
INVx3_ASAP7_75t_L g531 ( .A(n_422), .Y(n_531) );
OAI21x1_ASAP7_75t_L g532 ( .A1(n_406), .A2(n_374), .B(n_199), .Y(n_532) );
AND2x2_ASAP7_75t_L g533 ( .A(n_393), .B(n_374), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_391), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_422), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_396), .Y(n_536) );
OR2x2_ASAP7_75t_L g537 ( .A(n_396), .B(n_38), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_438), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_439), .B(n_39), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_426), .Y(n_540) );
INVx4_ASAP7_75t_L g541 ( .A(n_452), .Y(n_541) );
BUFx2_ASAP7_75t_L g542 ( .A(n_430), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_439), .B(n_42), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_429), .B(n_43), .Y(n_544) );
HB1xp67_ASAP7_75t_L g545 ( .A(n_441), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_426), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_441), .B(n_44), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_444), .B(n_45), .Y(n_548) );
INVx1_ASAP7_75t_L g549 ( .A(n_444), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_445), .Y(n_550) );
BUFx2_ASAP7_75t_L g551 ( .A(n_541), .Y(n_551) );
NOR2x1_ASAP7_75t_L g552 ( .A(n_541), .B(n_453), .Y(n_552) );
NOR2xp67_ASAP7_75t_L g553 ( .A(n_541), .B(n_445), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_461), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_457), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_468), .B(n_428), .Y(n_556) );
INVx2_ASAP7_75t_L g557 ( .A(n_457), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_464), .Y(n_558) );
INVx4_ASAP7_75t_L g559 ( .A(n_542), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_466), .Y(n_560) );
AND2x2_ASAP7_75t_L g561 ( .A(n_475), .B(n_428), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_483), .B(n_424), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_522), .B(n_448), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_483), .B(n_424), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_484), .B(n_424), .Y(n_566) );
INVx1_ASAP7_75t_L g567 ( .A(n_471), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_517), .B(n_448), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_469), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_469), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_488), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_484), .B(n_424), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_460), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_488), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_521), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_521), .Y(n_576) );
OR2x2_ASAP7_75t_L g577 ( .A(n_507), .B(n_451), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_538), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_512), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g581 ( .A(n_522), .B(n_408), .C(n_435), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_545), .Y(n_582) );
AND2x2_ASAP7_75t_L g583 ( .A(n_513), .B(n_451), .Y(n_583) );
AND2x2_ASAP7_75t_L g584 ( .A(n_470), .B(n_406), .Y(n_584) );
OR2x2_ASAP7_75t_L g585 ( .A(n_507), .B(n_423), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_545), .Y(n_586) );
INVx4_ASAP7_75t_L g587 ( .A(n_528), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_463), .B(n_406), .Y(n_588) );
INVx2_ASAP7_75t_L g589 ( .A(n_460), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_465), .B(n_449), .Y(n_590) );
INVx2_ASAP7_75t_SL g591 ( .A(n_502), .Y(n_591) );
OR2x2_ASAP7_75t_L g592 ( .A(n_455), .B(n_423), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_477), .B(n_449), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_489), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_533), .B(n_406), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_482), .B(n_443), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_476), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_533), .B(n_423), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_493), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_497), .B(n_423), .Y(n_600) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_462), .B(n_443), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_476), .Y(n_602) );
INVx1_ASAP7_75t_L g603 ( .A(n_496), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_513), .B(n_419), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_458), .B(n_419), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_523), .B(n_421), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_482), .B(n_442), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_458), .B(n_442), .Y(n_608) );
HB1xp67_ASAP7_75t_L g609 ( .A(n_520), .Y(n_609) );
NOR2x1_ASAP7_75t_L g610 ( .A(n_539), .B(n_450), .Y(n_610) );
INVx2_ASAP7_75t_L g611 ( .A(n_479), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_485), .B(n_421), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_456), .B(n_421), .Y(n_613) );
OR2x2_ASAP7_75t_L g614 ( .A(n_495), .B(n_421), .Y(n_614) );
AND2x2_ASAP7_75t_L g615 ( .A(n_485), .B(n_421), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_503), .B(n_450), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_528), .B(n_480), .Y(n_617) );
AND2x2_ASAP7_75t_L g618 ( .A(n_480), .B(n_420), .Y(n_618) );
NOR2xp67_ASAP7_75t_R g619 ( .A(n_454), .B(n_430), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_504), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_474), .B(n_419), .Y(n_621) );
INVx2_ASAP7_75t_L g622 ( .A(n_479), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_505), .Y(n_623) );
INVx4_ASAP7_75t_L g624 ( .A(n_456), .Y(n_624) );
INVx2_ASAP7_75t_SL g625 ( .A(n_491), .Y(n_625) );
INVx2_ASAP7_75t_L g626 ( .A(n_492), .Y(n_626) );
INVx2_ASAP7_75t_L g627 ( .A(n_492), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_508), .B(n_420), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_510), .Y(n_629) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_514), .B(n_420), .Y(n_630) );
OR2x2_ASAP7_75t_L g631 ( .A(n_473), .B(n_420), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_525), .A2(n_420), .B(n_400), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_515), .Y(n_633) );
BUFx3_ASAP7_75t_L g634 ( .A(n_490), .Y(n_634) );
OR2x2_ASAP7_75t_L g635 ( .A(n_478), .B(n_400), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_459), .B(n_400), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_549), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_534), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_524), .B(n_400), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_486), .B(n_400), .Y(n_640) );
OR2x2_ASAP7_75t_L g641 ( .A(n_520), .B(n_46), .Y(n_641) );
INVx2_ASAP7_75t_L g642 ( .A(n_494), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_494), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_536), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_474), .B(n_57), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_511), .B(n_60), .Y(n_646) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_472), .B(n_61), .Y(n_647) );
NAND4xp25_ASAP7_75t_L g648 ( .A(n_487), .B(n_62), .C(n_63), .D(n_64), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_520), .Y(n_649) );
AND2x2_ASAP7_75t_L g650 ( .A(n_481), .B(n_66), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_554), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_621), .A2(n_481), .B1(n_511), .B2(n_499), .C(n_509), .Y(n_652) );
AND2x2_ASAP7_75t_L g653 ( .A(n_600), .B(n_486), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_621), .B(n_531), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_556), .B(n_486), .Y(n_655) );
NAND4xp25_ASAP7_75t_L g656 ( .A(n_581), .B(n_516), .C(n_519), .D(n_544), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_605), .B(n_550), .Y(n_657) );
HB1xp67_ASAP7_75t_L g658 ( .A(n_575), .Y(n_658) );
NOR2x1_ASAP7_75t_L g659 ( .A(n_559), .B(n_548), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_605), .B(n_550), .Y(n_660) );
INVx2_ASAP7_75t_L g661 ( .A(n_575), .Y(n_661) );
INVxp67_ASAP7_75t_L g662 ( .A(n_591), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_558), .Y(n_663) );
INVx1_ASAP7_75t_SL g664 ( .A(n_551), .Y(n_664) );
AND2x4_ASAP7_75t_L g665 ( .A(n_587), .B(n_509), .Y(n_665) );
AND2x4_ASAP7_75t_L g666 ( .A(n_587), .B(n_509), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_560), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_564), .Y(n_668) );
NAND2x1_ASAP7_75t_L g669 ( .A(n_587), .B(n_531), .Y(n_669) );
NOR2x1_ASAP7_75t_L g670 ( .A(n_559), .B(n_548), .Y(n_670) );
INVx2_ASAP7_75t_SL g671 ( .A(n_591), .Y(n_671) );
INVx2_ASAP7_75t_L g672 ( .A(n_625), .Y(n_672) );
AND2x2_ASAP7_75t_L g673 ( .A(n_566), .B(n_518), .Y(n_673) );
INVx2_ASAP7_75t_L g674 ( .A(n_625), .Y(n_674) );
INVx2_ASAP7_75t_L g675 ( .A(n_577), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_567), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_559), .A2(n_526), .B1(n_527), .B2(n_490), .Y(n_677) );
NAND2x1_ASAP7_75t_L g678 ( .A(n_553), .B(n_531), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_580), .Y(n_679) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_604), .B(n_529), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_604), .B(n_529), .Y(n_681) );
AND2x2_ASAP7_75t_L g682 ( .A(n_566), .B(n_490), .Y(n_682) );
INVxp67_ASAP7_75t_SL g683 ( .A(n_609), .Y(n_683) );
AND2x2_ASAP7_75t_L g684 ( .A(n_572), .B(n_500), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_594), .Y(n_685) );
INVx2_ASAP7_75t_L g686 ( .A(n_555), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_624), .B(n_547), .Y(n_687) );
NOR2xp67_ASAP7_75t_L g688 ( .A(n_624), .B(n_501), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_568), .B(n_500), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_599), .Y(n_690) );
OR2x2_ASAP7_75t_L g691 ( .A(n_583), .B(n_535), .Y(n_691) );
NOR2xp33_ASAP7_75t_L g692 ( .A(n_592), .B(n_500), .Y(n_692) );
INVxp67_ASAP7_75t_L g693 ( .A(n_617), .Y(n_693) );
NOR3xp33_ASAP7_75t_L g694 ( .A(n_648), .B(n_543), .C(n_547), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_603), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_620), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_623), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_569), .B(n_546), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_629), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_624), .B(n_546), .Y(n_700) );
AND2x2_ASAP7_75t_L g701 ( .A(n_572), .B(n_540), .Y(n_701) );
OR2x2_ASAP7_75t_L g702 ( .A(n_583), .B(n_540), .Y(n_702) );
INVx2_ASAP7_75t_L g703 ( .A(n_555), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_633), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_563), .B(n_535), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_634), .Y(n_706) );
AND2x2_ASAP7_75t_L g707 ( .A(n_562), .B(n_506), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_637), .Y(n_708) );
AND2x2_ASAP7_75t_L g709 ( .A(n_562), .B(n_506), .Y(n_709) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_570), .B(n_498), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_634), .B(n_498), .Y(n_711) );
INVx1_ASAP7_75t_SL g712 ( .A(n_584), .Y(n_712) );
AND2x4_ASAP7_75t_L g713 ( .A(n_618), .B(n_532), .Y(n_713) );
INVx2_ASAP7_75t_L g714 ( .A(n_557), .Y(n_714) );
AND2x2_ASAP7_75t_L g715 ( .A(n_565), .B(n_532), .Y(n_715) );
NAND4xp25_ASAP7_75t_L g716 ( .A(n_645), .B(n_530), .C(n_537), .D(n_74), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_571), .B(n_69), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_561), .B(n_72), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_638), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_574), .B(n_75), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_565), .B(n_77), .Y(n_721) );
INVxp33_ASAP7_75t_L g722 ( .A(n_619), .Y(n_722) );
AND2x2_ASAP7_75t_L g723 ( .A(n_588), .B(n_78), .Y(n_723) );
AND2x2_ASAP7_75t_L g724 ( .A(n_595), .B(n_79), .Y(n_724) );
AND2x4_ASAP7_75t_L g725 ( .A(n_688), .B(n_586), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_711), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_675), .B(n_576), .Y(n_727) );
O2A1O1Ixp33_ASAP7_75t_L g728 ( .A1(n_722), .A2(n_650), .B(n_645), .C(n_646), .Y(n_728) );
OAI21xp5_ASAP7_75t_SL g729 ( .A1(n_656), .A2(n_552), .B(n_601), .Y(n_729) );
OAI22xp33_ASAP7_75t_L g730 ( .A1(n_656), .A2(n_610), .B1(n_590), .B2(n_608), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_679), .B(n_578), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_712), .B(n_606), .Y(n_732) );
AND2x2_ASAP7_75t_L g733 ( .A(n_712), .B(n_639), .Y(n_733) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_716), .A2(n_650), .B1(n_647), .B2(n_630), .Y(n_734) );
NAND2xp33_ASAP7_75t_SL g735 ( .A(n_669), .B(n_609), .Y(n_735) );
AND2x2_ASAP7_75t_L g736 ( .A(n_682), .B(n_598), .Y(n_736) );
NOR2xp33_ASAP7_75t_L g737 ( .A(n_662), .B(n_585), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_684), .B(n_630), .Y(n_738) );
AND2x2_ASAP7_75t_L g739 ( .A(n_655), .B(n_640), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_651), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_659), .A2(n_632), .B1(n_607), .B2(n_596), .Y(n_741) );
NAND2xp5_ASAP7_75t_L g742 ( .A(n_705), .B(n_582), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_716), .A2(n_647), .B1(n_593), .B2(n_579), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_663), .Y(n_744) );
AOI22x1_ASAP7_75t_SL g745 ( .A1(n_664), .A2(n_649), .B1(n_644), .B2(n_611), .Y(n_745) );
NOR2xp33_ASAP7_75t_L g746 ( .A(n_671), .B(n_635), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_667), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_711), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_693), .B(n_615), .Y(n_749) );
OR2x2_ASAP7_75t_L g750 ( .A(n_680), .B(n_631), .Y(n_750) );
INVx1_ASAP7_75t_L g751 ( .A(n_668), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_676), .Y(n_752) );
INVxp67_ASAP7_75t_L g753 ( .A(n_658), .Y(n_753) );
AO22x1_ASAP7_75t_L g754 ( .A1(n_670), .A2(n_612), .B1(n_616), .B2(n_643), .Y(n_754) );
AOI22xp5_ASAP7_75t_L g755 ( .A1(n_652), .A2(n_636), .B1(n_632), .B2(n_643), .Y(n_755) );
AOI22xp5_ASAP7_75t_L g756 ( .A1(n_715), .A2(n_557), .B1(n_627), .B2(n_626), .Y(n_756) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_664), .B(n_614), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_661), .B(n_642), .Y(n_758) );
INVx1_ASAP7_75t_L g759 ( .A(n_685), .Y(n_759) );
AND2x2_ASAP7_75t_L g760 ( .A(n_701), .B(n_613), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_680), .B(n_642), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_690), .Y(n_762) );
INVx1_ASAP7_75t_L g763 ( .A(n_695), .Y(n_763) );
OAI221xp5_ASAP7_75t_L g764 ( .A1(n_677), .A2(n_613), .B1(n_628), .B2(n_627), .C(n_626), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_681), .B(n_602), .Y(n_765) );
OAI322xp33_ASAP7_75t_L g766 ( .A1(n_654), .A2(n_602), .A3(n_622), .B1(n_573), .B2(n_611), .C1(n_589), .C2(n_597), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_687), .A2(n_613), .B(n_641), .Y(n_767) );
NOR2xp33_ASAP7_75t_L g768 ( .A(n_731), .B(n_672), .Y(n_768) );
INVx2_ASAP7_75t_SL g769 ( .A(n_732), .Y(n_769) );
AOI22xp5_ASAP7_75t_L g770 ( .A1(n_730), .A2(n_692), .B1(n_689), .B2(n_674), .Y(n_770) );
AOI322xp5_ASAP7_75t_L g771 ( .A1(n_730), .A2(n_706), .A3(n_673), .B1(n_707), .B2(n_709), .C1(n_683), .C2(n_681), .Y(n_771) );
OAI21xp5_ASAP7_75t_SL g772 ( .A1(n_729), .A2(n_706), .B(n_666), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_743), .A2(n_697), .B1(n_699), .B2(n_696), .C(n_704), .Y(n_773) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_743), .A2(n_665), .B1(n_666), .B2(n_678), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g775 ( .A1(n_734), .A2(n_708), .B1(n_660), .B2(n_657), .C(n_719), .Y(n_775) );
AOI222xp33_ASAP7_75t_L g776 ( .A1(n_734), .A2(n_657), .B1(n_660), .B2(n_710), .C1(n_698), .C2(n_718), .Y(n_776) );
OAI32xp33_ASAP7_75t_L g777 ( .A1(n_735), .A2(n_694), .A3(n_700), .B1(n_702), .B2(n_691), .Y(n_777) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_741), .A2(n_713), .B1(n_721), .B2(n_665), .Y(n_778) );
AOI21xp5_ASAP7_75t_L g779 ( .A1(n_754), .A2(n_698), .B(n_710), .Y(n_779) );
AOI21xp33_ASAP7_75t_L g780 ( .A1(n_728), .A2(n_720), .B(n_717), .Y(n_780) );
INVx1_ASAP7_75t_L g781 ( .A(n_742), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_740), .Y(n_782) );
AOI21xp5_ASAP7_75t_L g783 ( .A1(n_767), .A2(n_713), .B(n_720), .Y(n_783) );
AOI22xp33_ASAP7_75t_SL g784 ( .A1(n_745), .A2(n_723), .B1(n_724), .B2(n_653), .Y(n_784) );
OAI22x1_ASAP7_75t_L g785 ( .A1(n_725), .A2(n_714), .B1(n_703), .B2(n_686), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_744), .Y(n_786) );
NOR2xp33_ASAP7_75t_L g787 ( .A(n_731), .B(n_717), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_753), .B(n_622), .Y(n_788) );
AOI21xp33_ASAP7_75t_SL g789 ( .A1(n_728), .A2(n_597), .B(n_589), .Y(n_789) );
AOI22xp5_ASAP7_75t_L g790 ( .A1(n_737), .A2(n_573), .B1(n_172), .B2(n_250), .Y(n_790) );
OAI21xp5_ASAP7_75t_L g791 ( .A1(n_771), .A2(n_767), .B(n_753), .Y(n_791) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_776), .A2(n_764), .B1(n_755), .B2(n_746), .Y(n_792) );
AOI211xp5_ASAP7_75t_L g793 ( .A1(n_777), .A2(n_766), .B(n_725), .C(n_757), .Y(n_793) );
AO21x1_ASAP7_75t_L g794 ( .A1(n_772), .A2(n_751), .B(n_763), .Y(n_794) );
NOR2x1_ASAP7_75t_L g795 ( .A(n_774), .B(n_747), .Y(n_795) );
NOR3xp33_ASAP7_75t_L g796 ( .A(n_773), .B(n_762), .C(n_759), .Y(n_796) );
NOR3xp33_ASAP7_75t_L g797 ( .A(n_775), .B(n_752), .C(n_727), .Y(n_797) );
A2O1A1Ixp33_ASAP7_75t_L g798 ( .A1(n_789), .A2(n_756), .B(n_760), .C(n_749), .Y(n_798) );
A2O1A1Ixp33_ASAP7_75t_L g799 ( .A1(n_784), .A2(n_733), .B(n_726), .C(n_748), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_785), .A2(n_758), .B(n_761), .Y(n_800) );
NOR4xp25_ASAP7_75t_L g801 ( .A(n_778), .B(n_765), .C(n_750), .D(n_739), .Y(n_801) );
NAND3xp33_ASAP7_75t_L g802 ( .A(n_776), .B(n_738), .C(n_736), .Y(n_802) );
NAND3xp33_ASAP7_75t_L g803 ( .A(n_791), .B(n_770), .C(n_783), .Y(n_803) );
UNKNOWN g804 ( );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_799), .A2(n_779), .B(n_780), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_797), .B(n_781), .Y(n_806) );
NAND4xp25_ASAP7_75t_L g807 ( .A(n_793), .B(n_790), .C(n_787), .D(n_768), .Y(n_807) );
NAND3xp33_ASAP7_75t_SL g808 ( .A(n_794), .B(n_788), .C(n_786), .Y(n_808) );
NAND2xp33_ASAP7_75t_L g809 ( .A(n_803), .B(n_795), .Y(n_809) );
NOR2x1_ASAP7_75t_L g810 ( .A(n_808), .B(n_802), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_806), .Y(n_811) );
NOR3xp33_ASAP7_75t_L g812 ( .A(n_804), .B(n_798), .C(n_796), .Y(n_812) );
NOR2x1_ASAP7_75t_L g813 ( .A(n_809), .B(n_807), .Y(n_813) );
NOR4xp25_ASAP7_75t_L g814 ( .A(n_811), .B(n_782), .C(n_805), .D(n_801), .Y(n_814) );
AND3x2_ASAP7_75t_L g815 ( .A(n_812), .B(n_800), .C(n_769), .Y(n_815) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_813), .A2(n_810), .B1(n_172), .B2(n_250), .Y(n_816) );
NOR2xp33_ASAP7_75t_SL g817 ( .A(n_815), .B(n_172), .Y(n_817) );
NOR4xp75_ASAP7_75t_L g818 ( .A(n_817), .B(n_814), .C(n_82), .D(n_84), .Y(n_818) );
AND2x2_ASAP7_75t_L g819 ( .A(n_816), .B(n_80), .Y(n_819) );
NAND2xp5_ASAP7_75t_L g820 ( .A(n_819), .B(n_85), .Y(n_820) );
OAI21xp5_ASAP7_75t_L g821 ( .A1(n_820), .A2(n_818), .B(n_88), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_821), .B(n_87), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_822), .A2(n_89), .B(n_90), .Y(n_823) );
XNOR2x1_ASAP7_75t_L g824 ( .A(n_823), .B(n_93), .Y(n_824) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_824), .A2(n_100), .B1(n_94), .B2(n_95), .Y(n_825) );
endmodule