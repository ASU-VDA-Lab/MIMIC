module fake_netlist_1_3610_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
BUFx3_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
INVx3_ASAP7_75t_L g4 ( .A(n_2), .Y(n_4) );
OAI21x1_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B(n_1), .Y(n_5) );
OAI21x1_ASAP7_75t_SL g6 ( .A1(n_4), .A2(n_0), .B(n_2), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
OAI221xp5_ASAP7_75t_SL g9 ( .A1(n_8), .A2(n_3), .B1(n_5), .B2(n_6), .C(n_4), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
CKINVDCx20_ASAP7_75t_R g11 ( .A(n_10), .Y(n_11) );
endmodule