module fake_jpeg_2622_n_349 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_349);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_349;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

HB1xp67_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

BUFx4f_ASAP7_75t_SL g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_11),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_41),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_42),
.Y(n_116)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_43),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_44),
.Y(n_122)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_15),
.B(n_13),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_47),
.B(n_33),
.Y(n_102)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

INVx11_ASAP7_75t_L g110 ( 
.A(n_48),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_49),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_30),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_50),
.A2(n_61),
.B1(n_17),
.B2(n_35),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

INVx6_ASAP7_75t_L g123 ( 
.A(n_52),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_26),
.B(n_13),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_53),
.B(n_67),
.Y(n_94)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_26),
.B(n_38),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_55),
.B(n_64),
.Y(n_90)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx8_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_30),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_0),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_16),
.B(n_2),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_65),
.B(n_71),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_66),
.Y(n_105)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_16),
.B(n_2),
.Y(n_67)
);

INVx13_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_68),
.Y(n_106)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_19),
.Y(n_69)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_19),
.Y(n_70)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_16),
.B(n_4),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_72),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_16),
.B(n_4),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_34),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_19),
.B(n_5),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_27),
.C(n_35),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_30),
.Y(n_76)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_23),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_75),
.A2(n_22),
.B1(n_23),
.B2(n_20),
.Y(n_77)
);

AOI22x1_ASAP7_75t_L g165 ( 
.A1(n_77),
.A2(n_95),
.B1(n_97),
.B2(n_117),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_20),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_82),
.B(n_112),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_57),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_89),
.B(n_108),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_69),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_107),
.B1(n_118),
.B2(n_39),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_76),
.A2(n_74),
.B1(n_59),
.B2(n_42),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_41),
.A2(n_22),
.B1(n_23),
.B2(n_32),
.Y(n_97)
);

NAND2x1_ASAP7_75t_SL g161 ( 
.A(n_98),
.B(n_104),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_33),
.B1(n_37),
.B2(n_32),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_109),
.B1(n_54),
.B2(n_48),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_102),
.B(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_103),
.B(n_119),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_46),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_67),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_45),
.B(n_18),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_62),
.B(n_18),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_81),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_44),
.A2(n_17),
.B1(n_29),
.B2(n_27),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_58),
.A2(n_29),
.B1(n_34),
.B2(n_39),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_70),
.B(n_49),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_121),
.B(n_100),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_63),
.B(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_104),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_78),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_126),
.B(n_129),
.Y(n_202)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_94),
.A2(n_68),
.B(n_60),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_127),
.B(n_141),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g128 ( 
.A(n_120),
.Y(n_128)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_128),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_96),
.Y(n_129)
);

AO22x1_ASAP7_75t_SL g130 ( 
.A1(n_77),
.A2(n_63),
.B1(n_52),
.B2(n_51),
.Y(n_130)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_130),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_132),
.B(n_153),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_66),
.B1(n_43),
.B2(n_39),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_133),
.A2(n_149),
.B1(n_153),
.B2(n_140),
.Y(n_187)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_134),
.Y(n_181)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_78),
.Y(n_135)
);

INVx11_ASAP7_75t_L g178 ( 
.A(n_135),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_136),
.Y(n_183)
);

INVx5_ASAP7_75t_L g137 ( 
.A(n_106),
.Y(n_137)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_121),
.Y(n_138)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_138),
.Y(n_173)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_139),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_90),
.B(n_92),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_106),
.Y(n_144)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_144),
.Y(n_185)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_93),
.Y(n_145)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_145),
.Y(n_193)
);

AO22x1_ASAP7_75t_SL g146 ( 
.A1(n_82),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_146)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_117),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_147),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_112),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_148),
.B(n_151),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_98),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_149)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_78),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_88),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_152),
.B(n_154),
.Y(n_180)
);

A2O1A1Ixp33_ASAP7_75t_L g153 ( 
.A1(n_113),
.A2(n_9),
.B(n_83),
.C(n_81),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_79),
.B(n_87),
.C(n_114),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_155),
.B(n_162),
.Y(n_195)
);

OA22x2_ASAP7_75t_L g156 ( 
.A1(n_79),
.A2(n_87),
.B1(n_105),
.B2(n_88),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_158),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_115),
.A2(n_122),
.B1(n_86),
.B2(n_116),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_160),
.B1(n_158),
.B2(n_165),
.Y(n_175)
);

OR2x6_ASAP7_75t_L g158 ( 
.A(n_120),
.B(n_114),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_96),
.A2(n_101),
.B(n_80),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_159),
.A2(n_164),
.B(n_133),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g160 ( 
.A1(n_86),
.A2(n_122),
.B1(n_116),
.B2(n_110),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_161),
.Y(n_201)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_84),
.Y(n_163)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_163),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_80),
.A2(n_84),
.B(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_166),
.B(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_110),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_168),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_123),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_90),
.B(n_92),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_125),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_175),
.A2(n_170),
.B1(n_189),
.B2(n_207),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_179),
.B(n_196),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_182),
.B(n_156),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_138),
.A2(n_150),
.B1(n_166),
.B2(n_165),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_150),
.A2(n_165),
.B1(n_130),
.B2(n_154),
.Y(n_189)
);

BUFx2_ASAP7_75t_SL g191 ( 
.A(n_135),
.Y(n_191)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_191),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_154),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g197 ( 
.A1(n_130),
.A2(n_168),
.B1(n_158),
.B2(n_156),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_152),
.B1(n_128),
.B2(n_139),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_137),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_199),
.B(n_129),
.Y(n_226)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_134),
.Y(n_203)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_203),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_131),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_204),
.B(n_207),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_205),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_155),
.B(n_158),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_158),
.B(n_161),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_144),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_179),
.B(n_161),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_209),
.B(n_181),
.C(n_192),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_212),
.A2(n_213),
.B(n_237),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g213 ( 
.A1(n_208),
.A2(n_164),
.B(n_159),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_156),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_214),
.A2(n_183),
.B(n_190),
.Y(n_249)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_176),
.Y(n_215)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_215),
.Y(n_256)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_176),
.Y(n_216)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_216),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_174),
.B(n_143),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_217),
.B(n_223),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_219),
.B1(n_239),
.B2(n_177),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_201),
.B(n_128),
.Y(n_220)
);

NAND2xp33_ASAP7_75t_SL g255 ( 
.A(n_220),
.B(n_235),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_188),
.B(n_142),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_221),
.B(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_222),
.B(n_228),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_204),
.B(n_145),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_226),
.Y(n_248)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

OA21x2_ASAP7_75t_SL g254 ( 
.A1(n_229),
.A2(n_181),
.B(n_185),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_202),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_231),
.B(n_234),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_173),
.B(n_202),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_232),
.B(n_233),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_170),
.A2(n_206),
.B1(n_182),
.B2(n_194),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g235 ( 
.A(n_177),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_173),
.B(n_195),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_236),
.B(n_240),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_196),
.A2(n_206),
.B(n_187),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_200),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_238),
.B(n_193),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_175),
.A2(n_183),
.B1(n_194),
.B2(n_177),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_206),
.B(n_186),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_227),
.B(n_198),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_253),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_243),
.A2(n_250),
.B1(n_220),
.B2(n_229),
.Y(n_278)
);

OAI32xp33_ASAP7_75t_L g244 ( 
.A1(n_227),
.A2(n_198),
.A3(n_186),
.B1(n_193),
.B2(n_203),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_246),
.B(n_263),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_249),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_224),
.A2(n_190),
.B1(n_171),
.B2(n_199),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g252 ( 
.A1(n_212),
.A2(n_171),
.B1(n_192),
.B2(n_178),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_252),
.A2(n_214),
.B1(n_218),
.B2(n_215),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_254),
.A2(n_264),
.B(n_266),
.Y(n_285)
);

BUFx5_ASAP7_75t_L g258 ( 
.A(n_230),
.Y(n_258)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_258),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_185),
.Y(n_261)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_261),
.B(n_220),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_221),
.B(n_172),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_240),
.A2(n_172),
.B(n_178),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_226),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_232),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_213),
.A2(n_237),
.B(n_220),
.Y(n_266)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_235),
.A2(n_214),
.B(n_212),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_267),
.A2(n_223),
.B(n_216),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_246),
.B(n_225),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_268),
.B(n_271),
.Y(n_293)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_236),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_270),
.B(n_283),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_245),
.B(n_238),
.Y(n_271)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_274),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_286),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_247),
.A2(n_212),
.B1(n_211),
.B2(n_233),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_277),
.A2(n_278),
.B1(n_288),
.B2(n_261),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_245),
.B(n_217),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_279),
.B(n_287),
.Y(n_303)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_241),
.Y(n_281)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_281),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_209),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_284),
.B(n_244),
.Y(n_297)
);

OAI322xp33_ASAP7_75t_L g287 ( 
.A1(n_262),
.A2(n_210),
.A3(n_222),
.B1(n_228),
.B2(n_230),
.C1(n_265),
.C2(n_257),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_243),
.A2(n_210),
.B1(n_247),
.B2(n_257),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_283),
.C(n_253),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_290),
.B(n_275),
.C(n_286),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_282),
.A2(n_267),
.B1(n_250),
.B2(n_249),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_300),
.B1(n_285),
.B2(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_248),
.Y(n_295)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_295),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_282),
.A2(n_251),
.B1(n_252),
.B2(n_259),
.Y(n_296)
);

XNOR2x1_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_275),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_277),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_280),
.B(n_266),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_299),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_284),
.B(n_261),
.Y(n_299)
);

OAI321xp33_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_251),
.A3(n_255),
.B1(n_263),
.B2(n_259),
.C(n_256),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_281),
.B(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_302),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_306),
.B(n_316),
.Y(n_328)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_318),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_314),
.C(n_290),
.Y(n_325)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_317),
.Y(n_322)
);

AOI21x1_ASAP7_75t_SL g312 ( 
.A1(n_289),
.A2(n_285),
.B(n_264),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_312),
.A2(n_296),
.B(n_255),
.Y(n_323)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_313),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_301),
.B(n_272),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_304),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_315),
.A2(n_289),
.B1(n_291),
.B2(n_294),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_310),
.A2(n_297),
.B1(n_303),
.B2(n_272),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_323),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_325),
.A2(n_314),
.B(n_309),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_311),
.A2(n_298),
.B(n_273),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_326),
.B(n_292),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_316),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g330 ( 
.A(n_327),
.B(n_308),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_329),
.B(n_331),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_321),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_328),
.B(n_307),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_333),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_322),
.B(n_256),
.Y(n_333)
);

AOI31xp33_ASAP7_75t_SL g335 ( 
.A1(n_320),
.A2(n_312),
.A3(n_318),
.B(n_292),
.Y(n_335)
);

INVx1_ASAP7_75t_SL g341 ( 
.A(n_335),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_336),
.B(n_325),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_338),
.A2(n_341),
.B1(n_337),
.B2(n_319),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_339),
.A2(n_323),
.B1(n_273),
.B2(n_324),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_340),
.A2(n_322),
.B1(n_334),
.B2(n_333),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g346 ( 
.A1(n_342),
.A2(n_343),
.B(n_344),
.Y(n_346)
);

AOI211x1_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_324),
.B(n_338),
.C(n_299),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g347 ( 
.A1(n_345),
.A2(n_254),
.B(n_260),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_346),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_348),
.B(n_260),
.Y(n_349)
);


endmodule