module fake_jpeg_19212_n_209 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_209);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_209;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_130;
wire n_99;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_5),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_11),
.B(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

INVxp33_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_0),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_35),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_32),
.Y(n_41)
);

INVx5_ASAP7_75t_L g32 ( 
.A(n_16),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_7),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_34),
.Y(n_44)
);

BUFx2_ASAP7_75t_R g34 ( 
.A(n_25),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_36),
.B(n_17),
.Y(n_49)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_29),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_42),
.B(n_49),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_26),
.B1(n_19),
.B2(n_15),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_47),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_26),
.B1(n_19),
.B2(n_15),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_25),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_36),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_54),
.B(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_55),
.B(n_66),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_40),
.A2(n_34),
.B1(n_32),
.B2(n_24),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_56),
.A2(n_57),
.B1(n_65),
.B2(n_73),
.Y(n_92)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_32),
.B1(n_20),
.B2(n_24),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_28),
.B1(n_24),
.B2(n_20),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_58),
.A2(n_72),
.B1(n_48),
.B2(n_69),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_49),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_46),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_51),
.Y(n_60)
);

OR2x2_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_31),
.Y(n_61)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_61),
.A2(n_46),
.B1(n_39),
.B2(n_25),
.Y(n_83)
);

AOI32xp33_ASAP7_75t_L g64 ( 
.A1(n_44),
.A2(n_33),
.A3(n_37),
.B1(n_32),
.B2(n_18),
.Y(n_64)
);

AOI21xp33_ASAP7_75t_L g79 ( 
.A1(n_64),
.A2(n_47),
.B(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_48),
.A2(n_20),
.B1(n_17),
.B2(n_28),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_42),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_67),
.Y(n_78)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_45),
.B(n_35),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_74),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_L g71 ( 
.A1(n_45),
.A2(n_37),
.B1(n_36),
.B2(n_35),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_39),
.B1(n_38),
.B2(n_30),
.Y(n_89)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_72),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_18),
.B1(n_27),
.B2(n_28),
.Y(n_73)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_81),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_89),
.B1(n_90),
.B2(n_96),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_27),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_82),
.A2(n_88),
.B1(n_63),
.B2(n_87),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_53),
.Y(n_102)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_53),
.Y(n_85)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_85),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_97),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_60),
.A2(n_39),
.B1(n_30),
.B2(n_38),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_52),
.A2(n_67),
.B1(n_66),
.B2(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_64),
.B(n_23),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_91),
.B(n_95),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_93),
.Y(n_120)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_53),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_30),
.B1(n_38),
.B2(n_50),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_73),
.B(n_23),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_80),
.B(n_61),
.Y(n_98)
);

AOI221xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_8),
.B1(n_11),
.B2(n_13),
.C(n_3),
.Y(n_134)
);

OAI32xp33_ASAP7_75t_L g100 ( 
.A1(n_94),
.A2(n_70),
.A3(n_55),
.B1(n_62),
.B2(n_61),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_100),
.B(n_102),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_62),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_103),
.B(n_105),
.Y(n_138)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_56),
.B(n_57),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_86),
.A2(n_63),
.B1(n_65),
.B2(n_59),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_106),
.A2(n_118),
.B1(n_76),
.B2(n_95),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_90),
.B(n_92),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_113),
.C(n_75),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_22),
.Y(n_141)
);

A2O1A1O1Ixp25_ASAP7_75t_L g111 ( 
.A1(n_83),
.A2(n_84),
.B(n_92),
.C(n_87),
.D(n_78),
.Y(n_111)
);

A2O1A1O1Ixp25_ASAP7_75t_L g127 ( 
.A1(n_111),
.A2(n_83),
.B(n_85),
.C(n_22),
.D(n_77),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_115),
.B1(n_75),
.B2(n_93),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_38),
.C(n_50),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_88),
.Y(n_114)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_114),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_89),
.A2(n_22),
.B1(n_16),
.B2(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_116),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_84),
.B(n_25),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_117),
.B(n_77),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_86),
.A2(n_22),
.B1(n_23),
.B2(n_2),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_96),
.B(n_7),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g139 ( 
.A(n_119),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_101),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_121),
.B(n_122),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_123),
.A2(n_133),
.B1(n_114),
.B2(n_115),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_124),
.B(n_130),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_127),
.B(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g129 ( 
.A(n_107),
.B(n_9),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_129),
.B(n_132),
.Y(n_143)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_113),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_131),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_SL g135 ( 
.A(n_110),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_99),
.B(n_93),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_137),
.Y(n_142)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_140),
.Y(n_157)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_119),
.Y(n_165)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_105),
.B(n_104),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_147),
.A2(n_156),
.B(n_108),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_129),
.B(n_103),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_100),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_150),
.A2(n_151),
.B1(n_135),
.B2(n_122),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_138),
.A2(n_99),
.B1(n_102),
.B2(n_105),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_131),
.C(n_136),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_155),
.B(n_117),
.C(n_140),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_136),
.A2(n_111),
.B(n_104),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_159),
.B(n_166),
.C(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_160),
.B(n_161),
.Y(n_172)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_163),
.B1(n_164),
.B2(n_170),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_142),
.A2(n_125),
.B1(n_133),
.B2(n_127),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_144),
.A2(n_125),
.B1(n_139),
.B2(n_121),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_165),
.B(n_167),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_154),
.B(n_124),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_168),
.A2(n_6),
.B1(n_12),
.B2(n_4),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_128),
.C(n_126),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_151),
.A2(n_126),
.B1(n_1),
.B2(n_2),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_153),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_171),
.Y(n_175)
);

AOI322xp5_ASAP7_75t_SL g173 ( 
.A1(n_159),
.A2(n_146),
.A3(n_156),
.B1(n_148),
.B2(n_143),
.C1(n_157),
.C2(n_152),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_173),
.B(n_180),
.Y(n_187)
);

AOI322xp5_ASAP7_75t_L g174 ( 
.A1(n_162),
.A2(n_146),
.A3(n_143),
.B1(n_152),
.B2(n_150),
.C1(n_158),
.C2(n_8),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_174),
.B(n_170),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_158),
.C(n_8),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_177),
.B(n_181),
.C(n_163),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_6),
.C(n_12),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_179),
.A2(n_168),
.B1(n_161),
.B2(n_160),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_182),
.A2(n_189),
.B1(n_181),
.B2(n_187),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_186),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_178),
.B(n_164),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_184),
.A2(n_176),
.B(n_5),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_176),
.B(n_10),
.C(n_12),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_175),
.B(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_188),
.B(n_190),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_172),
.A2(n_180),
.B(n_177),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_172),
.B(n_4),
.Y(n_190)
);

HB1xp67_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_191),
.B(n_184),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_194),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_197),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_198),
.B(n_200),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_11),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_199),
.A2(n_191),
.B1(n_192),
.B2(n_200),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_202),
.B(n_13),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_204),
.B(n_205),
.Y(n_206)
);

AOI21x1_ASAP7_75t_L g205 ( 
.A1(n_201),
.A2(n_0),
.B(n_1),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_206),
.B(n_203),
.C(n_202),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_207),
.B(n_1),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g209 ( 
.A(n_208),
.B(n_1),
.Y(n_209)
);


endmodule