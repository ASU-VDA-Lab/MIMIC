module fake_jpeg_5466_n_14 (n_3, n_2, n_1, n_0, n_4, n_14);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_14;

wire n_13;
wire n_11;
wire n_10;
wire n_12;
wire n_8;
wire n_9;
wire n_6;
wire n_5;
wire n_7;

INVx5_ASAP7_75t_L g5 ( 
.A(n_2),
.Y(n_5)
);

NOR2xp33_ASAP7_75t_SL g6 ( 
.A(n_3),
.B(n_4),
.Y(n_6)
);

OAI21xp5_ASAP7_75t_L g7 ( 
.A1(n_6),
.A2(n_5),
.B(n_1),
.Y(n_7)
);

MAJIxp5_ASAP7_75t_L g11 ( 
.A(n_7),
.B(n_5),
.C(n_0),
.Y(n_11)
);

OAI22xp5_ASAP7_75t_L g8 ( 
.A1(n_6),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_8),
.B(n_9),
.Y(n_12)
);

INVx13_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

AOI321xp33_ASAP7_75t_SL g10 ( 
.A1(n_7),
.A2(n_5),
.A3(n_6),
.B1(n_3),
.B2(n_4),
.C(n_0),
.Y(n_10)
);

XOR2x2_ASAP7_75t_L g13 ( 
.A(n_10),
.B(n_11),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_12),
.B1(n_11),
.B2(n_5),
.Y(n_14)
);


endmodule