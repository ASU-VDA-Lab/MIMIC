module fake_jpeg_3140_n_74 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_74);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_74;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_10;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_44;
wire n_28;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_43;
wire n_29;
wire n_50;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_1),
.B(n_6),
.Y(n_9)
);

BUFx8_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

INVx11_ASAP7_75t_SL g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_1),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx6_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_9),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_13),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g29 ( 
.A(n_21),
.B(n_25),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_11),
.B(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_13),
.B(n_5),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_24),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_16),
.B(n_7),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_10),
.B(n_19),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_12),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_18),
.C(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_30),
.B(n_37),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_24),
.Y(n_32)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_20),
.B(n_14),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_44),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_30),
.A2(n_26),
.B1(n_15),
.B2(n_17),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_41),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_37),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_33),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_25),
.B1(n_34),
.B2(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_48),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_42),
.B(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_54),
.B(n_31),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_39),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_56),
.B(n_44),
.C(n_46),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_52),
.Y(n_57)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVxp33_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_59),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_49),
.C(n_58),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_60),
.Y(n_65)
);

OA21x2_ASAP7_75t_SL g69 ( 
.A1(n_65),
.A2(n_66),
.B(n_40),
.Y(n_69)
);

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_61),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_64),
.B1(n_53),
.B2(n_40),
.Y(n_68)
);

NOR3xp33_ASAP7_75t_L g70 ( 
.A(n_68),
.B(n_53),
.C(n_38),
.Y(n_70)
);

OA21x2_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_15),
.B(n_22),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g72 ( 
.A1(n_70),
.A2(n_71),
.B(n_17),
.Y(n_72)
);

BUFx24_ASAP7_75t_SL g73 ( 
.A(n_72),
.Y(n_73)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_26),
.Y(n_74)
);


endmodule