module fake_jpeg_24088_n_105 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_105);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_105;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx10_ASAP7_75t_L g11 ( 
.A(n_10),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_SL g14 ( 
.A(n_2),
.Y(n_14)
);

AND2x2_ASAP7_75t_SL g15 ( 
.A(n_3),
.B(n_8),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_1),
.B(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx8_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_9),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_22),
.Y(n_24)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_24),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_22),
.Y(n_25)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp67_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_0),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_26),
.B(n_15),
.Y(n_42)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_27),
.B(n_31),
.Y(n_36)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_32),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_34),
.B(n_12),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_27),
.B(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_37),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_SL g38 ( 
.A1(n_32),
.A2(n_15),
.B(n_14),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_26),
.C(n_12),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_21),
.Y(n_47)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_23),
.Y(n_62)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_49),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_47),
.B(n_48),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_38),
.B(n_25),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_35),
.A2(n_31),
.B1(n_16),
.B2(n_28),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_50),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_32),
.C(n_28),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_43),
.C(n_39),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_43),
.B(n_17),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

OAI22x1_ASAP7_75t_L g54 ( 
.A1(n_42),
.A2(n_30),
.B1(n_29),
.B2(n_25),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_57),
.B1(n_45),
.B2(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_55),
.Y(n_60)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_0),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_33),
.A2(n_21),
.B1(n_17),
.B2(n_18),
.Y(n_57)
);

INVxp67_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_58),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_35),
.A2(n_16),
.B1(n_19),
.B2(n_20),
.Y(n_59)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_59),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_62),
.B(n_68),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_63),
.A2(n_58),
.B(n_55),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_41),
.B(n_39),
.Y(n_65)
);

AO21x1_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_71),
.B(n_24),
.Y(n_76)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_73),
.Y(n_84)
);

NAND3xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_54),
.C(n_44),
.Y(n_73)
);

OAI21xp33_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_51),
.B(n_3),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_74),
.A2(n_81),
.B(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_75),
.Y(n_83)
);

AOI221xp5_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_79),
.B1(n_69),
.B2(n_67),
.C(n_24),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_60),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_78),
.Y(n_82)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_63),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_80),
.Y(n_85)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

XOR2x2_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_62),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_SL g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_88),
.A2(n_81),
.B1(n_74),
.B2(n_77),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_90),
.B(n_93),
.C(n_82),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_86),
.A2(n_79),
.B1(n_61),
.B2(n_30),
.Y(n_91)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_84),
.A2(n_29),
.B1(n_19),
.B2(n_20),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_83),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g93 ( 
.A1(n_87),
.A2(n_20),
.B(n_1),
.C(n_5),
.D(n_6),
.Y(n_93)
);

XNOR2x1_ASAP7_75t_L g94 ( 
.A(n_89),
.B(n_85),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_85),
.B(n_93),
.Y(n_99)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_97),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_95),
.B(n_96),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_101),
.A2(n_102),
.B1(n_98),
.B2(n_7),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_100),
.B(n_4),
.Y(n_102)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_6),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_8),
.Y(n_105)
);


endmodule