module fake_jpeg_29147_n_322 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_322);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_322;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_1),
.B(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_7),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_6),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_12),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_15),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_8),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_47),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_4),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_48),
.B(n_50),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_25),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g113 ( 
.A(n_49),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_16),
.B(n_40),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_17),
.B(n_4),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_51),
.B(n_86),
.Y(n_136)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_4),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_63),
.Y(n_106)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_58),
.B(n_59),
.Y(n_104)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_20),
.B(n_5),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_60),
.B(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_39),
.A2(n_5),
.B1(n_6),
.B2(n_9),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_61),
.A2(n_88),
.B1(n_89),
.B2(n_41),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_62),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_5),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_24),
.Y(n_64)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_65),
.Y(n_126)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_21),
.B(n_44),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_21),
.B(n_44),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_68),
.B(n_71),
.Y(n_109)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_69),
.Y(n_107)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_70),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_23),
.B(n_14),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

INVx5_ASAP7_75t_L g127 ( 
.A(n_72),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_23),
.B(n_14),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_77),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx5_ASAP7_75t_L g129 ( 
.A(n_74),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_37),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_43),
.Y(n_76)
);

BUFx12f_ASAP7_75t_L g124 ( 
.A(n_76),
.Y(n_124)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_9),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_78),
.B(n_83),
.Y(n_122)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_79),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_25),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g94 ( 
.A(n_80),
.Y(n_94)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_81),
.Y(n_134)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

CKINVDCx9p33_ASAP7_75t_R g121 ( 
.A(n_82),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_45),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_45),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_84),
.B(n_85),
.Y(n_133)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_32),
.Y(n_86)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_87),
.Y(n_96)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_26),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_53),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_91),
.B(n_102),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_82),
.B1(n_70),
.B2(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_92),
.A2(n_95),
.B1(n_110),
.B2(n_111),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_46),
.A2(n_29),
.B1(n_27),
.B2(n_39),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_54),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_103),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_69),
.A2(n_41),
.B1(n_28),
.B2(n_18),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_62),
.A2(n_29),
.B1(n_38),
.B2(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_41),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_112),
.B(n_118),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_65),
.B(n_19),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_88),
.A2(n_28),
.B1(n_38),
.B2(n_19),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_119),
.A2(n_132),
.B1(n_112),
.B2(n_96),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_72),
.B(n_18),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_106),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_87),
.B(n_34),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_128),
.B(n_130),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_83),
.B(n_34),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_74),
.A2(n_36),
.B1(n_28),
.B2(n_12),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_75),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_94),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_121),
.A2(n_76),
.B1(n_83),
.B2(n_28),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_138),
.A2(n_146),
.B1(n_150),
.B2(n_160),
.Y(n_174)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_124),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_139),
.Y(n_184)
);

OA22x2_ASAP7_75t_L g140 ( 
.A1(n_125),
.A2(n_61),
.B1(n_10),
.B2(n_11),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_153),
.B1(n_127),
.B2(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_SL g141 ( 
.A(n_113),
.Y(n_141)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_141),
.Y(n_201)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

INVx11_ASAP7_75t_L g144 ( 
.A(n_93),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g181 ( 
.A(n_144),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_10),
.B1(n_11),
.B2(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_159),
.Y(n_178)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_125),
.Y(n_148)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_148),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_149),
.B(n_155),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_136),
.A2(n_133),
.B1(n_114),
.B2(n_118),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_113),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_151),
.B(n_156),
.Y(n_172)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_114),
.Y(n_152)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_152),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_107),
.Y(n_154)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_154),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_106),
.B(n_123),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_104),
.B(n_117),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_122),
.B(n_107),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g197 ( 
.A1(n_157),
.A2(n_158),
.B(n_164),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_97),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_116),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_120),
.A2(n_131),
.B1(n_100),
.B2(n_99),
.Y(n_160)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_109),
.B(n_108),
.Y(n_163)
);

NAND3xp33_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_94),
.C(n_101),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_96),
.A2(n_97),
.B(n_116),
.Y(n_164)
);

INVx4_ASAP7_75t_SL g165 ( 
.A(n_93),
.Y(n_165)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_105),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_166),
.B(n_168),
.Y(n_187)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_90),
.B(n_98),
.C(n_126),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_98),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_169),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_127),
.A2(n_129),
.B1(n_126),
.B2(n_124),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_171),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_94),
.B(n_124),
.Y(n_175)
);

OR2x2_ASAP7_75t_L g205 ( 
.A(n_175),
.B(n_186),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_160),
.B1(n_140),
.B2(n_169),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_182),
.B(n_191),
.Y(n_209)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_152),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_183),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_161),
.A2(n_101),
.B1(n_99),
.B2(n_100),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_170),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVxp33_ASAP7_75t_L g220 ( 
.A(n_190),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_163),
.B(n_137),
.Y(n_191)
);

BUFx2_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_193),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_161),
.B(n_149),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_158),
.C(n_141),
.Y(n_207)
);

AOI32xp33_ASAP7_75t_L g196 ( 
.A1(n_168),
.A2(n_157),
.A3(n_155),
.B1(n_150),
.B2(n_140),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_199),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_SL g199 ( 
.A(n_156),
.B(n_157),
.Y(n_199)
);

AO22x2_ASAP7_75t_L g202 ( 
.A1(n_190),
.A2(n_140),
.B1(n_145),
.B2(n_148),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_202),
.B(n_223),
.Y(n_238)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_195),
.Y(n_203)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_203),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_216),
.B1(n_217),
.B2(n_200),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_192),
.B(n_162),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_210),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_207),
.B(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_186),
.B(n_158),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_208),
.B(n_177),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_192),
.B(n_165),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_198),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_221),
.Y(n_241)
);

BUFx6f_ASAP7_75t_L g215 ( 
.A(n_180),
.Y(n_215)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_179),
.A2(n_139),
.B1(n_144),
.B2(n_194),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_174),
.A2(n_187),
.B1(n_200),
.B2(n_197),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_175),
.C(n_178),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_172),
.B(n_176),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_198),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_222),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_184),
.B(n_188),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_177),
.B(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_225),
.Y(n_260)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_210),
.A2(n_206),
.B(n_205),
.C(n_220),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_226),
.A2(n_202),
.B(n_218),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_231),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_205),
.A2(n_201),
.B(n_188),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_229),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_224),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_234),
.B(n_235),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_209),
.B(n_208),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_203),
.Y(n_236)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_212),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_239),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_212),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_217),
.B(n_189),
.Y(n_240)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_240),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_219),
.A2(n_201),
.B(n_184),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_243),
.Y(n_261)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_215),
.Y(n_244)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_244),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_204),
.B1(n_216),
.B2(n_238),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_238),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_230),
.B(n_211),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_249),
.B(n_251),
.C(n_254),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_218),
.B1(n_202),
.B2(n_207),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_L g263 ( 
.A1(n_250),
.A2(n_225),
.B(n_227),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_242),
.B(n_202),
.Y(n_251)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_252),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_202),
.C(n_180),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_226),
.B(n_183),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_243),
.B(n_173),
.C(n_214),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_262),
.A2(n_263),
.B1(n_271),
.B2(n_241),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_248),
.B(n_234),
.Y(n_264)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_264),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_246),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_236),
.Y(n_277)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_257),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_258),
.A2(n_250),
.B(n_254),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g289 ( 
.A1(n_269),
.A2(n_274),
.B(n_276),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_256),
.B1(n_247),
.B2(n_258),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_253),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_231),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_272),
.B(n_275),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_259),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_260),
.B(n_230),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_251),
.Y(n_276)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_277),
.Y(n_297)
);

A2O1A1Ixp33_ASAP7_75t_L g278 ( 
.A1(n_266),
.A2(n_226),
.B(n_229),
.C(n_261),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_278),
.B(n_281),
.Y(n_295)
);

XNOR2x1_ASAP7_75t_L g279 ( 
.A(n_273),
.B(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_279),
.B(n_284),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_265),
.B(n_249),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_273),
.B(n_241),
.C(n_235),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_283),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_232),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_274),
.B(n_232),
.C(n_214),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_285),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_276),
.B(n_173),
.C(n_239),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_286),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_264),
.B(n_237),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_287),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_280),
.A2(n_263),
.B1(n_271),
.B2(n_262),
.Y(n_291)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_291),
.Y(n_301)
);

BUFx24_ASAP7_75t_SL g293 ( 
.A(n_281),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_293),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g298 ( 
.A(n_278),
.Y(n_298)
);

NOR3xp33_ASAP7_75t_SL g303 ( 
.A(n_298),
.B(n_275),
.C(n_272),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_290),
.A2(n_289),
.B(n_266),
.Y(n_300)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_300),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_284),
.C(n_285),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_302),
.B(n_303),
.Y(n_311)
);

AND2x4_ASAP7_75t_L g304 ( 
.A(n_295),
.B(n_279),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_304),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_296),
.A2(n_269),
.B1(n_282),
.B2(n_286),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_305),
.A2(n_294),
.B1(n_292),
.B2(n_270),
.Y(n_307)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_307),
.B(n_299),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_301),
.A2(n_297),
.B1(n_267),
.B2(n_268),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_310),
.Y(n_315)
);

AOI322xp5_ASAP7_75t_L g312 ( 
.A1(n_308),
.A2(n_303),
.A3(n_304),
.B1(n_306),
.B2(n_302),
.C1(n_288),
.C2(n_244),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_312),
.A2(n_313),
.B(n_314),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_233),
.Y(n_314)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_315),
.A2(n_309),
.B(n_304),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_316),
.B(n_309),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_318),
.A2(n_317),
.B(n_233),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_319),
.A2(n_181),
.B(n_215),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_320),
.A2(n_181),
.B1(n_212),
.B2(n_193),
.Y(n_321)
);

OR2x2_ASAP7_75t_L g322 ( 
.A(n_321),
.B(n_181),
.Y(n_322)
);


endmodule