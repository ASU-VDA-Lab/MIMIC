module fake_ariane_1574_n_934 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_934);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_934;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_913;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_878;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_908;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_906;
wire n_416;
wire n_283;
wire n_919;
wire n_525;
wire n_187;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_817;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_924;
wire n_927;
wire n_781;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_634;
wire n_391;
wire n_349;
wire n_756;
wire n_466;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_897;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_891;
wire n_737;
wire n_885;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_917;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_905;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_898;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_926;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_900;
wire n_883;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_801;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_818;
wire n_500;
wire n_665;
wire n_731;
wire n_336;
wire n_754;
wire n_779;
wire n_871;
wire n_315;
wire n_903;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_879;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_320;
wire n_309;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_721;
wire n_600;
wire n_481;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_928;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_901;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_894;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_677;
wire n_614;
wire n_604;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_874;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_694;
wire n_884;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_921;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_929;
wire n_206;
wire n_352;
wire n_538;
wire n_899;
wire n_920;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_455;
wire n_429;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_887;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_904;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_715;
wire n_512;
wire n_889;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_321;
wire n_221;
wire n_911;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_877;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_181;
wire n_723;
wire n_617;
wire n_658;
wire n_616;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_683;
wire n_601;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_907;
wire n_235;
wire n_881;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_910;
wire n_290;
wire n_527;
wire n_747;
wire n_741;
wire n_772;
wire n_847;
wire n_371;
wire n_845;
wire n_888;
wire n_199;
wire n_918;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_708;
wire n_308;
wire n_551;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_922;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_851;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_890;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_896;
wire n_409;
wire n_930;
wire n_519;
wire n_902;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_872;
wire n_933;
wire n_916;
wire n_254;
wire n_596;
wire n_912;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_915;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_544;
wire n_540;
wire n_216;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_179;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_895;
wire n_659;
wire n_583;
wire n_509;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_875;
wire n_669;
wire n_785;
wire n_827;
wire n_931;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_880;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_873;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_925;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_892;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_923;
wire n_250;
wire n_932;
wire n_773;
wire n_882;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_909;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_893;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_886;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

CKINVDCx14_ASAP7_75t_R g177 ( 
.A(n_2),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_112),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_56),
.Y(n_179)
);

BUFx2_ASAP7_75t_L g180 ( 
.A(n_90),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_58),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_110),
.Y(n_182)
);

BUFx10_ASAP7_75t_L g183 ( 
.A(n_43),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_100),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_143),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_49),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_87),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_72),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_82),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_101),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_36),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_148),
.Y(n_193)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_103),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_16),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_22),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_0),
.Y(n_197)
);

BUFx8_ASAP7_75t_SL g198 ( 
.A(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_60),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_106),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_70),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_16),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_76),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_129),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_131),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_14),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_120),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_64),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_126),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_108),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_111),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_40),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_149),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_65),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_119),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_61),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_116),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_7),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_33),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_134),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_136),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_104),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_96),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_46),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_160),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_26),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_63),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_151),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_137),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_53),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_94),
.Y(n_234)
);

BUFx2_ASAP7_75t_L g235 ( 
.A(n_133),
.Y(n_235)
);

INVx2_ASAP7_75t_SL g236 ( 
.A(n_109),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_22),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_170),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_39),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_113),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_132),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_125),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_48),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_138),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_150),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_144),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g248 ( 
.A(n_23),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_145),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_92),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_165),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_10),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_172),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_5),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_3),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_127),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_169),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_57),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_163),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_97),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_93),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_105),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_121),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_23),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_154),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_88),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_86),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_153),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_107),
.Y(n_269)
);

INVx1_ASAP7_75t_SL g270 ( 
.A(n_102),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_175),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_176),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_114),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_66),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_10),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_25),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_166),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_117),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_71),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_177),
.Y(n_280)
);

INVx5_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_177),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_252),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_252),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_244),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_248),
.B(n_0),
.Y(n_287)
);

INVx3_ASAP7_75t_L g288 ( 
.A(n_252),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_180),
.B(n_235),
.Y(n_289)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_244),
.Y(n_290)
);

AND2x4_ASAP7_75t_L g291 ( 
.A(n_243),
.B(n_1),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_207),
.B(n_1),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_220),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_259),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_244),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_241),
.B(n_31),
.Y(n_297)
);

INVx5_ASAP7_75t_L g298 ( 
.A(n_271),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_184),
.B(n_2),
.Y(n_299)
);

INVx3_ASAP7_75t_L g300 ( 
.A(n_252),
.Y(n_300)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

BUFx3_ASAP7_75t_L g302 ( 
.A(n_259),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_194),
.B(n_3),
.Y(n_303)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_189),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_254),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_191),
.B(n_4),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g307 ( 
.A(n_198),
.B(n_32),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_192),
.Y(n_309)
);

INVx5_ASAP7_75t_L g310 ( 
.A(n_271),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_195),
.Y(n_311)
);

BUFx8_ASAP7_75t_SL g312 ( 
.A(n_196),
.Y(n_312)
);

BUFx6f_ASAP7_75t_L g313 ( 
.A(n_194),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g314 ( 
.A(n_232),
.Y(n_314)
);

INVx5_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_199),
.B(n_4),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_203),
.B(n_5),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_204),
.B(n_6),
.Y(n_318)
);

INVx5_ASAP7_75t_L g319 ( 
.A(n_183),
.Y(n_319)
);

INVx5_ASAP7_75t_L g320 ( 
.A(n_183),
.Y(n_320)
);

INVx3_ASAP7_75t_L g321 ( 
.A(n_188),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_208),
.Y(n_322)
);

INVx5_ASAP7_75t_L g323 ( 
.A(n_188),
.Y(n_323)
);

AND2x4_ASAP7_75t_L g324 ( 
.A(n_211),
.B(n_6),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g325 ( 
.A(n_263),
.B(n_7),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_255),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_214),
.B(n_8),
.Y(n_327)
);

INVx2_ASAP7_75t_L g328 ( 
.A(n_224),
.Y(n_328)
);

INVx2_ASAP7_75t_SL g329 ( 
.A(n_264),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_228),
.B(n_8),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_234),
.B(n_9),
.Y(n_331)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_211),
.B(n_9),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_253),
.B(n_11),
.Y(n_334)
);

HB1xp67_ASAP7_75t_L g335 ( 
.A(n_197),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_313),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g337 ( 
.A(n_292),
.B(n_202),
.Y(n_337)
);

AO22x2_ASAP7_75t_L g338 ( 
.A1(n_293),
.A2(n_270),
.B1(n_216),
.B2(n_279),
.Y(n_338)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_288),
.Y(n_339)
);

AND2x4_ASAP7_75t_L g340 ( 
.A(n_321),
.B(n_260),
.Y(n_340)
);

OR2x2_ASAP7_75t_L g341 ( 
.A(n_321),
.B(n_206),
.Y(n_341)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_293),
.A2(n_276),
.B1(n_237),
.B2(n_266),
.Y(n_342)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_286),
.Y(n_343)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_SL g345 ( 
.A1(n_297),
.A2(n_274),
.B1(n_261),
.B2(n_267),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_321),
.B(n_186),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_289),
.A2(n_325),
.B1(n_287),
.B2(n_282),
.Y(n_347)
);

AO22x2_ASAP7_75t_L g348 ( 
.A1(n_287),
.A2(n_268),
.B1(n_223),
.B2(n_229),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_313),
.Y(n_349)
);

AO22x2_ASAP7_75t_L g350 ( 
.A1(n_325),
.A2(n_291),
.B1(n_324),
.B2(n_303),
.Y(n_350)
);

OAI22xp33_ASAP7_75t_L g351 ( 
.A1(n_307),
.A2(n_275),
.B1(n_190),
.B2(n_187),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_319),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_280),
.A2(n_200),
.B1(n_277),
.B2(n_273),
.Y(n_353)
);

OAI22xp33_ASAP7_75t_L g354 ( 
.A1(n_280),
.A2(n_278),
.B1(n_272),
.B2(n_269),
.Y(n_354)
);

OAI22xp33_ASAP7_75t_L g355 ( 
.A1(n_282),
.A2(n_265),
.B1(n_262),
.B2(n_258),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g356 ( 
.A1(n_306),
.A2(n_317),
.B1(n_327),
.B2(n_318),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_319),
.B(n_178),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_R g358 ( 
.A1(n_299),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_12),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_311),
.A2(n_257),
.B1(n_256),
.B2(n_251),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_313),
.Y(n_361)
);

AO22x2_ASAP7_75t_L g362 ( 
.A1(n_291),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_362)
);

HB1xp67_ASAP7_75t_L g363 ( 
.A(n_285),
.Y(n_363)
);

OAI22xp33_ASAP7_75t_SL g364 ( 
.A1(n_330),
.A2(n_250),
.B1(n_249),
.B2(n_247),
.Y(n_364)
);

OR2x6_ASAP7_75t_L g365 ( 
.A(n_329),
.B(n_15),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g366 ( 
.A1(n_291),
.A2(n_246),
.B1(n_245),
.B2(n_242),
.Y(n_366)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_319),
.B(n_320),
.Y(n_367)
);

OAI22xp33_ASAP7_75t_L g368 ( 
.A1(n_319),
.A2(n_240),
.B1(n_239),
.B2(n_238),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_319),
.B(n_179),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_320),
.B(n_181),
.Y(n_370)
);

AND2x6_ASAP7_75t_L g371 ( 
.A(n_303),
.B(n_34),
.Y(n_371)
);

INVx2_ASAP7_75t_L g372 ( 
.A(n_288),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_312),
.A2(n_233),
.B1(n_231),
.B2(n_230),
.Y(n_373)
);

OR2x2_ASAP7_75t_L g374 ( 
.A(n_329),
.B(n_17),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_320),
.B(n_182),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_303),
.A2(n_324),
.B1(n_333),
.B2(n_334),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_300),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_313),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_L g379 ( 
.A1(n_324),
.A2(n_227),
.B1(n_226),
.B2(n_225),
.Y(n_379)
);

OAI22xp33_ASAP7_75t_L g380 ( 
.A1(n_320),
.A2(n_222),
.B1(n_221),
.B2(n_219),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_300),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_333),
.A2(n_218),
.B1(n_217),
.B2(n_215),
.Y(n_382)
);

OAI22xp33_ASAP7_75t_L g383 ( 
.A1(n_320),
.A2(n_213),
.B1(n_212),
.B2(n_210),
.Y(n_383)
);

CKINVDCx6p67_ASAP7_75t_R g384 ( 
.A(n_323),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_300),
.Y(n_385)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_323),
.A2(n_209),
.B1(n_205),
.B2(n_201),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_283),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_285),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_283),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_284),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_323),
.B(n_185),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_284),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_290),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_295),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_393),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_351),
.B(n_316),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_354),
.B(n_355),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_353),
.Y(n_398)
);

INVx4_ASAP7_75t_L g399 ( 
.A(n_384),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_339),
.Y(n_400)
);

AND2x4_ASAP7_75t_L g401 ( 
.A(n_388),
.B(n_323),
.Y(n_401)
);

CKINVDCx16_ASAP7_75t_R g402 ( 
.A(n_346),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_323),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_350),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_337),
.B(n_295),
.Y(n_405)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_343),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_344),
.Y(n_407)
);

INVx2_ASAP7_75t_SL g408 ( 
.A(n_341),
.Y(n_408)
);

XOR2x2_ASAP7_75t_L g409 ( 
.A(n_373),
.B(n_312),
.Y(n_409)
);

BUFx8_ASAP7_75t_L g410 ( 
.A(n_359),
.Y(n_410)
);

AND2x4_ASAP7_75t_L g411 ( 
.A(n_388),
.B(n_302),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_372),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_363),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_348),
.B(n_338),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_377),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_381),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_385),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_348),
.B(n_338),
.Y(n_418)
);

INVx2_ASAP7_75t_L g419 ( 
.A(n_336),
.Y(n_419)
);

OR2x2_ASAP7_75t_SL g420 ( 
.A(n_358),
.B(n_294),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_394),
.B(n_302),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_336),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_394),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_356),
.B(n_314),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g425 ( 
.A(n_382),
.B(n_314),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_349),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_349),
.Y(n_427)
);

NOR2xp67_ASAP7_75t_L g428 ( 
.A(n_360),
.B(n_315),
.Y(n_428)
);

NAND2x1p5_ASAP7_75t_L g429 ( 
.A(n_374),
.B(n_304),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_361),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_379),
.B(n_340),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_387),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_350),
.B(n_305),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_361),
.Y(n_434)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_347),
.B(n_326),
.Y(n_435)
);

AND2x6_ASAP7_75t_L g436 ( 
.A(n_367),
.B(n_304),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g437 ( 
.A(n_340),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_366),
.B(n_314),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_378),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_365),
.Y(n_440)
);

CKINVDCx16_ASAP7_75t_R g441 ( 
.A(n_365),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_375),
.B(n_315),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_375),
.B(n_315),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_378),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_389),
.Y(n_445)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_369),
.B(n_326),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_371),
.B(n_332),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_390),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_392),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_370),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_392),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_343),
.Y(n_452)
);

BUFx2_ASAP7_75t_L g453 ( 
.A(n_362),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

AND2x2_ASAP7_75t_L g455 ( 
.A(n_362),
.B(n_326),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_371),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_371),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_371),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_352),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_391),
.Y(n_460)
);

AND2x2_ASAP7_75t_L g461 ( 
.A(n_357),
.B(n_309),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_345),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_342),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_386),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_368),
.B(n_380),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_383),
.B(n_332),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g467 ( 
.A(n_358),
.B(n_309),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g468 ( 
.A(n_364),
.B(n_193),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_393),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_393),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_354),
.B(n_315),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_449),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_433),
.B(n_322),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_451),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_404),
.B(n_322),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_408),
.B(n_315),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_422),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_396),
.B(n_331),
.Y(n_478)
);

BUFx6f_ASAP7_75t_SL g479 ( 
.A(n_399),
.Y(n_479)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_456),
.A2(n_328),
.B(n_301),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_419),
.Y(n_481)
);

AND2x2_ASAP7_75t_L g482 ( 
.A(n_404),
.B(n_435),
.Y(n_482)
);

OAI21xp5_ASAP7_75t_L g483 ( 
.A1(n_457),
.A2(n_328),
.B(n_301),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_455),
.B(n_290),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_427),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_413),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_426),
.Y(n_487)
);

INVx2_ASAP7_75t_SL g488 ( 
.A(n_411),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_430),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_434),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_439),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_332),
.Y(n_492)
);

BUFx3_ASAP7_75t_L g493 ( 
.A(n_411),
.Y(n_493)
);

AND2x2_ASAP7_75t_L g494 ( 
.A(n_405),
.B(n_290),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_406),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_402),
.Y(n_496)
);

BUFx4f_ASAP7_75t_L g497 ( 
.A(n_436),
.Y(n_497)
);

BUFx6f_ASAP7_75t_L g498 ( 
.A(n_406),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_301),
.Y(n_499)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_437),
.B(n_332),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_436),
.Y(n_501)
);

AND2x2_ASAP7_75t_L g502 ( 
.A(n_429),
.B(n_332),
.Y(n_502)
);

INVx2_ASAP7_75t_SL g503 ( 
.A(n_401),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_444),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_429),
.B(n_17),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_431),
.B(n_18),
.Y(n_506)
);

INVx2_ASAP7_75t_L g507 ( 
.A(n_395),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_431),
.B(n_18),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_396),
.B(n_281),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_421),
.B(n_446),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_458),
.A2(n_298),
.B(n_281),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_421),
.B(n_286),
.Y(n_512)
);

BUFx3_ASAP7_75t_L g513 ( 
.A(n_436),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_453),
.B(n_19),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g515 ( 
.A(n_465),
.B(n_281),
.Y(n_515)
);

BUFx6f_ASAP7_75t_L g516 ( 
.A(n_406),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_462),
.B(n_403),
.Y(n_517)
);

AND3x1_ASAP7_75t_SL g518 ( 
.A(n_420),
.B(n_463),
.C(n_441),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_403),
.B(n_286),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_409),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_469),
.Y(n_521)
);

AND2x2_ASAP7_75t_SL g522 ( 
.A(n_438),
.B(n_286),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_424),
.B(n_19),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_436),
.Y(n_524)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_450),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_470),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_465),
.B(n_281),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_436),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_464),
.B(n_20),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_432),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_423),
.B(n_296),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_448),
.Y(n_533)
);

INVxp67_ASAP7_75t_L g534 ( 
.A(n_424),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_440),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_425),
.B(n_20),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_400),
.Y(n_537)
);

HB1xp67_ASAP7_75t_L g538 ( 
.A(n_401),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_432),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_423),
.B(n_21),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_398),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_407),
.Y(n_542)
);

AND2x2_ASAP7_75t_SL g543 ( 
.A(n_447),
.B(n_296),
.Y(n_543)
);

BUFx6f_ASAP7_75t_L g544 ( 
.A(n_452),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_412),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_397),
.B(n_21),
.Y(n_546)
);

INVxp67_ASAP7_75t_L g547 ( 
.A(n_410),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_454),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_399),
.B(n_24),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_447),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_415),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g552 ( 
.A(n_460),
.B(n_416),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_410),
.Y(n_553)
);

INVx4_ASAP7_75t_L g554 ( 
.A(n_417),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_428),
.Y(n_555)
);

INVx4_ASAP7_75t_L g556 ( 
.A(n_459),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_466),
.B(n_471),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_474),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_474),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_517),
.B(n_466),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_524),
.Y(n_561)
);

OR2x2_ASAP7_75t_L g562 ( 
.A(n_486),
.B(n_418),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_553),
.B(n_442),
.Y(n_563)
);

AND2x2_ASAP7_75t_L g564 ( 
.A(n_482),
.B(n_414),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_517),
.B(n_443),
.Y(n_565)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_496),
.Y(n_566)
);

AND2x6_ASAP7_75t_L g567 ( 
.A(n_501),
.B(n_296),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_490),
.Y(n_568)
);

NOR2x1_ASAP7_75t_L g569 ( 
.A(n_493),
.B(n_468),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_479),
.Y(n_570)
);

AND2x4_ASAP7_75t_L g571 ( 
.A(n_482),
.B(n_25),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_490),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

HB1xp67_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_491),
.Y(n_575)
);

BUFx8_ASAP7_75t_SL g576 ( 
.A(n_553),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_510),
.B(n_26),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_524),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_499),
.B(n_27),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_485),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_478),
.B(n_27),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_499),
.B(n_28),
.Y(n_582)
);

INVx3_ASAP7_75t_L g583 ( 
.A(n_524),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g584 ( 
.A(n_529),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_521),
.Y(n_585)
);

INVx5_ASAP7_75t_L g586 ( 
.A(n_524),
.Y(n_586)
);

INVxp67_ASAP7_75t_L g587 ( 
.A(n_538),
.Y(n_587)
);

AND2x4_ASAP7_75t_L g588 ( 
.A(n_493),
.B(n_28),
.Y(n_588)
);

AND2x4_ASAP7_75t_L g589 ( 
.A(n_488),
.B(n_29),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_506),
.B(n_29),
.Y(n_590)
);

AND2x2_ASAP7_75t_L g591 ( 
.A(n_475),
.B(n_30),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g592 ( 
.A(n_506),
.B(n_30),
.Y(n_592)
);

AND2x2_ASAP7_75t_L g593 ( 
.A(n_475),
.B(n_296),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

NAND2x1p5_ASAP7_75t_L g595 ( 
.A(n_497),
.B(n_310),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_521),
.Y(n_596)
);

OR2x6_ASAP7_75t_L g597 ( 
.A(n_547),
.B(n_308),
.Y(n_597)
);

BUFx6f_ASAP7_75t_L g598 ( 
.A(n_528),
.Y(n_598)
);

OR2x6_ASAP7_75t_L g599 ( 
.A(n_529),
.B(n_308),
.Y(n_599)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_536),
.B(n_281),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_536),
.B(n_298),
.Y(n_601)
);

BUFx6f_ASAP7_75t_L g602 ( 
.A(n_528),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_528),
.Y(n_603)
);

NOR2xp67_ASAP7_75t_L g604 ( 
.A(n_531),
.B(n_35),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_488),
.B(n_37),
.Y(n_605)
);

INVx3_ASAP7_75t_L g606 ( 
.A(n_528),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_528),
.Y(n_608)
);

OR2x6_ASAP7_75t_L g609 ( 
.A(n_529),
.B(n_308),
.Y(n_609)
);

NAND2xp5_ASAP7_75t_L g610 ( 
.A(n_508),
.B(n_308),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_485),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_495),
.Y(n_612)
);

BUFx3_ASAP7_75t_L g613 ( 
.A(n_541),
.Y(n_613)
);

OR2x6_ASAP7_75t_L g614 ( 
.A(n_501),
.B(n_38),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_508),
.B(n_298),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_489),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_477),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_489),
.Y(n_618)
);

AND2x2_ASAP7_75t_L g619 ( 
.A(n_473),
.B(n_298),
.Y(n_619)
);

OR2x6_ASAP7_75t_L g620 ( 
.A(n_513),
.B(n_41),
.Y(n_620)
);

BUFx6f_ASAP7_75t_L g621 ( 
.A(n_495),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_531),
.B(n_298),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_473),
.B(n_310),
.Y(n_623)
);

OR2x6_ASAP7_75t_L g624 ( 
.A(n_513),
.B(n_42),
.Y(n_624)
);

NAND2x1p5_ASAP7_75t_L g625 ( 
.A(n_586),
.B(n_497),
.Y(n_625)
);

NAND2x1p5_ASAP7_75t_L g626 ( 
.A(n_586),
.B(n_497),
.Y(n_626)
);

BUFx6f_ASAP7_75t_L g627 ( 
.A(n_612),
.Y(n_627)
);

BUFx6f_ASAP7_75t_L g628 ( 
.A(n_612),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_576),
.Y(n_629)
);

INVx1_ASAP7_75t_SL g630 ( 
.A(n_566),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_613),
.Y(n_631)
);

AOI22xp33_ASAP7_75t_L g632 ( 
.A1(n_581),
.A2(n_546),
.B1(n_522),
.B2(n_523),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g633 ( 
.A(n_565),
.B(n_534),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_560),
.B(n_539),
.Y(n_634)
);

INVxp67_ASAP7_75t_L g635 ( 
.A(n_566),
.Y(n_635)
);

INVx4_ASAP7_75t_L g636 ( 
.A(n_586),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_560),
.B(n_539),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_565),
.B(n_515),
.Y(n_638)
);

CKINVDCx20_ASAP7_75t_R g639 ( 
.A(n_570),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_607),
.B(n_546),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_612),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_621),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g644 ( 
.A(n_584),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_588),
.Y(n_645)
);

INVx1_ASAP7_75t_SL g646 ( 
.A(n_571),
.Y(n_646)
);

NOR2xp33_ASAP7_75t_L g647 ( 
.A(n_587),
.B(n_535),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_568),
.Y(n_648)
);

NAND2x1p5_ASAP7_75t_L g649 ( 
.A(n_598),
.B(n_503),
.Y(n_649)
);

AOI22xp33_ASAP7_75t_L g650 ( 
.A1(n_581),
.A2(n_522),
.B1(n_584),
.B2(n_523),
.Y(n_650)
);

CKINVDCx11_ASAP7_75t_R g651 ( 
.A(n_563),
.Y(n_651)
);

INVx5_ASAP7_75t_L g652 ( 
.A(n_567),
.Y(n_652)
);

BUFx2_ASAP7_75t_L g653 ( 
.A(n_571),
.Y(n_653)
);

BUFx4f_ASAP7_75t_L g654 ( 
.A(n_563),
.Y(n_654)
);

AND2x4_ASAP7_75t_L g655 ( 
.A(n_563),
.B(n_503),
.Y(n_655)
);

BUFx12f_ASAP7_75t_L g656 ( 
.A(n_597),
.Y(n_656)
);

AOI22xp5_ASAP7_75t_L g657 ( 
.A1(n_588),
.A2(n_522),
.B1(n_505),
.B2(n_514),
.Y(n_657)
);

BUFx12f_ASAP7_75t_L g658 ( 
.A(n_597),
.Y(n_658)
);

NAND2x1p5_ASAP7_75t_L g659 ( 
.A(n_598),
.B(n_602),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_572),
.Y(n_660)
);

INVx5_ASAP7_75t_L g661 ( 
.A(n_567),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_585),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_596),
.Y(n_663)
);

INVx2_ASAP7_75t_SL g664 ( 
.A(n_597),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_617),
.Y(n_665)
);

BUFx2_ASAP7_75t_L g666 ( 
.A(n_587),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_564),
.B(n_514),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_573),
.Y(n_668)
);

BUFx8_ASAP7_75t_L g669 ( 
.A(n_589),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_589),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_575),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_558),
.B(n_484),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_580),
.Y(n_673)
);

AO21x2_ASAP7_75t_L g674 ( 
.A1(n_610),
.A2(n_519),
.B(n_483),
.Y(n_674)
);

INVx6_ASAP7_75t_L g675 ( 
.A(n_598),
.Y(n_675)
);

BUFx3_ASAP7_75t_L g676 ( 
.A(n_614),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_559),
.Y(n_677)
);

INVx2_ASAP7_75t_SL g678 ( 
.A(n_569),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_611),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_605),
.Y(n_680)
);

INVx4_ASAP7_75t_L g681 ( 
.A(n_602),
.Y(n_681)
);

BUFx12f_ASAP7_75t_L g682 ( 
.A(n_614),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_652),
.Y(n_683)
);

INVx6_ASAP7_75t_L g684 ( 
.A(n_669),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_633),
.B(n_591),
.Y(n_685)
);

NAND2xp33_ASAP7_75t_SL g686 ( 
.A(n_634),
.B(n_590),
.Y(n_686)
);

BUFx2_ASAP7_75t_L g687 ( 
.A(n_641),
.Y(n_687)
);

BUFx3_ASAP7_75t_L g688 ( 
.A(n_631),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_636),
.Y(n_689)
);

CKINVDCx11_ASAP7_75t_R g690 ( 
.A(n_639),
.Y(n_690)
);

CKINVDCx11_ASAP7_75t_R g691 ( 
.A(n_629),
.Y(n_691)
);

INVx4_ASAP7_75t_L g692 ( 
.A(n_636),
.Y(n_692)
);

INVx2_ASAP7_75t_SL g693 ( 
.A(n_654),
.Y(n_693)
);

INVx3_ASAP7_75t_L g694 ( 
.A(n_675),
.Y(n_694)
);

BUFx3_ASAP7_75t_L g695 ( 
.A(n_654),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_651),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_655),
.Y(n_697)
);

INVx1_ASAP7_75t_SL g698 ( 
.A(n_630),
.Y(n_698)
);

INVx1_ASAP7_75t_SL g699 ( 
.A(n_630),
.Y(n_699)
);

INVx11_ASAP7_75t_L g700 ( 
.A(n_669),
.Y(n_700)
);

INVx1_ASAP7_75t_L g701 ( 
.A(n_662),
.Y(n_701)
);

OAI22xp33_ASAP7_75t_SL g702 ( 
.A1(n_657),
.A2(n_646),
.B1(n_680),
.B2(n_592),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_666),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_663),
.Y(n_704)
);

CKINVDCx20_ASAP7_75t_R g705 ( 
.A(n_647),
.Y(n_705)
);

BUFx10_ASAP7_75t_L g706 ( 
.A(n_675),
.Y(n_706)
);

AOI22xp33_ASAP7_75t_L g707 ( 
.A1(n_632),
.A2(n_592),
.B1(n_590),
.B2(n_579),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_673),
.Y(n_708)
);

AOI22xp33_ASAP7_75t_L g709 ( 
.A1(n_632),
.A2(n_599),
.B1(n_609),
.B2(n_582),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_635),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_667),
.B(n_505),
.Y(n_711)
);

INVx4_ASAP7_75t_L g712 ( 
.A(n_675),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_653),
.Y(n_713)
);

AND2x4_ASAP7_75t_L g714 ( 
.A(n_655),
.B(n_561),
.Y(n_714)
);

AOI22xp33_ASAP7_75t_L g715 ( 
.A1(n_650),
.A2(n_599),
.B1(n_609),
.B2(n_526),
.Y(n_715)
);

OAI22xp5_ASAP7_75t_SL g716 ( 
.A1(n_646),
.A2(n_541),
.B1(n_520),
.B2(n_535),
.Y(n_716)
);

INVx1_ASAP7_75t_SL g717 ( 
.A(n_645),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_665),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_677),
.Y(n_719)
);

AOI22xp33_ASAP7_75t_L g720 ( 
.A1(n_650),
.A2(n_599),
.B1(n_609),
.B2(n_507),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_633),
.B(n_494),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_668),
.Y(n_722)
);

INVx6_ASAP7_75t_L g723 ( 
.A(n_656),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_648),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_679),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_660),
.Y(n_726)
);

INVx4_ASAP7_75t_L g727 ( 
.A(n_627),
.Y(n_727)
);

OAI22xp33_ASAP7_75t_R g728 ( 
.A1(n_638),
.A2(n_562),
.B1(n_518),
.B2(n_520),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_671),
.Y(n_729)
);

BUFx3_ASAP7_75t_L g730 ( 
.A(n_658),
.Y(n_730)
);

BUFx3_ASAP7_75t_L g731 ( 
.A(n_627),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_634),
.Y(n_732)
);

AOI22xp33_ASAP7_75t_L g733 ( 
.A1(n_638),
.A2(n_507),
.B1(n_526),
.B2(n_527),
.Y(n_733)
);

INVx4_ASAP7_75t_SL g734 ( 
.A(n_683),
.Y(n_734)
);

AOI22xp33_ASAP7_75t_L g735 ( 
.A1(n_707),
.A2(n_682),
.B1(n_640),
.B2(n_670),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_707),
.A2(n_685),
.B1(n_711),
.B2(n_686),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_716),
.A2(n_678),
.B1(n_676),
.B2(n_640),
.Y(n_737)
);

AOI22xp33_ASAP7_75t_L g738 ( 
.A1(n_702),
.A2(n_533),
.B1(n_530),
.B2(n_616),
.Y(n_738)
);

AOI22xp33_ASAP7_75t_L g739 ( 
.A1(n_728),
.A2(n_533),
.B1(n_530),
.B2(n_618),
.Y(n_739)
);

OAI22xp5_ASAP7_75t_L g740 ( 
.A1(n_721),
.A2(n_635),
.B1(n_577),
.B2(n_644),
.Y(n_740)
);

HB1xp67_ASAP7_75t_L g741 ( 
.A(n_732),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_708),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_708),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_687),
.Y(n_744)
);

BUFx5_ASAP7_75t_L g745 ( 
.A(n_731),
.Y(n_745)
);

OAI22xp5_ASAP7_75t_L g746 ( 
.A1(n_705),
.A2(n_577),
.B1(n_644),
.B2(n_620),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_698),
.B(n_637),
.Y(n_747)
);

HB1xp67_ASAP7_75t_L g748 ( 
.A(n_732),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_699),
.B(n_637),
.Y(n_749)
);

OAI22xp5_ASAP7_75t_L g750 ( 
.A1(n_705),
.A2(n_620),
.B1(n_624),
.B2(n_614),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_690),
.Y(n_751)
);

AOI22xp33_ASAP7_75t_SL g752 ( 
.A1(n_684),
.A2(n_620),
.B1(n_624),
.B2(n_549),
.Y(n_752)
);

OAI222xp33_ASAP7_75t_L g753 ( 
.A1(n_709),
.A2(n_624),
.B1(n_672),
.B2(n_509),
.C1(n_557),
.C2(n_610),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_709),
.A2(n_472),
.B1(n_545),
.B2(n_551),
.Y(n_754)
);

BUFx6f_ASAP7_75t_L g755 ( 
.A(n_683),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_710),
.B(n_549),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_SL g757 ( 
.A1(n_684),
.A2(n_664),
.B1(n_556),
.B2(n_605),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_701),
.Y(n_758)
);

OAI22xp5_ASAP7_75t_L g759 ( 
.A1(n_703),
.A2(n_540),
.B1(n_556),
.B2(n_487),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_704),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_718),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_700),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_725),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_719),
.Y(n_764)
);

INVx1_ASAP7_75t_L g765 ( 
.A(n_722),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_724),
.Y(n_766)
);

AND2x2_ASAP7_75t_L g767 ( 
.A(n_713),
.B(n_540),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_726),
.Y(n_768)
);

AOI22xp33_ASAP7_75t_SL g769 ( 
.A1(n_684),
.A2(n_600),
.B1(n_601),
.B2(n_672),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_706),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_715),
.A2(n_479),
.B1(n_556),
.B2(n_494),
.Y(n_771)
);

AOI22xp33_ASAP7_75t_L g772 ( 
.A1(n_715),
.A2(n_537),
.B1(n_545),
.B2(n_504),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_725),
.Y(n_773)
);

AND2x2_ASAP7_75t_L g774 ( 
.A(n_717),
.B(n_593),
.Y(n_774)
);

AOI22xp33_ASAP7_75t_L g775 ( 
.A1(n_720),
.A2(n_554),
.B1(n_542),
.B2(n_481),
.Y(n_775)
);

BUFx4f_ASAP7_75t_SL g776 ( 
.A(n_688),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_729),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_729),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_733),
.A2(n_554),
.B1(n_697),
.B2(n_481),
.Y(n_779)
);

AOI22xp33_ASAP7_75t_L g780 ( 
.A1(n_733),
.A2(n_481),
.B1(n_500),
.B2(n_619),
.Y(n_780)
);

BUFx12f_ASAP7_75t_L g781 ( 
.A(n_690),
.Y(n_781)
);

BUFx4f_ASAP7_75t_SL g782 ( 
.A(n_695),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_697),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_695),
.A2(n_500),
.B1(n_623),
.B2(n_502),
.Y(n_784)
);

OAI22xp5_ASAP7_75t_SL g785 ( 
.A1(n_696),
.A2(n_555),
.B1(n_552),
.B2(n_649),
.Y(n_785)
);

AOI222xp33_ASAP7_75t_L g786 ( 
.A1(n_730),
.A2(n_479),
.B1(n_476),
.B2(n_604),
.C1(n_484),
.C2(n_502),
.Y(n_786)
);

AOI22xp33_ASAP7_75t_L g787 ( 
.A1(n_750),
.A2(n_723),
.B1(n_714),
.B2(n_730),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_736),
.A2(n_692),
.B1(n_723),
.B2(n_689),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_736),
.A2(n_723),
.B1(n_714),
.B2(n_693),
.Y(n_789)
);

AOI22xp33_ASAP7_75t_L g790 ( 
.A1(n_746),
.A2(n_714),
.B1(n_615),
.B2(n_550),
.Y(n_790)
);

OAI222xp33_ASAP7_75t_L g791 ( 
.A1(n_752),
.A2(n_615),
.B1(n_712),
.B2(n_649),
.C1(n_727),
.C2(n_492),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_SL g792 ( 
.A1(n_740),
.A2(n_683),
.B1(n_661),
.B2(n_652),
.Y(n_792)
);

AOI22xp33_ASAP7_75t_L g793 ( 
.A1(n_752),
.A2(n_550),
.B1(n_543),
.B2(n_544),
.Y(n_793)
);

AOI22xp33_ASAP7_75t_SL g794 ( 
.A1(n_757),
.A2(n_683),
.B1(n_661),
.B2(n_652),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_758),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_766),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_747),
.B(n_731),
.Y(n_797)
);

AND2x2_ASAP7_75t_SL g798 ( 
.A(n_741),
.B(n_712),
.Y(n_798)
);

AOI22xp33_ASAP7_75t_SL g799 ( 
.A1(n_759),
.A2(n_661),
.B1(n_543),
.B2(n_567),
.Y(n_799)
);

BUFx2_ASAP7_75t_L g800 ( 
.A(n_744),
.Y(n_800)
);

AOI22xp33_ASAP7_75t_L g801 ( 
.A1(n_735),
.A2(n_550),
.B1(n_544),
.B2(n_594),
.Y(n_801)
);

OAI22xp5_ASAP7_75t_L g802 ( 
.A1(n_769),
.A2(n_689),
.B1(n_694),
.B2(n_727),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_735),
.A2(n_550),
.B1(n_544),
.B2(n_561),
.Y(n_803)
);

AOI22xp33_ASAP7_75t_L g804 ( 
.A1(n_772),
.A2(n_550),
.B1(n_674),
.B2(n_691),
.Y(n_804)
);

AOI22xp33_ASAP7_75t_L g805 ( 
.A1(n_738),
.A2(n_544),
.B1(n_603),
.B2(n_578),
.Y(n_805)
);

OAI22xp5_ASAP7_75t_L g806 ( 
.A1(n_771),
.A2(n_737),
.B1(n_776),
.B2(n_784),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_749),
.B(n_627),
.Y(n_807)
);

OAI211xp5_ASAP7_75t_L g808 ( 
.A1(n_756),
.A2(n_691),
.B(n_532),
.C(n_548),
.Y(n_808)
);

OAI221xp5_ASAP7_75t_SL g809 ( 
.A1(n_739),
.A2(n_512),
.B1(n_548),
.B2(n_606),
.C(n_603),
.Y(n_809)
);

OA21x2_ASAP7_75t_L g810 ( 
.A1(n_753),
.A2(n_480),
.B(n_622),
.Y(n_810)
);

AOI22xp33_ASAP7_75t_L g811 ( 
.A1(n_754),
.A2(n_772),
.B1(n_786),
.B2(n_774),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_SL g812 ( 
.A1(n_785),
.A2(n_567),
.B1(n_602),
.B2(n_608),
.Y(n_812)
);

OA21x2_ASAP7_75t_L g813 ( 
.A1(n_753),
.A2(n_768),
.B(n_765),
.Y(n_813)
);

AOI22xp33_ASAP7_75t_L g814 ( 
.A1(n_767),
.A2(n_578),
.B1(n_583),
.B2(n_594),
.Y(n_814)
);

OAI221xp5_ASAP7_75t_L g815 ( 
.A1(n_779),
.A2(n_548),
.B1(n_583),
.B2(n_606),
.C(n_681),
.Y(n_815)
);

BUFx2_ASAP7_75t_SL g816 ( 
.A(n_762),
.Y(n_816)
);

AOI221xp5_ASAP7_75t_L g817 ( 
.A1(n_760),
.A2(n_622),
.B1(n_628),
.B2(n_643),
.C(n_642),
.Y(n_817)
);

AOI22xp33_ASAP7_75t_L g818 ( 
.A1(n_775),
.A2(n_674),
.B1(n_608),
.B2(n_681),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_780),
.A2(n_628),
.B1(n_643),
.B2(n_642),
.Y(n_819)
);

AOI22xp33_ASAP7_75t_L g820 ( 
.A1(n_741),
.A2(n_642),
.B1(n_621),
.B2(n_498),
.Y(n_820)
);

AOI22xp33_ASAP7_75t_L g821 ( 
.A1(n_748),
.A2(n_621),
.B1(n_498),
.B2(n_495),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_761),
.B(n_706),
.Y(n_822)
);

AOI22xp33_ASAP7_75t_L g823 ( 
.A1(n_748),
.A2(n_516),
.B1(n_495),
.B2(n_498),
.Y(n_823)
);

NAND3xp33_ASAP7_75t_L g824 ( 
.A(n_783),
.B(n_516),
.C(n_498),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_764),
.B(n_706),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_745),
.B(n_659),
.Y(n_826)
);

AOI221x1_ASAP7_75t_L g827 ( 
.A1(n_770),
.A2(n_516),
.B1(n_498),
.B2(n_495),
.C(n_511),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_742),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_807),
.B(n_745),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_SL g830 ( 
.A(n_798),
.B(n_745),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_798),
.B(n_745),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_800),
.B(n_745),
.Y(n_832)
);

OAI22xp5_ASAP7_75t_L g833 ( 
.A1(n_789),
.A2(n_776),
.B1(n_782),
.B2(n_751),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_795),
.Y(n_834)
);

OAI21xp33_ASAP7_75t_L g835 ( 
.A1(n_808),
.A2(n_770),
.B(n_755),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_797),
.B(n_745),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_787),
.B(n_796),
.Y(n_837)
);

INVx2_ASAP7_75t_L g838 ( 
.A(n_828),
.Y(n_838)
);

NAND3xp33_ASAP7_75t_L g839 ( 
.A(n_817),
.B(n_825),
.C(n_822),
.Y(n_839)
);

OAI21xp5_ASAP7_75t_SL g840 ( 
.A1(n_806),
.A2(n_781),
.B(n_782),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_813),
.B(n_790),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_787),
.B(n_755),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_789),
.B(n_743),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_788),
.B(n_802),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_804),
.B(n_763),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_826),
.B(n_773),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_804),
.B(n_777),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_811),
.A2(n_659),
.B1(n_625),
.B2(n_626),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_SL g849 ( 
.A(n_792),
.B(n_734),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_818),
.B(n_778),
.Y(n_850)
);

AND2x2_ASAP7_75t_L g851 ( 
.A(n_816),
.B(n_734),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_SL g852 ( 
.A1(n_812),
.A2(n_626),
.B(n_625),
.Y(n_852)
);

NAND3xp33_ASAP7_75t_L g853 ( 
.A(n_809),
.B(n_516),
.C(n_310),
.Y(n_853)
);

NAND3xp33_ASAP7_75t_L g854 ( 
.A(n_814),
.B(n_516),
.C(n_310),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_820),
.B(n_819),
.Y(n_855)
);

OAI22xp5_ASAP7_75t_SL g856 ( 
.A1(n_799),
.A2(n_595),
.B1(n_45),
.B2(n_47),
.Y(n_856)
);

OAI221xp5_ASAP7_75t_L g857 ( 
.A1(n_793),
.A2(n_595),
.B1(n_310),
.B2(n_52),
.C(n_54),
.Y(n_857)
);

AND2x2_ASAP7_75t_L g858 ( 
.A(n_810),
.B(n_821),
.Y(n_858)
);

AND2x2_ASAP7_75t_L g859 ( 
.A(n_810),
.B(n_44),
.Y(n_859)
);

OA21x2_ASAP7_75t_L g860 ( 
.A1(n_827),
.A2(n_50),
.B(n_55),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_832),
.B(n_810),
.Y(n_861)
);

NAND4xp75_ASAP7_75t_L g862 ( 
.A(n_849),
.B(n_791),
.C(n_794),
.D(n_803),
.Y(n_862)
);

AND2x2_ASAP7_75t_L g863 ( 
.A(n_834),
.B(n_823),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_836),
.B(n_824),
.Y(n_864)
);

AND2x2_ASAP7_75t_L g865 ( 
.A(n_841),
.B(n_801),
.Y(n_865)
);

OAI211xp5_ASAP7_75t_L g866 ( 
.A1(n_844),
.A2(n_815),
.B(n_805),
.C(n_67),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_841),
.B(n_59),
.Y(n_867)
);

HB1xp67_ASAP7_75t_L g868 ( 
.A(n_829),
.Y(n_868)
);

AND2x2_ASAP7_75t_L g869 ( 
.A(n_858),
.B(n_62),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_L g870 ( 
.A(n_840),
.B(n_68),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_846),
.B(n_69),
.Y(n_871)
);

NAND4xp75_ASAP7_75t_L g872 ( 
.A(n_849),
.B(n_73),
.C(n_74),
.D(n_75),
.Y(n_872)
);

INVx2_ASAP7_75t_L g873 ( 
.A(n_838),
.Y(n_873)
);

NAND3xp33_ASAP7_75t_L g874 ( 
.A(n_839),
.B(n_77),
.C(n_78),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_858),
.B(n_79),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_844),
.B(n_80),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_837),
.B(n_81),
.Y(n_877)
);

XNOR2xp5_ASAP7_75t_L g878 ( 
.A(n_876),
.B(n_833),
.Y(n_878)
);

NOR3xp33_ASAP7_75t_SL g879 ( 
.A(n_870),
.B(n_835),
.C(n_831),
.Y(n_879)
);

OAI31xp33_ASAP7_75t_L g880 ( 
.A1(n_866),
.A2(n_853),
.A3(n_859),
.B(n_856),
.Y(n_880)
);

OR2x2_ASAP7_75t_L g881 ( 
.A(n_868),
.B(n_847),
.Y(n_881)
);

NOR2x1_ASAP7_75t_L g882 ( 
.A(n_864),
.B(n_830),
.Y(n_882)
);

NOR4xp25_ASAP7_75t_L g883 ( 
.A(n_876),
.B(n_859),
.C(n_855),
.D(n_857),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_861),
.B(n_851),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_877),
.Y(n_885)
);

AND2x4_ASAP7_75t_L g886 ( 
.A(n_863),
.B(n_830),
.Y(n_886)
);

NAND4xp75_ASAP7_75t_SL g887 ( 
.A(n_870),
.B(n_860),
.C(n_842),
.D(n_845),
.Y(n_887)
);

XNOR2xp5_ASAP7_75t_L g888 ( 
.A(n_862),
.B(n_831),
.Y(n_888)
);

NOR3xp33_ASAP7_75t_L g889 ( 
.A(n_874),
.B(n_848),
.C(n_854),
.Y(n_889)
);

XNOR2x1_ASAP7_75t_L g890 ( 
.A(n_888),
.B(n_867),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_884),
.B(n_861),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_881),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_886),
.Y(n_893)
);

INVxp67_ASAP7_75t_L g894 ( 
.A(n_882),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_886),
.Y(n_895)
);

XNOR2x1_ASAP7_75t_L g896 ( 
.A(n_885),
.B(n_867),
.Y(n_896)
);

OA22x2_ASAP7_75t_L g897 ( 
.A1(n_892),
.A2(n_878),
.B1(n_865),
.B2(n_869),
.Y(n_897)
);

AOI22xp5_ASAP7_75t_L g898 ( 
.A1(n_890),
.A2(n_883),
.B1(n_865),
.B2(n_889),
.Y(n_898)
);

OA22x2_ASAP7_75t_L g899 ( 
.A1(n_893),
.A2(n_875),
.B1(n_887),
.B2(n_863),
.Y(n_899)
);

AOI22x1_ASAP7_75t_L g900 ( 
.A1(n_894),
.A2(n_875),
.B1(n_880),
.B2(n_879),
.Y(n_900)
);

OA22x2_ASAP7_75t_L g901 ( 
.A1(n_895),
.A2(n_852),
.B1(n_880),
.B2(n_873),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_891),
.B(n_873),
.Y(n_902)
);

OA22x2_ASAP7_75t_L g903 ( 
.A1(n_896),
.A2(n_845),
.B1(n_843),
.B2(n_850),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_898),
.A2(n_872),
.B1(n_860),
.B2(n_871),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_900),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_897),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_902),
.Y(n_907)
);

AOI22xp5_ASAP7_75t_L g908 ( 
.A1(n_904),
.A2(n_901),
.B1(n_903),
.B2(n_899),
.Y(n_908)
);

AOI22xp5_ASAP7_75t_L g909 ( 
.A1(n_904),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_909)
);

AOI221xp5_ASAP7_75t_L g910 ( 
.A1(n_908),
.A2(n_906),
.B1(n_905),
.B2(n_907),
.C(n_95),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_909),
.Y(n_911)
);

OAI21xp5_ASAP7_75t_SL g912 ( 
.A1(n_910),
.A2(n_98),
.B(n_99),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_911),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_913),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_912),
.Y(n_915)
);

NAND4xp25_ASAP7_75t_L g916 ( 
.A(n_914),
.B(n_115),
.C(n_118),
.D(n_122),
.Y(n_916)
);

AND3x1_ASAP7_75t_L g917 ( 
.A(n_915),
.B(n_123),
.C(n_124),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_SL g918 ( 
.A(n_915),
.B(n_128),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_914),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_919),
.Y(n_920)
);

AND2x2_ASAP7_75t_L g921 ( 
.A(n_917),
.B(n_130),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_916),
.Y(n_922)
);

INVxp33_ASAP7_75t_SL g923 ( 
.A(n_918),
.Y(n_923)
);

OAI22xp5_ASAP7_75t_L g924 ( 
.A1(n_920),
.A2(n_139),
.B1(n_140),
.B2(n_141),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_922),
.A2(n_142),
.B1(n_146),
.B2(n_147),
.Y(n_925)
);

HB1xp67_ASAP7_75t_L g926 ( 
.A(n_921),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_923),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_926),
.Y(n_928)
);

AO22x2_ASAP7_75t_L g929 ( 
.A1(n_928),
.A2(n_925),
.B1(n_927),
.B2(n_924),
.Y(n_929)
);

INVx1_ASAP7_75t_L g930 ( 
.A(n_929),
.Y(n_930)
);

AOI22xp5_ASAP7_75t_L g931 ( 
.A1(n_930),
.A2(n_158),
.B1(n_159),
.B2(n_161),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_931),
.Y(n_932)
);

AOI221xp5_ASAP7_75t_L g933 ( 
.A1(n_932),
.A2(n_162),
.B1(n_164),
.B2(n_167),
.C(n_168),
.Y(n_933)
);

AOI211xp5_ASAP7_75t_L g934 ( 
.A1(n_933),
.A2(n_171),
.B(n_173),
.C(n_174),
.Y(n_934)
);


endmodule