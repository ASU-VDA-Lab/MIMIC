module fake_jpeg_7865_n_80 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_80);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx3_ASAP7_75t_L g9 ( 
.A(n_8),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_8),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx10_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

AND2x2_ASAP7_75t_L g18 ( 
.A(n_13),
.B(n_0),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_18),
.B(n_21),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

NOR2xp67_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_10),
.B(n_1),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_23),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_10),
.B(n_1),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_16),
.B1(n_9),
.B2(n_13),
.Y(n_25)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_36),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

AND2x6_ASAP7_75t_L g34 ( 
.A(n_24),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_18),
.Y(n_35)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_29),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_43),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_42),
.Y(n_50)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_44),
.A2(n_27),
.B1(n_28),
.B2(n_26),
.Y(n_45)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_38),
.A2(n_32),
.B1(n_28),
.B2(n_16),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_48),
.B(n_49),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_28),
.B1(n_9),
.B2(n_26),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_42),
.A2(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g54 ( 
.A1(n_51),
.A2(n_52),
.B1(n_50),
.B2(n_40),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_47),
.A2(n_7),
.B(n_6),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_5),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_54),
.B(n_59),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_52),
.B(n_51),
.Y(n_56)
);

XOR2xp5_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_58),
.Y(n_62)
);

MAJx2_ASAP7_75t_L g58 ( 
.A(n_49),
.B(n_19),
.C(n_12),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_46),
.Y(n_59)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_55),
.Y(n_63)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_57),
.A2(n_40),
.B1(n_44),
.B2(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_64),
.A2(n_65),
.B1(n_14),
.B2(n_3),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_57),
.B(n_7),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_62),
.B(n_19),
.C(n_14),
.Y(n_67)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_67),
.A2(n_64),
.B(n_14),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_68),
.B(n_2),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g70 ( 
.A1(n_67),
.A2(n_60),
.B(n_63),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_70),
.B(n_72),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_69),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_74),
.B(n_69),
.C(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_66),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_75),
.B(n_2),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_76),
.A2(n_77),
.B1(n_73),
.B2(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_78),
.B(n_3),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_4),
.Y(n_80)
);


endmodule